module kick_lookup(index, out);
	input logic unsigned [9:0] index;
	output logic signed [23:0] out;
	always_comb begin
		case(index)
			0: out = 0;
			1: out = 0;
			2: out = 77;
			3: out = 914;
			4: out = 1259;
			5: out = 1129;
			6: out = 1227;
			7: out = 1250;
			8: out = 1690;
			9: out = 2049;
			10: out = 2614;
			11: out = 3196;
			12: out = 3209;
			13: out = 2814;
			14: out = 2952;
			15: out = 2987;
			16: out = 3182;
			17: out = 2991;
			18: out = 2665;
			19: out = 2916;
			20: out = 3069;
			21: out = 3236;
			22: out = 3568;
			23: out = 4049;
			24: out = 4561;
			25: out = 5004;
			26: out = 5163;
			27: out = 5576;
			28: out = 6078;
			29: out = 6479;
			30: out = 6577;
			31: out = 6093;
			32: out = 6316;
			33: out = 6766;
			34: out = 7091;
			35: out = 7179;
			36: out = 6881;
			37: out = 7284;
			38: out = 7359;
			39: out = 7263;
			40: out = 6789;
			41: out = 6113;
			42: out = 5706;
			43: out = 5508;
			44: out = 5283;
			45: out = 5504;
			46: out = 5395;
			47: out = 4820;
			48: out = 5057;
			49: out = 5415;
			50: out = 5331;
			51: out = 5240;
			52: out = 5497;
			53: out = 6365;
			54: out = 7033;
			55: out = 7398;
			56: out = 7415;
			57: out = 6813;
			58: out = 7024;
			59: out = 8134;
			60: out = 9756;
			61: out = 11347;
			62: out = 13079;
			63: out = 13755;
			64: out = 14459;
			65: out = 15902;
			66: out = 17206;
			67: out = 18245;
			68: out = 19484;
			69: out = 20343;
			70: out = 22086;
			71: out = 23148;
			72: out = 24088;
			73: out = 24673;
			74: out = 27450;
			75: out = 32241;
			76: out = 32312;
			77: out = 32412;
			78: out = 32277;
			79: out = 32268;
			80: out = 32112;
			81: out = 32109;
			82: out = 32054;
			83: out = 32095;
			84: out = 32061;
			85: out = 32071;
			86: out = 32022;
			87: out = 32007;
			88: out = 31955;
			89: out = 31934;
			90: out = 31899;
			91: out = 31886;
			92: out = 31859;
			93: out = 31846;
			94: out = 31819;
			95: out = 31799;
			96: out = 31768;
			97: out = 31745;
			98: out = 31716;
			99: out = 31697;
			100: out = 31670;
			101: out = 31651;
			102: out = 31629;
			103: out = 31608;
			104: out = 31578;
			105: out = 31561;
			106: out = 31529;
			107: out = 31508;
			108: out = 31474;
			109: out = 31468;
			110: out = 31418;
			111: out = 31448;
			112: out = 31120;
			113: out = 29390;
			114: out = 27954;
			115: out = 26486;
			116: out = 24857;
			117: out = 23719;
			118: out = 23311;
			119: out = 22864;
			120: out = 22038;
			121: out = 20778;
			122: out = 19947;
			123: out = 19314;
			124: out = 18218;
			125: out = 16569;
			126: out = 15098;
			127: out = 13522;
			128: out = 11622;
			129: out = 9757;
			130: out = 8423;
			131: out = 7616;
			132: out = 6324;
			133: out = 4719;
			134: out = 3594;
			135: out = 2124;
			136: out = 696;
			137: out = -1233;
			138: out = -3194;
			139: out = -4759;
			140: out = -6732;
			141: out = -8771;
			142: out = -10236;
			143: out = -11293;
			144: out = -12712;
			145: out = -13700;
			146: out = -14622;
			147: out = -15701;
			148: out = -16357;
			149: out = -16888;
			150: out = -17982;
			151: out = -18931;
			152: out = -20442;
			153: out = -21982;
			154: out = -22929;
			155: out = -23588;
			156: out = -24487;
			157: out = -26078;
			158: out = -26746;
			159: out = -27695;
			160: out = -28912;
			161: out = -30039;
			162: out = -31472;
			163: out = -32488;
			164: out = -32561;
			165: out = -32584;
			166: out = -32568;
			167: out = -32552;
			168: out = -32521;
			169: out = -32502;
			170: out = -32481;
			171: out = -32453;
			172: out = -32432;
			173: out = -32422;
			174: out = -32406;
			175: out = -32378;
			176: out = -32354;
			177: out = -32330;
			178: out = -32309;
			179: out = -32284;
			180: out = -32262;
			181: out = -32239;
			182: out = -32213;
			183: out = -32188;
			184: out = -32161;
			185: out = -32137;
			186: out = -32113;
			187: out = -32087;
			188: out = -32061;
			189: out = -32040;
			190: out = -32014;
			191: out = -31988;
			192: out = -31963;
			193: out = -31934;
			194: out = -31915;
			195: out = -31885;
			196: out = -31859;
			197: out = -31834;
			198: out = -31803;
			199: out = -31780;
			200: out = -31750;
			201: out = -31723;
			202: out = -31688;
			203: out = -31651;
			204: out = -31614;
			205: out = -31593;
			206: out = -31562;
			207: out = -31484;
			208: out = -31410;
			209: out = -31306;
			210: out = -31208;
			211: out = -30225;
			212: out = -28673;
			213: out = -27786;
			214: out = -27365;
			215: out = -27601;
			216: out = -26871;
			217: out = -26122;
			218: out = -25663;
			219: out = -25265;
			220: out = -25403;
			221: out = -25399;
			222: out = -24890;
			223: out = -24273;
			224: out = -23297;
			225: out = -22252;
			226: out = -21821;
			227: out = -20717;
			228: out = -19508;
			229: out = -18571;
			230: out = -17368;
			231: out = -15866;
			232: out = -14095;
			233: out = -12471;
			234: out = -11637;
			235: out = -10356;
			236: out = -9140;
			237: out = -8465;
			238: out = -7235;
			239: out = -5327;
			240: out = -3197;
			241: out = -1314;
			242: out = -18;
			243: out = 1442;
			244: out = 2533;
			245: out = 3724;
			246: out = 4529;
			247: out = 5256;
			248: out = 6175;
			249: out = 6624;
			250: out = 7403;
			251: out = 8586;
			252: out = 10067;
			253: out = 11296;
			254: out = 12911;
			255: out = 14708;
			256: out = 15980;
			257: out = 17581;
			258: out = 19083;
			259: out = 19600;
			260: out = 20281;
			261: out = 21026;
			262: out = 22206;
			263: out = 22879;
			264: out = 23240;
			265: out = 23527;
			266: out = 23929;
			267: out = 24252;
			268: out = 24488;
			269: out = 25015;
			270: out = 25683;
			271: out = 26441;
			272: out = 27362;
			273: out = 28418;
			274: out = 29351;
			275: out = 30164;
			276: out = 31668;
			277: out = 32602;
			278: out = 32522;
			279: out = 32546;
			280: out = 32481;
			281: out = 32480;
			282: out = 32441;
			283: out = 32432;
			284: out = 32396;
			285: out = 32380;
			286: out = 32342;
			287: out = 32326;
			288: out = 32294;
			289: out = 32272;
			290: out = 32243;
			291: out = 32225;
			292: out = 32196;
			293: out = 32178;
			294: out = 32150;
			295: out = 32130;
			296: out = 32101;
			297: out = 32079;
			298: out = 32054;
			299: out = 32030;
			300: out = 31999;
			301: out = 31991;
			302: out = 31399;
			303: out = 30454;
			304: out = 29814;
			305: out = 29212;
			306: out = 28529;
			307: out = 27545;
			308: out = 26983;
			309: out = 26769;
			310: out = 26189;
			311: out = 25787;
			312: out = 25692;
			313: out = 25190;
			314: out = 24878;
			315: out = 24723;
			316: out = 24339;
			317: out = 23942;
			318: out = 23258;
			319: out = 23055;
			320: out = 22692;
			321: out = 22060;
			322: out = 21214;
			323: out = 20405;
			324: out = 19372;
			325: out = 18327;
			326: out = 18001;
			327: out = 18124;
			328: out = 18178;
			329: out = 17829;
			330: out = 16739;
			331: out = 16616;
			332: out = 16173;
			333: out = 15443;
			334: out = 14611;
			335: out = 12840;
			336: out = 11296;
			337: out = 10020;
			338: out = 9240;
			339: out = 8645;
			340: out = 8592;
			341: out = 7623;
			342: out = 6889;
			343: out = 6696;
			344: out = 5284;
			345: out = 3906;
			346: out = 3111;
			347: out = 1958;
			348: out = 1232;
			349: out = -12;
			350: out = -1469;
			351: out = -3460;
			352: out = -4886;
			353: out = -6034;
			354: out = -7059;
			355: out = -8312;
			356: out = -9846;
			357: out = -10606;
			358: out = -11587;
			359: out = -12976;
			360: out = -14380;
			361: out = -15710;
			362: out = -16427;
			363: out = -17070;
			364: out = -18116;
			365: out = -19354;
			366: out = -19721;
			367: out = -20015;
			368: out = -20700;
			369: out = -22087;
			370: out = -22764;
			371: out = -23157;
			372: out = -24121;
			373: out = -24895;
			374: out = -25752;
			375: out = -26109;
			376: out = -26445;
			377: out = -26669;
			378: out = -27551;
			379: out = -28250;
			380: out = -29308;
			381: out = -30791;
			382: out = -31996;
			383: out = -32215;
			384: out = -32199;
			385: out = -32195;
			386: out = -32158;
			387: out = -32125;
			388: out = -32122;
			389: out = -32107;
			390: out = -32062;
			391: out = -32050;
			392: out = -32035;
			393: out = -32031;
			394: out = -32008;
			395: out = -31986;
			396: out = -31955;
			397: out = -31931;
			398: out = -31923;
			399: out = -31909;
			400: out = -31885;
			401: out = -31866;
			402: out = -31851;
			403: out = -31824;
			404: out = -31797;
			405: out = -31762;
			406: out = -31732;
			407: out = -31699;
			408: out = -31661;
			409: out = -31651;
			410: out = -31622;
			411: out = -31596;
			412: out = -31564;
			413: out = -31547;
			414: out = -31493;
			415: out = -31457;
			416: out = -31398;
			417: out = -31326;
			418: out = -31285;
			419: out = -31313;
			420: out = -31144;
			421: out = -30928;
			422: out = -30468;
			423: out = -29738;
			424: out = -28786;
			425: out = -28204;
			426: out = -28043;
			427: out = -27188;
			428: out = -27072;
			429: out = -26828;
			430: out = -26715;
			431: out = -26560;
			432: out = -26226;
			433: out = -26457;
			434: out = -26475;
			435: out = -26519;
			436: out = -26579;
			437: out = -26357;
			438: out = -25668;
			439: out = -24707;
			440: out = -23476;
			441: out = -22629;
			442: out = -22401;
			443: out = -21742;
			444: out = -20624;
			445: out = -20059;
			446: out = -19592;
			447: out = -18833;
			448: out = -17889;
			449: out = -17455;
			450: out = -16861;
			451: out = -16162;
			452: out = -16220;
			453: out = -16225;
			454: out = -15662;
			455: out = -14746;
			456: out = -13886;
			457: out = -13030;
			458: out = -12905;
			459: out = -12495;
			460: out = -11318;
			461: out = -10708;
			462: out = -9819;
			463: out = -9198;
			464: out = -8723;
			465: out = -8037;
			466: out = -7316;
			467: out = -6301;
			468: out = -5202;
			469: out = -4294;
			470: out = -3527;
			471: out = -2914;
			472: out = -1557;
			473: out = -560;
			474: out = 586;
			475: out = 1489;
			476: out = 2459;
			477: out = 3331;
			478: out = 3981;
			479: out = 5039;
			480: out = 5527;
			481: out = 5948;
			482: out = 6281;
			483: out = 7087;
			484: out = 7832;
			485: out = 8640;
			486: out = 9436;
			487: out = 10230;
			488: out = 11282;
			489: out = 12419;
			490: out = 13353;
			491: out = 14083;
			492: out = 14702;
			493: out = 15470;
			494: out = 16350;
			495: out = 17166;
			496: out = 17850;
			497: out = 18021;
			498: out = 18250;
			499: out = 18901;
			500: out = 20041;
			501: out = 21332;
			502: out = 22932;
			503: out = 23898;
			504: out = 24693;
			505: out = 25711;
			506: out = 26368;
			507: out = 26366;
			508: out = 26560;
			509: out = 27468;
			510: out = 27987;
			511: out = 28714;
			512: out = 29029;
			513: out = 29419;
			514: out = 29741;
			515: out = 30041;
			516: out = 30251;
			517: out = 30355;
			518: out = 30675;
			519: out = 31389;
			520: out = 32429;
			521: out = 32765;
			522: out = 32727;
			523: out = 32708;
			524: out = 32679;
			525: out = 32656;
			526: out = 32629;
			527: out = 32603;
			528: out = 32582;
			529: out = 32556;
			530: out = 32529;
			531: out = 32504;
			532: out = 32479;
			533: out = 32453;
			534: out = 32431;
			535: out = 32406;
			536: out = 32383;
			537: out = 32358;
			538: out = 32334;
			539: out = 32307;
			540: out = 32289;
			541: out = 32262;
			542: out = 32238;
			543: out = 32214;
			544: out = 32189;
			545: out = 32157;
			546: out = 32141;
			547: out = 32110;
			548: out = 32098;
			549: out = 32058;
			550: out = 32064;
			551: out = 31906;
			552: out = 31343;
			553: out = 30948;
			554: out = 29988;
			555: out = 29410;
			556: out = 28658;
			557: out = 28195;
			558: out = 27623;
			559: out = 27114;
			560: out = 26841;
			561: out = 26308;
			562: out = 25907;
			563: out = 25774;
			564: out = 25576;
			565: out = 25416;
			566: out = 25355;
			567: out = 24836;
			568: out = 24311;
			569: out = 24102;
			570: out = 23805;
			571: out = 23119;
			572: out = 22031;
			573: out = 21377;
			574: out = 20845;
			575: out = 20254;
			576: out = 19618;
			577: out = 19263;
			578: out = 19133;
			579: out = 18831;
			580: out = 18304;
			581: out = 17650;
			582: out = 17222;
			583: out = 16948;
			584: out = 15896;
			585: out = 14876;
			586: out = 14297;
			587: out = 13519;
			588: out = 12664;
			589: out = 12206;
			590: out = 12004;
			591: out = 11771;
			592: out = 11362;
			593: out = 10584;
			594: out = 10054;
			595: out = 9968;
			596: out = 9401;
			597: out = 8888;
			598: out = 8339;
			599: out = 7352;
			600: out = 6280;
			601: out = 5744;
			602: out = 5379;
			603: out = 4925;
			604: out = 4229;
			605: out = 3485;
			606: out = 2493;
			607: out = 1716;
			608: out = 1229;
			609: out = 1046;
			610: out = 566;
			611: out = -293;
			612: out = -1329;
			613: out = -2360;
			614: out = -3338;
			615: out = -4325;
			616: out = -4862;
			617: out = -5642;
			618: out = -6585;
			619: out = -7524;
			620: out = -8205;
			621: out = -9011;
			622: out = -10146;
			623: out = -11061;
			624: out = -12193;
			625: out = -13149;
			626: out = -13981;
			627: out = -14828;
			628: out = -15226;
			629: out = -16109;
			630: out = -17018;
			631: out = -17698;
			632: out = -18221;
			633: out = -18755;
			634: out = -19289;
			635: out = -20043;
			636: out = -20249;
			637: out = -20475;
			638: out = -20972;
			639: out = -21693;
			640: out = -22653;
			641: out = -23529;
			642: out = -24197;
			643: out = -24727;
			644: out = -25328;
			645: out = -25912;
			646: out = -26254;
			647: out = -26609;
			648: out = -26945;
			649: out = -27428;
			650: out = -27747;
			651: out = -28054;
			652: out = -28369;
			653: out = -28653;
			654: out = -28716;
			655: out = -28853;
			656: out = -29324;
			657: out = -29235;
			658: out = -29574;
			659: out = -30446;
			660: out = -30874;
			661: out = -30487;
			662: out = -30100;
			663: out = -29728;
			664: out = -29739;
			665: out = -30414;
			666: out = -30745;
			667: out = -30390;
			668: out = -30481;
			669: out = -30721;
			670: out = -31424;
			671: out = -31716;
			672: out = -31698;
			673: out = -31757;
			674: out = -31739;
			675: out = -31718;
			676: out = -31655;
			677: out = -31597;
			678: out = -31490;
			679: out = -31399;
			680: out = -31388;
			681: out = -31371;
			682: out = -31373;
			683: out = -31405;
			684: out = -31363;
			685: out = -31225;
			686: out = -31144;
			687: out = -31035;
			688: out = -30607;
			689: out = -30372;
			690: out = -30081;
			691: out = -29283;
			692: out = -28871;
			693: out = -28677;
			694: out = -28202;
			695: out = -27635;
			696: out = -27226;
			697: out = -26738;
			698: out = -26596;
			699: out = -26748;
			700: out = -26401;
			701: out = -26085;
			702: out = -25731;
			703: out = -25361;
			704: out = -25104;
			705: out = -24668;
			706: out = -24493;
			707: out = -24423;
			708: out = -24681;
			709: out = -24488;
			710: out = -24275;
			711: out = -23992;
			712: out = -23898;
			713: out = -23727;
			714: out = -23603;
			715: out = -23452;
			716: out = -23277;
			717: out = -22639;
			718: out = -22177;
			719: out = -21911;
			720: out = -21378;
			721: out = -20832;
			722: out = -20550;
			723: out = -19921;
			724: out = -18943;
			725: out = -18067;
			726: out = -17361;
			727: out = -16990;
			728: out = -16700;
			729: out = -16289;
			730: out = -15849;
			731: out = -15610;
			732: out = -15422;
			733: out = -14997;
			734: out = -14755;
			735: out = -14767;
			736: out = -14646;
			737: out = -14232;
			738: out = -13792;
			739: out = -13219;
			740: out = -12879;
			741: out = -11952;
			742: out = -11246;
			743: out = -11118;
			744: out = -10507;
			745: out = -10319;
			746: out = -10445;
			747: out = -10184;
			748: out = -9526;
			749: out = -9003;
			750: out = -8194;
			751: out = -7508;
			752: out = -7139;
			753: out = -6767;
			754: out = -6300;
			755: out = -6061;
			756: out = -5638;
			757: out = -5355;
			758: out = -5460;
			759: out = -5059;
			760: out = -4659;
			761: out = -4098;
			762: out = -3402;
			763: out = -2655;
			764: out = -1993;
			765: out = -1226;
			766: out = -369;
			767: out = 333;
			768: out = 823;
			769: out = 1287;
			770: out = 1442;
			771: out = 1959;
			772: out = 2450;
			773: out = 2734;
			774: out = 3319;
			775: out = 4099;
			776: out = 4885;
			777: out = 5557;
			778: out = 6241;
			779: out = 6776;
			780: out = 7214;
			781: out = 8090;
			782: out = 8636;
			783: out = 9118;
			784: out = 9390;
			785: out = 10030;
			786: out = 10799;
			787: out = 11010;
			788: out = 11307;
			789: out = 11520;
			790: out = 12008;
			791: out = 12518;
			792: out = 13037;
			793: out = 13498;
			794: out = 13662;
			795: out = 13998;
			796: out = 14326;
			797: out = 14887;
			798: out = 15338;
			799: out = 15588;
			800: out = 15761;
			801: out = 16394;
			802: out = 17143;
			803: out = 17807;
			804: out = 18576;
			805: out = 18847;
			806: out = 19023;
			807: out = 19707;
			808: out = 20391;
			809: out = 21177;
			810: out = 22042;
			811: out = 22492;
			812: out = 22512;
			813: out = 22971;
			814: out = 23782;
			815: out = 24125;
			816: out = 24664;
			817: out = 24635;
			818: out = 24695;
			819: out = 25024;
			820: out = 25025;
			821: out = 25167;
			822: out = 25381;
			823: out = 25804;
			824: out = 26348;
			825: out = 26701;
			826: out = 26971;
			827: out = 27296;
			828: out = 27576;
			829: out = 27592;
			830: out = 27743;
			831: out = 28109;
			832: out = 28649;
			833: out = 29026;
			834: out = 29415;
			835: out = 29805;
			836: out = 30042;
			837: out = 30348;
			838: out = 30713;
			839: out = 31018;
			840: out = 31368;
			841: out = 31434;
			842: out = 31519;
			843: out = 31637;
			844: out = 31613;
			845: out = 31516;
			846: out = 31428;
			847: out = 31218;
			848: out = 31104;
			849: out = 30775;
			850: out = 30596;
			851: out = 30468;
			852: out = 30282;
			853: out = 30323;
			854: out = 30300;
			855: out = 29982;
			856: out = 29682;
			857: out = 29525;
			858: out = 29623;
			859: out = 29468;
			860: out = 29331;
			861: out = 29250;
			862: out = 28969;
			863: out = 28639;
			864: out = 28403;
			865: out = 28333;
			866: out = 28027;
			867: out = 27628;
			868: out = 27032;
			869: out = 26803;
			870: out = 26587;
			871: out = 26346;
			872: out = 25982;
			873: out = 25603;
			874: out = 25471;
			875: out = 25119;
			876: out = 24680;
			877: out = 24248;
			878: out = 24068;
			879: out = 24002;
			880: out = 23742;
			881: out = 23201;
			882: out = 22588;
			883: out = 22254;
			884: out = 21842;
			885: out = 21634;
			886: out = 21308;
			887: out = 21048;
			888: out = 20849;
			889: out = 20319;
			890: out = 19942;
			891: out = 19440;
			892: out = 19003;
			893: out = 18662;
			894: out = 18324;
			895: out = 18072;
			896: out = 17571;
			897: out = 16972;
			898: out = 16551;
			899: out = 16071;
			900: out = 15591;
			901: out = 15316;
			902: out = 15105;
			903: out = 14645;
			904: out = 14335;
			905: out = 14033;
			906: out = 13766;
			907: out = 13457;
			908: out = 13101;
			909: out = 12541;
			910: out = 12196;
			911: out = 12032;
			912: out = 11828;
			913: out = 11535;
			914: out = 11243;
			915: out = 10772;
			916: out = 10187;
			917: out = 9875;
			918: out = 9915;
			919: out = 9933;
			920: out = 9865;
			921: out = 9708;
			922: out = 9141;
			923: out = 8632;
			924: out = 8369;
			925: out = 8362;
			926: out = 8396;
			927: out = 8115;
			928: out = 7566;
			929: out = 6960;
			930: out = 6665;
			931: out = 6551;
			932: out = 6482;
			933: out = 6134;
			934: out = 5464;
			935: out = 5001;
			936: out = 4651;
			937: out = 4290;
			938: out = 4071;
			939: out = 3636;
			940: out = 2968;
			941: out = 2356;
			942: out = 1744;
			943: out = 1406;
			944: out = 1087;
			945: out = 682;
			946: out = 226;
			947: out = -469;
			948: out = -1187;
			949: out = -1824;
			950: out = -2273;
			951: out = -2923;
			952: out = -3633;
			953: out = -4227;
			954: out = -4680;
			955: out = -5216;
			956: out = -5880;
			957: out = -6618;
			958: out = -7338;
			959: out = -7979;
			960: out = -8893;
			961: out = -9843;
			962: out = -10517;
			963: out = -11145;
			964: out = -11778;
			965: out = -12372;
			966: out = -12800;
			967: out = -13278;
			968: out = -13863;
			969: out = -14344;
			970: out = -14876;
			971: out = -15414;
			972: out = -15936;
			973: out = -16256;
			974: out = -16683;
			975: out = -17102;
			976: out = -17568;
			977: out = -17957;
			978: out = -18295;
			979: out = -18734;
			980: out = -19162;
			981: out = -19621;
			982: out = -20186;
			983: out = -20561;
			984: out = -20687;
			985: out = -20738;
			986: out = -20883;
			987: out = -21362;
			988: out = -21615;
			989: out = -21650;
			990: out = -21984;
			991: out = -22215;
			992: out = -22504;
			993: out = -22855;
			994: out = -23067;
			995: out = -23187;
			996: out = -23498;
			997: out = -23698;
			998: out = -23763;
			999: out = -24143;
			1000: out = -24208;
			1001: out = -24501;
			1002: out = -24738;
			1003: out = -24954;
			1004: out = -25423;
			1005: out = -25830;
			1006: out = -26164;
			1007: out = -26499;
			1008: out = -26753;
			1009: out = -26990;
			1010: out = -27172;
			1011: out = -27159;
			1012: out = -27244;
			1013: out = -27348;
			1014: out = -27312;
			1015: out = -27292;
			1016: out = -27397;
			1017: out = -27420;
			1018: out = -27438;
			1019: out = -27719;
			1020: out = -28007;
			1021: out = -27969;
			1022: out = -27875;
			1023: out = -27989;
			1024: out = -27981;
			1025: out = -27909;
			1026: out = -28231;
			1027: out = -28311;
			1028: out = -28311;
			1029: out = -28245;
			1030: out = -28281;
			1031: out = -28444;
			1032: out = -28484;
			1033: out = -28619;
			1034: out = -28841;
			1035: out = -28880;
			1036: out = -28803;
			1037: out = -28646;
			1038: out = -28373;
			1039: out = -28358;
			1040: out = -28503;
			1041: out = -28196;
			1042: out = -27942;
			1043: out = -27802;
			1044: out = -27687;
			1045: out = -27532;
			1046: out = -27271;
			1047: out = -27243;
			1048: out = -27119;
			1049: out = -27036;
			1050: out = -26781;
			1051: out = -26369;
			1052: out = -26085;
			1053: out = -25717;
			1054: out = -25568;
			1055: out = -25429;
			1056: out = -25220;
			1057: out = -25067;
			1058: out = -24942;
			1059: out = -24690;
			1060: out = -24537;
			1061: out = -24203;
			1062: out = -23887;
			1063: out = -23645;
			1064: out = -23428;
			1065: out = -23283;
			1066: out = -22940;
			1067: out = -22538;
			1068: out = -22071;
			1069: out = -21565;
			1070: out = -21082;
			1071: out = -20823;
			1072: out = -20494;
			1073: out = -20114;
			1074: out = -19904;
			1075: out = -19772;
			1076: out = -19640;
			1077: out = -19374;
			1078: out = -18950;
			1079: out = -18659;
			1080: out = -18451;
			1081: out = -18410;
			1082: out = -18216;
			1083: out = -18113;
			1084: out = -18045;
			1085: out = -17918;
			1086: out = -17719;
			1087: out = -17458;
			1088: out = -17257;
			1089: out = -17058;
			1090: out = -16706;
			1091: out = -16407;
			1092: out = -16254;
			1093: out = -16080;
			1094: out = -15846;
			1095: out = -15641;
			1096: out = -15511;
			1097: out = -15214;
			1098: out = -14778;
			1099: out = -14493;
			1100: out = -14245;
			1101: out = -14011;
			1102: out = -13546;
			1103: out = -13063;
			1104: out = -12607;
			1105: out = -12210;
			1106: out = -11808;
			1107: out = -11433;
			1108: out = -11144;
			1109: out = -10849;
			1110: out = -10480;
			1111: out = -10241;
			1112: out = -10027;
			1113: out = -9795;
			1114: out = -9388;
			1115: out = -9068;
			1116: out = -8818;
			1117: out = -8649;
			1118: out = -8576;
			1119: out = -8334;
			1120: out = -7969;
			1121: out = -7744;
			1122: out = -7445;
			1123: out = -7099;
			1124: out = -6882;
			1125: out = -6630;
			1126: out = -6172;
			1127: out = -6098;
			1128: out = -5890;
			1129: out = -5650;
			1130: out = -5562;
			1131: out = -5492;
			1132: out = -5379;
			1133: out = -5092;
			1134: out = -4862;
			1135: out = -4705;
			1136: out = -4481;
			1137: out = -4328;
			1138: out = -4063;
			1139: out = -3754;
			1140: out = -3386;
			1141: out = -3046;
			1142: out = -2766;
			1143: out = -2506;
			1144: out = -2151;
			1145: out = -1745;
			1146: out = -1439;
			1147: out = -1045;
			1148: out = -756;
			1149: out = -384;
			1150: out = 49;
			1151: out = 472;
			1152: out = 798;
			1153: out = 1135;
			1154: out = 1444;
			1155: out = 1737;
			1156: out = 1939;
			1157: out = 2054;
			1158: out = 2368;
			1159: out = 2765;
			1160: out = 3190;
			1161: out = 3667;
			1162: out = 4246;
			1163: out = 4738;
			1164: out = 5202;
			1165: out = 5686;
			1166: out = 6242;
			1167: out = 6492;
			1168: out = 6834;
			1169: out = 7362;
			1170: out = 7729;
			1171: out = 8039;
			1172: out = 8468;
			1173: out = 8998;
			1174: out = 9319;
			1175: out = 9661;
			1176: out = 10126;
			1177: out = 10420;
			1178: out = 10758;
			1179: out = 11080;
			1180: out = 11344;
			1181: out = 11745;
			1182: out = 11950;
			1183: out = 12118;
			1184: out = 12446;
			1185: out = 12761;
			1186: out = 13122;
			1187: out = 13497;
			1188: out = 13878;
			1189: out = 14356;
			1190: out = 14686;
			1191: out = 14914;
			1192: out = 15129;
			1193: out = 15352;
			1194: out = 15625;
			1195: out = 15871;
			1196: out = 16275;
			1197: out = 16597;
			1198: out = 16853;
			1199: out = 17059;
			1200: out = 17468;
			1201: out = 17771;
			1202: out = 17968;
			1203: out = 18142;
			1204: out = 18380;
			1205: out = 18703;
			1206: out = 18996;
			1207: out = 19282;
			1208: out = 19446;
			1209: out = 19749;
			1210: out = 19976;
			1211: out = 20165;
			1212: out = 20357;
			1213: out = 20509;
			1214: out = 20751;
			1215: out = 20981;
			1216: out = 21237;
			1217: out = 21462;
			1218: out = 21772;
			1219: out = 22051;
			1220: out = 22175;
			1221: out = 22333;
			1222: out = 22572;
			1223: out = 22899;
			1224: out = 23211;
			1225: out = 23484;
			1226: out = 23573;
			1227: out = 23721;
			1228: out = 24050;
			1229: out = 24360;
			1230: out = 24655;
			1231: out = 24827;
			1232: out = 24948;
			1233: out = 25028;
			1234: out = 25196;
			1235: out = 25324;
			1236: out = 25549;
			1237: out = 25809;
			1238: out = 25987;
			1239: out = 26161;
			1240: out = 26295;
			1241: out = 26314;
			1242: out = 26410;
			1243: out = 26659;
			1244: out = 26758;
			1245: out = 26856;
			1246: out = 26951;
			1247: out = 27058;
			1248: out = 27155;
			1249: out = 27310;
			1250: out = 27493;
			1251: out = 27685;
			1252: out = 27872;
			1253: out = 27896;
			1254: out = 27831;
			1255: out = 27850;
			1256: out = 27872;
			1257: out = 27910;
			1258: out = 27892;
			1259: out = 27739;
			1260: out = 27597;
			1261: out = 27603;
			1262: out = 27576;
			1263: out = 27515;
			1264: out = 27329;
			1265: out = 27114;
			1266: out = 26974;
			1267: out = 26763;
			1268: out = 26517;
			1269: out = 26360;
			1270: out = 26181;
			1271: out = 26024;
			1272: out = 25912;
			1273: out = 25762;
			1274: out = 25540;
			1275: out = 25325;
			1276: out = 25244;
			1277: out = 25065;
			1278: out = 24772;
			1279: out = 24512;
			1280: out = 24352;
			1281: out = 24163;
			1282: out = 24059;
			1283: out = 23964;
			1284: out = 23808;
			1285: out = 23628;
			1286: out = 23400;
			1287: out = 23145;
			1288: out = 22833;
			1289: out = 22583;
			1290: out = 22345;
			1291: out = 22094;
			1292: out = 21735;
			1293: out = 21402;
			1294: out = 21182;
			1295: out = 20949;
			1296: out = 20700;
			1297: out = 20475;
			1298: out = 20219;
			1299: out = 19999;
			1300: out = 19807;
			1301: out = 19605;
			1302: out = 19357;
			1303: out = 19068;
			1304: out = 18822;
			1305: out = 18492;
			1306: out = 18160;
			1307: out = 17926;
			1308: out = 17716;
			1309: out = 17497;
			1310: out = 17353;
			1311: out = 17193;
			1312: out = 17008;
			1313: out = 16831;
			1314: out = 16666;
			1315: out = 16409;
			1316: out = 16102;
			1317: out = 15841;
			1318: out = 15626;
			1319: out = 15476;
			1320: out = 15304;
			1321: out = 15069;
			1322: out = 14770;
			1323: out = 14554;
			1324: out = 14353;
			1325: out = 14103;
			1326: out = 13828;
			1327: out = 13553;
			1328: out = 13357;
			1329: out = 13193;
			1330: out = 12994;
			1331: out = 12788;
			1332: out = 12489;
			1333: out = 12222;
			1334: out = 11914;
			1335: out = 11572;
			1336: out = 11267;
			1337: out = 10960;
			1338: out = 10619;
			1339: out = 10344;
			1340: out = 10087;
			1341: out = 9782;
			1342: out = 9495;
			1343: out = 9226;
			1344: out = 9014;
			1345: out = 8812;
			1346: out = 8625;
			1347: out = 8373;
			1348: out = 8121;
			1349: out = 7899;
			1350: out = 7692;
			1351: out = 7522;
			1352: out = 7304;
			1353: out = 7131;
			1354: out = 6862;
			1355: out = 6573;
			1356: out = 6392;
			1357: out = 6192;
			1358: out = 5949;
			1359: out = 5748;
			1360: out = 5519;
			1361: out = 5199;
			1362: out = 4965;
			1363: out = 4758;
			1364: out = 4613;
			1365: out = 4442;
			1366: out = 4139;
			1367: out = 3862;
			1368: out = 3607;
			1369: out = 3376;
			1370: out = 3179;
			1371: out = 3034;
			1372: out = 2885;
			1373: out = 2683;
			1374: out = 2393;
			1375: out = 2119;
			1376: out = 1863;
			1377: out = 1593;
			1378: out = 1330;
			1379: out = 1134;
			1380: out = 990;
			1381: out = 826;
			1382: out = 631;
			1383: out = 391;
			1384: out = 73;
			1385: out = -238;
			1386: out = -487;
			1387: out = -705;
			1388: out = -984;
			1389: out = -1283;
			1390: out = -1522;
			1391: out = -1711;
			1392: out = -1946;
			1393: out = -2161;
			1394: out = -2450;
			1395: out = -2871;
			1396: out = -3217;
			1397: out = -3528;
			1398: out = -3892;
			1399: out = -4250;
			1400: out = -4602;
			1401: out = -4911;
			1402: out = -5163;
			1403: out = -5470;
			1404: out = -5868;
			1405: out = -6294;
			1406: out = -6554;
			1407: out = -6848;
			1408: out = -7205;
			1409: out = -7622;
			1410: out = -8074;
			1411: out = -8481;
			1412: out = -8906;
			1413: out = -9390;
			1414: out = -9781;
			1415: out = -10109;
			1416: out = -10492;
			1417: out = -10835;
			1418: out = -11197;
			1419: out = -11599;
			1420: out = -12017;
			1421: out = -12367;
			1422: out = -12644;
			1423: out = -12908;
			1424: out = -13184;
			1425: out = -13534;
			1426: out = -13886;
			1427: out = -14179;
			1428: out = -14464;
			1429: out = -14797;
			1430: out = -15124;
			1431: out = -15477;
			1432: out = -15818;
			1433: out = -16123;
			1434: out = -16355;
			1435: out = -16588;
			1436: out = -16855;
			1437: out = -17090;
			1438: out = -17357;
			1439: out = -17602;
			1440: out = -17874;
			1441: out = -18172;
			1442: out = -18437;
			1443: out = -18635;
			1444: out = -18870;
			1445: out = -19112;
			1446: out = -19249;
			1447: out = -19412;
			1448: out = -19598;
			1449: out = -19784;
			1450: out = -19992;
			1451: out = -20174;
			1452: out = -20312;
			1453: out = -20510;
			1454: out = -20759;
			1455: out = -20971;
			1456: out = -21078;
			1457: out = -21188;
			1458: out = -21361;
			1459: out = -21573;
			1460: out = -21737;
			1461: out = -21861;
			1462: out = -22040;
			1463: out = -22189;
			1464: out = -22297;
			1465: out = -22465;
			1466: out = -22598;
			1467: out = -22692;
			1468: out = -22824;
			1469: out = -22939;
			1470: out = -23058;
			1471: out = -23113;
			1472: out = -23162;
			1473: out = -23227;
			1474: out = -23292;
			1475: out = -23372;
			1476: out = -23468;
			1477: out = -23541;
			1478: out = -23539;
			1479: out = -23558;
			1480: out = -23589;
			1481: out = -23652;
			1482: out = -23751;
			1483: out = -23843;
			1484: out = -23866;
			1485: out = -23894;
			1486: out = -23913;
			1487: out = -23960;
			1488: out = -24034;
			1489: out = -24063;
			1490: out = -24103;
			1491: out = -24171;
			1492: out = -24191;
			1493: out = -24247;
			1494: out = -24300;
			1495: out = -24318;
			1496: out = -24289;
			1497: out = -24190;
			1498: out = -24237;
			1499: out = -24292;
			1500: out = -24291;
			1501: out = -24379;
			1502: out = -24481;
			1503: out = -24531;
			1504: out = -24499;
			1505: out = -24441;
			1506: out = -24426;
			1507: out = -24461;
			1508: out = -24464;
			1509: out = -24462;
			1510: out = -24521;
			1511: out = -24593;
			1512: out = -24609;
			1513: out = -24579;
			1514: out = -24533;
			1515: out = -24462;
			1516: out = -24375;
			1517: out = -24344;
			1518: out = -24335;
			1519: out = -24236;
			1520: out = -24087;
			1521: out = -23941;
			1522: out = -23826;
			1523: out = -23740;
			1524: out = -23621;
			1525: out = -23479;
			1526: out = -23351;
			1527: out = -23198;
			1528: out = -23045;
			1529: out = -22961;
			1530: out = -22858;
			1531: out = -22718;
			1532: out = -22545;
			1533: out = -22366;
			1534: out = -22189;
			1535: out = -22009;
			1536: out = -21847;
			1537: out = -21676;
			1538: out = -21461;
			1539: out = -21266;
			1540: out = -21100;
			1541: out = -20922;
			1542: out = -20727;
			1543: out = -20513;
			1544: out = -20299;
			1545: out = -20048;
			1546: out = -19820;
			1547: out = -19554;
			1548: out = -19313;
			1549: out = -19113;
			1550: out = -18925;
			1551: out = -18740;
			1552: out = -18485;
			1553: out = -18201;
			1554: out = -17941;
			1555: out = -17722;
			1556: out = -17507;
			1557: out = -17303;
			1558: out = -17086;
			1559: out = -16856;
			1560: out = -16648;
			1561: out = -16458;
			1562: out = -16279;
			1563: out = -16080;
			1564: out = -15843;
			1565: out = -15618;
			1566: out = -15413;
			1567: out = -15264;
			1568: out = -15127;
			1569: out = -14942;
			1570: out = -14747;
			1571: out = -14550;
			1572: out = -14376;
			1573: out = -14183;
			1574: out = -13966;
			1575: out = -13763;
			1576: out = -13567;
			1577: out = -13370;
			1578: out = -13235;
			1579: out = -13090;
			1580: out = -12911;
			1581: out = -12761;
			1582: out = -12596;
			1583: out = -12417;
			1584: out = -12230;
			1585: out = -12057;
			1586: out = -11899;
			1587: out = -11755;
			1588: out = -11609;
			1589: out = -11479;
			1590: out = -11346;
			1591: out = -11189;
			1592: out = -10994;
			1593: out = -10775;
			1594: out = -10608;
			1595: out = -10458;
			1596: out = -10296;
			1597: out = -10138;
			1598: out = -9969;
			1599: out = -9745;
			1600: out = -9520;
			1601: out = -9286;
			1602: out = -9053;
			1603: out = -8841;
			1604: out = -8619;
			1605: out = -8387;
			1606: out = -8160;
			1607: out = -7966;
			1608: out = -7772;
			1609: out = -7551;
			1610: out = -7319;
			1611: out = -7107;
			1612: out = -6936;
			1613: out = -6766;
			1614: out = -6570;
			1615: out = -6376;
			1616: out = -6187;
			1617: out = -6000;
			1618: out = -5813;
			1619: out = -5665;
			1620: out = -5521;
			1621: out = -5351;
			1622: out = -5175;
			1623: out = -4987;
			1624: out = -4821;
			1625: out = -4644;
			1626: out = -4454;
			1627: out = -4286;
			1628: out = -4140;
			1629: out = -3997;
			1630: out = -3829;
			1631: out = -3655;
			1632: out = -3472;
			1633: out = -3309;
			1634: out = -3137;
			1635: out = -2956;
			1636: out = -2807;
			1637: out = -2624;
			1638: out = -2407;
			1639: out = -2208;
			1640: out = -2043;
			1641: out = -1882;
			1642: out = -1709;
			1643: out = -1559;
			1644: out = -1399;
			1645: out = -1223;
			1646: out = -1063;
			1647: out = -920;
			1648: out = -760;
			1649: out = -611;
			1650: out = -458;
			1651: out = -288;
			1652: out = -93;
			1653: out = 107;
			1654: out = 280;
			1655: out = 420;
			1656: out = 575;
			1657: out = 752;
			1658: out = 945;
			1659: out = 1135;
			1660: out = 1268;
			1661: out = 1395;
			1662: out = 1565;
			1663: out = 1761;
			1664: out = 1960;
			1665: out = 2170;
			1666: out = 2379;
			1667: out = 2609;
			1668: out = 2838;
			1669: out = 3049;
			1670: out = 3269;
			1671: out = 3482;
			1672: out = 3704;
			1673: out = 3934;
			1674: out = 4180;
			1675: out = 4436;
			1676: out = 4681;
			1677: out = 4929;
			1678: out = 5176;
			1679: out = 5418;
			1680: out = 5665;
			1681: out = 5929;
			1682: out = 6203;
			1683: out = 6505;
			1684: out = 6749;
			1685: out = 6994;
			1686: out = 7263;
			1687: out = 7539;
			1688: out = 7802;
			1689: out = 8031;
			1690: out = 8248;
			1691: out = 8481;
			1692: out = 8725;
			1693: out = 8974;
			1694: out = 9211;
			1695: out = 9463;
			1696: out = 9704;
			1697: out = 9917;
			1698: out = 10171;
			1699: out = 10396;
			1700: out = 10601;
			1701: out = 10819;
			1702: out = 11065;
			1703: out = 11298;
			1704: out = 11528;
			1705: out = 11729;
			1706: out = 11926;
			1707: out = 12128;
			1708: out = 12322;
			1709: out = 12506;
			1710: out = 12705;
			1711: out = 12907;
			1712: out = 13094;
			1713: out = 13302;
			1714: out = 13495;
			1715: out = 13704;
			1716: out = 13899;
			1717: out = 14094;
			1718: out = 14295;
			1719: out = 14498;
			1720: out = 14695;
			1721: out = 14882;
			1722: out = 15039;
			1723: out = 15207;
			1724: out = 15412;
			1725: out = 15619;
			1726: out = 15813;
			1727: out = 15960;
			1728: out = 16103;
			1729: out = 16261;
			1730: out = 16418;
			1731: out = 16581;
			1732: out = 16734;
			1733: out = 16860;
			1734: out = 16999;
			1735: out = 17152;
			1736: out = 17292;
			1737: out = 17436;
			1738: out = 17585;
			1739: out = 17727;
			1740: out = 17852;
			1741: out = 17995;
			1742: out = 18107;
			1743: out = 18224;
			1744: out = 18367;
			1745: out = 18510;
			1746: out = 18632;
			1747: out = 18751;
			1748: out = 18887;
			1749: out = 19018;
			1750: out = 19125;
			1751: out = 19245;
			1752: out = 19365;
			1753: out = 19483;
			1754: out = 19611;
			1755: out = 19735;
			1756: out = 19878;
			1757: out = 19987;
			1758: out = 20127;
			1759: out = 20241;
			1760: out = 20370;
			1761: out = 20482;
			1762: out = 20582;
			1763: out = 20676;
			1764: out = 20766;
			1765: out = 20875;
			1766: out = 20976;
			1767: out = 21076;
			1768: out = 21191;
			1769: out = 21280;
			1770: out = 21368;
			1771: out = 21475;
			1772: out = 21569;
			1773: out = 21662;
			1774: out = 21730;
			1775: out = 21818;
			1776: out = 21901;
			1777: out = 22000;
			1778: out = 22079;
			1779: out = 22174;
			1780: out = 22242;
			1781: out = 22327;
			1782: out = 22410;
			1783: out = 22488;
			1784: out = 22569;
			1785: out = 22639;
			1786: out = 22715;
			1787: out = 22778;
			1788: out = 22868;
			1789: out = 22950;
			1790: out = 23010;
			1791: out = 23059;
			1792: out = 23119;
			1793: out = 23166;
			1794: out = 23202;
			1795: out = 23233;
			1796: out = 23271;
			1797: out = 23307;
			1798: out = 23321;
			1799: out = 23350;
			1800: out = 23334;
			1801: out = 23336;
			1802: out = 23326;
			1803: out = 23328;
			1804: out = 23278;
			1805: out = 23239;
			1806: out = 23165;
			1807: out = 23084;
			1808: out = 23041;
			1809: out = 22938;
			1810: out = 22840;
			1811: out = 22766;
			1812: out = 22678;
			1813: out = 22524;
			1814: out = 22427;
			1815: out = 22334;
			1816: out = 22205;
			1817: out = 22040;
			1818: out = 21911;
			1819: out = 21798;
			1820: out = 21656;
			1821: out = 21508;
			1822: out = 21369;
			1823: out = 21235;
			1824: out = 21056;
			1825: out = 20954;
			1826: out = 20771;
			1827: out = 20574;
			1828: out = 20422;
			1829: out = 20264;
			1830: out = 20104;
			1831: out = 19929;
			1832: out = 19752;
			1833: out = 19575;
			1834: out = 19390;
			1835: out = 19209;
			1836: out = 19035;
			1837: out = 18876;
			1838: out = 18675;
			1839: out = 18498;
			1840: out = 18323;
			1841: out = 18118;
			1842: out = 17970;
			1843: out = 17778;
			1844: out = 17607;
			1845: out = 17424;
			1846: out = 17249;
			1847: out = 17081;
			1848: out = 16909;
			1849: out = 16725;
			1850: out = 16539;
			1851: out = 16346;
			1852: out = 16165;
			1853: out = 15984;
			1854: out = 15824;
			1855: out = 15647;
			1856: out = 15447;
			1857: out = 15275;
			1858: out = 15122;
			1859: out = 14952;
			1860: out = 14779;
			1861: out = 14637;
			1862: out = 14476;
			1863: out = 14291;
			1864: out = 14118;
			1865: out = 13949;
			1866: out = 13795;
			1867: out = 13615;
			1868: out = 13474;
			1869: out = 13254;
			1870: out = 13048;
			1871: out = 12940;
			1872: out = 12797;
			1873: out = 12652;
			1874: out = 12513;
			1875: out = 12345;
			1876: out = 12194;
			1877: out = 12027;
			1878: out = 11879;
			1879: out = 11753;
			1880: out = 11575;
			1881: out = 11447;
			1882: out = 11307;
			1883: out = 11169;
			1884: out = 11038;
			1885: out = 10892;
			1886: out = 10764;
			1887: out = 10617;
			1888: out = 10495;
			1889: out = 10361;
			1890: out = 10229;
			1891: out = 10114;
			1892: out = 9979;
			1893: out = 9862;
			1894: out = 9723;
			1895: out = 9603;
			1896: out = 9491;
			1897: out = 9341;
			1898: out = 9227;
			1899: out = 9120;
			1900: out = 9014;
			1901: out = 8878;
			1902: out = 8766;
			1903: out = 8632;
			1904: out = 8528;
			1905: out = 8408;
			1906: out = 8292;
			1907: out = 8177;
			1908: out = 8069;
			1909: out = 7972;
			1910: out = 7875;
			1911: out = 7783;
			1912: out = 7666;
			1913: out = 7546;
			1914: out = 7439;
			1915: out = 7261;
			1916: out = 7036;
			1917: out = 6820;
			1918: out = 6620;
			1919: out = 6400;
			1920: out = 6198;
			1921: out = 5974;
			1922: out = 5816;
			1923: out = 5625;
			1924: out = 5412;
			1925: out = 5236;
			1926: out = 5042;
			1927: out = 4850;
			1928: out = 4664;
			1929: out = 4503;
			1930: out = 4333;
			1931: out = 4161;
			1932: out = 3988;
			1933: out = 3813;
			1934: out = 3649;
			1935: out = 3488;
			1936: out = 3346;
			1937: out = 3198;
			1938: out = 3056;
			1939: out = 2877;
			1940: out = 2711;
			1941: out = 2592;
			1942: out = 2409;
			1943: out = 2246;
			1944: out = 2110;
			1945: out = 1974;
			1946: out = 1812;
			1947: out = 1667;
			1948: out = 1531;
			1949: out = 1387;
			1950: out = 1226;
			1951: out = 1081;
			1952: out = 949;
			1953: out = 793;
			1954: out = 713;
			1955: out = 562;
			1956: out = 412;
			1957: out = 276;
			1958: out = 113;
			1959: out = -39;
			1960: out = -176;
			1961: out = -333;
			1962: out = -465;
			1963: out = -585;
			1964: out = -736;
			1965: out = -868;
			1966: out = -1012;
			1967: out = -1140;
			1968: out = -1271;
			1969: out = -1416;
			1970: out = -1568;
			1971: out = -1673;
			1972: out = -1808;
			1973: out = -1950;
			1974: out = -2083;
			1975: out = -2230;
			1976: out = -2346;
			1977: out = -2518;
			1978: out = -2655;
			1979: out = -2803;
			1980: out = -2950;
			1981: out = -3104;
			1982: out = -3247;
			1983: out = -3401;
			1984: out = -3552;
			1985: out = -3713;
			1986: out = -3851;
			1987: out = -3989;
			1988: out = -4173;
			1989: out = -4323;
			1990: out = -4503;
			1991: out = -4670;
			1992: out = -4857;
			1993: out = -5014;
			1994: out = -5199;
			1995: out = -5401;
			1996: out = -5582;
			1997: out = -5783;
			1998: out = -5963;
			1999: out = -6180;
			2000: out = -6363;
			2001: out = -6576;
			2002: out = -6786;
			2003: out = -7001;
			2004: out = -7226;
			2005: out = -7446;
			2006: out = -7655;
			2007: out = -7884;
			2008: out = -8125;
			2009: out = -8334;
			2010: out = -8578;
			2011: out = -8809;
			2012: out = -9056;
			2013: out = -9310;
			2014: out = -9531;
			2015: out = -9770;
			2016: out = -10012;
			2017: out = -10264;
			2018: out = -10510;
			2019: out = -10759;
			2020: out = -10989;
			2021: out = -11235;
			2022: out = -11474;
			2023: out = -11702;
			2024: out = -11952;
			2025: out = -12172;
			2026: out = -12424;
			2027: out = -12657;
			2028: out = -12872;
			2029: out = -13092;
			2030: out = -13314;
			2031: out = -13542;
			2032: out = -13759;
			2033: out = -13957;
			2034: out = -14155;
			2035: out = -14374;
			2036: out = -14561;
			2037: out = -14752;
			2038: out = -14942;
			2039: out = -15141;
			2040: out = -15320;
			2041: out = -15517;
			2042: out = -15700;
			2043: out = -15850;
			2044: out = -16040;
			2045: out = -16207;
			2046: out = -16363;
			2047: out = -16525;
			2048: out = -16689;
			2049: out = -16823;
			2050: out = -16994;
			2051: out = -17136;
			2052: out = -17277;
			2053: out = -17419;
			2054: out = -17546;
			2055: out = -17718;
			2056: out = -17839;
			2057: out = -17948;
			2058: out = -18074;
			2059: out = -18166;
			2060: out = -18278;
			2061: out = -18385;
			2062: out = -18473;
			2063: out = -18592;
			2064: out = -18718;
			2065: out = -18793;
			2066: out = -18900;
			2067: out = -18977;
			2068: out = -19061;
			2069: out = -19171;
			2070: out = -19232;
			2071: out = -19328;
			2072: out = -19407;
			2073: out = -19488;
			2074: out = -19568;
			2075: out = -19650;
			2076: out = -19716;
			2077: out = -19769;
			2078: out = -19828;
			2079: out = -19891;
			2080: out = -19959;
			2081: out = -20011;
			2082: out = -20070;
			2083: out = -20131;
			2084: out = -20155;
			2085: out = -20239;
			2086: out = -20271;
			2087: out = -20336;
			2088: out = -20363;
			2089: out = -20399;
			2090: out = -20437;
			2091: out = -20477;
			2092: out = -20494;
			2093: out = -20535;
			2094: out = -20576;
			2095: out = -20585;
			2096: out = -20620;
			2097: out = -20650;
			2098: out = -20658;
			2099: out = -20691;
			2100: out = -20712;
			2101: out = -20729;
			2102: out = -20738;
			2103: out = -20750;
			2104: out = -20774;
			2105: out = -20766;
			2106: out = -20789;
			2107: out = -20809;
			2108: out = -20801;
			2109: out = -20824;
			2110: out = -20824;
			2111: out = -20819;
			2112: out = -20841;
			2113: out = -20829;
			2114: out = -20830;
			2115: out = -20853;
			2116: out = -20852;
			2117: out = -20842;
			2118: out = -20828;
			2119: out = -20818;
			2120: out = -20830;
			2121: out = -20819;
			2122: out = -20811;
			2123: out = -20800;
			2124: out = -20783;
			2125: out = -20780;
			2126: out = -20760;
			2127: out = -20740;
			2128: out = -20746;
			2129: out = -20715;
			2130: out = -20695;
			2131: out = -20668;
			2132: out = -20668;
			2133: out = -20644;
			2134: out = -20603;
			2135: out = -20567;
			2136: out = -20546;
			2137: out = -20517;
			2138: out = -20478;
			2139: out = -20451;
			2140: out = -20376;
			2141: out = -20320;
			2142: out = -20310;
			2143: out = -20262;
			2144: out = -20214;
			2145: out = -20180;
			2146: out = -20125;
			2147: out = -20086;
			2148: out = -20016;
			2149: out = -19962;
			2150: out = -19888;
			2151: out = -19812;
			2152: out = -19755;
			2153: out = -19661;
			2154: out = -19600;
			2155: out = -19520;
			2156: out = -19419;
			2157: out = -19344;
			2158: out = -19230;
			2159: out = -19135;
			2160: out = -19056;
			2161: out = -18955;
			2162: out = -18846;
			2163: out = -18715;
			2164: out = -18611;
			2165: out = -18477;
			2166: out = -18357;
			2167: out = -18234;
			2168: out = -18108;
			2169: out = -17962;
			2170: out = -17806;
			2171: out = -17685;
			2172: out = -17533;
			2173: out = -17397;
			2174: out = -17226;
			2175: out = -17080;
			2176: out = -16918;
			2177: out = -16761;
			2178: out = -16601;
			2179: out = -16446;
			2180: out = -16254;
			2181: out = -16101;
			2182: out = -15930;
			2183: out = -15763;
			2184: out = -15623;
			2185: out = -15438;
			2186: out = -15259;
			2187: out = -15100;
			2188: out = -14929;
			2189: out = -14749;
			2190: out = -14595;
			2191: out = -14420;
			2192: out = -14245;
			2193: out = -14073;
			2194: out = -13924;
			2195: out = -13764;
			2196: out = -13594;
			2197: out = -13437;
			2198: out = -13272;
			2199: out = -13097;
			2200: out = -12921;
			2201: out = -12774;
			2202: out = -12613;
			2203: out = -12450;
			2204: out = -12308;
			2205: out = -12138;
			2206: out = -11996;
			2207: out = -11851;
			2208: out = -11686;
			2209: out = -11546;
			2210: out = -11377;
			2211: out = -11247;
			2212: out = -11087;
			2213: out = -10954;
			2214: out = -10804;
			2215: out = -10653;
			2216: out = -10527;
			2217: out = -10361;
			2218: out = -10244;
			2219: out = -10103;
			2220: out = -9971;
			2221: out = -9852;
			2222: out = -9689;
			2223: out = -9570;
			2224: out = -9435;
			2225: out = -9290;
			2226: out = -9168;
			2227: out = -9046;
			2228: out = -8915;
			2229: out = -8794;
			2230: out = -8669;
			2231: out = -8542;
			2232: out = -8431;
			2233: out = -8324;
			2234: out = -8185;
			2235: out = -8064;
			2236: out = -7953;
			2237: out = -7817;
			2238: out = -7717;
			2239: out = -7601;
			2240: out = -7504;
			2241: out = -7389;
			2242: out = -7295;
			2243: out = -7187;
			2244: out = -7074;
			2245: out = -6953;
			2246: out = -6882;
			2247: out = -6788;
			2248: out = -6675;
			2249: out = -6586;
			2250: out = -6431;
			2251: out = -6261;
			2252: out = -6102;
			2253: out = -5942;
			2254: out = -5778;
			2255: out = -5621;
			2256: out = -5464;
			2257: out = -5331;
			2258: out = -5167;
			2259: out = -5014;
			2260: out = -4873;
			2261: out = -4722;
			2262: out = -4564;
			2263: out = -4443;
			2264: out = -4300;
			2265: out = -4151;
			2266: out = -4014;
			2267: out = -3895;
			2268: out = -3741;
			2269: out = -3628;
			2270: out = -3511;
			2271: out = -3368;
			2272: out = -3251;
			2273: out = -3125;
			2274: out = -3001;
			2275: out = -2885;
			2276: out = -2759;
			2277: out = -2648;
			2278: out = -2515;
			2279: out = -2395;
			2280: out = -2301;
			2281: out = -2184;
			2282: out = -2077;
			2283: out = -1957;
			2284: out = -1863;
			2285: out = -1736;
			2286: out = -1627;
			2287: out = -1534;
			2288: out = -1411;
			2289: out = -1309;
			2290: out = -1182;
			2291: out = -1094;
			2292: out = -999;
			2293: out = -894;
			2294: out = -800;
			2295: out = -667;
			2296: out = -563;
			2297: out = -455;
			2298: out = -337;
			2299: out = -241;
			2300: out = -138;
			2301: out = -41;
			2302: out = 65;
			2303: out = 171;
			2304: out = 268;
			2305: out = 353;
			2306: out = 463;
			2307: out = 583;
			2308: out = 684;
			2309: out = 808;
			2310: out = 905;
			2311: out = 1004;
			2312: out = 1138;
			2313: out = 1220;
			2314: out = 1336;
			2315: out = 1450;
			2316: out = 1530;
			2317: out = 1660;
			2318: out = 1719;
			2319: out = 1815;
			2320: out = 1957;
			2321: out = 2073;
			2322: out = 2214;
			2323: out = 2323;
			2324: out = 2446;
			2325: out = 2563;
			2326: out = 2714;
			2327: out = 2836;
			2328: out = 2965;
			2329: out = 3091;
			2330: out = 3225;
			2331: out = 3363;
			2332: out = 3494;
			2333: out = 3641;
			2334: out = 3769;
			2335: out = 3923;
			2336: out = 4085;
			2337: out = 4230;
			2338: out = 4395;
			2339: out = 4569;
			2340: out = 4705;
			2341: out = 4870;
			2342: out = 5031;
			2343: out = 5220;
			2344: out = 5369;
			2345: out = 5532;
			2346: out = 5716;
			2347: out = 5901;
			2348: out = 6071;
			2349: out = 6256;
			2350: out = 6433;
			2351: out = 6597;
			2352: out = 6790;
			2353: out = 6963;
			2354: out = 7155;
			2355: out = 7328;
			2356: out = 7524;
			2357: out = 7682;
			2358: out = 7849;
			2359: out = 8053;
			2360: out = 8220;
			2361: out = 8387;
			2362: out = 8583;
			2363: out = 8752;
			2364: out = 8917;
			2365: out = 9098;
			2366: out = 9266;
			2367: out = 9427;
			2368: out = 9588;
			2369: out = 9758;
			2370: out = 9915;
			2371: out = 10104;
			2372: out = 10264;
			2373: out = 10412;
			2374: out = 10563;
			2375: out = 10739;
			2376: out = 10876;
			2377: out = 11037;
			2378: out = 11192;
			2379: out = 11339;
			2380: out = 11473;
			2381: out = 11614;
			2382: out = 11770;
			2383: out = 11913;
			2384: out = 12048;
			2385: out = 12182;
			2386: out = 12307;
			2387: out = 12450;
			2388: out = 12563;
			2389: out = 12720;
			2390: out = 12855;
			2391: out = 12955;
			2392: out = 13086;
			2393: out = 13207;
			2394: out = 13333;
			2395: out = 13445;
			2396: out = 13614;
			2397: out = 13709;
			2398: out = 13836;
			2399: out = 13946;
			2400: out = 14067;
			2401: out = 14171;
			2402: out = 14333;
			2403: out = 14458;
			2404: out = 14548;
			2405: out = 14659;
			2406: out = 14736;
			2407: out = 14842;
			2408: out = 14940;
			2409: out = 15033;
			2410: out = 15126;
			2411: out = 15242;
			2412: out = 15340;
			2413: out = 15450;
			2414: out = 15523;
			2415: out = 15629;
			2416: out = 15723;
			2417: out = 15822;
			2418: out = 15902;
			2419: out = 16015;
			2420: out = 16101;
			2421: out = 16177;
			2422: out = 16270;
			2423: out = 16363;
			2424: out = 16447;
			2425: out = 16544;
			2426: out = 16615;
			2427: out = 16706;
			2428: out = 16777;
			2429: out = 16864;
			2430: out = 16935;
			2431: out = 17015;
			2432: out = 17091;
			2433: out = 17173;
			2434: out = 17239;
			2435: out = 17319;
			2436: out = 17393;
			2437: out = 17468;
			2438: out = 17548;
			2439: out = 17615;
			2440: out = 17700;
			2441: out = 17769;
			2442: out = 17829;
			2443: out = 17893;
			2444: out = 17969;
			2445: out = 18060;
			2446: out = 18113;
			2447: out = 18194;
			2448: out = 18244;
			2449: out = 18327;
			2450: out = 18388;
			2451: out = 18456;
			2452: out = 18532;
			2453: out = 18587;
			2454: out = 18633;
			2455: out = 18718;
			2456: out = 18774;
			2457: out = 18825;
			2458: out = 18896;
			2459: out = 18935;
			2460: out = 19012;
			2461: out = 19061;
			2462: out = 19121;
			2463: out = 19173;
			2464: out = 19234;
			2465: out = 19259;
			2466: out = 19263;
			2467: out = 19257;
			2468: out = 19283;
			2469: out = 19323;
			2470: out = 19336;
			2471: out = 19368;
			2472: out = 19389;
			2473: out = 19416;
			2474: out = 19365;
			2475: out = 19305;
			2476: out = 19258;
			2477: out = 19238;
			2478: out = 19237;
			2479: out = 19248;
			2480: out = 19194;
			2481: out = 19159;
			2482: out = 19156;
			2483: out = 19169;
			2484: out = 19156;
			2485: out = 19157;
			2486: out = 19187;
			2487: out = 19105;
			2488: out = 19085;
			2489: out = 19045;
			2490: out = 19035;
			2491: out = 19037;
			2492: out = 19045;
			2493: out = 19049;
			2494: out = 19009;
			2495: out = 18894;
			2496: out = 18858;
			2497: out = 18825;
			2498: out = 18821;
			2499: out = 18834;
			2500: out = 18788;
			2501: out = 18728;
			2502: out = 18647;
			2503: out = 18600;
			2504: out = 18533;
			2505: out = 18565;
			2506: out = 18503;
			2507: out = 18429;
			2508: out = 18392;
			2509: out = 18348;
			2510: out = 18351;
			2511: out = 18280;
			2512: out = 18181;
			2513: out = 18125;
			2514: out = 18040;
			2515: out = 18014;
			2516: out = 17937;
			2517: out = 17822;
			2518: out = 17777;
			2519: out = 17693;
			2520: out = 17613;
			2521: out = 17533;
			2522: out = 17437;
			2523: out = 17360;
			2524: out = 17247;
			2525: out = 17154;
			2526: out = 17036;
			2527: out = 16901;
			2528: out = 16825;
			2529: out = 16725;
			2530: out = 16591;
			2531: out = 16505;
			2532: out = 16399;
			2533: out = 16261;
			2534: out = 16186;
			2535: out = 16040;
			2536: out = 15898;
			2537: out = 15805;
			2538: out = 15631;
			2539: out = 15528;
			2540: out = 15428;
			2541: out = 15274;
			2542: out = 15164;
			2543: out = 15045;
			2544: out = 14925;
			2545: out = 14770;
			2546: out = 14631;
			2547: out = 14509;
			2548: out = 14348;
			2549: out = 14253;
			2550: out = 14142;
			2551: out = 14003;
			2552: out = 13858;
			2553: out = 13681;
			2554: out = 13576;
			2555: out = 13438;
			2556: out = 13314;
			2557: out = 13213;
			2558: out = 13073;
			2559: out = 12972;
			2560: out = 12829;
			2561: out = 12670;
			2562: out = 12546;
			2563: out = 12380;
			2564: out = 12238;
			2565: out = 12142;
			2566: out = 12031;
			2567: out = 11883;
			2568: out = 11775;
			2569: out = 11659;
			2570: out = 11536;
			2571: out = 11384;
			2572: out = 11273;
			2573: out = 11155;
			2574: out = 11012;
			2575: out = 10909;
			2576: out = 10751;
			2577: out = 10648;
			2578: out = 10524;
			2579: out = 10398;
			2580: out = 10281;
			2581: out = 10180;
			2582: out = 10079;
			2583: out = 9947;
			2584: out = 9828;
			2585: out = 9714;
			2586: out = 9604;
			2587: out = 9481;
			2588: out = 9389;
			2589: out = 9321;
			2590: out = 9189;
			2591: out = 9065;
			2592: out = 8943;
			2593: out = 8841;
			2594: out = 8732;
			2595: out = 8619;
			2596: out = 8523;
			2597: out = 8404;
			2598: out = 8301;
			2599: out = 8206;
			2600: out = 8107;
			2601: out = 8022;
			2602: out = 7922;
			2603: out = 7824;
			2604: out = 7729;
			2605: out = 7645;
			2606: out = 7555;
			2607: out = 7468;
			2608: out = 7344;
			2609: out = 7268;
			2610: out = 7186;
			2611: out = 7092;
			2612: out = 6992;
			2613: out = 6908;
			2614: out = 6824;
			2615: out = 6718;
			2616: out = 6635;
			2617: out = 6582;
			2618: out = 6510;
			2619: out = 6411;
			2620: out = 6314;
			2621: out = 6217;
			2622: out = 6135;
			2623: out = 6072;
			2624: out = 5989;
			2625: out = 5913;
			2626: out = 5825;
			2627: out = 5738;
			2628: out = 5662;
			2629: out = 5575;
			2630: out = 5531;
			2631: out = 5459;
			2632: out = 5385;
			2633: out = 5295;
			2634: out = 5213;
			2635: out = 5154;
			2636: out = 5087;
			2637: out = 5008;
			2638: out = 4947;
			2639: out = 4874;
			2640: out = 4807;
			2641: out = 4731;
			2642: out = 4685;
			2643: out = 4602;
			2644: out = 4467;
			2645: out = 4325;
			2646: out = 4152;
			2647: out = 3992;
			2648: out = 3853;
			2649: out = 3711;
			2650: out = 3556;
			2651: out = 3387;
			2652: out = 3251;
			2653: out = 3105;
			2654: out = 2983;
			2655: out = 2843;
			2656: out = 2699;
			2657: out = 2575;
			2658: out = 2436;
			2659: out = 2330;
			2660: out = 2192;
			2661: out = 2068;
			2662: out = 1935;
			2663: out = 1825;
			2664: out = 1712;
			2665: out = 1575;
			2666: out = 1490;
			2667: out = 1344;
			2668: out = 1248;
			2669: out = 1118;
			2670: out = 1025;
			2671: out = 903;
			2672: out = 775;
			2673: out = 680;
			2674: out = 573;
			2675: out = 443;
			2676: out = 342;
			2677: out = 229;
			2678: out = 128;
			2679: out = 27;
			2680: out = -83;
			2681: out = -199;
			2682: out = -280;
			2683: out = -386;
			2684: out = -489;
			2685: out = -586;
			2686: out = -671;
			2687: out = -783;
			2688: out = -894;
			2689: out = -995;
			2690: out = -1093;
			2691: out = -1192;
			2692: out = -1288;
			2693: out = -1375;
			2694: out = -1456;
			2695: out = -1567;
			2696: out = -1631;
			2697: out = -1759;
			2698: out = -1880;
			2699: out = -1948;
			2700: out = -2060;
			2701: out = -2152;
			2702: out = -2265;
			2703: out = -2362;
			2704: out = -2474;
			2705: out = -2571;
			2706: out = -2645;
			2707: out = -2760;
			2708: out = -2859;
			2709: out = -2988;
			2710: out = -3081;
			2711: out = -3170;
			2712: out = -3274;
			2713: out = -3373;
			2714: out = -3486;
			2715: out = -3578;
			2716: out = -3691;
			2717: out = -3787;
			2718: out = -3891;
			2719: out = -3985;
			2720: out = -4083;
			2721: out = -4199;
			2722: out = -4316;
			2723: out = -4411;
			2724: out = -4521;
			2725: out = -4641;
			2726: out = -4758;
			2727: out = -4855;
			2728: out = -4982;
			2729: out = -5086;
			2730: out = -5220;
			2731: out = -5333;
			2732: out = -5466;
			2733: out = -5604;
			2734: out = -5720;
			2735: out = -5838;
			2736: out = -5980;
			2737: out = -6119;
			2738: out = -6267;
			2739: out = -6384;
			2740: out = -6529;
			2741: out = -6678;
			2742: out = -6807;
			2743: out = -6943;
			2744: out = -7115;
			2745: out = -7262;
			2746: out = -7412;
			2747: out = -7589;
			2748: out = -7753;
			2749: out = -7902;
			2750: out = -8077;
			2751: out = -8219;
			2752: out = -8409;
			2753: out = -8577;
			2754: out = -8745;
			2755: out = -8938;
			2756: out = -9129;
			2757: out = -9282;
			2758: out = -9439;
			2759: out = -9623;
			2760: out = -9830;
			2761: out = -10024;
			2762: out = -10186;
			2763: out = -10387;
			2764: out = -10563;
			2765: out = -10737;
			2766: out = -10947;
			2767: out = -11160;
			2768: out = -11343;
			2769: out = -11475;
			2770: out = -11666;
			2771: out = -11841;
			2772: out = -12003;
			2773: out = -12179;
			2774: out = -12351;
			2775: out = -12520;
			2776: out = -12688;
			2777: out = -12838;
			2778: out = -13011;
			2779: out = -13181;
			2780: out = -13321;
			2781: out = -13468;
			2782: out = -13621;
			2783: out = -13772;
			2784: out = -13901;
			2785: out = -14062;
			2786: out = -14182;
			2787: out = -14334;
			2788: out = -14458;
			2789: out = -14595;
			2790: out = -14738;
			2791: out = -14845;
			2792: out = -14979;
			2793: out = -15107;
			2794: out = -15220;
			2795: out = -15318;
			2796: out = -15441;
			2797: out = -15550;
			2798: out = -15673;
			2799: out = -15765;
			2800: out = -15863;
			2801: out = -15969;
			2802: out = -16061;
			2803: out = -16163;
			2804: out = -16251;
			2805: out = -16344;
			2806: out = -16414;
			2807: out = -16511;
			2808: out = -16600;
			2809: out = -16682;
			2810: out = -16752;
			2811: out = -16831;
			2812: out = -16907;
			2813: out = -16977;
			2814: out = -17053;
			2815: out = -17120;
			2816: out = -17159;
			2817: out = -17236;
			2818: out = -17285;
			2819: out = -17370;
			2820: out = -17403;
			2821: out = -17459;
			2822: out = -17534;
			2823: out = -17574;
			2824: out = -17642;
			2825: out = -17661;
			2826: out = -17705;
			2827: out = -17763;
			2828: out = -17807;
			2829: out = -17841;
			2830: out = -17878;
			2831: out = -17898;
			2832: out = -17919;
			2833: out = -17974;
			2834: out = -18009;
			2835: out = -18035;
			2836: out = -18062;
			2837: out = -18078;
			2838: out = -18084;
			2839: out = -18132;
			2840: out = -18170;
			2841: out = -18161;
			2842: out = -18182;
			2843: out = -18202;
			2844: out = -18218;
			2845: out = -18234;
			2846: out = -18256;
			2847: out = -18267;
			2848: out = -18266;
			2849: out = -18280;
			2850: out = -18290;
			2851: out = -18250;
			2852: out = -18274;
			2853: out = -18289;
			2854: out = -18292;
			2855: out = -18320;
			2856: out = -18326;
			2857: out = -18337;
			2858: out = -18326;
			2859: out = -18315;
			2860: out = -18320;
			2861: out = -18321;
			2862: out = -18317;
			2863: out = -18337;
			2864: out = -18305;
			2865: out = -18310;
			2866: out = -18289;
			2867: out = -18291;
			2868: out = -18297;
			2869: out = -18278;
			2870: out = -18268;
			2871: out = -18276;
			2872: out = -18244;
			2873: out = -18221;
			2874: out = -18225;
			2875: out = -18205;
			2876: out = -18192;
			2877: out = -18171;
			2878: out = -18134;
			2879: out = -18118;
			2880: out = -18129;
			2881: out = -18087;
			2882: out = -18077;
			2883: out = -18045;
			2884: out = -18026;
			2885: out = -17993;
			2886: out = -17966;
			2887: out = -17940;
			2888: out = -17911;
			2889: out = -17865;
			2890: out = -17840;
			2891: out = -17806;
			2892: out = -17807;
			2893: out = -17761;
			2894: out = -17719;
			2895: out = -17701;
			2896: out = -17647;
			2897: out = -17630;
			2898: out = -17583;
			2899: out = -17559;
			2900: out = -17531;
			2901: out = -17498;
			2902: out = -17461;
			2903: out = -17425;
			2904: out = -17393;
			2905: out = -17342;
			2906: out = -17309;
			2907: out = -17258;
			2908: out = -17214;
			2909: out = -17176;
			2910: out = -17102;
			2911: out = -17080;
			2912: out = -17003;
			2913: out = -16967;
			2914: out = -16896;
			2915: out = -16853;
			2916: out = -16789;
			2917: out = -16724;
			2918: out = -16663;
			2919: out = -16587;
			2920: out = -16523;
			2921: out = -16453;
			2922: out = -16376;
			2923: out = -16297;
			2924: out = -16207;
			2925: out = -16139;
			2926: out = -16047;
			2927: out = -15967;
			2928: out = -15878;
			2929: out = -15763;
			2930: out = -15683;
			2931: out = -15562;
			2932: out = -15482;
			2933: out = -15367;
			2934: out = -15270;
			2935: out = -15150;
			2936: out = -15042;
			2937: out = -14930;
			2938: out = -14813;
			2939: out = -14710;
			2940: out = -14576;
			2941: out = -14449;
			2942: out = -14312;
			2943: out = -14198;
			2944: out = -14089;
			2945: out = -13943;
			2946: out = -13804;
			2947: out = -13682;
			2948: out = -13551;
			2949: out = -13413;
			2950: out = -13273;
			2951: out = -13148;
			2952: out = -13033;
			2953: out = -12879;
			2954: out = -12737;
			2955: out = -12588;
			2956: out = -12449;
			2957: out = -12319;
			2958: out = -12162;
			2959: out = -12021;
			2960: out = -11887;
			2961: out = -11757;
			2962: out = -11613;
			2963: out = -11468;
			2964: out = -11347;
			2965: out = -11201;
			2966: out = -11067;
			2967: out = -10947;
			2968: out = -10806;
			2969: out = -10666;
			2970: out = -10545;
			2971: out = -10404;
			2972: out = -10266;
			2973: out = -10152;
			2974: out = -10014;
			2975: out = -9888;
			2976: out = -9763;
			2977: out = -9636;
			2978: out = -9527;
			2979: out = -9399;
			2980: out = -9260;
			2981: out = -9140;
			2982: out = -9016;
			2983: out = -8889;
			2984: out = -8789;
			2985: out = -8654;
			2986: out = -8550;
			2987: out = -8430;
			2988: out = -8305;
			2989: out = -8184;
			2990: out = -8089;
			2991: out = -7967;
			2992: out = -7853;
			2993: out = -7732;
			2994: out = -7615;
			2995: out = -7512;
			2996: out = -7403;
			2997: out = -7298;
			2998: out = -7197;
			2999: out = -7066;
			3000: out = -6974;
			3001: out = -6871;
			3002: out = -6779;
			3003: out = -6682;
			3004: out = -6570;
			3005: out = -6482;
			3006: out = -6379;
			3007: out = -6278;
			3008: out = -6198;
			3009: out = -6108;
			3010: out = -6012;
			3011: out = -5919;
			3012: out = -5834;
			3013: out = -5746;
			3014: out = -5666;
			3015: out = -5576;
			3016: out = -5495;
			3017: out = -5397;
			3018: out = -5316;
			3019: out = -5234;
			3020: out = -5153;
			3021: out = -5079;
			3022: out = -4998;
			3023: out = -4886;
			3024: out = -4826;
			3025: out = -4759;
			3026: out = -4655;
			3027: out = -4601;
			3028: out = -4510;
			3029: out = -4438;
			3030: out = -4357;
			3031: out = -4256;
			3032: out = -4114;
			3033: out = -3991;
			3034: out = -3850;
			3035: out = -3725;
			3036: out = -3620;
			3037: out = -3472;
			3038: out = -3347;
			3039: out = -3246;
			3040: out = -3133;
			3041: out = -3032;
			3042: out = -2912;
			3043: out = -2809;
			3044: out = -2719;
			3045: out = -2608;
			3046: out = -2512;
			3047: out = -2397;
			3048: out = -2293;
			3049: out = -2192;
			3050: out = -2089;
			3051: out = -1994;
			3052: out = -1914;
			3053: out = -1802;
			3054: out = -1719;
			3055: out = -1638;
			3056: out = -1531;
			3057: out = -1435;
			3058: out = -1340;
			3059: out = -1246;
			3060: out = -1169;
			3061: out = -1074;
			3062: out = -993;
			3063: out = -909;
			3064: out = -829;
			3065: out = -759;
			3066: out = -647;
			3067: out = -577;
			3068: out = -495;
			3069: out = -411;
			3070: out = -333;
			3071: out = -267;
			3072: out = -175;
			3073: out = -97;
			3074: out = -6;
			3075: out = 68;
			3076: out = 140;
			3077: out = 195;
			3078: out = 300;
			3079: out = 356;
			3080: out = 463;
			3081: out = 528;
			3082: out = 596;
			3083: out = 665;
			3084: out = 719;
			3085: out = 820;
			3086: out = 885;
			3087: out = 947;
			3088: out = 1031;
			3089: out = 1083;
			3090: out = 1167;
			3091: out = 1231;
			3092: out = 1298;
			3093: out = 1380;
			3094: out = 1444;
			3095: out = 1505;
			3096: out = 1582;
			3097: out = 1651;
			3098: out = 1755;
			3099: out = 1802;
			3100: out = 1861;
			3101: out = 1961;
			3102: out = 2042;
			3103: out = 2112;
			3104: out = 2191;
			3105: out = 2279;
			3106: out = 2355;
			3107: out = 2439;
			3108: out = 2514;
			3109: out = 2618;
			3110: out = 2681;
			3111: out = 2756;
			3112: out = 2848;
			3113: out = 2951;
			3114: out = 3025;
			3115: out = 3118;
			3116: out = 3210;
			3117: out = 3280;
			3118: out = 3376;
			3119: out = 3489;
			3120: out = 3575;
			3121: out = 3679;
			3122: out = 3779;
			3123: out = 3876;
			3124: out = 3977;
			3125: out = 4066;
			3126: out = 4178;
			3127: out = 4286;
			3128: out = 4379;
			3129: out = 4491;
			3130: out = 4602;
			3131: out = 4727;
			3132: out = 4840;
			3133: out = 4966;
			3134: out = 5090;
			3135: out = 5215;
			3136: out = 5338;
			3137: out = 5463;
			3138: out = 5571;
			3139: out = 5696;
			3140: out = 5830;
			3141: out = 5965;
			3142: out = 6107;
			3143: out = 6216;
			3144: out = 6364;
			3145: out = 6499;
			3146: out = 6616;
			3147: out = 6753;
			3148: out = 6882;
			3149: out = 7025;
			3150: out = 7144;
			3151: out = 7268;
			3152: out = 7412;
			3153: out = 7530;
			3154: out = 7670;
			3155: out = 7790;
			3156: out = 7934;
			3157: out = 8040;
			3158: out = 8168;
			3159: out = 8304;
			3160: out = 8421;
			3161: out = 8546;
			3162: out = 8679;
			3163: out = 8786;
			3164: out = 8900;
			3165: out = 9037;
			3166: out = 9149;
			3167: out = 9264;
			3168: out = 9382;
			3169: out = 9488;
			3170: out = 9602;
			3171: out = 9717;
			3172: out = 9812;
			3173: out = 9935;
			3174: out = 10023;
			3175: out = 10137;
			3176: out = 10244;
			3177: out = 10349;
			3178: out = 10463;
			3179: out = 10553;
			3180: out = 10652;
			3181: out = 10748;
			3182: out = 10858;
			3183: out = 10940;
			3184: out = 11060;
			3185: out = 11120;
			3186: out = 11229;
			3187: out = 11310;
			3188: out = 11405;
			3189: out = 11496;
			3190: out = 11578;
			3191: out = 11670;
			3192: out = 11741;
			3193: out = 11829;
			3194: out = 11919;
			3195: out = 12000;
			3196: out = 12085;
			3197: out = 12152;
			3198: out = 12225;
			3199: out = 12320;
			3200: out = 12383;
			3201: out = 12465;
			3202: out = 12542;
			3203: out = 12616;
			3204: out = 12676;
			3205: out = 12765;
			3206: out = 12840;
			3207: out = 12917;
			3208: out = 12978;
			3209: out = 13054;
			3210: out = 13124;
			3211: out = 13189;
			3212: out = 13246;
			3213: out = 13318;
			3214: out = 13389;
			3215: out = 13440;
			3216: out = 13518;
			3217: out = 13557;
			3218: out = 13611;
			3219: out = 13686;
			3220: out = 13746;
			3221: out = 13789;
			3222: out = 13860;
			3223: out = 13866;
			3224: out = 13935;
			3225: out = 13979;
			3226: out = 14050;
			3227: out = 14109;
			3228: out = 14172;
			3229: out = 14232;
			3230: out = 14288;
			3231: out = 14317;
			3232: out = 14387;
			3233: out = 14424;
			3234: out = 14485;
			3235: out = 14542;
			3236: out = 14575;
			3237: out = 14616;
			3238: out = 14676;
			3239: out = 14725;
			3240: out = 14772;
			3241: out = 14820;
			3242: out = 14863;
			3243: out = 14911;
			3244: out = 14952;
			3245: out = 15025;
			3246: out = 15043;
			3247: out = 15101;
			3248: out = 15120;
			3249: out = 15184;
			3250: out = 15203;
			3251: out = 15254;
			3252: out = 15284;
			3253: out = 15321;
			3254: out = 15351;
			3255: out = 15390;
			3256: out = 15425;
			3257: out = 15473;
			3258: out = 15481;
			3259: out = 15476;
			3260: out = 15484;
			3261: out = 15492;
			3262: out = 15475;
			3263: out = 15481;
			3264: out = 15437;
			3265: out = 15370;
			3266: out = 15361;
			3267: out = 15397;
			3268: out = 15405;
			3269: out = 15389;
			3270: out = 15376;
			3271: out = 15322;
			3272: out = 15309;
			3273: out = 15302;
			3274: out = 15293;
			3275: out = 15255;
			3276: out = 15267;
			3277: out = 15245;
			3278: out = 15259;
			3279: out = 15275;
			3280: out = 15240;
			3281: out = 15220;
			3282: out = 15224;
			3283: out = 15151;
			3284: out = 15145;
			3285: out = 15145;
			3286: out = 15132;
			3287: out = 15108;
			3288: out = 15114;
			3289: out = 15124;
			3290: out = 15104;
			3291: out = 15059;
			3292: out = 15021;
			3293: out = 15041;
			3294: out = 15012;
			3295: out = 15002;
			3296: out = 15046;
			3297: out = 15041;
			3298: out = 15002;
			3299: out = 14983;
			3300: out = 14895;
			3301: out = 14907;
			3302: out = 14909;
			3303: out = 14895;
			3304: out = 14891;
			3305: out = 14909;
			3306: out = 14855;
			3307: out = 14834;
			3308: out = 14845;
			3309: out = 14841;
			3310: out = 14792;
			3311: out = 14753;
			3312: out = 14743;
			3313: out = 14679;
			3314: out = 14689;
			3315: out = 14607;
			3316: out = 14565;
			3317: out = 14587;
			3318: out = 14525;
			3319: out = 14489;
			3320: out = 14477;
			3321: out = 14455;
			3322: out = 14450;
			3323: out = 14344;
			3324: out = 14282;
			3325: out = 14242;
			3326: out = 14209;
			3327: out = 14177;
			3328: out = 14111;
			3329: out = 14062;
			3330: out = 14033;
			3331: out = 13934;
			3332: out = 13873;
			3333: out = 13841;
			3334: out = 13772;
			3335: out = 13651;
			3336: out = 13614;
			3337: out = 13559;
			3338: out = 13468;
			3339: out = 13388;
			3340: out = 13333;
			3341: out = 13260;
			3342: out = 13136;
			3343: out = 13083;
			3344: out = 13037;
			3345: out = 12912;
			3346: out = 12789;
			3347: out = 12707;
			3348: out = 12598;
			3349: out = 12527;
			3350: out = 12441;
			3351: out = 12362;
			3352: out = 12257;
			3353: out = 12180;
			3354: out = 12086;
			3355: out = 12016;
			3356: out = 11896;
			3357: out = 11794;
			3358: out = 11681;
			3359: out = 11552;
			3360: out = 11476;
			3361: out = 11390;
			3362: out = 11278;
			3363: out = 11178;
			3364: out = 11058;
			3365: out = 10979;
			3366: out = 10896;
			3367: out = 10778;
			3368: out = 10668;
			3369: out = 10546;
			3370: out = 10468;
			3371: out = 10368;
			3372: out = 10269;
			3373: out = 10190;
			3374: out = 10079;
			3375: out = 9954;
			3376: out = 9850;
			3377: out = 9747;
			3378: out = 9654;
			3379: out = 9543;
			3380: out = 9437;
			3381: out = 9356;
			3382: out = 9266;
			3383: out = 9141;
			3384: out = 9058;
			3385: out = 8962;
			3386: out = 8865;
			3387: out = 8752;
			3388: out = 8642;
			3389: out = 8540;
			3390: out = 8470;
			3391: out = 8374;
			3392: out = 8267;
			3393: out = 8174;
			3394: out = 8085;
			3395: out = 7973;
			3396: out = 7880;
			3397: out = 7831;
			3398: out = 7726;
			3399: out = 7625;
			3400: out = 7538;
			3401: out = 7432;
			3402: out = 7363;
			3403: out = 7256;
			3404: out = 7183;
			3405: out = 7108;
			3406: out = 7007;
			3407: out = 6915;
			3408: out = 6845;
			3409: out = 6751;
			3410: out = 6621;
			3411: out = 6542;
			3412: out = 6481;
			3413: out = 6407;
			3414: out = 6331;
			3415: out = 6255;
			3416: out = 6194;
			3417: out = 6101;
			3418: out = 6027;
			3419: out = 5955;
			3420: out = 5866;
			3421: out = 5782;
			3422: out = 5709;
			3423: out = 5641;
			3424: out = 5559;
			3425: out = 5500;
			3426: out = 5437;
			3427: out = 5327;
			3428: out = 5288;
			3429: out = 5226;
			3430: out = 5191;
			3431: out = 5107;
			3432: out = 5040;
			3433: out = 4952;
			3434: out = 4895;
			3435: out = 4822;
			3436: out = 4766;
			3437: out = 4710;
			3438: out = 4641;
			3439: out = 4600;
			3440: out = 4529;
			3441: out = 4485;
			3442: out = 4416;
			3443: out = 4339;
			3444: out = 4272;
			3445: out = 4201;
			3446: out = 4160;
			3447: out = 4089;
			3448: out = 4050;
			3449: out = 4001;
			3450: out = 3912;
			3451: out = 3864;
			3452: out = 3819;
			3453: out = 3758;
			3454: out = 3716;
			3455: out = 3645;
			3456: out = 3594;
			3457: out = 3525;
			3458: out = 3481;
			3459: out = 3424;
			3460: out = 3386;
			3461: out = 3323;
			3462: out = 3290;
			3463: out = 3210;
			3464: out = 3200;
			3465: out = 3133;
			3466: out = 3102;
			3467: out = 3051;
			3468: out = 2997;
			3469: out = 2952;
			3470: out = 2914;
			3471: out = 2882;
			3472: out = 2827;
			3473: out = 2741;
			3474: out = 2625;
			3475: out = 2514;
			3476: out = 2404;
			3477: out = 2299;
			3478: out = 2182;
			3479: out = 2080;
			3480: out = 1963;
			3481: out = 1871;
			3482: out = 1741;
			3483: out = 1643;
			3484: out = 1567;
			3485: out = 1468;
			3486: out = 1351;
			3487: out = 1240;
			3488: out = 1169;
			3489: out = 1070;
			3490: out = 967;
			3491: out = 880;
			3492: out = 786;
			3493: out = 675;
			3494: out = 624;
			3495: out = 547;
			3496: out = 434;
			3497: out = 347;
			3498: out = 251;
			3499: out = 160;
			3500: out = 67;
			3501: out = -19;
			3502: out = -112;
			3503: out = -196;
			3504: out = -274;
			3505: out = -347;
			3506: out = -413;
			3507: out = -496;
			3508: out = -597;
			3509: out = -670;
			3510: out = -747;
			3511: out = -818;
			3512: out = -884;
			3513: out = -941;
			3514: out = -1030;
			3515: out = -1095;
			3516: out = -1152;
			3517: out = -1236;
			3518: out = -1308;
			3519: out = -1368;
			3520: out = -1450;
			3521: out = -1500;
			3522: out = -1592;
			3523: out = -1640;
			3524: out = -1724;
			3525: out = -1797;
			3526: out = -1863;
			3527: out = -1946;
			3528: out = -2010;
			3529: out = -2066;
			3530: out = -2157;
			3531: out = -2215;
			3532: out = -2280;
			3533: out = -2357;
			3534: out = -2416;
			3535: out = -2488;
			3536: out = -2570;
			3537: out = -2630;
			3538: out = -2697;
			3539: out = -2760;
			3540: out = -2819;
			3541: out = -2898;
			3542: out = -2981;
			3543: out = -3042;
			3544: out = -3110;
			3545: out = -3176;
			3546: out = -3245;
			3547: out = -3310;
			3548: out = -3393;
			3549: out = -3451;
			3550: out = -3518;
			3551: out = -3567;
			3552: out = -3661;
			3553: out = -3720;
			3554: out = -3807;
			3555: out = -3876;
			3556: out = -3950;
			3557: out = -4027;
			3558: out = -4095;
			3559: out = -4171;
			3560: out = -4250;
			3561: out = -4339;
			3562: out = -4409;
			3563: out = -4504;
			3564: out = -4589;
			3565: out = -4685;
			3566: out = -4750;
			3567: out = -4845;
			3568: out = -4926;
			3569: out = -5031;
			3570: out = -5136;
			3571: out = -5205;
			3572: out = -5323;
			3573: out = -5415;
			3574: out = -5499;
			3575: out = -5603;
			3576: out = -5714;
			3577: out = -5831;
			3578: out = -5933;
			3579: out = -6026;
			3580: out = -6132;
			3581: out = -6241;
			3582: out = -6362;
			3583: out = -6469;
			3584: out = -6593;
			3585: out = -6701;
			3586: out = -6846;
			3587: out = -6952;
			3588: out = -7084;
			3589: out = -7202;
			3590: out = -7323;
			3591: out = -7465;
			3592: out = -7571;
			3593: out = -7710;
			3594: out = -7846;
			3595: out = -7995;
			3596: out = -8118;
			3597: out = -8237;
			3598: out = -8390;
			3599: out = -8523;
			3600: out = -8654;
			3601: out = -8790;
			3602: out = -8924;
			3603: out = -9055;
			3604: out = -9201;
			3605: out = -9323;
			3606: out = -9467;
			3607: out = -9604;
			3608: out = -9717;
			3609: out = -9881;
			3610: out = -9984;
			3611: out = -10107;
			3612: out = -10248;
			3613: out = -10360;
			3614: out = -10477;
			3615: out = -10600;
			3616: out = -10720;
			3617: out = -10832;
			3618: out = -10936;
			3619: out = -11072;
			3620: out = -11197;
			3621: out = -11304;
			3622: out = -11414;
			3623: out = -11506;
			3624: out = -11615;
			3625: out = -11730;
			3626: out = -11822;
			3627: out = -11945;
			3628: out = -12030;
			3629: out = -12128;
			3630: out = -12221;
			3631: out = -12325;
			3632: out = -12410;
			3633: out = -12502;
			3634: out = -12571;
			3635: out = -12667;
			3636: out = -12738;
			3637: out = -12810;
			3638: out = -12904;
			3639: out = -12967;
			3640: out = -13045;
			3641: out = -13118;
			3642: out = -13189;
			3643: out = -13260;
			3644: out = -13333;
			3645: out = -13388;
			3646: out = -13435;
			3647: out = -13509;
			3648: out = -13563;
			3649: out = -13611;
			3650: out = -13678;
			3651: out = -13732;
			3652: out = -13766;
			3653: out = -13817;
			3654: out = -13874;
			3655: out = -13917;
			3656: out = -13976;
			3657: out = -14017;
			3658: out = -14050;
			3659: out = -14078;
			3660: out = -14109;
			3661: out = -14166;
			3662: out = -14199;
			3663: out = -14240;
			3664: out = -14264;
			3665: out = -14295;
			3666: out = -14334;
			3667: out = -14359;
			3668: out = -14403;
			3669: out = -14422;
			3670: out = -14446;
			3671: out = -14469;
			3672: out = -14521;
			3673: out = -14579;
			3674: out = -14575;
			3675: out = -14571;
			3676: out = -14595;
			3677: out = -14606;
			3678: out = -14601;
			3679: out = -14629;
			3680: out = -14633;
			3681: out = -14641;
			3682: out = -14674;
			3683: out = -14652;
			3684: out = -14692;
			3685: out = -14689;
			3686: out = -14707;
			3687: out = -14695;
			3688: out = -14717;
			3689: out = -14694;
			3690: out = -14701;
			3691: out = -14712;
			3692: out = -14714;
			3693: out = -14717;
			3694: out = -14730;
			3695: out = -14713;
			3696: out = -14719;
			3697: out = -14719;
			3698: out = -14711;
			3699: out = -14726;
			3700: out = -14705;
			3701: out = -14705;
			3702: out = -14701;
			3703: out = -14696;
			3704: out = -14675;
			3705: out = -14671;
			3706: out = -14650;
			3707: out = -14654;
			3708: out = -14644;
			3709: out = -14642;
			3710: out = -14616;
			3711: out = -14609;
			3712: out = -14591;
			3713: out = -14584;
			3714: out = -14585;
			3715: out = -14562;
			3716: out = -14563;
			3717: out = -14535;
			3718: out = -14520;
			3719: out = -14508;
			3720: out = -14502;
			3721: out = -14481;
			3722: out = -14463;
			3723: out = -14437;
			3724: out = -14421;
			3725: out = -14404;
			3726: out = -14362;
			3727: out = -14378;
			3728: out = -14336;
			3729: out = -14307;
			3730: out = -14276;
			3731: out = -14268;
			3732: out = -14226;
			3733: out = -14201;
			3734: out = -14205;
			3735: out = -14156;
			3736: out = -14135;
			3737: out = -14119;
			3738: out = -14085;
			3739: out = -14052;
			3740: out = -14035;
			3741: out = -14002;
			3742: out = -13986;
			3743: out = -13969;
			3744: out = -13929;
			3745: out = -13899;
			3746: out = -13865;
			3747: out = -13820;
			3748: out = -13799;
			3749: out = -13760;
			3750: out = -13729;
			3751: out = -13709;
			3752: out = -13663;
			3753: out = -13614;
			3754: out = -13593;
			3755: out = -13560;
			3756: out = -13519;
			3757: out = -13437;
			3758: out = -13396;
			3759: out = -13368;
			3760: out = -13332;
			3761: out = -13285;
			3762: out = -13258;
			3763: out = -13199;
			3764: out = -13153;
			3765: out = -13098;
			3766: out = -13032;
			3767: out = -12979;
			3768: out = -12929;
			3769: out = -12875;
			3770: out = -12808;
			3771: out = -12747;
			3772: out = -12698;
			3773: out = -12627;
			3774: out = -12569;
			3775: out = -12495;
			3776: out = -12426;
			3777: out = -12348;
			3778: out = -12264;
			3779: out = -12219;
			3780: out = -12132;
			3781: out = -12041;
			3782: out = -11977;
			3783: out = -11895;
			3784: out = -11804;
			3785: out = -11730;
			3786: out = -11625;
			3787: out = -11553;
			3788: out = -11448;
			3789: out = -11343;
			3790: out = -11262;
			3791: out = -11155;
			3792: out = -11068;
			3793: out = -10950;
			3794: out = -10872;
			3795: out = -10779;
			3796: out = -10666;
			3797: out = -10566;
			3798: out = -10456;
			3799: out = -10368;
			3800: out = -10251;
			3801: out = -10144;
			3802: out = -10049;
			3803: out = -9934;
			3804: out = -9829;
			3805: out = -9728;
			3806: out = -9616;
			3807: out = -9503;
			3808: out = -9414;
			3809: out = -9306;
			3810: out = -9189;
			3811: out = -9074;
			3812: out = -8978;
			3813: out = -8858;
			3814: out = -8765;
			3815: out = -8656;
			3816: out = -8535;
			3817: out = -8434;
			3818: out = -8331;
			3819: out = -8250;
			3820: out = -8120;
			3821: out = -8041;
			3822: out = -7934;
			3823: out = -7825;
			3824: out = -7724;
			3825: out = -7626;
			3826: out = -7524;
			3827: out = -7421;
			3828: out = -7334;
			3829: out = -7222;
			3830: out = -7149;
			3831: out = -7050;
			3832: out = -6944;
			3833: out = -6852;
			3834: out = -6746;
			3835: out = -6669;
			3836: out = -6561;
			3837: out = -6489;
			3838: out = -6387;
			3839: out = -6310;
			3840: out = -6220;
			3841: out = -6138;
			3842: out = -6040;
			3843: out = -5959;
			3844: out = -5866;
			3845: out = -5781;
			3846: out = -5705;
			3847: out = -5617;
			3848: out = -5522;
			3849: out = -5464;
			3850: out = -5369;
			3851: out = -5283;
			3852: out = -5203;
			3853: out = -5137;
			3854: out = -5068;
			3855: out = -4968;
			3856: out = -4901;
			3857: out = -4852;
			3858: out = -4790;
			3859: out = -4703;
			3860: out = -4616;
			3861: out = -4563;
			3862: out = -4479;
			3863: out = -4407;
			3864: out = -4333;
			3865: out = -4274;
			3866: out = -4197;
			3867: out = -4134;
			3868: out = -4052;
			3869: out = -3996;
			3870: out = -3942;
			3871: out = -3875;
			3872: out = -3812;
			3873: out = -3743;
			3874: out = -3689;
			3875: out = -3608;
			3876: out = -3558;
			3877: out = -3504;
			3878: out = -3451;
			3879: out = -3377;
			3880: out = -3323;
			3881: out = -3276;
			3882: out = -3213;
			3883: out = -3166;
			3884: out = -3098;
			3885: out = -3062;
			3886: out = -2999;
			3887: out = -2897;
			3888: out = -2813;
			3889: out = -2713;
			3890: out = -2622;
			3891: out = -2525;
			3892: out = -2441;
			3893: out = -2344;
			3894: out = -2270;
			3895: out = -2159;
			3896: out = -2080;
			3897: out = -1997;
			3898: out = -1903;
			3899: out = -1829;
			3900: out = -1756;
			3901: out = -1673;
			3902: out = -1575;
			3903: out = -1517;
			3904: out = -1427;
			3905: out = -1371;
			3906: out = -1284;
			3907: out = -1209;
			3908: out = -1146;
			3909: out = -1062;
			3910: out = -993;
			3911: out = -926;
			3912: out = -854;
			3913: out = -787;
			3914: out = -723;
			3915: out = -641;
			3916: out = -590;
			3917: out = -534;
			3918: out = -475;
			3919: out = -387;
			3920: out = -330;
			3921: out = -258;
			3922: out = -208;
			3923: out = -146;
			3924: out = -86;
			3925: out = -41;
			3926: out = 32;
			3927: out = 90;
			3928: out = 136;
			3929: out = 205;
			3930: out = 265;
			3931: out = 317;
			3932: out = 391;
			3933: out = 438;
			3934: out = 470;
			3935: out = 538;
			3936: out = 600;
			3937: out = 655;
			3938: out = 723;
			3939: out = 762;
			3940: out = 820;
			3941: out = 869;
			3942: out = 926;
			3943: out = 1000;
			3944: out = 1057;
			3945: out = 1093;
			3946: out = 1151;
			3947: out = 1194;
			3948: out = 1247;
			3949: out = 1294;
			3950: out = 1344;
			3951: out = 1394;
			3952: out = 1459;
			3953: out = 1518;
			3954: out = 1556;
			3955: out = 1627;
			3956: out = 1674;
			3957: out = 1730;
			3958: out = 1778;
			3959: out = 1847;
			3960: out = 1888;
			3961: out = 1949;
			3962: out = 2006;
			3963: out = 2060;
			3964: out = 2112;
			3965: out = 2185;
			3966: out = 2246;
			3967: out = 2294;
			3968: out = 2339;
			3969: out = 2415;
			3970: out = 2465;
			3971: out = 2525;
			3972: out = 2600;
			3973: out = 2648;
			3974: out = 2726;
			3975: out = 2784;
			3976: out = 2850;
			3977: out = 2921;
			3978: out = 2994;
			3979: out = 3057;
			3980: out = 3117;
			3981: out = 3194;
			3982: out = 3281;
			3983: out = 3358;
			3984: out = 3430;
			3985: out = 3519;
			3986: out = 3594;
			3987: out = 3661;
			3988: out = 3753;
			3989: out = 3856;
			3990: out = 3932;
			3991: out = 4028;
			3992: out = 4116;
			3993: out = 4207;
			3994: out = 4291;
			3995: out = 4391;
			3996: out = 4479;
			3997: out = 4569;
			3998: out = 4660;
			3999: out = 4764;
			4000: out = 4855;
			4001: out = 4952;
			4002: out = 5049;
			4003: out = 5156;
			4004: out = 5246;
			4005: out = 5342;
			4006: out = 5441;
			4007: out = 5541;
			4008: out = 5639;
			4009: out = 5738;
			4010: out = 5850;
			4011: out = 5946;
			4012: out = 6025;
			4013: out = 6134;
			4014: out = 6237;
			4015: out = 6332;
			4016: out = 6444;
			4017: out = 6540;
			4018: out = 6635;
			4019: out = 6727;
			4020: out = 6826;
			4021: out = 6936;
			4022: out = 7018;
			4023: out = 7105;
			4024: out = 7179;
			4025: out = 7300;
			4026: out = 7383;
			4027: out = 7487;
			4028: out = 7580;
			4029: out = 7655;
			4030: out = 7740;
			4031: out = 7838;
			4032: out = 7913;
			4033: out = 7980;
			4034: out = 8079;
			4035: out = 8155;
			4036: out = 8249;
			4037: out = 8319;
			4038: out = 8421;
			4039: out = 8482;
			4040: out = 8561;
			4041: out = 8653;
			4042: out = 8714;
			4043: out = 8789;
			4044: out = 8874;
			4045: out = 8943;
			4046: out = 9020;
			4047: out = 9091;
			4048: out = 9162;
			4049: out = 9238;
			4050: out = 9303;
			4051: out = 9367;
			4052: out = 9433;
			4053: out = 9495;
			4054: out = 9562;
			4055: out = 9629;
			4056: out = 9693;
			4057: out = 9764;
			4058: out = 9828;
			4059: out = 9884;
			4060: out = 9937;
			4061: out = 10020;
			4062: out = 10068;
			4063: out = 10148;
			4064: out = 10192;
			4065: out = 10240;
			4066: out = 10310;
			4067: out = 10348;
			4068: out = 10421;
			4069: out = 10456;
			4070: out = 10524;
			4071: out = 10570;
			4072: out = 10636;
			4073: out = 10678;
			4074: out = 10726;
			4075: out = 10757;
			4076: out = 10828;
			4077: out = 10867;
			4078: out = 10921;
			4079: out = 10975;
			4080: out = 11019;
			4081: out = 11057;
			4082: out = 11101;
			4083: out = 11161;
			4084: out = 11201;
			4085: out = 11249;
			4086: out = 11287;
			4087: out = 11321;
			4088: out = 11363;
			4089: out = 11408;
			4090: out = 11460;
			4091: out = 11508;
			4092: out = 11547;
			4093: out = 11595;
			4094: out = 11616;
			4095: out = 11666;
			4096: out = 11708;
			4097: out = 11745;
			4098: out = 11776;
			4099: out = 11811;
			4100: out = 11856;
			4101: out = 11908;
			4102: out = 11943;
			4103: out = 11979;
			4104: out = 12013;
			4105: out = 12047;
			4106: out = 12085;
			4107: out = 12127;
			4108: out = 12163;
			4109: out = 12202;
			4110: out = 12220;
			4111: out = 12255;
			4112: out = 12307;
			4113: out = 12324;
			4114: out = 12369;
			4115: out = 12388;
			4116: out = 12415;
			4117: out = 12441;
			4118: out = 12442;
			4119: out = 12467;
			4120: out = 12489;
			4121: out = 12476;
			4122: out = 12435;
			4123: out = 12470;
			4124: out = 12452;
			4125: out = 12398;
			4126: out = 12403;
			4127: out = 12421;
			4128: out = 12421;
			4129: out = 12430;
			4130: out = 12419;
			4131: out = 12358;
			4132: out = 12380;
			4133: out = 12375;
			4134: out = 12378;
			4135: out = 12353;
			4136: out = 12344;
			4137: out = 12329;
			4138: out = 12278;
			4139: out = 12241;
			4140: out = 12246;
			4141: out = 12223;
			4142: out = 12210;
			4143: out = 12243;
			4144: out = 12248;
			4145: out = 12219;
			4146: out = 12163;
			4147: out = 12165;
			4148: out = 12169;
			4149: out = 12149;
			4150: out = 12174;
			4151: out = 12162;
			4152: out = 12108;
			4153: out = 12113;
			4154: out = 12110;
			4155: out = 12106;
			4156: out = 12144;
			4157: out = 12122;
			4158: out = 12047;
			4159: out = 12041;
			4160: out = 12012;
			4161: out = 12053;
			4162: out = 12052;
			4163: out = 12019;
			4164: out = 12020;
			4165: out = 12042;
			4166: out = 12044;
			4167: out = 12007;
			4168: out = 11965;
			4169: out = 11964;
			4170: out = 11919;
			4171: out = 11938;
			4172: out = 11953;
			4173: out = 11960;
			4174: out = 11955;
			4175: out = 11938;
			4176: out = 11927;
			4177: out = 11925;
			4178: out = 11893;
			4179: out = 11854;
			4180: out = 11835;
			4181: out = 11865;
			4182: out = 11791;
			4183: out = 11719;
			4184: out = 11711;
			4185: out = 11665;
			4186: out = 11659;
			4187: out = 11686;
			4188: out = 11692;
			4189: out = 11636;
			4190: out = 11619;
			4191: out = 11547;
			4192: out = 11517;
			4193: out = 11516;
			4194: out = 11480;
			4195: out = 11445;
			4196: out = 11439;
			4197: out = 11373;
			4198: out = 11359;
			4199: out = 11293;
			4200: out = 11213;
			4201: out = 11205;
			4202: out = 11199;
			4203: out = 11130;
			4204: out = 11026;
			4205: out = 11011;
			4206: out = 10979;
			4207: out = 10931;
			4208: out = 10864;
			4209: out = 10824;
			4210: out = 10779;
			4211: out = 10708;
			4212: out = 10601;
			4213: out = 10542;
			4214: out = 10489;
			4215: out = 10409;
			4216: out = 10345;
			4217: out = 10296;
			4218: out = 10233;
			4219: out = 10168;
			4220: out = 10108;
			4221: out = 10041;
			4222: out = 9959;
			4223: out = 9867;
			4224: out = 9789;
			4225: out = 9735;
			4226: out = 9636;
			4227: out = 9572;
			4228: out = 9476;
			4229: out = 9414;
			4230: out = 9351;
			4231: out = 9274;
			4232: out = 9187;
			4233: out = 9103;
			4234: out = 9023;
			4235: out = 8935;
			4236: out = 8870;
			4237: out = 8784;
			4238: out = 8710;
			4239: out = 8608;
			4240: out = 8547;
			4241: out = 8465;
			4242: out = 8365;
			4243: out = 8297;
			4244: out = 8234;
			4245: out = 8173;
			4246: out = 8048;
			4247: out = 7984;
			4248: out = 7909;
			4249: out = 7816;
			4250: out = 7729;
			4251: out = 7654;
			4252: out = 7586;
			4253: out = 7507;
			4254: out = 7434;
			4255: out = 7369;
			4256: out = 7282;
			4257: out = 7205;
			4258: out = 7129;
			4259: out = 7044;
			4260: out = 6974;
			4261: out = 6873;
			4262: out = 6791;
			4263: out = 6735;
			4264: out = 6660;
			4265: out = 6590;
			4266: out = 6498;
			4267: out = 6417;
			4268: out = 6356;
			4269: out = 6297;
			4270: out = 6233;
			4271: out = 6156;
			4272: out = 6081;
			4273: out = 5997;
			4274: out = 5918;
			4275: out = 5876;
			4276: out = 5808;
			4277: out = 5742;
			4278: out = 5664;
			4279: out = 5602;
			4280: out = 5528;
			4281: out = 5445;
			4282: out = 5394;
			4283: out = 5328;
			4284: out = 5253;
			4285: out = 5189;
			4286: out = 5128;
			4287: out = 5070;
			4288: out = 5000;
			4289: out = 4969;
			4290: out = 4888;
			4291: out = 4834;
			4292: out = 4769;
			4293: out = 4700;
			4294: out = 4652;
			4295: out = 4586;
			4296: out = 4507;
			4297: out = 4444;
			4298: out = 4388;
			4299: out = 4361;
			4300: out = 4280;
			4301: out = 4225;
			4302: out = 4176;
			4303: out = 4123;
			4304: out = 4065;
			4305: out = 4032;
			4306: out = 3958;
			4307: out = 3890;
			4308: out = 3833;
			4309: out = 3769;
			4310: out = 3752;
			4311: out = 3706;
			4312: out = 3643;
			4313: out = 3622;
			4314: out = 3568;
			4315: out = 3506;
			4316: out = 3459;
			4317: out = 3403;
			4318: out = 3366;
			4319: out = 3316;
			4320: out = 3286;
			4321: out = 3233;
			4322: out = 3180;
			4323: out = 3140;
			4324: out = 3103;
			4325: out = 3048;
			4326: out = 2996;
			4327: out = 2968;
			4328: out = 2933;
			4329: out = 2877;
			4330: out = 2844;
			4331: out = 2802;
			4332: out = 2737;
			4333: out = 2712;
			4334: out = 2673;
			4335: out = 2648;
			4336: out = 2607;
			4337: out = 2558;
			4338: out = 2527;
			4339: out = 2476;
			4340: out = 2446;
			4341: out = 2426;
			4342: out = 2376;
			4343: out = 2352;
			4344: out = 2294;
			4345: out = 2281;
			4346: out = 2247;
			4347: out = 2186;
			4348: out = 2134;
			4349: out = 2029;
			4350: out = 1950;
			4351: out = 1851;
			4352: out = 1772;
			4353: out = 1665;
			4354: out = 1584;
			4355: out = 1489;
			4356: out = 1417;
			4357: out = 1328;
			4358: out = 1228;
			4359: out = 1154;
			4360: out = 1058;
			4361: out = 974;
			4362: out = 895;
			4363: out = 831;
			4364: out = 749;
			4365: out = 669;
			4366: out = 616;
			4367: out = 527;
			4368: out = 448;
			4369: out = 386;
			4370: out = 303;
			4371: out = 246;
			4372: out = 154;
			4373: out = 89;
			4374: out = 31;
			4375: out = -38;
			4376: out = -95;
			4377: out = -161;
			4378: out = -238;
			4379: out = -321;
			4380: out = -358;
			4381: out = -423;
			4382: out = -496;
			4383: out = -545;
			4384: out = -619;
			4385: out = -682;
			4386: out = -748;
			4387: out = -799;
			4388: out = -859;
			4389: out = -913;
			4390: out = -968;
			4391: out = -1019;
			4392: out = -1056;
			4393: out = -1120;
			4394: out = -1192;
			4395: out = -1260;
			4396: out = -1321;
			4397: out = -1377;
			4398: out = -1447;
			4399: out = -1500;
			4400: out = -1546;
			4401: out = -1591;
			4402: out = -1659;
			4403: out = -1713;
			4404: out = -1759;
			4405: out = -1809;
			4406: out = -1870;
			4407: out = -1912;
			4408: out = -1969;
			4409: out = -2025;
			4410: out = -2077;
			4411: out = -2147;
			4412: out = -2194;
			4413: out = -2234;
			4414: out = -2311;
			4415: out = -2356;
			4416: out = -2406;
			4417: out = -2453;
			4418: out = -2509;
			4419: out = -2559;
			4420: out = -2607;
			4421: out = -2651;
			4422: out = -2718;
			4423: out = -2775;
			4424: out = -2812;
			4425: out = -2872;
			4426: out = -2931;
			4427: out = -2995;
			4428: out = -3034;
			4429: out = -3084;
			4430: out = -3143;
			4431: out = -3198;
			4432: out = -3256;
			4433: out = -3319;
			4434: out = -3389;
			4435: out = -3452;
			4436: out = -3509;
			4437: out = -3596;
			4438: out = -3655;
			4439: out = -3718;
			4440: out = -3787;
			4441: out = -3852;
			4442: out = -3913;
			4443: out = -3992;
			4444: out = -4060;
			4445: out = -4143;
			4446: out = -4223;
			4447: out = -4279;
			4448: out = -4369;
			4449: out = -4446;
			4450: out = -4516;
			4451: out = -4585;
			4452: out = -4684;
			4453: out = -4743;
			4454: out = -4821;
			4455: out = -4913;
			4456: out = -4994;
			4457: out = -5074;
			4458: out = -5173;
			4459: out = -5253;
			4460: out = -5346;
			4461: out = -5452;
			4462: out = -5532;
			4463: out = -5624;
			4464: out = -5722;
			4465: out = -5815;
			4466: out = -5907;
			4467: out = -6015;
			4468: out = -6128;
			4469: out = -6213;
			4470: out = -6308;
			4471: out = -6412;
			4472: out = -6525;
			4473: out = -6631;
			4474: out = -6746;
			4475: out = -6843;
			4476: out = -6935;
			4477: out = -7048;
			4478: out = -7158;
			4479: out = -7281;
			4480: out = -7381;
			4481: out = -7495;
			4482: out = -7605;
			4483: out = -7720;
			4484: out = -7835;
			4485: out = -7942;
			4486: out = -8051;
			4487: out = -8167;
			4488: out = -8254;
			4489: out = -8362;
			4490: out = -8455;
			4491: out = -8573;
			4492: out = -8663;
			4493: out = -8774;
			4494: out = -8874;
			4495: out = -8950;
			4496: out = -9043;
			4497: out = -9139;
			4498: out = -9231;
			4499: out = -9313;
			4500: out = -9402;
			4501: out = -9476;
			4502: out = -9552;
			4503: out = -9628;
			4504: out = -9706;
			4505: out = -9780;
			4506: out = -9878;
			4507: out = -9939;
			4508: out = -10032;
			4509: out = -10108;
			4510: out = -10171;
			4511: out = -10252;
			4512: out = -10309;
			4513: out = -10397;
			4514: out = -10452;
			4515: out = -10522;
			4516: out = -10577;
			4517: out = -10649;
			4518: out = -10703;
			4519: out = -10766;
			4520: out = -10818;
			4521: out = -10889;
			4522: out = -10918;
			4523: out = -10980;
			4524: out = -11039;
			4525: out = -11090;
			4526: out = -11120;
			4527: out = -11196;
			4528: out = -11225;
			4529: out = -11252;
			4530: out = -11315;
			4531: out = -11354;
			4532: out = -11401;
			4533: out = -11427;
			4534: out = -11462;
			4535: out = -11491;
			4536: out = -11539;
			4537: out = -11577;
			4538: out = -11590;
			4539: out = -11631;
			4540: out = -11649;
			4541: out = -11682;
			4542: out = -11719;
			4543: out = -11742;
			4544: out = -11772;
			4545: out = -11781;
			4546: out = -11806;
			4547: out = -11835;
			4548: out = -11864;
			4549: out = -11870;
			4550: out = -11890;
			4551: out = -11907;
			4552: out = -11915;
			4553: out = -11919;
			4554: out = -11957;
			4555: out = -11958;
			4556: out = -11970;
			4557: out = -11969;
			4558: out = -12007;
			4559: out = -11997;
			4560: out = -12014;
			4561: out = -12014;
			4562: out = -12020;
			4563: out = -12010;
			4564: out = -12036;
			4565: out = -12036;
			4566: out = -12036;
			4567: out = -12047;
			4568: out = -12051;
			4569: out = -12055;
			4570: out = -12091;
			4571: out = -12079;
			4572: out = -12073;
			4573: out = -12064;
			4574: out = -12059;
			4575: out = -12068;
			4576: out = -12043;
			4577: out = -12049;
			4578: out = -12043;
			4579: out = -12041;
			4580: out = -12039;
			4581: out = -12021;
			4582: out = -12028;
			4583: out = -12023;
			4584: out = -12012;
			4585: out = -12013;
			4586: out = -11989;
			4587: out = -11984;
			4588: out = -11971;
			4589: out = -11973;
			4590: out = -11968;
			4591: out = -11943;
			4592: out = -11936;
			4593: out = -11919;
			4594: out = -11908;
			4595: out = -11891;
			4596: out = -11887;
			4597: out = -11849;
			4598: out = -11847;
			4599: out = -11835;
			4600: out = -11825;
			4601: out = -11812;
			4602: out = -11785;
			4603: out = -11764;
			4604: out = -11756;
			4605: out = -11732;
			4606: out = -11707;
			4607: out = -11707;
			4608: out = -11684;
			4609: out = -11652;
			4610: out = -11650;
			4611: out = -11623;
			4612: out = -11613;
			4613: out = -11587;
			4614: out = -11559;
			4615: out = -11554;
			4616: out = -11511;
			4617: out = -11493;
			4618: out = -11473;
			4619: out = -11448;
			4620: out = -11420;
			4621: out = -11406;
			4622: out = -11363;
			4623: out = -11343;
			4624: out = -11330;
			4625: out = -11303;
			4626: out = -11254;
			4627: out = -11236;
			4628: out = -11216;
			4629: out = -11180;
			4630: out = -11150;
			4631: out = -11134;
			4632: out = -11112;
			4633: out = -11075;
			4634: out = -11032;
			4635: out = -11032;
			4636: out = -10982;
			4637: out = -10943;
			4638: out = -10924;
			4639: out = -10889;
			4640: out = -10837;
			4641: out = -10818;
			4642: out = -10775;
			4643: out = -10738;
			4644: out = -10702;
			4645: out = -10662;
			4646: out = -10618;
			4647: out = -10585;
			4648: out = -10537;
			4649: out = -10489;
			4650: out = -10431;
			4651: out = -10411;
			4652: out = -10340;
			4653: out = -10302;
			4654: out = -10231;
			4655: out = -10175;
			4656: out = -10142;
			4657: out = -10079;
			4658: out = -10024;
			4659: out = -9965;
			4660: out = -9919;
			4661: out = -9838;
			4662: out = -9793;
			4663: out = -9700;
			4664: out = -9653;
			4665: out = -9586;
			4666: out = -9519;
			4667: out = -9445;
			4668: out = -9371;
			4669: out = -9300;
			4670: out = -9221;
			4671: out = -9151;
			4672: out = -9079;
			4673: out = -9002;
			4674: out = -8920;
			4675: out = -8834;
			4676: out = -8762;
			4677: out = -8676;
			4678: out = -8589;
			4679: out = -8512;
			4680: out = -8404;
			4681: out = -8345;
			4682: out = -8256;
			4683: out = -8152;
			4684: out = -8084;
			4685: out = -7986;
			4686: out = -7901;
			4687: out = -7815;
			4688: out = -7740;
			4689: out = -7646;
			4690: out = -7555;
			4691: out = -7482;
			4692: out = -7380;
			4693: out = -7298;
			4694: out = -7214;
			4695: out = -7139;
			4696: out = -7045;
			4697: out = -6971;
			4698: out = -6862;
			4699: out = -6800;
			4700: out = -6718;
			4701: out = -6628;
			4702: out = -6553;
			4703: out = -6445;
			4704: out = -6398;
			4705: out = -6302;
			4706: out = -6222;
			4707: out = -6135;
			4708: out = -6048;
			4709: out = -5973;
			4710: out = -5895;
			4711: out = -5830;
			4712: out = -5748;
			4713: out = -5664;
			4714: out = -5583;
			4715: out = -5510;
			4716: out = -5427;
			4717: out = -5357;
			4718: out = -5283;
			4719: out = -5199;
			4720: out = -5129;
			4721: out = -5061;
			4722: out = -4978;
			4723: out = -4916;
			4724: out = -4831;
			4725: out = -4766;
			4726: out = -4693;
			4727: out = -4611;
			4728: out = -4574;
			4729: out = -4483;
			4730: out = -4423;
			4731: out = -4360;
			4732: out = -4293;
			4733: out = -4227;
			4734: out = -4172;
			4735: out = -4109;
			4736: out = -4045;
			4737: out = -3982;
			4738: out = -3917;
			4739: out = -3868;
			4740: out = -3805;
			4741: out = -3742;
			4742: out = -3681;
			4743: out = -3626;
			4744: out = -3571;
			4745: out = -3517;
			4746: out = -3453;
			4747: out = -3413;
			4748: out = -3343;
			4749: out = -3290;
			4750: out = -3250;
			4751: out = -3178;
			4752: out = -3144;
			4753: out = -3078;
			4754: out = -3035;
			4755: out = -2991;
			4756: out = -2950;
			4757: out = -2888;
			4758: out = -2834;
			4759: out = -2796;
			4760: out = -2738;
			4761: out = -2682;
			4762: out = -2642;
			4763: out = -2605;
			4764: out = -2561;
			4765: out = -2503;
			4766: out = -2465;
			4767: out = -2421;
			4768: out = -2382;
			4769: out = -2339;
			4770: out = -2276;
			4771: out = -2206;
			4772: out = -2134;
			4773: out = -2044;
			4774: out = -1980;
			4775: out = -1889;
			4776: out = -1823;
			4777: out = -1754;
			4778: out = -1682;
			4779: out = -1615;
			4780: out = -1552;
			4781: out = -1474;
			4782: out = -1406;
			4783: out = -1351;
			4784: out = -1279;
			4785: out = -1225;
			4786: out = -1153;
			4787: out = -1102;
			4788: out = -1036;
			4789: out = -973;
			4790: out = -915;
			4791: out = -847;
			4792: out = -802;
			4793: out = -740;
			4794: out = -680;
			4795: out = -635;
			4796: out = -577;
			4797: out = -516;
			4798: out = -469;
			4799: out = -411;
			4800: out = -348;
			4801: out = -306;
			4802: out = -264;
			4803: out = -210;
			4804: out = -147;
			4805: out = -102;
			4806: out = -61;
			4807: out = -19;
			4808: out = 27;
			4809: out = 88;
			4810: out = 125;
			4811: out = 167;
			4812: out = 227;
			4813: out = 270;
			4814: out = 317;
			4815: out = 349;
			4816: out = 401;
			4817: out = 438;
			4818: out = 490;
			4819: out = 529;
			4820: out = 574;
			4821: out = 625;
			4822: out = 669;
			4823: out = 707;
			4824: out = 756;
			4825: out = 796;
			4826: out = 835;
			4827: out = 890;
			4828: out = 920;
			4829: out = 961;
			4830: out = 1000;
			4831: out = 1047;
			4832: out = 1092;
			4833: out = 1133;
			4834: out = 1185;
			4835: out = 1213;
			4836: out = 1276;
			4837: out = 1291;
			4838: out = 1350;
			4839: out = 1390;
			4840: out = 1436;
			4841: out = 1485;
			4842: out = 1536;
			4843: out = 1571;
			4844: out = 1607;
			4845: out = 1648;
			4846: out = 1697;
			4847: out = 1724;
			4848: out = 1774;
			4849: out = 1823;
			4850: out = 1859;
			4851: out = 1925;
			4852: out = 1953;
			4853: out = 2014;
			4854: out = 2051;
			4855: out = 2105;
			4856: out = 2152;
			4857: out = 2198;
			4858: out = 2245;
			4859: out = 2293;
			4860: out = 2338;
			4861: out = 2397;
			4862: out = 2448;
			4863: out = 2514;
			4864: out = 2564;
			4865: out = 2628;
			4866: out = 2690;
			4867: out = 2756;
			4868: out = 2805;
			4869: out = 2873;
			4870: out = 2933;
			4871: out = 2994;
			4872: out = 3069;
			4873: out = 3129;
			4874: out = 3199;
			4875: out = 3276;
			4876: out = 3340;
			4877: out = 3404;
			4878: out = 3472;
			4879: out = 3556;
			4880: out = 3618;
			4881: out = 3676;
			4882: out = 3771;
			4883: out = 3842;
			4884: out = 3926;
			4885: out = 3994;
			4886: out = 4096;
			4887: out = 4151;
			4888: out = 4234;
			4889: out = 4318;
			4890: out = 4401;
			4891: out = 4463;
			4892: out = 4560;
			4893: out = 4631;
			4894: out = 4714;
			4895: out = 4795;
			4896: out = 4884;
			4897: out = 4963;
			4898: out = 5046;
			4899: out = 5118;
			4900: out = 5201;
			4901: out = 5285;
			4902: out = 5356;
			4903: out = 5442;
			4904: out = 5522;
			4905: out = 5583;
			4906: out = 5681;
			4907: out = 5763;
			4908: out = 5832;
			4909: out = 5919;
			4910: out = 5982;
			4911: out = 6061;
			4912: out = 6125;
			4913: out = 6206;
			4914: out = 6282;
			4915: out = 6346;
			4916: out = 6423;
			4917: out = 6470;
			4918: out = 6554;
			4919: out = 6621;
			4920: out = 6692;
			4921: out = 6741;
			4922: out = 6819;
			4923: out = 6883;
			4924: out = 6940;
			4925: out = 7014;
			4926: out = 7071;
			4927: out = 7146;
			4928: out = 7188;
			4929: out = 7252;
			4930: out = 7320;
			4931: out = 7368;
			4932: out = 7432;
			4933: out = 7482;
			4934: out = 7548;
			4935: out = 7613;
			4936: out = 7669;
			4937: out = 7718;
			4938: out = 7797;
			4939: out = 7834;
			4940: out = 7894;
			4941: out = 7941;
			4942: out = 8010;
			4943: out = 8060;
			4944: out = 8115;
			4945: out = 8158;
			4946: out = 8228;
			4947: out = 8260;
			4948: out = 8333;
			4949: out = 8361;
			4950: out = 8408;
			4951: out = 8458;
			4952: out = 8497;
			4953: out = 8550;
			4954: out = 8590;
			4955: out = 8630;
			4956: out = 8661;
			4957: out = 8717;
			4958: out = 8757;
			4959: out = 8796;
			4960: out = 8843;
			4961: out = 8864;
			4962: out = 8921;
			4963: out = 8944;
			4964: out = 8990;
			4965: out = 9045;
			4966: out = 9068;
			4967: out = 9098;
			4968: out = 9150;
			4969: out = 9193;
			4970: out = 9231;
			4971: out = 9271;
			4972: out = 9308;
			4973: out = 9352;
			4974: out = 9377;
			4975: out = 9409;
			4976: out = 9459;
			4977: out = 9484;
			4978: out = 9527;
			4979: out = 9543;
			4980: out = 9597;
			4981: out = 9635;
			4982: out = 9659;
			4983: out = 9692;
			4984: out = 9730;
			4985: out = 9765;
			4986: out = 9781;
			4987: out = 9816;
			4988: out = 9850;
			4989: out = 9882;
			4990: out = 9907;
			4991: out = 9934;
			4992: out = 9977;
			4993: out = 9996;
			4994: out = 10019;
			4995: out = 10055;
			4996: out = 10085;
			4997: out = 10104;
			4998: out = 10134;
			4999: out = 10157;
			5000: out = 10182;
			5001: out = 10216;
			5002: out = 10227;
			5003: out = 10244;
			5004: out = 10267;
			5005: out = 10285;
			5006: out = 10281;
			5007: out = 10265;
			5008: out = 10280;
			5009: out = 10231;
			5010: out = 10233;
			5011: out = 10272;
			5012: out = 10246;
			5013: out = 10229;
			5014: out = 10180;
			5015: out = 10192;
			5016: out = 10148;
			5017: out = 10159;
			5018: out = 10173;
			5019: out = 10151;
			5020: out = 10157;
			5021: out = 10131;
			5022: out = 10125;
			5023: out = 10106;
			5024: out = 10143;
			5025: out = 10124;
			5026: out = 10091;
			5027: out = 10114;
			5028: out = 10094;
			5029: out = 10111;
			5030: out = 10123;
			5031: out = 10090;
			5032: out = 10102;
			5033: out = 10084;
			5034: out = 10087;
			5035: out = 10074;
			5036: out = 10065;
			5037: out = 10054;
			5038: out = 10053;
			5039: out = 10025;
			5040: out = 10031;
			5041: out = 10025;
			5042: out = 10028;
			5043: out = 10036;
			5044: out = 10004;
			5045: out = 10021;
			5046: out = 9995;
			5047: out = 10009;
			5048: out = 10002;
			5049: out = 9970;
			5050: out = 9937;
			5051: out = 9941;
			5052: out = 9952;
			5053: out = 9974;
			5054: out = 9967;
			5055: out = 9984;
			5056: out = 9976;
			5057: out = 9941;
			5058: out = 9937;
			5059: out = 9927;
			5060: out = 9915;
			5061: out = 9895;
			5062: out = 9856;
			5063: out = 9829;
			5064: out = 9831;
			5065: out = 9820;
			5066: out = 9791;
			5067: out = 9748;
			5068: out = 9747;
			5069: out = 9745;
			5070: out = 9757;
			5071: out = 9746;
			5072: out = 9730;
			5073: out = 9701;
			5074: out = 9627;
			5075: out = 9655;
			5076: out = 9594;
			5077: out = 9590;
			5078: out = 9574;
			5079: out = 9528;
			5080: out = 9529;
			5081: out = 9487;
			5082: out = 9486;
			5083: out = 9451;
			5084: out = 9439;
			5085: out = 9412;
			5086: out = 9399;
			5087: out = 9333;
			5088: out = 9294;
			5089: out = 9247;
			5090: out = 9185;
			5091: out = 9168;
			5092: out = 9125;
			5093: out = 9059;
			5094: out = 9011;
			5095: out = 8990;
			5096: out = 8914;
			5097: out = 8890;
			5098: out = 8836;
			5099: out = 8782;
			5100: out = 8716;
			5101: out = 8659;
			5102: out = 8631;
			5103: out = 8583;
			5104: out = 8548;
			5105: out = 8478;
			5106: out = 8423;
			5107: out = 8362;
			5108: out = 8296;
			5109: out = 8237;
			5110: out = 8186;
			5111: out = 8124;
			5112: out = 8074;
			5113: out = 8000;
			5114: out = 7910;
			5115: out = 7852;
			5116: out = 7775;
			5117: out = 7722;
			5118: out = 7686;
			5119: out = 7587;
			5120: out = 7519;
			5121: out = 7465;
			5122: out = 7369;
			5123: out = 7315;
			5124: out = 7285;
			5125: out = 7205;
			5126: out = 7136;
			5127: out = 7080;
			5128: out = 6987;
			5129: out = 6938;
			5130: out = 6864;
			5131: out = 6795;
			5132: out = 6744;
			5133: out = 6694;
			5134: out = 6619;
			5135: out = 6554;
			5136: out = 6483;
			5137: out = 6429;
			5138: out = 6353;
			5139: out = 6279;
			5140: out = 6240;
			5141: out = 6158;
			5142: out = 6060;
			5143: out = 6021;
			5144: out = 5965;
			5145: out = 5910;
			5146: out = 5830;
			5147: out = 5781;
			5148: out = 5722;
			5149: out = 5638;
			5150: out = 5577;
			5151: out = 5550;
			5152: out = 5477;
			5153: out = 5400;
			5154: out = 5349;
			5155: out = 5284;
			5156: out = 5231;
			5157: out = 5172;
			5158: out = 5104;
			5159: out = 5050;
			5160: out = 4988;
			5161: out = 4938;
			5162: out = 4882;
			5163: out = 4852;
			5164: out = 4769;
			5165: out = 4710;
			5166: out = 4653;
			5167: out = 4619;
			5168: out = 4527;
			5169: out = 4470;
			5170: out = 4429;
			5171: out = 4372;
			5172: out = 4326;
			5173: out = 4286;
			5174: out = 4229;
			5175: out = 4183;
			5176: out = 4107;
			5177: out = 4080;
			5178: out = 4014;
			5179: out = 3969;
			5180: out = 3910;
			5181: out = 3872;
			5182: out = 3802;
			5183: out = 3765;
			5184: out = 3726;
			5185: out = 3678;
			5186: out = 3630;
			5187: out = 3580;
			5188: out = 3543;
			5189: out = 3501;
			5190: out = 3450;
			5191: out = 3391;
			5192: out = 3343;
			5193: out = 3334;
			5194: out = 3269;
			5195: out = 3213;
			5196: out = 3190;
			5197: out = 3139;
			5198: out = 3087;
			5199: out = 3063;
			5200: out = 3038;
			5201: out = 2976;
			5202: out = 2939;
			5203: out = 2896;
			5204: out = 2834;
			5205: out = 2803;
			5206: out = 2768;
			5207: out = 2742;
			5208: out = 2694;
			5209: out = 2679;
			5210: out = 2651;
			5211: out = 2602;
			5212: out = 2561;
			5213: out = 2524;
			5214: out = 2502;
			5215: out = 2469;
			5216: out = 2429;
			5217: out = 2383;
			5218: out = 2347;
			5219: out = 2325;
			5220: out = 2266;
			5221: out = 2240;
			5222: out = 2202;
			5223: out = 2180;
			5224: out = 2147;
			5225: out = 2108;
			5226: out = 2073;
			5227: out = 2051;
			5228: out = 2037;
			5229: out = 1982;
			5230: out = 1962;
			5231: out = 1918;
			5232: out = 1878;
			5233: out = 1867;
			5234: out = 1835;
			5235: out = 1816;
			5236: out = 1796;
			5237: out = 1729;
			5238: out = 1650;
			5239: out = 1576;
			5240: out = 1493;
			5241: out = 1425;
			5242: out = 1345;
			5243: out = 1260;
			5244: out = 1204;
			5245: out = 1115;
			5246: out = 1061;
			5247: out = 985;
			5248: out = 925;
			5249: out = 862;
			5250: out = 787;
			5251: out = 720;
			5252: out = 654;
			5253: out = 596;
			5254: out = 537;
			5255: out = 475;
			5256: out = 416;
			5257: out = 372;
			5258: out = 304;
			5259: out = 239;
			5260: out = 202;
			5261: out = 151;
			5262: out = 96;
			5263: out = 31;
			5264: out = -32;
			5265: out = -91;
			5266: out = -148;
			5267: out = -211;
			5268: out = -257;
			5269: out = -302;
			5270: out = -365;
			5271: out = -411;
			5272: out = -469;
			5273: out = -521;
			5274: out = -566;
			5275: out = -626;
			5276: out = -680;
			5277: out = -735;
			5278: out = -787;
			5279: out = -833;
			5280: out = -886;
			5281: out = -927;
			5282: out = -978;
			5283: out = -1033;
			5284: out = -1081;
			5285: out = -1125;
			5286: out = -1175;
			5287: out = -1221;
			5288: out = -1269;
			5289: out = -1294;
			5290: out = -1314;
			5291: out = -1394;
			5292: out = -1429;
			5293: out = -1477;
			5294: out = -1529;
			5295: out = -1582;
			5296: out = -1617;
			5297: out = -1664;
			5298: out = -1699;
			5299: out = -1728;
			5300: out = -1800;
			5301: out = -1817;
			5302: out = -1870;
			5303: out = -1914;
			5304: out = -1956;
			5305: out = -1991;
			5306: out = -2051;
			5307: out = -2105;
			5308: out = -2149;
			5309: out = -2173;
			5310: out = -2227;
			5311: out = -2261;
			5312: out = -2309;
			5313: out = -2372;
			5314: out = -2417;
			5315: out = -2459;
			5316: out = -2498;
			5317: out = -2547;
			5318: out = -2618;
			5319: out = -2652;
			5320: out = -2705;
			5321: out = -2752;
			5322: out = -2796;
			5323: out = -2841;
			5324: out = -2903;
			5325: out = -2962;
			5326: out = -3019;
			5327: out = -3059;
			5328: out = -3111;
			5329: out = -3177;
			5330: out = -3228;
			5331: out = -3281;
			5332: out = -3350;
			5333: out = -3382;
			5334: out = -3458;
			5335: out = -3509;
			5336: out = -3572;
			5337: out = -3631;
			5338: out = -3696;
			5339: out = -3756;
			5340: out = -3820;
			5341: out = -3895;
			5342: out = -3963;
			5343: out = -4024;
			5344: out = -4090;
			5345: out = -4159;
			5346: out = -4225;
			5347: out = -4291;
			5348: out = -4381;
			5349: out = -4445;
			5350: out = -4519;
			5351: out = -4578;
			5352: out = -4682;
			5353: out = -4770;
			5354: out = -4831;
			5355: out = -4914;
			5356: out = -5003;
			5357: out = -5080;
			5358: out = -5166;
			5359: out = -5260;
			5360: out = -5342;
			5361: out = -5436;
			5362: out = -5510;
			5363: out = -5603;
			5364: out = -5711;
			5365: out = -5803;
			5366: out = -5875;
			5367: out = -5980;
			5368: out = -6071;
			5369: out = -6145;
			5370: out = -6235;
			5371: out = -6328;
			5372: out = -6411;
			5373: out = -6507;
			5374: out = -6583;
			5375: out = -6688;
			5376: out = -6758;
			5377: out = -6861;
			5378: out = -6949;
			5379: out = -7032;
			5380: out = -7128;
			5381: out = -7203;
			5382: out = -7292;
			5383: out = -7378;
			5384: out = -7449;
			5385: out = -7527;
			5386: out = -7604;
			5387: out = -7673;
			5388: out = -7740;
			5389: out = -7827;
			5390: out = -7874;
			5391: out = -7959;
			5392: out = -8022;
			5393: out = -8093;
			5394: out = -8161;
			5395: out = -8226;
			5396: out = -8292;
			5397: out = -8335;
			5398: out = -8397;
			5399: out = -8461;
			5400: out = -8515;
			5401: out = -8581;
			5402: out = -8644;
			5403: out = -8682;
			5404: out = -8746;
			5405: out = -8793;
			5406: out = -8846;
			5407: out = -8883;
			5408: out = -8940;
			5409: out = -8986;
			5410: out = -9027;
			5411: out = -9085;
			5412: out = -9118;
			5413: out = -9168;
			5414: out = -9196;
			5415: out = -9240;
			5416: out = -9280;
			5417: out = -9322;
			5418: out = -9352;
			5419: out = -9393;
			5420: out = -9400;
			5421: out = -9453;
			5422: out = -9476;
			5423: out = -9518;
			5424: out = -9538;
			5425: out = -9559;
			5426: out = -9595;
			5427: out = -9619;
			5428: out = -9643;
			5429: out = -9681;
			5430: out = -9690;
			5431: out = -9707;
			5432: out = -9726;
			5433: out = -9743;
			5434: out = -9772;
			5435: out = -9779;
			5436: out = -9796;
			5437: out = -9816;
			5438: out = -9829;
			5439: out = -9832;
			5440: out = -9860;
			5441: out = -9865;
			5442: out = -9867;
			5443: out = -9895;
			5444: out = -9895;
			5445: out = -9897;
			5446: out = -9924;
			5447: out = -9920;
			5448: out = -9936;
			5449: out = -9934;
			5450: out = -9936;
			5451: out = -9960;
			5452: out = -9977;
			5453: out = -9957;
			5454: out = -9967;
			5455: out = -9965;
			5456: out = -9959;
			5457: out = -9971;
			5458: out = -9972;
			5459: out = -9967;
			5460: out = -9961;
			5461: out = -9972;
			5462: out = -9968;
			5463: out = -9955;
			5464: out = -9962;
			5465: out = -9958;
			5466: out = -9952;
			5467: out = -9974;
			5468: out = -9968;
			5469: out = -9948;
			5470: out = -9943;
			5471: out = -9935;
			5472: out = -9911;
			5473: out = -9910;
			5474: out = -9903;
			5475: out = -9898;
			5476: out = -9885;
			5477: out = -9873;
			5478: out = -9865;
			5479: out = -9856;
			5480: out = -9847;
			5481: out = -9836;
			5482: out = -9839;
			5483: out = -9814;
			5484: out = -9806;
			5485: out = -9791;
			5486: out = -9783;
			5487: out = -9764;
			5488: out = -9749;
			5489: out = -9737;
			5490: out = -9728;
			5491: out = -9701;
			5492: out = -9686;
			5493: out = -9683;
			5494: out = -9657;
			5495: out = -9646;
			5496: out = -9625;
			5497: out = -9607;
			5498: out = -9591;
			5499: out = -9567;
			5500: out = -9566;
			5501: out = -9528;
			5502: out = -9529;
			5503: out = -9494;
			5504: out = -9492;
			5505: out = -9473;
			5506: out = -9456;
			5507: out = -9426;
			5508: out = -9401;
			5509: out = -9389;
			5510: out = -9361;
			5511: out = -9351;
			5512: out = -9333;
			5513: out = -9304;
			5514: out = -9271;
			5515: out = -9267;
			5516: out = -9235;
			5517: out = -9233;
			5518: out = -9186;
			5519: out = -9163;
			5520: out = -9143;
			5521: out = -9114;
			5522: out = -9085;
			5523: out = -9054;
			5524: out = -9053;
			5525: out = -9011;
			5526: out = -8972;
			5527: out = -8958;
			5528: out = -8943;
			5529: out = -8880;
			5530: out = -8871;
			5531: out = -8817;
			5532: out = -8799;
			5533: out = -8771;
			5534: out = -8729;
			5535: out = -8708;
			5536: out = -8656;
			5537: out = -8622;
			5538: out = -8599;
			5539: out = -8557;
			5540: out = -8521;
			5541: out = -8470;
			5542: out = -8431;
			5543: out = -8388;
			5544: out = -8338;
			5545: out = -8303;
			5546: out = -8266;
			5547: out = -8215;
			5548: out = -8158;
			5549: out = -8120;
			5550: out = -8059;
			5551: out = -8013;
			5552: out = -7956;
			5553: out = -7896;
			5554: out = -7835;
			5555: out = -7782;
			5556: out = -7731;
			5557: out = -7659;
			5558: out = -7623;
			5559: out = -7555;
			5560: out = -7497;
			5561: out = -7428;
			5562: out = -7375;
			5563: out = -7315;
			5564: out = -7244;
			5565: out = -7174;
			5566: out = -7119;
			5567: out = -7035;
			5568: out = -6967;
			5569: out = -6902;
			5570: out = -6832;
			5571: out = -6759;
			5572: out = -6690;
			5573: out = -6615;
			5574: out = -6535;
			5575: out = -6483;
			5576: out = -6398;
			5577: out = -6332;
			5578: out = -6266;
			5579: out = -6189;
			5580: out = -6121;
			5581: out = -6043;
			5582: out = -5973;
			5583: out = -5902;
			5584: out = -5842;
			5585: out = -5770;
			5586: out = -5701;
			5587: out = -5622;
			5588: out = -5558;
			5589: out = -5501;
			5590: out = -5425;
			5591: out = -5363;
			5592: out = -5294;
			5593: out = -5231;
			5594: out = -5158;
			5595: out = -5090;
			5596: out = -5039;
			5597: out = -4949;
			5598: out = -4898;
			5599: out = -4832;
			5600: out = -4766;
			5601: out = -4710;
			5602: out = -4634;
			5603: out = -4566;
			5604: out = -4505;
			5605: out = -4447;
			5606: out = -4375;
			5607: out = -4322;
			5608: out = -4269;
			5609: out = -4207;
			5610: out = -4137;
			5611: out = -4077;
			5612: out = -4027;
			5613: out = -3970;
			5614: out = -3901;
			5615: out = -3851;
			5616: out = -3790;
			5617: out = -3746;
			5618: out = -3675;
			5619: out = -3626;
			5620: out = -3577;
			5621: out = -3504;
			5622: out = -3461;
			5623: out = -3417;
			5624: out = -3356;
			5625: out = -3307;
			5626: out = -3256;
			5627: out = -3203;
			5628: out = -3148;
			5629: out = -3099;
			5630: out = -3061;
			5631: out = -3010;
			5632: out = -2953;
			5633: out = -2905;
			5634: out = -2864;
			5635: out = -2813;
			5636: out = -2781;
			5637: out = -2728;
			5638: out = -2682;
			5639: out = -2631;
			5640: out = -2596;
			5641: out = -2554;
			5642: out = -2510;
			5643: out = -2467;
			5644: out = -2436;
			5645: out = -2384;
			5646: out = -2344;
			5647: out = -2309;
			5648: out = -2266;
			5649: out = -2228;
			5650: out = -2193;
			5651: out = -2155;
			5652: out = -2126;
			5653: out = -2081;
			5654: out = -2058;
			5655: out = -2007;
			5656: out = -1970;
			5657: out = -1936;
			5658: out = -1900;
			5659: out = -1865;
			5660: out = -1813;
			5661: out = -1745;
			5662: out = -1682;
			5663: out = -1613;
			5664: out = -1566;
			5665: out = -1495;
			5666: out = -1442;
			5667: out = -1386;
			5668: out = -1314;
			5669: out = -1269;
			5670: out = -1203;
			5671: out = -1152;
			5672: out = -1095;
			5673: out = -1038;
			5674: out = -989;
			5675: out = -927;
			5676: out = -900;
			5677: out = -829;
			5678: out = -780;
			5679: out = -742;
			5680: out = -680;
			5681: out = -643;
			5682: out = -595;
			5683: out = -551;
			5684: out = -499;
			5685: out = -448;
			5686: out = -411;
			5687: out = -380;
			5688: out = -329;
			5689: out = -279;
			5690: out = -242;
			5691: out = -195;
			5692: out = -152;
			5693: out = -108;
			5694: out = -80;
			5695: out = -44;
			5696: out = 3;
			5697: out = 39;
			5698: out = 100;
			5699: out = 112;
			5700: out = 163;
			5701: out = 205;
			5702: out = 231;
			5703: out = 278;
			5704: out = 317;
			5705: out = 354;
			5706: out = 382;
			5707: out = 432;
			5708: out = 462;
			5709: out = 510;
			5710: out = 533;
			5711: out = 560;
			5712: out = 596;
			5713: out = 634;
			5714: out = 682;
			5715: out = 694;
			5716: out = 760;
			5717: out = 774;
			5718: out = 813;
			5719: out = 837;
			5720: out = 880;
			5721: out = 903;
			5722: out = 945;
			5723: out = 983;
			5724: out = 1006;
			5725: out = 1056;
			5726: out = 1090;
			5727: out = 1110;
			5728: out = 1143;
			5729: out = 1199;
			5730: out = 1216;
			5731: out = 1245;
			5732: out = 1299;
			5733: out = 1317;
			5734: out = 1358;
			5735: out = 1386;
			5736: out = 1427;
			5737: out = 1484;
			5738: out = 1513;
			5739: out = 1555;
			5740: out = 1590;
			5741: out = 1612;
			5742: out = 1662;
			5743: out = 1693;
			5744: out = 1723;
			5745: out = 1755;
			5746: out = 1811;
			5747: out = 1853;
			5748: out = 1885;
			5749: out = 1942;
			5750: out = 1981;
			5751: out = 2026;
			5752: out = 2068;
			5753: out = 2120;
			5754: out = 2152;
			5755: out = 2216;
			5756: out = 2266;
			5757: out = 2294;
			5758: out = 2356;
			5759: out = 2412;
			5760: out = 2467;
			5761: out = 2510;
			5762: out = 2561;
			5763: out = 2613;
			5764: out = 2665;
			5765: out = 2729;
			5766: out = 2782;
			5767: out = 2848;
			5768: out = 2903;
			5769: out = 2959;
			5770: out = 3028;
			5771: out = 3074;
			5772: out = 3139;
			5773: out = 3208;
			5774: out = 3260;
			5775: out = 3321;
			5776: out = 3390;
			5777: out = 3463;
			5778: out = 3528;
			5779: out = 3594;
			5780: out = 3651;
			5781: out = 3718;
			5782: out = 3785;
			5783: out = 3860;
			5784: out = 3909;
			5785: out = 3980;
			5786: out = 4040;
			5787: out = 4113;
			5788: out = 4186;
			5789: out = 4245;
			5790: out = 4323;
			5791: out = 4375;
			5792: out = 4441;
			5793: out = 4505;
			5794: out = 4570;
			5795: out = 4633;
			5796: out = 4693;
			5797: out = 4747;
			5798: out = 4809;
			5799: out = 4885;
			5800: out = 4944;
			5801: out = 4996;
			5802: out = 5067;
			5803: out = 5109;
			5804: out = 5173;
			5805: out = 5213;
			5806: out = 5291;
			5807: out = 5347;
			5808: out = 5397;
			5809: out = 5438;
			5810: out = 5520;
			5811: out = 5560;
			5812: out = 5617;
			5813: out = 5675;
			5814: out = 5728;
			5815: out = 5767;
			5816: out = 5828;
			5817: out = 5870;
			5818: out = 5943;
			5819: out = 5973;
			5820: out = 6017;
			5821: out = 6061;
			5822: out = 6136;
			5823: out = 6186;
			5824: out = 6218;
			5825: out = 6276;
			5826: out = 6315;
			5827: out = 6352;
			5828: out = 6406;
			5829: out = 6439;
			5830: out = 6483;
			5831: out = 6527;
			5832: out = 6571;
			5833: out = 6624;
			5834: out = 6652;
			5835: out = 6706;
			5836: out = 6746;
			5837: out = 6770;
			5838: out = 6826;
			5839: out = 6850;
			5840: out = 6891;
			5841: out = 6949;
			5842: out = 6950;
			5843: out = 7011;
			5844: out = 7048;
			5845: out = 7080;
			5846: out = 7117;
			5847: out = 7160;
			5848: out = 7195;
			5849: out = 7214;
			5850: out = 7259;
			5851: out = 7300;
			5852: out = 7339;
			5853: out = 7355;
			5854: out = 7402;
			5855: out = 7422;
			5856: out = 7468;
			5857: out = 7491;
			5858: out = 7522;
			5859: out = 7559;
			5860: out = 7575;
			5861: out = 7609;
			5862: out = 7648;
			5863: out = 7687;
			5864: out = 7706;
			5865: out = 7741;
			5866: out = 7766;
			5867: out = 7790;
			5868: out = 7823;
			5869: out = 7856;
			5870: out = 7879;
			5871: out = 7908;
			5872: out = 7934;
			5873: out = 7973;
			5874: out = 7978;
			5875: out = 8022;
			5876: out = 8062;
			5877: out = 8076;
			5878: out = 8095;
			5879: out = 8123;
			5880: out = 8149;
			5881: out = 8180;
			5882: out = 8195;
			5883: out = 8209;
			5884: out = 8246;
			5885: out = 8275;
			5886: out = 8304;
			5887: out = 8326;
			5888: out = 8346;
			5889: out = 8375;
			5890: out = 8382;
			5891: out = 8386;
			5892: out = 8427;
			5893: out = 8442;
			5894: out = 8428;
			5895: out = 8450;
			5896: out = 8467;
			5897: out = 8438;
			5898: out = 8427;
			5899: out = 8432;
			5900: out = 8405;
			5901: out = 8406;
			5902: out = 8427;
			5903: out = 8402;
			5904: out = 8444;
			5905: out = 8414;
			5906: out = 8417;
			5907: out = 8403;
			5908: out = 8368;
			5909: out = 8387;
			5910: out = 8398;
			5911: out = 8381;
			5912: out = 8372;
			5913: out = 8379;
			5914: out = 8360;
			5915: out = 8377;
			5916: out = 8304;
			5917: out = 8323;
			5918: out = 8349;
			5919: out = 8347;
			5920: out = 8332;
			5921: out = 8323;
			5922: out = 8331;
			5923: out = 8326;
			5924: out = 8292;
			5925: out = 8287;
			5926: out = 8275;
			5927: out = 8262;
			5928: out = 8269;
			5929: out = 8300;
			5930: out = 8272;
			5931: out = 8274;
			5932: out = 8281;
			5933: out = 8260;
			5934: out = 8266;
			5935: out = 8292;
			5936: out = 8218;
			5937: out = 8242;
			5938: out = 8198;
			5939: out = 8217;
			5940: out = 8238;
			5941: out = 8210;
			5942: out = 8226;
			5943: out = 8264;
			5944: out = 8248;
			5945: out = 8194;
			5946: out = 8185;
			5947: out = 8196;
			5948: out = 8159;
			5949: out = 8125;
			5950: out = 8147;
			5951: out = 8113;
			5952: out = 8102;
			5953: out = 8114;
			5954: out = 8106;
			5955: out = 8113;
			5956: out = 8113;
			5957: out = 8098;
			5958: out = 8076;
			5959: out = 8074;
			5960: out = 8080;
			5961: out = 8075;
			5962: out = 8010;
			5963: out = 8022;
			5964: out = 7998;
			5965: out = 8001;
			5966: out = 7977;
			5967: out = 7951;
			5968: out = 7914;
			5969: out = 7894;
			5970: out = 7894;
			5971: out = 7863;
			5972: out = 7849;
			5973: out = 7834;
			5974: out = 7843;
			5975: out = 7771;
			5976: out = 7737;
			5977: out = 7713;
			5978: out = 7681;
			5979: out = 7671;
			5980: out = 7637;
			5981: out = 7609;
			5982: out = 7580;
			5983: out = 7512;
			5984: out = 7504;
			5985: out = 7463;
			5986: out = 7396;
			5987: out = 7374;
			5988: out = 7332;
			5989: out = 7278;
			5990: out = 7251;
			5991: out = 7201;
			5992: out = 7146;
			5993: out = 7116;
			5994: out = 7069;
			5995: out = 7066;
			5996: out = 6960;
			5997: out = 6928;
			5998: out = 6870;
			5999: out = 6833;
			6000: out = 6826;
			6001: out = 6761;
			6002: out = 6702;
			6003: out = 6646;
			6004: out = 6602;
			6005: out = 6530;
			6006: out = 6470;
			6007: out = 6450;
			6008: out = 6376;
			6009: out = 6344;
			6010: out = 6284;
			6011: out = 6235;
			6012: out = 6182;
			6013: out = 6125;
			6014: out = 6074;
			6015: out = 5997;
			6016: out = 5954;
			6017: out = 5895;
			6018: out = 5840;
			6019: out = 5785;
			6020: out = 5748;
			6021: out = 5673;
			6022: out = 5616;
			6023: out = 5569;
			6024: out = 5520;
			6025: out = 5465;
			6026: out = 5391;
			6027: out = 5361;
			6028: out = 5287;
			6029: out = 5239;
			6030: out = 5196;
			6031: out = 5132;
			6032: out = 5072;
			6033: out = 5047;
			6034: out = 4967;
			6035: out = 4927;
			6036: out = 4867;
			6037: out = 4820;
			6038: out = 4761;
			6039: out = 4704;
			6040: out = 4656;
			6041: out = 4605;
			6042: out = 4546;
			6043: out = 4523;
			6044: out = 4442;
			6045: out = 4400;
			6046: out = 4351;
			6047: out = 4305;
			6048: out = 4264;
			6049: out = 4206;
			6050: out = 4150;
			6051: out = 4119;
			6052: out = 4071;
			6053: out = 4029;
			6054: out = 3977;
			6055: out = 3918;
			6056: out = 3896;
			6057: out = 3819;
			6058: out = 3788;
			6059: out = 3742;
			6060: out = 3713;
			6061: out = 3633;
			6062: out = 3601;
			6063: out = 3575;
			6064: out = 3532;
			6065: out = 3473;
			6066: out = 3442;
			6067: out = 3404;
			6068: out = 3329;
			6069: out = 3305;
			6070: out = 3285;
			6071: out = 3228;
			6072: out = 3182;
			6073: out = 3142;
			6074: out = 3098;
			6075: out = 3078;
			6076: out = 3034;
			6077: out = 2992;
			6078: out = 2952;
			6079: out = 2928;
			6080: out = 2889;
			6081: out = 2864;
			6082: out = 2827;
			6083: out = 2764;
			6084: out = 2741;
			6085: out = 2681;
			6086: out = 2667;
			6087: out = 2630;
			6088: out = 2601;
			6089: out = 2563;
			6090: out = 2533;
			6091: out = 2486;
			6092: out = 2453;
			6093: out = 2421;
			6094: out = 2374;
			6095: out = 2346;
			6096: out = 2330;
			6097: out = 2289;
			6098: out = 2261;
			6099: out = 2243;
			6100: out = 2192;
			6101: out = 2155;
			6102: out = 2110;
			6103: out = 2087;
			6104: out = 2077;
			6105: out = 2044;
			6106: out = 2018;
			6107: out = 2010;
			6108: out = 1963;
			6109: out = 1948;
			6110: out = 1913;
			6111: out = 1904;
			6112: out = 1868;
			6113: out = 1817;
			6114: out = 1801;
			6115: out = 1773;
			6116: out = 1761;
			6117: out = 1746;
			6118: out = 1702;
			6119: out = 1701;
			6120: out = 1660;
			6121: out = 1634;
			6122: out = 1612;
			6123: out = 1595;
			6124: out = 1551;
			6125: out = 1533;
			6126: out = 1497;
			6127: out = 1437;
			6128: out = 1376;
			6129: out = 1300;
			6130: out = 1238;
			6131: out = 1179;
			6132: out = 1108;
			6133: out = 1054;
			6134: out = 1007;
			6135: out = 938;
			6136: out = 872;
			6137: out = 813;
			6138: out = 768;
			6139: out = 713;
			6140: out = 670;
			6141: out = 626;
			6142: out = 569;
			6143: out = 503;
			6144: out = 469;
			6145: out = 404;
			6146: out = 345;
			6147: out = 315;
			6148: out = 243;
			6149: out = 207;
			6150: out = 144;
			6151: out = 101;
			6152: out = 51;
			6153: out = 27;
			6154: out = -41;
			6155: out = -75;
			6156: out = -123;
			6157: out = -179;
			6158: out = -218;
			6159: out = -287;
			6160: out = -326;
			6161: out = -358;
			6162: out = -401;
			6163: out = -446;
			6164: out = -478;
			6165: out = -538;
			6166: out = -573;
			6167: out = -629;
			6168: out = -647;
			6169: out = -700;
			6170: out = -737;
			6171: out = -788;
			6172: out = -817;
			6173: out = -854;
			6174: out = -898;
			6175: out = -917;
			6176: out = -989;
			6177: out = -1003;
			6178: out = -1036;
			6179: out = -1108;
			6180: out = -1107;
			6181: out = -1163;
			6182: out = -1197;
			6183: out = -1243;
			6184: out = -1286;
			6185: out = -1303;
			6186: out = -1335;
			6187: out = -1368;
			6188: out = -1404;
			6189: out = -1444;
			6190: out = -1497;
			6191: out = -1511;
			6192: out = -1566;
			6193: out = -1616;
			6194: out = -1634;
			6195: out = -1676;
			6196: out = -1713;
			6197: out = -1736;
			6198: out = -1769;
			6199: out = -1824;
			6200: out = -1844;
			6201: out = -1890;
			6202: out = -1936;
			6203: out = -1967;
			6204: out = -1992;
			6205: out = -2050;
			6206: out = -2078;
			6207: out = -2125;
			6208: out = -2171;
			6209: out = -2199;
			6210: out = -2257;
			6211: out = -2289;
			6212: out = -2332;
			6213: out = -2377;
			6214: out = -2412;
			6215: out = -2462;
			6216: out = -2501;
			6217: out = -2554;
			6218: out = -2587;
			6219: out = -2646;
			6220: out = -2678;
			6221: out = -2724;
			6222: out = -2788;
			6223: out = -2841;
			6224: out = -2877;
			6225: out = -2921;
			6226: out = -2969;
			6227: out = -3015;
			6228: out = -3086;
			6229: out = -3126;
			6230: out = -3181;
			6231: out = -3238;
			6232: out = -3286;
			6233: out = -3336;
			6234: out = -3420;
			6235: out = -3466;
			6236: out = -3515;
			6237: out = -3596;
			6238: out = -3651;
			6239: out = -3698;
			6240: out = -3772;
			6241: out = -3837;
			6242: out = -3899;
			6243: out = -3960;
			6244: out = -4046;
			6245: out = -4108;
			6246: out = -4187;
			6247: out = -4247;
			6248: out = -4314;
			6249: out = -4379;
			6250: out = -4457;
			6251: out = -4521;
			6252: out = -4602;
			6253: out = -4680;
			6254: out = -4751;
			6255: out = -4813;
			6256: out = -4896;
			6257: out = -4969;
			6258: out = -5039;
			6259: out = -5118;
			6260: out = -5187;
			6261: out = -5261;
			6262: out = -5347;
			6263: out = -5410;
			6264: out = -5473;
			6265: out = -5559;
			6266: out = -5623;
			6267: out = -5689;
			6268: out = -5777;
			6269: out = -5842;
			6270: out = -5910;
			6271: out = -5966;
			6272: out = -6044;
			6273: out = -6105;
			6274: out = -6173;
			6275: out = -6239;
			6276: out = -6312;
			6277: out = -6363;
			6278: out = -6443;
			6279: out = -6502;
			6280: out = -6554;
			6281: out = -6623;
			6282: out = -6668;
			6283: out = -6736;
			6284: out = -6777;
			6285: out = -6829;
			6286: out = -6881;
			6287: out = -6941;
			6288: out = -6985;
			6289: out = -7032;
			6290: out = -7078;
			6291: out = -7128;
			6292: out = -7160;
			6293: out = -7216;
			6294: out = -7267;
			6295: out = -7282;
			6296: out = -7339;
			6297: out = -7383;
			6298: out = -7411;
			6299: out = -7463;
			6300: out = -7486;
			6301: out = -7531;
			6302: out = -7558;
			6303: out = -7601;
			6304: out = -7630;
			6305: out = -7659;
			6306: out = -7689;
			6307: out = -7728;
			6308: out = -7745;
			6309: out = -7778;
			6310: out = -7823;
			6311: out = -7838;
			6312: out = -7864;
			6313: out = -7874;
			6314: out = -7898;
			6315: out = -7926;
			6316: out = -7943;
			6317: out = -7971;
			6318: out = -7992;
			6319: out = -8001;
			6320: out = -8027;
			6321: out = -8042;
			6322: out = -8063;
			6323: out = -8076;
			6324: out = -8091;
			6325: out = -8092;
			6326: out = -8119;
			6327: out = -8128;
			6328: out = -8140;
			6329: out = -8151;
			6330: out = -8150;
			6331: out = -8178;
			6332: out = -8178;
			6333: out = -8186;
			6334: out = -8186;
			6335: out = -8206;
			6336: out = -8199;
			6337: out = -8209;
			6338: out = -8206;
			6339: out = -8226;
			6340: out = -8220;
			6341: out = -8225;
			6342: out = -8239;
			6343: out = -8241;
			6344: out = -8227;
			6345: out = -8244;
			6346: out = -8227;
			6347: out = -8242;
			6348: out = -8223;
			6349: out = -8253;
			6350: out = -8231;
			6351: out = -8225;
			6352: out = -8226;
			6353: out = -8228;
			6354: out = -8223;
			6355: out = -8233;
			6356: out = -8206;
			6357: out = -8211;
			6358: out = -8214;
			6359: out = -8198;
			6360: out = -8207;
			6361: out = -8189;
			6362: out = -8183;
			6363: out = -8180;
			6364: out = -8184;
			6365: out = -8183;
			6366: out = -8168;
			6367: out = -8149;
			6368: out = -8133;
			6369: out = -8137;
			6370: out = -8101;
			6371: out = -8103;
			6372: out = -8096;
			6373: out = -8074;
			6374: out = -8064;
			6375: out = -8066;
			6376: out = -8049;
			6377: out = -8038;
			6378: out = -8027;
			6379: out = -8009;
			6380: out = -8005;
			6381: out = -7970;
			6382: out = -7981;
			6383: out = -7969;
			6384: out = -7947;
			6385: out = -7943;
			6386: out = -7922;
			6387: out = -7907;
			6388: out = -7887;
			6389: out = -7885;
			6390: out = -7867;
			6391: out = -7855;
			6392: out = -7823;
			6393: out = -7822;
			6394: out = -7811;
			6395: out = -7795;
			6396: out = -7758;
			6397: out = -7753;
			6398: out = -7741;
			6399: out = -7704;
			6400: out = -7702;
			6401: out = -7683;
			6402: out = -7662;
			6403: out = -7646;
			6404: out = -7624;
			6405: out = -7593;
			6406: out = -7590;
			6407: out = -7568;
			6408: out = -7548;
			6409: out = -7523;
			6410: out = -7499;
			6411: out = -7471;
			6412: out = -7457;
			6413: out = -7433;
			6414: out = -7421;
			6415: out = -7388;
			6416: out = -7351;
			6417: out = -7342;
			6418: out = -7318;
			6419: out = -7290;
			6420: out = -7256;
			6421: out = -7237;
			6422: out = -7213;
			6423: out = -7186;
			6424: out = -7150;
			6425: out = -7127;
			6426: out = -7091;
			6427: out = -7056;
			6428: out = -7039;
			6429: out = -7000;
			6430: out = -6967;
			6431: out = -6947;
			6432: out = -6895;
			6433: out = -6869;
			6434: out = -6831;
			6435: out = -6791;
			6436: out = -6760;
			6437: out = -6717;
			6438: out = -6675;
			6439: out = -6644;
			6440: out = -6578;
			6441: out = -6558;
			6442: out = -6512;
			6443: out = -6452;
			6444: out = -6416;
			6445: out = -6369;
			6446: out = -6310;
			6447: out = -6276;
			6448: out = -6204;
			6449: out = -6154;
			6450: out = -6098;
			6451: out = -6061;
			6452: out = -6012;
			6453: out = -5950;
			6454: out = -5899;
			6455: out = -5849;
			6456: out = -5802;
			6457: out = -5736;
			6458: out = -5683;
			6459: out = -5619;
			6460: out = -5578;
			6461: out = -5508;
			6462: out = -5450;
			6463: out = -5392;
			6464: out = -5342;
			6465: out = -5285;
			6466: out = -5236;
			6467: out = -5164;
			6468: out = -5099;
			6469: out = -5051;
			6470: out = -5000;
			6471: out = -4940;
			6472: out = -4868;
			6473: out = -4822;
			6474: out = -4755;
			6475: out = -4707;
			6476: out = -4640;
			6477: out = -4588;
			6478: out = -4529;
			6479: out = -4479;
			6480: out = -4416;
			6481: out = -4363;
			6482: out = -4313;
			6483: out = -4252;
			6484: out = -4194;
			6485: out = -4132;
			6486: out = -4081;
			6487: out = -4015;
			6488: out = -3983;
			6489: out = -3912;
			6490: out = -3871;
			6491: out = -3800;
			6492: out = -3756;
			6493: out = -3702;
			6494: out = -3654;
			6495: out = -3604;
			6496: out = -3546;
			6497: out = -3496;
			6498: out = -3456;
			6499: out = -3404;
			6500: out = -3345;
			6501: out = -3305;
			6502: out = -3250;
			6503: out = -3213;
			6504: out = -3169;
			6505: out = -3116;
			6506: out = -3079;
			6507: out = -3028;
			6508: out = -2986;
			6509: out = -2937;
			6510: out = -2888;
			6511: out = -2856;
			6512: out = -2805;
			6513: out = -2764;
			6514: out = -2720;
			6515: out = -2683;
			6516: out = -2635;
			6517: out = -2599;
			6518: out = -2550;
			6519: out = -2522;
			6520: out = -2459;
			6521: out = -2438;
			6522: out = -2393;
			6523: out = -2353;
			6524: out = -2317;
			6525: out = -2270;
			6526: out = -2235;
			6527: out = -2205;
			6528: out = -2175;
			6529: out = -2133;
			6530: out = -2108;
			6531: out = -2065;
			6532: out = -2016;
			6533: out = -1993;
			6534: out = -1949;
			6535: out = -1931;
			6536: out = -1891;
			6537: out = -1861;
			6538: out = -1828;
			6539: out = -1811;
			6540: out = -1778;
			6541: out = -1737;
			6542: out = -1711;
			6543: out = -1673;
			6544: out = -1652;
			6545: out = -1624;
			6546: out = -1600;
			6547: out = -1554;
			6548: out = -1535;
			6549: out = -1523;
			6550: out = -1473;
			6551: out = -1421;
			6552: out = -1375;
			6553: out = -1312;
			6554: out = -1264;
			6555: out = -1206;
			6556: out = -1166;
			6557: out = -1104;
			6558: out = -1071;
			6559: out = -1023;
			6560: out = -978;
			6561: out = -928;
			6562: out = -884;
			6563: out = -857;
			6564: out = -795;
			6565: out = -767;
			6566: out = -711;
			6567: out = -676;
			6568: out = -636;
			6569: out = -605;
			6570: out = -562;
			6571: out = -528;
			6572: out = -483;
			6573: out = -446;
			6574: out = -406;
			6575: out = -382;
			6576: out = -346;
			6577: out = -303;
			6578: out = -271;
			6579: out = -240;
			6580: out = -203;
			6581: out = -174;
			6582: out = -126;
			6583: out = -107;
			6584: out = -56;
			6585: out = -43;
			6586: out = -1;
			6587: out = 19;
			6588: out = 60;
			6589: out = 96;
			6590: out = 126;
			6591: out = 147;
			6592: out = 183;
			6593: out = 218;
			6594: out = 246;
			6595: out = 277;
			6596: out = 312;
			6597: out = 342;
			6598: out = 364;
			6599: out = 395;
			6600: out = 423;
			6601: out = 456;
			6602: out = 489;
			6603: out = 501;
			6604: out = 545;
			6605: out = 562;
			6606: out = 594;
			6607: out = 635;
			6608: out = 647;
			6609: out = 672;
			6610: out = 709;
			6611: out = 736;
			6612: out = 759;
			6613: out = 789;
			6614: out = 809;
			6615: out = 841;
			6616: out = 856;
			6617: out = 895;
			6618: out = 922;
			6619: out = 957;
			6620: out = 975;
			6621: out = 1016;
			6622: out = 1037;
			6623: out = 1067;
			6624: out = 1098;
			6625: out = 1129;
			6626: out = 1143;
			6627: out = 1179;
			6628: out = 1219;
			6629: out = 1241;
			6630: out = 1290;
			6631: out = 1308;
			6632: out = 1344;
			6633: out = 1365;
			6634: out = 1417;
			6635: out = 1444;
			6636: out = 1480;
			6637: out = 1515;
			6638: out = 1539;
			6639: out = 1577;
			6640: out = 1608;
			6641: out = 1640;
			6642: out = 1664;
			6643: out = 1709;
			6644: out = 1753;
			6645: out = 1781;
			6646: out = 1824;
			6647: out = 1872;
			6648: out = 1908;
			6649: out = 1945;
			6650: out = 1992;
			6651: out = 2030;
			6652: out = 2063;
			6653: out = 2129;
			6654: out = 2163;
			6655: out = 2204;
			6656: out = 2253;
			6657: out = 2304;
			6658: out = 2361;
			6659: out = 2398;
			6660: out = 2440;
			6661: out = 2503;
			6662: out = 2547;
			6663: out = 2597;
			6664: out = 2658;
			6665: out = 2696;
			6666: out = 2760;
			6667: out = 2798;
			6668: out = 2855;
			6669: out = 2908;
			6670: out = 2960;
			6671: out = 3018;
			6672: out = 3075;
			6673: out = 3119;
			6674: out = 3180;
			6675: out = 3226;
			6676: out = 3296;
			6677: out = 3326;
			6678: out = 3392;
			6679: out = 3445;
			6680: out = 3499;
			6681: out = 3551;
			6682: out = 3602;
			6683: out = 3663;
			6684: out = 3701;
			6685: out = 3753;
			6686: out = 3811;
			6687: out = 3867;
			6688: out = 3914;
			6689: out = 3960;
			6690: out = 4010;
			6691: out = 4056;
			6692: out = 4127;
			6693: out = 4152;
			6694: out = 4203;
			6695: out = 4269;
			6696: out = 4292;
			6697: out = 4347;
			6698: out = 4400;
			6699: out = 4441;
			6700: out = 4489;
			6701: out = 4524;
			6702: out = 4574;
			6703: out = 4616;
			6704: out = 4669;
			6705: out = 4708;
			6706: out = 4760;
			6707: out = 4801;
			6708: out = 4845;
			6709: out = 4884;
			6710: out = 4925;
			6711: out = 4979;
			6712: out = 5000;
			6713: out = 5046;
			6714: out = 5082;
			6715: out = 5126;
			6716: out = 5174;
			6717: out = 5188;
			6718: out = 5249;
			6719: out = 5268;
			6720: out = 5312;
			6721: out = 5352;
			6722: out = 5370;
			6723: out = 5417;
			6724: out = 5442;
			6725: out = 5474;
			6726: out = 5516;
			6727: out = 5551;
			6728: out = 5565;
			6729: out = 5614;
			6730: out = 5633;
			6731: out = 5663;
			6732: out = 5714;
			6733: out = 5729;
			6734: out = 5761;
			6735: out = 5803;
			6736: out = 5841;
			6737: out = 5855;
			6738: out = 5890;
			6739: out = 5925;
			6740: out = 5942;
			6741: out = 5992;
			6742: out = 6002;
			6743: out = 6026;
			6744: out = 6067;
			6745: out = 6073;
			6746: out = 6118;
			6747: out = 6138;
			6748: out = 6169;
			6749: out = 6197;
			6750: out = 6216;
			6751: out = 6245;
			6752: out = 6270;
			6753: out = 6305;
			6754: out = 6318;
			6755: out = 6332;
			6756: out = 6379;
			6757: out = 6385;
			6758: out = 6420;
			6759: out = 6443;
			6760: out = 6468;
			6761: out = 6485;
			6762: out = 6509;
			6763: out = 6535;
			6764: out = 6557;
			6765: out = 6586;
			6766: out = 6590;
			6767: out = 6613;
			6768: out = 6657;
			6769: out = 6657;
			6770: out = 6690;
			6771: out = 6712;
			6772: out = 6739;
			6773: out = 6750;
			6774: out = 6773;
			6775: out = 6801;
			6776: out = 6810;
			6777: out = 6859;
			6778: out = 6835;
			6779: out = 6878;
			6780: out = 6896;
			6781: out = 6897;
			6782: out = 6926;
			6783: out = 6944;
			6784: out = 6959;
			6785: out = 6959;
			6786: out = 6957;
			6787: out = 6960;
			6788: out = 6970;
			6789: out = 6982;
			6790: out = 6954;
			6791: out = 6953;
			6792: out = 6940;
			6793: out = 6932;
			6794: out = 6925;
			6795: out = 6925;
			6796: out = 6929;
			6797: out = 6908;
			6798: out = 6917;
			6799: out = 6885;
			6800: out = 6889;
			6801: out = 6878;
			6802: out = 6844;
			6803: out = 6871;
			6804: out = 6861;
			6805: out = 6860;
			6806: out = 6873;
			6807: out = 6884;
			6808: out = 6881;
			6809: out = 6899;
			6810: out = 6874;
			6811: out = 6891;
			6812: out = 6870;
			6813: out = 6882;
			6814: out = 6873;
			6815: out = 6841;
			6816: out = 6836;
			6817: out = 6857;
			6818: out = 6813;
			6819: out = 6815;
			6820: out = 6833;
			6821: out = 6825;
			6822: out = 6795;
			6823: out = 6797;
			6824: out = 6783;
			6825: out = 6774;
			6826: out = 6769;
			6827: out = 6807;
			6828: out = 6794;
			6829: out = 6802;
			6830: out = 6759;
			6831: out = 6778;
			6832: out = 6783;
			6833: out = 6772;
			6834: out = 6779;
			6835: out = 6795;
			6836: out = 6781;
			6837: out = 6762;
			6838: out = 6749;
			6839: out = 6708;
			6840: out = 6741;
			6841: out = 6713;
			6842: out = 6722;
			6843: out = 6713;
			6844: out = 6705;
			6845: out = 6706;
			6846: out = 6693;
			6847: out = 6701;
			6848: out = 6687;
			6849: out = 6701;
			6850: out = 6693;
			6851: out = 6671;
			6852: out = 6616;
			6853: out = 6594;
			6854: out = 6595;
			6855: out = 6584;
			6856: out = 6557;
			6857: out = 6574;
			6858: out = 6556;
			6859: out = 6536;
			6860: out = 6505;
			6861: out = 6511;
			6862: out = 6507;
			6863: out = 6445;
			6864: out = 6445;
			6865: out = 6440;
			6866: out = 6410;
			6867: out = 6389;
			6868: out = 6344;
			6869: out = 6324;
			6870: out = 6323;
			6871: out = 6268;
			6872: out = 6254;
			6873: out = 6221;
			6874: out = 6187;
			6875: out = 6173;
			6876: out = 6166;
			6877: out = 6089;
			6878: out = 6074;
			6879: out = 6052;
			6880: out = 6012;
			6881: out = 5981;
			6882: out = 5942;
			6883: out = 5902;
			6884: out = 5861;
			6885: out = 5848;
			6886: out = 5806;
			6887: out = 5749;
			6888: out = 5710;
			6889: out = 5651;
			6890: out = 5616;
			6891: out = 5602;
			6892: out = 5548;
			6893: out = 5527;
			6894: out = 5472;
			6895: out = 5425;
			6896: out = 5389;
			6897: out = 5326;
			6898: out = 5309;
			6899: out = 5253;
			6900: out = 5214;
			6901: out = 5162;
			6902: out = 5111;
			6903: out = 5089;
			6904: out = 5025;
			6905: out = 5010;
			6906: out = 4952;
			6907: out = 4905;
			6908: out = 4858;
			6909: out = 4806;
			6910: out = 4765;
			6911: out = 4734;
			6912: out = 4683;
			6913: out = 4613;
			6914: out = 4592;
			6915: out = 4523;
			6916: out = 4491;
			6917: out = 4447;
			6918: out = 4399;
			6919: out = 4361;
			6920: out = 4332;
			6921: out = 4264;
			6922: out = 4225;
			6923: out = 4183;
			6924: out = 4159;
			6925: out = 4088;
			6926: out = 4052;
			6927: out = 4010;
			6928: out = 3958;
			6929: out = 3929;
			6930: out = 3865;
			6931: out = 3848;
			6932: out = 3795;
			6933: out = 3764;
			6934: out = 3716;
			6935: out = 3665;
			6936: out = 3633;
			6937: out = 3583;
			6938: out = 3529;
			6939: out = 3520;
			6940: out = 3466;
			6941: out = 3410;
			6942: out = 3377;
			6943: out = 3362;
			6944: out = 3310;
			6945: out = 3287;
			6946: out = 3236;
			6947: out = 3182;
			6948: out = 3160;
			6949: out = 3111;
			6950: out = 3101;
			6951: out = 3055;
			6952: out = 3020;
			6953: out = 2978;
			6954: out = 2951;
			6955: out = 2903;
			6956: out = 2881;
			6957: out = 2827;
			6958: out = 2803;
			6959: out = 2774;
			6960: out = 2737;
			6961: out = 2703;
			6962: out = 2682;
			6963: out = 2626;
			6964: out = 2607;
			6965: out = 2568;
			6966: out = 2528;
			6967: out = 2512;
			6968: out = 2491;
			6969: out = 2459;
			6970: out = 2409;
			6971: out = 2387;
			6972: out = 2361;
			6973: out = 2315;
			6974: out = 2290;
			6975: out = 2275;
			6976: out = 2238;
			6977: out = 2214;
			6978: out = 2183;
			6979: out = 2146;
			6980: out = 2123;
			6981: out = 2097;
			6982: out = 2073;
			6983: out = 2033;
			6984: out = 2020;
			6985: out = 1985;
			6986: out = 1959;
			6987: out = 1929;
			6988: out = 1890;
			6989: out = 1876;
			6990: out = 1859;
			6991: out = 1817;
			6992: out = 1808;
			6993: out = 1773;
			6994: out = 1758;
			6995: out = 1713;
			6996: out = 1700;
			6997: out = 1691;
			6998: out = 1657;
			6999: out = 1619;
			7000: out = 1607;
			7001: out = 1582;
			7002: out = 1569;
			7003: out = 1534;
			7004: out = 1510;
			7005: out = 1506;
			7006: out = 1459;
			7007: out = 1434;
			7008: out = 1425;
			7009: out = 1399;
			7010: out = 1388;
			7011: out = 1370;
			7012: out = 1359;
			7013: out = 1338;
			7014: out = 1319;
			7015: out = 1282;
			7016: out = 1258;
			7017: out = 1237;
			7018: out = 1176;
			7019: out = 1128;
			7020: out = 1087;
			7021: out = 1031;
			7022: out = 966;
			7023: out = 924;
			7024: out = 867;
			7025: out = 813;
			7026: out = 782;
			7027: out = 716;
			7028: out = 666;
			7029: out = 619;
			7030: out = 573;
			7031: out = 537;
			7032: out = 486;
			7033: out = 442;
			7034: out = 394;
			7035: out = 367;
			7036: out = 310;
			7037: out = 270;
			7038: out = 241;
			7039: out = 174;
			7040: out = 135;
			7041: out = 107;
			7042: out = 53;
			7043: out = 26;
			7044: out = -10;
			7045: out = -54;
			7046: out = -92;
			7047: out = -140;
			7048: out = -173;
			7049: out = -202;
			7050: out = -242;
			7051: out = -280;
			7052: out = -325;
			7053: out = -350;
			7054: out = -389;
			7055: out = -410;
			7056: out = -460;
			7057: out = -471;
			7058: out = -538;
			7059: out = -541;
			7060: out = -576;
			7061: out = -625;
			7062: out = -660;
			7063: out = -703;
			7064: out = -725;
			7065: out = -766;
			7066: out = -789;
			7067: out = -829;
			7068: out = -849;
			7069: out = -886;
			7070: out = -918;
			7071: out = -945;
			7072: out = -967;
			7073: out = -1007;
			7074: out = -1050;
			7075: out = -1080;
			7076: out = -1101;
			7077: out = -1142;
			7078: out = -1158;
			7079: out = -1184;
			7080: out = -1222;
			7081: out = -1257;
			7082: out = -1276;
			7083: out = -1317;
			7084: out = -1341;
			7085: out = -1373;
			7086: out = -1416;
			7087: out = -1433;
			7088: out = -1469;
			7089: out = -1498;
			7090: out = -1521;
			7091: out = -1555;
			7092: out = -1566;
			7093: out = -1604;
			7094: out = -1648;
			7095: out = -1673;
			7096: out = -1716;
			7097: out = -1750;
			7098: out = -1790;
			7099: out = -1825;
			7100: out = -1860;
			7101: out = -1888;
			7102: out = -1918;
			7103: out = -1960;
			7104: out = -1990;
			7105: out = -2017;
			7106: out = -2064;
			7107: out = -2090;
			7108: out = -2133;
			7109: out = -2159;
			7110: out = -2216;
			7111: out = -2249;
			7112: out = -2282;
			7113: out = -2322;
			7114: out = -2375;
			7115: out = -2397;
			7116: out = -2444;
			7117: out = -2478;
			7118: out = -2521;
			7119: out = -2572;
			7120: out = -2614;
			7121: out = -2649;
			7122: out = -2696;
			7123: out = -2747;
			7124: out = -2783;
			7125: out = -2827;
			7126: out = -2889;
			7127: out = -2923;
			7128: out = -2987;
			7129: out = -3010;
			7130: out = -3087;
			7131: out = -3121;
			7132: out = -3180;
			7133: out = -3247;
			7134: out = -3288;
			7135: out = -3357;
			7136: out = -3415;
			7137: out = -3465;
			7138: out = -3519;
			7139: out = -3589;
			7140: out = -3640;
			7141: out = -3707;
			7142: out = -3769;
			7143: out = -3815;
			7144: out = -3880;
			7145: out = -3932;
			7146: out = -4016;
			7147: out = -4069;
			7148: out = -4142;
			7149: out = -4186;
			7150: out = -4247;
			7151: out = -4313;
			7152: out = -4374;
			7153: out = -4435;
			7154: out = -4482;
			7155: out = -4565;
			7156: out = -4604;
			7157: out = -4670;
			7158: out = -4725;
			7159: out = -4791;
			7160: out = -4836;
			7161: out = -4882;
			7162: out = -4956;
			7163: out = -5003;
			7164: out = -5055;
			7165: out = -5107;
			7166: out = -5169;
			7167: out = -5216;
			7168: out = -5261;
			7169: out = -5315;
			7170: out = -5377;
			7171: out = -5411;
			7172: out = -5458;
			7173: out = -5515;
			7174: out = -5544;
			7175: out = -5617;
			7176: out = -5639;
			7177: out = -5681;
			7178: out = -5741;
			7179: out = -5750;
			7180: out = -5814;
			7181: out = -5852;
			7182: out = -5894;
			7183: out = -5920;
			7184: out = -5974;
			7185: out = -5995;
			7186: out = -6044;
			7187: out = -6078;
			7188: out = -6101;
			7189: out = -6150;
			7190: out = -6171;
			7191: out = -6184;
			7192: out = -6230;
			7193: out = -6253;
			7194: out = -6287;
			7195: out = -6306;
			7196: out = -6331;
			7197: out = -6360;
			7198: out = -6380;
			7199: out = -6416;
			7200: out = -6427;
			7201: out = -6445;
			7202: out = -6470;
			7203: out = -6471;
			7204: out = -6513;
			7205: out = -6517;
			7206: out = -6538;
			7207: out = -6552;
			7208: out = -6569;
			7209: out = -6584;
			7210: out = -6598;
			7211: out = -6629;
			7212: out = -6627;
			7213: out = -6637;
			7214: out = -6653;
			7215: out = -6665;
			7216: out = -6666;
			7217: out = -6689;
			7218: out = -6682;
			7219: out = -6713;
			7220: out = -6705;
			7221: out = -6720;
			7222: out = -6738;
			7223: out = -6735;
			7224: out = -6748;
			7225: out = -6749;
			7226: out = -6748;
			7227: out = -6764;
			7228: out = -6759;
			7229: out = -6767;
			7230: out = -6781;
			7231: out = -6771;
			7232: out = -6775;
			7233: out = -6784;
			7234: out = -6787;
			7235: out = -6782;
			7236: out = -6785;
			7237: out = -6782;
			7238: out = -6778;
			7239: out = -6771;
			7240: out = -6782;
			7241: out = -6775;
			7242: out = -6762;
			7243: out = -6767;
			7244: out = -6772;
			7245: out = -6761;
			7246: out = -6761;
			7247: out = -6769;
			7248: out = -6744;
			7249: out = -6740;
			7250: out = -6746;
			7251: out = -6730;
			7252: out = -6729;
			7253: out = -6715;
			7254: out = -6724;
			7255: out = -6710;
			7256: out = -6700;
			7257: out = -6714;
			7258: out = -6694;
			7259: out = -6681;
			7260: out = -6681;
			7261: out = -6666;
			7262: out = -6663;
			7263: out = -6647;
			7264: out = -6639;
			7265: out = -6643;
			7266: out = -6628;
			7267: out = -6611;
			7268: out = -6606;
			7269: out = -6604;
			7270: out = -6598;
			7271: out = -6589;
			7272: out = -6572;
			7273: out = -6561;
			7274: out = -6546;
			7275: out = -6546;
			7276: out = -6513;
			7277: out = -6512;
			7278: out = -6500;
			7279: out = -6488;
			7280: out = -6474;
			7281: out = -6455;
			7282: out = -6454;
			7283: out = -6431;
			7284: out = -6415;
			7285: out = -6409;
			7286: out = -6402;
			7287: out = -6375;
			7288: out = -6374;
			7289: out = -6340;
			7290: out = -6332;
			7291: out = -6311;
			7292: out = -6296;
			7293: out = -6276;
			7294: out = -6279;
			7295: out = -6245;
			7296: out = -6234;
			7297: out = -6226;
			7298: out = -6208;
			7299: out = -6184;
			7300: out = -6176;
			7301: out = -6157;
			7302: out = -6125;
			7303: out = -6118;
			7304: out = -6096;
			7305: out = -6083;
			7306: out = -6061;
			7307: out = -6045;
			7308: out = -6024;
			7309: out = -6007;
			7310: out = -5992;
			7311: out = -5966;
			7312: out = -5941;
			7313: out = -5923;
			7314: out = -5894;
			7315: out = -5870;
			7316: out = -5856;
			7317: out = -5824;
			7318: out = -5800;
			7319: out = -5771;
			7320: out = -5745;
			7321: out = -5722;
			7322: out = -5696;
			7323: out = -5658;
			7324: out = -5629;
			7325: out = -5610;
			7326: out = -5563;
			7327: out = -5535;
			7328: out = -5511;
			7329: out = -5465;
			7330: out = -5442;
			7331: out = -5401;
			7332: out = -5363;
			7333: out = -5338;
			7334: out = -5295;
			7335: out = -5261;
			7336: out = -5212;
			7337: out = -5176;
			7338: out = -5136;
			7339: out = -5095;
			7340: out = -5046;
			7341: out = -5014;
			7342: out = -4962;
			7343: out = -4916;
			7344: out = -4889;
			7345: out = -4834;
			7346: out = -4788;
			7347: out = -4749;
			7348: out = -4694;
			7349: out = -4654;
			7350: out = -4606;
			7351: out = -4554;
			7352: out = -4512;
			7353: out = -4458;
			7354: out = -4406;
			7355: out = -4357;
			7356: out = -4312;
			7357: out = -4263;
			7358: out = -4225;
			7359: out = -4174;
			7360: out = -4131;
			7361: out = -4079;
			7362: out = -4043;
			7363: out = -3984;
			7364: out = -3934;
			7365: out = -3898;
			7366: out = -3841;
			7367: out = -3795;
			7368: out = -3754;
			7369: out = -3693;
			7370: out = -3653;
			7371: out = -3614;
			7372: out = -3549;
			7373: out = -3530;
			7374: out = -3487;
			7375: out = -3432;
			7376: out = -3388;
			7377: out = -3328;
			7378: out = -3295;
			7379: out = -3249;
			7380: out = -3197;
			7381: out = -3158;
			7382: out = -3118;
			7383: out = -3070;
			7384: out = -3035;
			7385: out = -2998;
			7386: out = -2947;
			7387: out = -2893;
			7388: out = -2872;
			7389: out = -2813;
			7390: out = -2779;
			7391: out = -2742;
			7392: out = -2707;
			7393: out = -2668;
			7394: out = -2621;
			7395: out = -2580;
			7396: out = -2555;
			7397: out = -2504;
			7398: out = -2480;
			7399: out = -2440;
			7400: out = -2398;
			7401: out = -2356;
			7402: out = -2323;
			7403: out = -2298;
			7404: out = -2258;
			7405: out = -2221;
			7406: out = -2183;
			7407: out = -2154;
			7408: out = -2129;
			7409: out = -2088;
			7410: out = -2051;
			7411: out = -2021;
			7412: out = -1992;
			7413: out = -1950;
			7414: out = -1924;
			7415: out = -1903;
			7416: out = -1862;
			7417: out = -1832;
			7418: out = -1804;
			7419: out = -1776;
			7420: out = -1750;
			7421: out = -1714;
			7422: out = -1694;
			7423: out = -1655;
			7424: out = -1627;
			7425: out = -1600;
			7426: out = -1576;
			7427: out = -1543;
			7428: out = -1515;
			7429: out = -1500;
			7430: out = -1465;
			7431: out = -1454;
			7432: out = -1426;
			7433: out = -1385;
			7434: out = -1370;
			7435: out = -1336;
			7436: out = -1316;
			7437: out = -1290;
			7438: out = -1269;
			7439: out = -1253;
			7440: out = -1219;
			7441: out = -1182;
			7442: out = -1146;
			7443: out = -1094;
			7444: out = -1073;
			7445: out = -1016;
			7446: out = -979;
			7447: out = -938;
			7448: out = -895;
			7449: out = -865;
			7450: out = -832;
			7451: out = -790;
			7452: out = -761;
			7453: out = -720;
			7454: out = -682;
			7455: out = -663;
			7456: out = -623;
			7457: out = -581;
			7458: out = -546;
			7459: out = -519;
			7460: out = -482;
			7461: out = -442;
			7462: out = -429;
			7463: out = -388;
			7464: out = -352;
			7465: out = -325;
			7466: out = -290;
			7467: out = -269;
			7468: out = -231;
			7469: out = -210;
			7470: out = -174;
			7471: out = -159;
			7472: out = -128;
			7473: out = -97;
			7474: out = -65;
			7475: out = -41;
			7476: out = -15;
			7477: out = 8;
			7478: out = 29;
			7479: out = 66;
			7480: out = 79;
			7481: out = 120;
			7482: out = 138;
			7483: out = 151;
			7484: out = 182;
			7485: out = 211;
			7486: out = 228;
			7487: out = 256;
			7488: out = 288;
			7489: out = 304;
			7490: out = 337;
			7491: out = 356;
			7492: out = 379;
			7493: out = 399;
			7494: out = 436;
			7495: out = 435;
			7496: out = 470;
			7497: out = 489;
			7498: out = 522;
			7499: out = 546;
			7500: out = 559;
			7501: out = 581;
			7502: out = 608;
			7503: out = 633;
			7504: out = 644;
			7505: out = 676;
			7506: out = 691;
			7507: out = 722;
			7508: out = 742;
			7509: out = 753;
			7510: out = 790;
			7511: out = 806;
			7512: out = 834;
			7513: out = 845;
			7514: out = 886;
			7515: out = 896;
			7516: out = 932;
			7517: out = 955;
			7518: out = 975;
			7519: out = 991;
			7520: out = 1035;
			7521: out = 1036;
			7522: out = 1069;
			7523: out = 1098;
			7524: out = 1121;
			7525: out = 1156;
			7526: out = 1168;
			7527: out = 1205;
			7528: out = 1226;
			7529: out = 1255;
			7530: out = 1280;
			7531: out = 1309;
			7532: out = 1341;
			7533: out = 1365;
			7534: out = 1393;
			7535: out = 1435;
			7536: out = 1468;
			7537: out = 1497;
			7538: out = 1528;
			7539: out = 1569;
			7540: out = 1600;
			7541: out = 1630;
			7542: out = 1684;
			7543: out = 1693;
			7544: out = 1749;
			7545: out = 1771;
			7546: out = 1813;
			7547: out = 1849;
			7548: out = 1865;
			7549: out = 1924;
			7550: out = 1949;
			7551: out = 1995;
			7552: out = 2032;
			7553: out = 2081;
			7554: out = 2117;
			7555: out = 2173;
			7556: out = 2193;
			7557: out = 2243;
			7558: out = 2293;
			7559: out = 2332;
			7560: out = 2370;
			7561: out = 2422;
			7562: out = 2464;
			7563: out = 2505;
			7564: out = 2548;
			7565: out = 2605;
			7566: out = 2632;
			7567: out = 2690;
			7568: out = 2722;
			7569: out = 2779;
			7570: out = 2809;
			7571: out = 2862;
			7572: out = 2898;
			7573: out = 2945;
			7574: out = 2988;
			7575: out = 3024;
			7576: out = 3066;
			7577: out = 3119;
			7578: out = 3160;
			7579: out = 3191;
			7580: out = 3245;
			7581: out = 3279;
			7582: out = 3317;
			7583: out = 3363;
			7584: out = 3397;
			7585: out = 3438;
			7586: out = 3476;
			7587: out = 3517;
			7588: out = 3555;
			7589: out = 3598;
			7590: out = 3619;
			7591: out = 3672;
			7592: out = 3706;
			7593: out = 3746;
			7594: out = 3778;
			7595: out = 3814;
			7596: out = 3838;
			7597: out = 3885;
			7598: out = 3921;
			7599: out = 3958;
			7600: out = 3988;
			7601: out = 4028;
			7602: out = 4053;
			7603: out = 4079;
			7604: out = 4115;
			7605: out = 4154;
			7606: out = 4183;
			7607: out = 4206;
			7608: out = 4247;
			7609: out = 4280;
			7610: out = 4301;
			7611: out = 4335;
			7612: out = 4364;
			7613: out = 4395;
			7614: out = 4415;
			7615: out = 4456;
			7616: out = 4472;
			7617: out = 4509;
			7618: out = 4538;
			7619: out = 4553;
			7620: out = 4577;
			7621: out = 4617;
			7622: out = 4637;
			7623: out = 4664;
			7624: out = 4687;
			7625: out = 4725;
			7626: out = 4749;
			7627: out = 4770;
			7628: out = 4786;
			7629: out = 4814;
			7630: out = 4844;
			7631: out = 4868;
			7632: out = 4873;
			7633: out = 4912;
			7634: out = 4926;
			7635: out = 4954;
			7636: out = 4976;
			7637: out = 4994;
			7638: out = 5025;
			7639: out = 5040;
			7640: out = 5066;
			7641: out = 5083;
			7642: out = 5107;
			7643: out = 5127;
			7644: out = 5149;
			7645: out = 5170;
			7646: out = 5197;
			7647: out = 5204;
			7648: out = 5223;
			7649: out = 5252;
			7650: out = 5270;
			7651: out = 5285;
			7652: out = 5314;
			7653: out = 5330;
			7654: out = 5351;
			7655: out = 5365;
			7656: out = 5397;
			7657: out = 5406;
			7658: out = 5422;
			7659: out = 5440;
			7660: out = 5456;
			7661: out = 5474;
			7662: out = 5501;
			7663: out = 5522;
			7664: out = 5523;
			7665: out = 5551;
			7666: out = 5567;
			7667: out = 5576;
			7668: out = 5603;
			7669: out = 5622;
			7670: out = 5615;
			7671: out = 5628;
			7672: out = 5669;
			7673: out = 5665;
			7674: out = 5672;
			7675: out = 5692;
			7676: out = 5674;
			7677: out = 5699;
			7678: out = 5676;
			7679: out = 5702;
			7680: out = 5694;
			7681: out = 5708;
			7682: out = 5692;
			7683: out = 5700;
			7684: out = 5694;
			7685: out = 5686;
			7686: out = 5684;
			7687: out = 5678;
			7688: out = 5708;
			7689: out = 5679;
			7690: out = 5681;
			7691: out = 5677;
			7692: out = 5681;
			7693: out = 5648;
			7694: out = 5651;
			7695: out = 5658;
			7696: out = 5648;
			7697: out = 5628;
			7698: out = 5634;
			7699: out = 5625;
			7700: out = 5633;
			7701: out = 5592;
			7702: out = 5604;
			7703: out = 5634;
			7704: out = 5610;
			7705: out = 5616;
			7706: out = 5608;
			7707: out = 5647;
			7708: out = 5622;
			7709: out = 5610;
			7710: out = 5622;
			7711: out = 5617;
			7712: out = 5594;
			7713: out = 5600;
			7714: out = 5575;
			7715: out = 5557;
			7716: out = 5594;
			7717: out = 5575;
			7718: out = 5595;
			7719: out = 5550;
			7720: out = 5592;
			7721: out = 5576;
			7722: out = 5571;
			7723: out = 5588;
			7724: out = 5602;
			7725: out = 5601;
			7726: out = 5580;
			7727: out = 5591;
			7728: out = 5580;
			7729: out = 5576;
			7730: out = 5570;
			7731: out = 5542;
			7732: out = 5537;
			7733: out = 5552;
			7734: out = 5515;
			7735: out = 5518;
			7736: out = 5506;
			7737: out = 5530;
			7738: out = 5510;
			7739: out = 5518;
			7740: out = 5504;
			7741: out = 5492;
			7742: out = 5477;
			7743: out = 5468;
			7744: out = 5476;
			7745: out = 5469;
			7746: out = 5446;
			7747: out = 5436;
			7748: out = 5423;
			7749: out = 5416;
			7750: out = 5382;
			7751: out = 5381;
			7752: out = 5361;
			7753: out = 5345;
			7754: out = 5341;
			7755: out = 5327;
			7756: out = 5294;
			7757: out = 5278;
			7758: out = 5258;
			7759: out = 5239;
			7760: out = 5240;
			7761: out = 5211;
			7762: out = 5173;
			7763: out = 5172;
			7764: out = 5114;
			7765: out = 5105;
			7766: out = 5089;
			7767: out = 5048;
			7768: out = 5042;
			7769: out = 5015;
			7770: out = 4967;
			7771: out = 4933;
			7772: out = 4930;
			7773: out = 4880;
			7774: out = 4842;
			7775: out = 4833;
			7776: out = 4789;
			7777: out = 4755;
			7778: out = 4752;
			7779: out = 4696;
			7780: out = 4684;
			7781: out = 4629;
			7782: out = 4600;
			7783: out = 4573;
			7784: out = 4527;
			7785: out = 4505;
			7786: out = 4474;
			7787: out = 4447;
			7788: out = 4409;
			7789: out = 4357;
			7790: out = 4344;
			7791: out = 4299;
			7792: out = 4252;
			7793: out = 4227;
			7794: out = 4192;
			7795: out = 4147;
			7796: out = 4097;
			7797: out = 4049;
			7798: out = 4013;
			7799: out = 3992;
			7800: out = 3945;
			7801: out = 3910;
			7802: out = 3890;
			7803: out = 3856;
			7804: out = 3833;
			7805: out = 3779;
			7806: out = 3745;
			7807: out = 3710;
			7808: out = 3654;
			7809: out = 3647;
			7810: out = 3567;
			7811: out = 3544;
			7812: out = 3511;
			7813: out = 3477;
			7814: out = 3441;
			7815: out = 3405;
			7816: out = 3380;
			7817: out = 3339;
			7818: out = 3290;
			7819: out = 3274;
			7820: out = 3244;
			7821: out = 3186;
			7822: out = 3148;
			7823: out = 3121;
			7824: out = 3082;
			7825: out = 3055;
			7826: out = 3027;
			7827: out = 2975;
			7828: out = 2963;
			7829: out = 2914;
			7830: out = 2884;
			7831: out = 2850;
			7832: out = 2836;
			7833: out = 2793;
			7834: out = 2736;
			7835: out = 2748;
			7836: out = 2680;
			7837: out = 2678;
			7838: out = 2629;
			7839: out = 2598;
			7840: out = 2584;
			7841: out = 2546;
			7842: out = 2517;
			7843: out = 2499;
			7844: out = 2444;
			7845: out = 2432;
			7846: out = 2383;
			7847: out = 2359;
			7848: out = 2347;
			7849: out = 2309;
			7850: out = 2275;
			7851: out = 2264;
			7852: out = 2215;
			7853: out = 2191;
			7854: out = 2178;
			7855: out = 2151;
			7856: out = 2128;
			7857: out = 2080;
			7858: out = 2073;
			7859: out = 2027;
			7860: out = 2021;
			7861: out = 2004;
			7862: out = 1961;
			7863: out = 1945;
			7864: out = 1913;
			7865: out = 1887;
			7866: out = 1875;
			7867: out = 1838;
			7868: out = 1815;
			7869: out = 1789;
			7870: out = 1755;
			7871: out = 1754;
			7872: out = 1720;
			7873: out = 1697;
			7874: out = 1679;
			7875: out = 1664;
			7876: out = 1629;
			7877: out = 1622;
			7878: out = 1593;
			7879: out = 1577;
			7880: out = 1536;
			7881: out = 1521;
			7882: out = 1513;
			7883: out = 1490;
			7884: out = 1465;
			7885: out = 1451;
			7886: out = 1439;
			7887: out = 1405;
			7888: out = 1383;
			7889: out = 1385;
			7890: out = 1357;
			7891: out = 1329;
			7892: out = 1321;
			7893: out = 1292;
			7894: out = 1281;
			7895: out = 1272;
			7896: out = 1233;
			7897: out = 1233;
			7898: out = 1201;
			7899: out = 1188;
			7900: out = 1175;
			7901: out = 1156;
			7902: out = 1141;
			7903: out = 1132;
			7904: out = 1114;
			7905: out = 1094;
			7906: out = 1081;
			7907: out = 1057;
			7908: out = 1028;
			7909: out = 992;
			7910: out = 951;
			7911: out = 885;
			7912: out = 843;
			7913: out = 793;
			7914: out = 768;
			7915: out = 727;
			7916: out = 677;
			7917: out = 654;
			7918: out = 611;
			7919: out = 558;
			7920: out = 529;
			7921: out = 489;
			7922: out = 452;
			7923: out = 418;
			7924: out = 389;
			7925: out = 339;
			7926: out = 298;
			7927: out = 292;
			7928: out = 225;
			7929: out = 205;
			7930: out = 163;
			7931: out = 127;
			7932: out = 108;
			7933: out = 52;
			7934: out = 37;
			7935: out = -3;
			7936: out = -36;
			7937: out = -63;
			7938: out = -101;
			7939: out = -125;
			7940: out = -151;
			7941: out = -185;
			7942: out = -229;
			7943: out = -241;
			7944: out = -281;
			7945: out = -306;
			7946: out = -329;
			7947: out = -372;
			7948: out = -387;
			7949: out = -423;
			7950: out = -434;
			7951: out = -469;
			7952: out = -493;
			7953: out = -533;
			7954: out = -559;
			7955: out = -572;
			7956: out = -618;
			7957: out = -628;
			7958: out = -653;
			7959: out = -695;
			7960: out = -709;
			7961: out = -739;
			7962: out = -756;
			7963: out = -788;
			7964: out = -813;
			7965: out = -855;
			7966: out = -868;
			7967: out = -891;
			7968: out = -928;
			7969: out = -945;
			7970: out = -967;
			7971: out = -997;
			7972: out = -1016;
			7973: out = -1043;
			7974: out = -1063;
			7975: out = -1093;
			7976: out = -1121;
			7977: out = -1142;
			7978: out = -1186;
			7979: out = -1188;
			7980: out = -1226;
			7981: out = -1245;
			7982: out = -1269;
			7983: out = -1298;
			7984: out = -1328;
			7985: out = -1352;
			7986: out = -1374;
			7987: out = -1403;
			7988: out = -1438;
			7989: out = -1436;
			7990: out = -1464;
			7991: out = -1501;
			7992: out = -1536;
			7993: out = -1561;
			7994: out = -1598;
			7995: out = -1631;
			7996: out = -1659;
			7997: out = -1686;
			7998: out = -1717;
			7999: out = -1749;
			8000: out = -1765;
			8001: out = -1809;
			8002: out = -1839;
			8003: out = -1867;
			8004: out = -1900;
			8005: out = -1939;
			8006: out = -1983;
			8007: out = -2006;
			8008: out = -2034;
			8009: out = -2077;
			8010: out = -2110;
			8011: out = -2142;
			8012: out = -2196;
			8013: out = -2216;
			8014: out = -2263;
			8015: out = -2290;
			8016: out = -2346;
			8017: out = -2373;
			8018: out = -2422;
			8019: out = -2462;
			8020: out = -2501;
			8021: out = -2540;
			8022: out = -2597;
			8023: out = -2636;
			8024: out = -2669;
			8025: out = -2723;
			8026: out = -2758;
			8027: out = -2821;
			8028: out = -2860;
			8029: out = -2913;
			8030: out = -2969;
			8031: out = -3006;
			8032: out = -3045;
			8033: out = -3109;
			8034: out = -3151;
			8035: out = -3197;
			8036: out = -3255;
			8037: out = -3308;
			8038: out = -3353;
			8039: out = -3409;
			8040: out = -3470;
			8041: out = -3505;
			8042: out = -3572;
			8043: out = -3616;
			8044: out = -3666;
			8045: out = -3712;
			8046: out = -3757;
			8047: out = -3814;
			8048: out = -3862;
			8049: out = -3910;
			8050: out = -3974;
			8051: out = -4005;
			8052: out = -4062;
			8053: out = -4095;
			8054: out = -4147;
			8055: out = -4193;
			8056: out = -4234;
			8057: out = -4284;
			8058: out = -4329;
			8059: out = -4367;
			8060: out = -4393;
			8061: out = -4452;
			8062: out = -4488;
			8063: out = -4526;
			8064: out = -4553;
			8065: out = -4608;
			8066: out = -4628;
			8067: out = -4675;
			8068: out = -4713;
			8069: out = -4736;
			8070: out = -4774;
			8071: out = -4808;
			8072: out = -4829;
			8073: out = -4879;
			8074: out = -4886;
			8075: out = -4928;
			8076: out = -4956;
			8077: out = -4992;
			8078: out = -5004;
			8079: out = -5048;
			8080: out = -5067;
			8081: out = -5102;
			8082: out = -5126;
			8083: out = -5145;
			8084: out = -5160;
			8085: out = -5190;
			8086: out = -5214;
			8087: out = -5214;
			8088: out = -5253;
			8089: out = -5272;
			8090: out = -5284;
			8091: out = -5307;
			8092: out = -5328;
			8093: out = -5342;
			8094: out = -5361;
			8095: out = -5357;
			8096: out = -5389;
			8097: out = -5389;
			8098: out = -5418;
			8099: out = -5423;
			8100: out = -5425;
			8101: out = -5447;
			8102: out = -5454;
			8103: out = -5470;
			8104: out = -5484;
			8105: out = -5492;
			8106: out = -5496;
			8107: out = -5509;
			8108: out = -5500;
			8109: out = -5531;
			8110: out = -5515;
			8111: out = -5533;
			8112: out = -5548;
			8113: out = -5542;
			8114: out = -5550;
			8115: out = -5564;
			8116: out = -5562;
			8117: out = -5563;
			8118: out = -5567;
			8119: out = -5570;
			8120: out = -5581;
			8121: out = -5581;
			8122: out = -5577;
			8123: out = -5581;
			8124: out = -5577;
			8125: out = -5587;
			8126: out = -5596;
			8127: out = -5587;
			8128: out = -5591;
			8129: out = -5581;
			8130: out = -5588;
			8131: out = -5579;
			8132: out = -5580;
			8133: out = -5596;
			8134: out = -5563;
			8135: out = -5576;
			8136: out = -5569;
			8137: out = -5574;
			8138: out = -5572;
			8139: out = -5559;
			8140: out = -5563;
			8141: out = -5548;
			8142: out = -5554;
			8143: out = -5545;
			8144: out = -5534;
			8145: out = -5535;
			8146: out = -5527;
			8147: out = -5510;
			8148: out = -5517;
			8149: out = -5519;
			8150: out = -5495;
			8151: out = -5493;
			8152: out = -5505;
			8153: out = -5474;
			8154: out = -5474;
			8155: out = -5463;
			8156: out = -5453;
			8157: out = -5457;
			8158: out = -5441;
			8159: out = -5425;
			8160: out = -5421;
			8161: out = -5414;
			8162: out = -5406;
			8163: out = -5403;
			8164: out = -5398;
			8165: out = -5366;
			8166: out = -5376;
			8167: out = -5376;
			8168: out = -5354;
			8169: out = -5349;
			8170: out = -5329;
			8171: out = -5323;
			8172: out = -5314;
			8173: out = -5298;
			8174: out = -5284;
			8175: out = -5267;
			8176: out = -5259;
			8177: out = -5237;
			8178: out = -5226;
			8179: out = -5233;
			8180: out = -5204;
			8181: out = -5184;
			8182: out = -5181;
			8183: out = -5170;
			8184: out = -5149;
			8185: out = -5138;
			8186: out = -5126;
			8187: out = -5117;
			8188: out = -5090;
			8189: out = -5095;
			8190: out = -5073;
			8191: out = -5056;
			8192: out = -5044;
			8193: out = -5030;
			8194: out = -5011;
			8195: out = -4992;
			8196: out = -4982;
			8197: out = -4967;
			8198: out = -4955;
			8199: out = -4931;
			8200: out = -4907;
			8201: out = -4900;
			8202: out = -4881;
			8203: out = -4872;
			8204: out = -4842;
			8205: out = -4831;
			8206: out = -4807;
			8207: out = -4790;
			8208: out = -4756;
			8209: out = -4765;
			8210: out = -4715;
			8211: out = -4711;
			8212: out = -4673;
			8213: out = -4667;
			8214: out = -4642;
			8215: out = -4611;
			8216: out = -4589;
			8217: out = -4561;
			8218: out = -4538;
			8219: out = -4502;
			8220: out = -4487;
			8221: out = -4450;
			8222: out = -4420;
			8223: out = -4393;
			8224: out = -4359;
			8225: out = -4345;
			8226: out = -4312;
			8227: out = -4264;
			8228: out = -4250;
			8229: out = -4194;
			8230: out = -4171;
			8231: out = -4136;
			8232: out = -4104;
			8233: out = -4054;
			8234: out = -4039;
			8235: out = -3992;
			8236: out = -3954;
			8237: out = -3925;
			8238: out = -3891;
			8239: out = -3846;
			8240: out = -3813;
			8241: out = -3762;
			8242: out = -3736;
			8243: out = -3685;
			8244: out = -3652;
			8245: out = -3622;
			8246: out = -3564;
			8247: out = -3541;
			8248: out = -3510;
			8249: out = -3454;
			8250: out = -3428;
			8251: out = -3369;
			8252: out = -3335;
			8253: out = -3300;
			8254: out = -3256;
			8255: out = -3224;
			8256: out = -3186;
			8257: out = -3146;
			8258: out = -3109;
			8259: out = -3069;
			8260: out = -3027;
			8261: out = -2991;
			8262: out = -2954;
			8263: out = -2917;
			8264: out = -2878;
			8265: out = -2845;
			8266: out = -2795;
			8267: out = -2786;
			8268: out = -2722;
			8269: out = -2696;
			8270: out = -2661;
			8271: out = -2614;
			8272: out = -2593;
			8273: out = -2542;
			8274: out = -2517;
			8275: out = -2476;
			8276: out = -2446;
			8277: out = -2408;
			8278: out = -2377;
			8279: out = -2349;
			8280: out = -2302;
			8281: out = -2274;
			8282: out = -2245;
			8283: out = -2205;
			8284: out = -2188;
			8285: out = -2142;
			8286: out = -2110;
			8287: out = -2089;
			8288: out = -2048;
			8289: out = -2022;
			8290: out = -1983;
			8291: out = -1969;
			8292: out = -1931;
			8293: out = -1902;
			8294: out = -1874;
			8295: out = -1848;
			8296: out = -1816;
			8297: out = -1790;
			8298: out = -1753;
			8299: out = -1735;
			8300: out = -1703;
			8301: out = -1672;
			8302: out = -1655;
			8303: out = -1629;
			8304: out = -1592;
			8305: out = -1588;
			8306: out = -1547;
			8307: out = -1520;
			8308: out = -1495;
			8309: out = -1471;
			8310: out = -1457;
			8311: out = -1424;
			8312: out = -1410;
			8313: out = -1361;
			8314: out = -1364;
			8315: out = -1338;
			8316: out = -1300;
			8317: out = -1292;
			8318: out = -1268;
			8319: out = -1239;
			8320: out = -1221;
			8321: out = -1198;
			8322: out = -1178;
			8323: out = -1160;
			8324: out = -1131;
			8325: out = -1118;
			8326: out = -1106;
			8327: out = -1081;
			8328: out = -1052;
			8329: out = -1043;
			8330: out = -1016;
			8331: out = -995;
			8332: out = -972;
			8333: out = -948;
			8334: out = -907;
			8335: out = -872;
			8336: out = -848;
			8337: out = -803;
			8338: out = -780;
			8339: out = -754;
			8340: out = -704;
			8341: out = -688;
			8342: out = -655;
			8343: out = -628;
			8344: out = -595;
			8345: out = -565;
			8346: out = -549;
			8347: out = -510;
			8348: out = -488;
			8349: out = -455;
			8350: out = -432;
			8351: out = -398;
			8352: out = -393;
			8353: out = -360;
			8354: out = -336;
			8355: out = -305;
			8356: out = -286;
			8357: out = -252;
			8358: out = -225;
			8359: out = -216;
			8360: out = -176;
			8361: out = -156;
			8362: out = -145;
			8363: out = -119;
			8364: out = -81;
			8365: out = -72;
			8366: out = -41;
			8367: out = -30;
			8368: out = -14;
			8369: out = 9;
			8370: out = 50;
			8371: out = 46;
			8372: out = 75;
			8373: out = 105;
			8374: out = 114;
			8375: out = 138;
			8376: out = 162;
			8377: out = 176;
			8378: out = 194;
			8379: out = 225;
			8380: out = 231;
			8381: out = 262;
			8382: out = 274;
			8383: out = 303;
			8384: out = 301;
			8385: out = 341;
			8386: out = 350;
			8387: out = 364;
			8388: out = 395;
			8389: out = 404;
			8390: out = 428;
			8391: out = 443;
			8392: out = 462;
			8393: out = 484;
			8394: out = 491;
			8395: out = 522;
			8396: out = 538;
			8397: out = 550;
			8398: out = 573;
			8399: out = 582;
			8400: out = 614;
			8401: out = 630;
			8402: out = 645;
			8403: out = 653;
			8404: out = 685;
			8405: out = 702;
			8406: out = 726;
			8407: out = 731;
			8408: out = 762;
			8409: out = 771;
			8410: out = 800;
			8411: out = 821;
			8412: out = 836;
			8413: out = 866;
			8414: out = 871;
			8415: out = 906;
			8416: out = 921;
			8417: out = 940;
			8418: out = 969;
			8419: out = 983;
			8420: out = 1011;
			8421: out = 1035;
			8422: out = 1059;
			8423: out = 1073;
			8424: out = 1108;
			8425: out = 1121;
			8426: out = 1150;
			8427: out = 1173;
			8428: out = 1205;
			8429: out = 1233;
			8430: out = 1259;
			8431: out = 1290;
			8432: out = 1305;
			8433: out = 1344;
			8434: out = 1358;
			8435: out = 1398;
			8436: out = 1414;
			8437: out = 1461;
			8438: out = 1486;
			8439: out = 1523;
			8440: out = 1552;
			8441: out = 1576;
			8442: out = 1614;
			8443: out = 1640;
			8444: out = 1674;
			8445: out = 1693;
			8446: out = 1746;
			8447: out = 1769;
			8448: out = 1806;
			8449: out = 1847;
			8450: out = 1878;
			8451: out = 1913;
			8452: out = 1950;
			8453: out = 1990;
			8454: out = 2013;
			8455: out = 2053;
			8456: out = 2098;
			8457: out = 2124;
			8458: out = 2169;
			8459: out = 2197;
			8460: out = 2240;
			8461: out = 2265;
			8462: out = 2304;
			8463: out = 2346;
			8464: out = 2384;
			8465: out = 2406;
			8466: out = 2447;
			8467: out = 2479;
			8468: out = 2512;
			8469: out = 2554;
			8470: out = 2577;
			8471: out = 2618;
			8472: out = 2654;
			8473: out = 2683;
			8474: out = 2720;
			8475: out = 2762;
			8476: out = 2782;
			8477: out = 2815;
			8478: out = 2849;
			8479: out = 2882;
			8480: out = 2906;
			8481: out = 2950;
			8482: out = 2979;
			8483: out = 3008;
			8484: out = 3035;
			8485: out = 3071;
			8486: out = 3087;
			8487: out = 3127;
			8488: out = 3152;
			8489: out = 3166;
			8490: out = 3212;
			8491: out = 3227;
			8492: out = 3264;
			8493: out = 3296;
			8494: out = 3308;
			8495: out = 3345;
			8496: out = 3363;
			8497: out = 3393;
			8498: out = 3421;
			8499: out = 3441;
			8500: out = 3458;
			8501: out = 3489;
			8502: out = 3515;
			8503: out = 3529;
			8504: out = 3575;
			8505: out = 3583;
			8506: out = 3610;
			8507: out = 3640;
			8508: out = 3645;
			8509: out = 3682;
			8510: out = 3707;
			8511: out = 3717;
			8512: out = 3736;
			8513: out = 3762;
			8514: out = 3778;
			8515: out = 3816;
			8516: out = 3830;
			8517: out = 3849;
			8518: out = 3877;
			8519: out = 3880;
			8520: out = 3917;
			8521: out = 3932;
			8522: out = 3966;
			8523: out = 3980;
			8524: out = 3996;
			8525: out = 4018;
			8526: out = 4034;
			8527: out = 4042;
			8528: out = 4072;
			8529: out = 4076;
			8530: out = 4109;
			8531: out = 4122;
			8532: out = 4120;
			8533: out = 4159;
			8534: out = 4169;
			8535: out = 4185;
			8536: out = 4203;
			8537: out = 4225;
			8538: out = 4239;
			8539: out = 4255;
			8540: out = 4255;
			8541: out = 4290;
			8542: out = 4292;
			8543: out = 4317;
			8544: out = 4340;
			8545: out = 4356;
			8546: out = 4359;
			8547: out = 4382;
			8548: out = 4404;
			8549: out = 4405;
			8550: out = 4433;
			8551: out = 4439;
			8552: out = 4447;
			8553: out = 4479;
			8554: out = 4490;
			8555: out = 4497;
			8556: out = 4524;
			8557: out = 4528;
			8558: out = 4547;
			8559: out = 4552;
			8560: out = 4584;
			8561: out = 4586;
			8562: out = 4599;
			8563: out = 4604;
			8564: out = 4635;
			8565: out = 4631;
			8566: out = 4634;
			8567: out = 4655;
			8568: out = 4661;
			8569: out = 4656;
			8570: out = 4640;
			8571: out = 4657;
			8572: out = 4651;
			8573: out = 4633;
			8574: out = 4635;
			8575: out = 4658;
			8576: out = 4630;
			8577: out = 4632;
			8578: out = 4636;
			8579: out = 4629;
			8580: out = 4642;
			8581: out = 4625;
			8582: out = 4621;
			8583: out = 4617;
			8584: out = 4634;
			8585: out = 4636;
			8586: out = 4590;
			8587: out = 4607;
			8588: out = 4616;
			8589: out = 4617;
			8590: out = 4604;
			8591: out = 4618;
			8592: out = 4620;
			8593: out = 4612;
			8594: out = 4598;
			8595: out = 4623;
			8596: out = 4598;
			8597: out = 4596;
			8598: out = 4584;
			8599: out = 4594;
			8600: out = 4587;
			8601: out = 4584;
			8602: out = 4569;
			8603: out = 4588;
			8604: out = 4593;
			8605: out = 4574;
			8606: out = 4588;
			8607: out = 4593;
			8608: out = 4573;
			8609: out = 4585;
			8610: out = 4559;
			8611: out = 4563;
			8612: out = 4568;
			8613: out = 4573;
			8614: out = 4587;
			8615: out = 4575;
			8616: out = 4565;
			8617: out = 4562;
			8618: out = 4574;
			8619: out = 4578;
			8620: out = 4554;
			8621: out = 4553;
			8622: out = 4559;
			8623: out = 4546;
			8624: out = 4533;
			8625: out = 4531;
			8626: out = 4525;
			8627: out = 4522;
			8628: out = 4535;
			8629: out = 4529;
			8630: out = 4518;
			8631: out = 4493;
			8632: out = 4510;
			8633: out = 4503;
			8634: out = 4482;
			8635: out = 4497;
			8636: out = 4481;
			8637: out = 4499;
			8638: out = 4463;
			8639: out = 4446;
			8640: out = 4445;
			8641: out = 4447;
			8642: out = 4429;
			8643: out = 4423;
			8644: out = 4414;
			8645: out = 4404;
			8646: out = 4375;
			8647: out = 4369;
			8648: out = 4383;
			8649: out = 4347;
			8650: out = 4314;
			8651: out = 4317;
			8652: out = 4301;
			8653: out = 4270;
			8654: out = 4249;
			8655: out = 4234;
			8656: out = 4209;
			8657: out = 4183;
			8658: out = 4180;
			8659: out = 4166;
			8660: out = 4140;
			8661: out = 4120;
			8662: out = 4089;
			8663: out = 4066;
			8664: out = 4052;
			8665: out = 4027;
			8666: out = 3984;
			8667: out = 3959;
			8668: out = 3936;
			8669: out = 3921;
			8670: out = 3890;
			8671: out = 3861;
			8672: out = 3844;
			8673: out = 3808;
			8674: out = 3788;
			8675: out = 3746;
			8676: out = 3726;
			8677: out = 3693;
			8678: out = 3676;
			8679: out = 3640;
			8680: out = 3601;
			8681: out = 3574;
			8682: out = 3556;
			8683: out = 3520;
			8684: out = 3499;
			8685: out = 3448;
			8686: out = 3417;
			8687: out = 3394;
			8688: out = 3378;
			8689: out = 3339;
			8690: out = 3310;
			8691: out = 3278;
			8692: out = 3250;
			8693: out = 3227;
			8694: out = 3185;
			8695: out = 3148;
			8696: out = 3130;
			8697: out = 3090;
			8698: out = 3059;
			8699: out = 3047;
			8700: out = 3013;
			8701: out = 2994;
			8702: out = 2959;
			8703: out = 2924;
			8704: out = 2889;
			8705: out = 2842;
			8706: out = 2835;
			8707: out = 2800;
			8708: out = 2752;
			8709: out = 2754;
			8710: out = 2705;
			8711: out = 2691;
			8712: out = 2642;
			8713: out = 2630;
			8714: out = 2601;
			8715: out = 2558;
			8716: out = 2540;
			8717: out = 2514;
			8718: out = 2491;
			8719: out = 2451;
			8720: out = 2435;
			8721: out = 2400;
			8722: out = 2391;
			8723: out = 2346;
			8724: out = 2317;
			8725: out = 2292;
			8726: out = 2277;
			8727: out = 2231;
			8728: out = 2219;
			8729: out = 2183;
			8730: out = 2164;
			8731: out = 2136;
			8732: out = 2115;
			8733: out = 2092;
			8734: out = 2063;
			8735: out = 2049;
			8736: out = 2002;
			8737: out = 1992;
			8738: out = 1967;
			8739: out = 1947;
			8740: out = 1923;
			8741: out = 1903;
			8742: out = 1868;
			8743: out = 1850;
			8744: out = 1823;
			8745: out = 1812;
			8746: out = 1771;
			8747: out = 1754;
			8748: out = 1725;
			8749: out = 1713;
			8750: out = 1690;
			8751: out = 1677;
			8752: out = 1648;
			8753: out = 1630;
			8754: out = 1611;
			8755: out = 1586;
			8756: out = 1574;
			8757: out = 1555;
			8758: out = 1530;
			8759: out = 1506;
			8760: out = 1483;
			8761: out = 1465;
			8762: out = 1452;
			8763: out = 1415;
			8764: out = 1415;
			8765: out = 1375;
			8766: out = 1373;
			8767: out = 1350;
			8768: out = 1334;
			8769: out = 1310;
			8770: out = 1299;
			8771: out = 1265;
			8772: out = 1259;
			8773: out = 1235;
			8774: out = 1225;
			8775: out = 1206;
			8776: out = 1177;
			8777: out = 1169;
			8778: out = 1151;
			8779: out = 1150;
			8780: out = 1125;
			8781: out = 1106;
			8782: out = 1082;
			8783: out = 1077;
			8784: out = 1057;
			8785: out = 1047;
			8786: out = 1032;
			8787: out = 1015;
			8788: out = 1003;
			8789: out = 997;
			8790: out = 963;
			8791: out = 963;
			8792: out = 948;
			8793: out = 917;
			8794: out = 922;
			8795: out = 910;
			8796: out = 893;
			8797: out = 879;
			8798: out = 867;
			8799: out = 856;
			8800: out = 811;
			8801: out = 771;
			8802: out = 724;
			8803: out = 693;
			8804: out = 663;
			8805: out = 624;
			8806: out = 597;
			8807: out = 555;
			8808: out = 535;
			8809: out = 490;
			8810: out = 463;
			8811: out = 421;
			8812: out = 382;
			8813: out = 357;
			8814: out = 329;
			8815: out = 299;
			8816: out = 270;
			8817: out = 249;
			8818: out = 199;
			8819: out = 182;
			8820: out = 154;
			8821: out = 111;
			8822: out = 98;
			8823: out = 64;
			8824: out = 37;
			8825: out = 13;
			8826: out = -9;
			8827: out = -20;
			8828: out = -70;
			8829: out = -84;
			8830: out = -117;
			8831: out = -132;
			8832: out = -156;
			8833: out = -188;
			8834: out = -209;
			8835: out = -241;
			8836: out = -257;
			8837: out = -286;
			8838: out = -304;
			8839: out = -323;
			8840: out = -356;
			8841: out = -370;
			8842: out = -404;
			8843: out = -423;
			8844: out = -439;
			8845: out = -468;
			8846: out = -495;
			8847: out = -516;
			8848: out = -529;
			8849: out = -567;
			8850: out = -572;
			8851: out = -610;
			8852: out = -621;
			8853: out = -638;
			8854: out = -680;
			8855: out = -677;
			8856: out = -707;
			8857: out = -727;
			8858: out = -759;
			8859: out = -765;
			8860: out = -798;
			8861: out = -813;
			8862: out = -831;
			8863: out = -861;
			8864: out = -872;
			8865: out = -894;
			8866: out = -916;
			8867: out = -931;
			8868: out = -959;
			8869: out = -975;
			8870: out = -998;
			8871: out = -1014;
			8872: out = -1036;
			8873: out = -1055;
			8874: out = -1077;
			8875: out = -1109;
			8876: out = -1116;
			8877: out = -1154;
			8878: out = -1158;
			8879: out = -1187;
			8880: out = -1221;
			8881: out = -1235;
			8882: out = -1268;
			8883: out = -1284;
			8884: out = -1306;
			8885: out = -1330;
			8886: out = -1350;
			8887: out = -1361;
			8888: out = -1394;
			8889: out = -1418;
			8890: out = -1453;
			8891: out = -1477;
			8892: out = -1505;
			8893: out = -1527;
			8894: out = -1565;
			8895: out = -1579;
			8896: out = -1600;
			8897: out = -1646;
			8898: out = -1653;
			8899: out = -1687;
			8900: out = -1717;
			8901: out = -1755;
			8902: out = -1774;
			8903: out = -1802;
			8904: out = -1840;
			8905: out = -1865;
			8906: out = -1894;
			8907: out = -1933;
			8908: out = -1969;
			8909: out = -2001;
			8910: out = -2030;
			8911: out = -2051;
			8912: out = -2089;
			8913: out = -2125;
			8914: out = -2156;
			8915: out = -2204;
			8916: out = -2230;
			8917: out = -2270;
			8918: out = -2306;
			8919: out = -2356;
			8920: out = -2384;
			8921: out = -2433;
			8922: out = -2471;
			8923: out = -2511;
			8924: out = -2557;
			8925: out = -2595;
			8926: out = -2630;
			8927: out = -2675;
			8928: out = -2723;
			8929: out = -2750;
			8930: out = -2795;
			8931: out = -2847;
			8932: out = -2885;
			8933: out = -2929;
			8934: out = -2964;
			8935: out = -3004;
			8936: out = -3048;
			8937: out = -3096;
			8938: out = -3126;
			8939: out = -3170;
			8940: out = -3214;
			8941: out = -3246;
			8942: out = -3282;
			8943: out = -3335;
			8944: out = -3362;
			8945: out = -3391;
			8946: out = -3446;
			8947: out = -3471;
			8948: out = -3499;
			8949: out = -3545;
			8950: out = -3584;
			8951: out = -3618;
			8952: out = -3640;
			8953: out = -3681;
			8954: out = -3725;
			8955: out = -3745;
			8956: out = -3779;
			8957: out = -3808;
			8958: out = -3835;
			8959: out = -3875;
			8960: out = -3890;
			8961: out = -3925;
			8962: out = -3963;
			8963: out = -3969;
			8964: out = -4010;
			8965: out = -4024;
			8966: out = -4059;
			8967: out = -4080;
			8968: out = -4096;
			8969: out = -4119;
			8970: out = -4149;
			8971: out = -4157;
			8972: out = -4178;
			8973: out = -4205;
			8974: out = -4228;
			8975: out = -4226;
			8976: out = -4265;
			8977: out = -4267;
			8978: out = -4298;
			8979: out = -4303;
			8980: out = -4343;
			8981: out = -4330;
			8982: out = -4363;
			8983: out = -4375;
			8984: out = -4381;
			8985: out = -4392;
			8986: out = -4400;
			8987: out = -4427;
			8988: out = -4434;
			8989: out = -4441;
			8990: out = -4453;
			8991: out = -4465;
			8992: out = -4475;
			8993: out = -4480;
			8994: out = -4490;
			8995: out = -4502;
			8996: out = -4513;
			8997: out = -4517;
			8998: out = -4523;
			8999: out = -4528;
			9000: out = -4523;
			9001: out = -4546;
			9002: out = -4542;
			9003: out = -4540;
			9004: out = -4559;
			9005: out = -4545;
			9006: out = -4557;
			9007: out = -4578;
			9008: out = -4562;
			9009: out = -4576;
			9010: out = -4562;
			9011: out = -4581;
			9012: out = -4575;
			9013: out = -4583;
			9014: out = -4570;
			9015: out = -4590;
			9016: out = -4571;
			9017: out = -4583;
			9018: out = -4581;
			9019: out = -4577;
			9020: out = -4590;
			9021: out = -4574;
			9022: out = -4571;
			9023: out = -4583;
			9024: out = -4574;
			9025: out = -4559;
			9026: out = -4583;
			9027: out = -4563;
			9028: out = -4554;
			9029: out = -4571;
			9030: out = -4564;
			9031: out = -4547;
			9032: out = -4558;
			9033: out = -4547;
			9034: out = -4546;
			9035: out = -4534;
			9036: out = -4531;
			9037: out = -4535;
			9038: out = -4526;
			9039: out = -4518;
			9040: out = -4507;
			9041: out = -4516;
			9042: out = -4507;
			9043: out = -4497;
			9044: out = -4491;
			9045: out = -4480;
			9046: out = -4491;
			9047: out = -4471;
			9048: out = -4460;
			9049: out = -4456;
			9050: out = -4455;
			9051: out = -4434;
			9052: out = -4435;
			9053: out = -4431;
			9054: out = -4422;
			9055: out = -4412;
			9056: out = -4405;
			9057: out = -4388;
			9058: out = -4383;
			9059: out = -4379;
			9060: out = -4370;
			9061: out = -4357;
			9062: out = -4357;
			9063: out = -4333;
			9064: out = -4345;
			9065: out = -4336;
			9066: out = -4310;
			9067: out = -4310;
			9068: out = -4289;
			9069: out = -4288;
			9070: out = -4269;
			9071: out = -4259;
			9072: out = -4254;
			9073: out = -4239;
			9074: out = -4223;
			9075: out = -4208;
			9076: out = -4205;
			9077: out = -4203;
			9078: out = -4184;
			9079: out = -4174;
			9080: out = -4172;
			9081: out = -4152;
			9082: out = -4145;
			9083: out = -4122;
			9084: out = -4117;
			9085: out = -4107;
			9086: out = -4096;
			9087: out = -4077;
			9088: out = -4064;
			9089: out = -4048;
			9090: out = -4040;
			9091: out = -4021;
			9092: out = -4010;
			9093: out = -3998;
			9094: out = -3982;
			9095: out = -3958;
			9096: out = -3953;
			9097: out = -3937;
			9098: out = -3915;
			9099: out = -3907;
			9100: out = -3886;
			9101: out = -3866;
			9102: out = -3850;
			9103: out = -3828;
			9104: out = -3804;
			9105: out = -3791;
			9106: out = -3771;
			9107: out = -3750;
			9108: out = -3731;
			9109: out = -3716;
			9110: out = -3691;
			9111: out = -3666;
			9112: out = -3647;
			9113: out = -3615;
			9114: out = -3595;
			9115: out = -3567;
			9116: out = -3549;
			9117: out = -3518;
			9118: out = -3493;
			9119: out = -3466;
			9120: out = -3442;
			9121: out = -3414;
			9122: out = -3390;
			9123: out = -3354;
			9124: out = -3324;
			9125: out = -3300;
			9126: out = -3268;
			9127: out = -3234;
			9128: out = -3212;
			9129: out = -3179;
			9130: out = -3144;
			9131: out = -3116;
			9132: out = -3094;
			9133: out = -3051;
			9134: out = -3027;
			9135: out = -2985;
			9136: out = -2960;
			9137: out = -2926;
			9138: out = -2897;
			9139: out = -2856;
			9140: out = -2836;
			9141: out = -2797;
			9142: out = -2767;
			9143: out = -2738;
			9144: out = -2700;
			9145: out = -2680;
			9146: out = -2642;
			9147: out = -2601;
			9148: out = -2571;
			9149: out = -2540;
			9150: out = -2493;
			9151: out = -2484;
			9152: out = -2441;
			9153: out = -2422;
			9154: out = -2383;
			9155: out = -2352;
			9156: out = -2333;
			9157: out = -2288;
			9158: out = -2269;
			9159: out = -2229;
			9160: out = -2211;
			9161: out = -2167;
			9162: out = -2147;
			9163: out = -2108;
			9164: out = -2091;
			9165: out = -2061;
			9166: out = -2029;
			9167: out = -2000;
			9168: out = -1980;
			9169: out = -1947;
			9170: out = -1911;
			9171: out = -1889;
			9172: out = -1862;
			9173: out = -1840;
			9174: out = -1806;
			9175: out = -1780;
			9176: out = -1765;
			9177: out = -1724;
			9178: out = -1708;
			9179: out = -1685;
			9180: out = -1650;
			9181: out = -1628;
			9182: out = -1608;
			9183: out = -1571;
			9184: out = -1553;
			9185: out = -1543;
			9186: out = -1509;
			9187: out = -1486;
			9188: out = -1466;
			9189: out = -1435;
			9190: out = -1417;
			9191: out = -1398;
			9192: out = -1369;
			9193: out = -1357;
			9194: out = -1326;
			9195: out = -1309;
			9196: out = -1298;
			9197: out = -1259;
			9198: out = -1255;
			9199: out = -1227;
			9200: out = -1205;
			9201: out = -1190;
			9202: out = -1157;
			9203: out = -1152;
			9204: out = -1131;
			9205: out = -1102;
			9206: out = -1086;
			9207: out = -1089;
			9208: out = -1046;
			9209: out = -1043;
			9210: out = -1003;
			9211: out = -1011;
			9212: out = -979;
			9213: out = -955;
			9214: out = -956;
			9215: out = -931;
			9216: out = -920;
			9217: out = -890;
			9218: out = -885;
			9219: out = -860;
			9220: out = -854;
			9221: out = -824;
			9222: out = -822;
			9223: out = -806;
			9224: out = -776;
			9225: out = -741;
			9226: out = -725;
			9227: out = -693;
			9228: out = -661;
			9229: out = -642;
			9230: out = -613;
			9231: out = -593;
			9232: out = -570;
			9233: out = -539;
			9234: out = -518;
			9235: out = -501;
			9236: out = -457;
			9237: out = -450;
			9238: out = -423;
			9239: out = -405;
			9240: out = -372;
			9241: out = -360;
			9242: out = -346;
			9243: out = -316;
			9244: out = -289;
			9245: out = -286;
			9246: out = -261;
			9247: out = -227;
			9248: out = -218;
			9249: out = -200;
			9250: out = -193;
			9251: out = -149;
			9252: out = -148;
			9253: out = -126;
			9254: out = -101;
			9255: out = -80;
			9256: out = -70;
			9257: out = -43;
			9258: out = -38;
			9259: out = -9;
			9260: out = 5;
			9261: out = 21;
			9262: out = 34;
			9263: out = 64;
			9264: out = 74;
			9265: out = 89;
			9266: out = 105;
			9267: out = 112;
			9268: out = 134;
			9269: out = 161;
			9270: out = 159;
			9271: out = 187;
			9272: out = 204;
			9273: out = 200;
			9274: out = 227;
			9275: out = 254;
			9276: out = 252;
			9277: out = 274;
			9278: out = 293;
			9279: out = 310;
			9280: out = 316;
			9281: out = 333;
			9282: out = 353;
			9283: out = 359;
			9284: out = 372;
			9285: out = 401;
			9286: out = 403;
			9287: out = 434;
			9288: out = 434;
			9289: out = 447;
			9290: out = 476;
			9291: out = 480;
			9292: out = 502;
			9293: out = 519;
			9294: out = 531;
			9295: out = 529;
			9296: out = 566;
			9297: out = 571;
			9298: out = 586;
			9299: out = 605;
			9300: out = 622;
			9301: out = 633;
			9302: out = 663;
			9303: out = 665;
			9304: out = 693;
			9305: out = 703;
			9306: out = 711;
			9307: out = 739;
			9308: out = 755;
			9309: out = 771;
			9310: out = 785;
			9311: out = 815;
			9312: out = 821;
			9313: out = 849;
			9314: out = 856;
			9315: out = 885;
			9316: out = 901;
			9317: out = 917;
			9318: out = 951;
			9319: out = 954;
			9320: out = 980;
			9321: out = 1000;
			9322: out = 1034;
			9323: out = 1043;
			9324: out = 1066;
			9325: out = 1096;
			9326: out = 1113;
			9327: out = 1140;
			9328: out = 1165;
			9329: out = 1188;
			9330: out = 1204;
			9331: out = 1239;
			9332: out = 1259;
			9333: out = 1295;
			9334: out = 1310;
			9335: out = 1354;
			9336: out = 1363;
			9337: out = 1405;
			9338: out = 1424;
			9339: out = 1460;
			9340: out = 1475;
			9341: out = 1507;
			9342: out = 1535;
			9343: out = 1563;
			9344: out = 1598;
			9345: out = 1622;
			9346: out = 1657;
			9347: out = 1683;
			9348: out = 1710;
			9349: out = 1742;
			9350: out = 1771;
			9351: out = 1796;
			9352: out = 1835;
			9353: out = 1855;
			9354: out = 1902;
			9355: out = 1914;
			9356: out = 1946;
			9357: out = 1981;
			9358: out = 2001;
			9359: out = 2028;
			9360: out = 2067;
			9361: out = 2091;
			9362: out = 2114;
			9363: out = 2152;
			9364: out = 2168;
			9365: out = 2200;
			9366: out = 2223;
			9367: out = 2254;
			9368: out = 2275;
			9369: out = 2309;
			9370: out = 2325;
			9371: out = 2368;
			9372: out = 2381;
			9373: out = 2399;
			9374: out = 2442;
			9375: out = 2450;
			9376: out = 2481;
			9377: out = 2498;
			9378: out = 2535;
			9379: out = 2553;
			9380: out = 2574;
			9381: out = 2605;
			9382: out = 2621;
			9383: out = 2641;
			9384: out = 2670;
			9385: out = 2688;
			9386: out = 2714;
			9387: out = 2726;
			9388: out = 2752;
			9389: out = 2784;
			9390: out = 2787;
			9391: out = 2811;
			9392: out = 2831;
			9393: out = 2856;
			9394: out = 2871;
			9395: out = 2901;
			9396: out = 2916;
			9397: out = 2932;
			9398: out = 2953;
			9399: out = 2971;
			9400: out = 2984;
			9401: out = 3012;
			9402: out = 3024;
			9403: out = 3049;
			9404: out = 3063;
			9405: out = 3070;
			9406: out = 3102;
			9407: out = 3115;
			9408: out = 3134;
			9409: out = 3145;
			9410: out = 3172;
			9411: out = 3170;
			9412: out = 3211;
			9413: out = 3209;
			9414: out = 3229;
			9415: out = 3241;
			9416: out = 3262;
			9417: out = 3276;
			9418: out = 3292;
			9419: out = 3312;
			9420: out = 3326;
			9421: out = 3343;
			9422: out = 3354;
			9423: out = 3371;
			9424: out = 3376;
			9425: out = 3404;
			9426: out = 3411;
			9427: out = 3426;
			9428: out = 3433;
			9429: out = 3453;
			9430: out = 3469;
			9431: out = 3488;
			9432: out = 3483;
			9433: out = 3513;
			9434: out = 3522;
			9435: out = 3528;
			9436: out = 3552;
			9437: out = 3559;
			9438: out = 3584;
			9439: out = 3581;
			9440: out = 3600;
			9441: out = 3620;
			9442: out = 3622;
			9443: out = 3638;
			9444: out = 3646;
			9445: out = 3658;
			9446: out = 3677;
			9447: out = 3687;
			9448: out = 3693;
			9449: out = 3708;
			9450: out = 3719;
			9451: out = 3736;
			9452: out = 3735;
			9453: out = 3760;
			9454: out = 3770;
			9455: out = 3769;
			9456: out = 3780;
			9457: out = 3793;
			9458: out = 3795;
			9459: out = 3812;
			9460: out = 3813;
			9461: out = 3818;
			9462: out = 3809;
			9463: out = 3788;
			9464: out = 3792;
			9465: out = 3772;
			9466: out = 3787;
			9467: out = 3773;
			9468: out = 3791;
			9469: out = 3792;
			9470: out = 3782;
			9471: out = 3803;
			9472: out = 3773;
			9473: out = 3779;
			9474: out = 3779;
			9475: out = 3794;
			9476: out = 3765;
			9477: out = 3776;
			9478: out = 3772;
			9479: out = 3783;
			9480: out = 3775;
			9481: out = 3775;
			9482: out = 3767;
			9483: out = 3777;
			9484: out = 3777;
			9485: out = 3761;
			9486: out = 3755;
			9487: out = 3762;
			9488: out = 3757;
			9489: out = 3734;
			9490: out = 3748;
			9491: out = 3738;
			9492: out = 3756;
			9493: out = 3744;
			9494: out = 3758;
			9495: out = 3742;
			9496: out = 3745;
			9497: out = 3732;
			9498: out = 3733;
			9499: out = 3747;
			9500: out = 3728;
			9501: out = 3725;
			9502: out = 3745;
			9503: out = 3725;
			9504: out = 3745;
			9505: out = 3705;
			9506: out = 3712;
			9507: out = 3721;
			9508: out = 3736;
			9509: out = 3699;
			9510: out = 3723;
			9511: out = 3719;
			9512: out = 3729;
			9513: out = 3709;
			9514: out = 3698;
			9515: out = 3706;
			9516: out = 3708;
			9517: out = 3707;
			9518: out = 3666;
			9519: out = 3695;
			9520: out = 3686;
			9521: out = 3688;
			9522: out = 3664;
			9523: out = 3667;
			9524: out = 3665;
			9525: out = 3654;
			9526: out = 3674;
			9527: out = 3667;
			9528: out = 3675;
			9529: out = 3641;
			9530: out = 3648;
			9531: out = 3610;
			9532: out = 3607;
			9533: out = 3620;
			9534: out = 3599;
			9535: out = 3579;
			9536: out = 3569;
			9537: out = 3577;
			9538: out = 3544;
			9539: out = 3559;
			9540: out = 3529;
			9541: out = 3521;
			9542: out = 3516;
			9543: out = 3491;
			9544: out = 3495;
			9545: out = 3471;
			9546: out = 3464;
			9547: out = 3461;
			9548: out = 3442;
			9549: out = 3413;
			9550: out = 3395;
			9551: out = 3364;
			9552: out = 3347;
			9553: out = 3333;
			9554: out = 3316;
			9555: out = 3292;
			9556: out = 3274;
			9557: out = 3263;
			9558: out = 3240;
			9559: out = 3225;
			9560: out = 3201;
			9561: out = 3190;
			9562: out = 3160;
			9563: out = 3145;
			9564: out = 3117;
			9565: out = 3078;
			9566: out = 3071;
			9567: out = 3054;
			9568: out = 3032;
			9569: out = 3000;
			9570: out = 2983;
			9571: out = 2954;
			9572: out = 2929;
			9573: out = 2900;
			9574: out = 2869;
			9575: out = 2861;
			9576: out = 2823;
			9577: out = 2806;
			9578: out = 2784;
			9579: out = 2758;
			9580: out = 2751;
			9581: out = 2704;
			9582: out = 2689;
			9583: out = 2654;
			9584: out = 2649;
			9585: out = 2607;
			9586: out = 2588;
			9587: out = 2559;
			9588: out = 2539;
			9589: out = 2501;
			9590: out = 2481;
			9591: out = 2471;
			9592: out = 2446;
			9593: out = 2408;
			9594: out = 2397;
			9595: out = 2360;
			9596: out = 2350;
			9597: out = 2321;
			9598: out = 2297;
			9599: out = 2279;
			9600: out = 2262;
			9601: out = 2214;
			9602: out = 2195;
			9603: out = 2186;
			9604: out = 2137;
			9605: out = 2124;
			9606: out = 2102;
			9607: out = 2081;
			9608: out = 2051;
			9609: out = 2050;
			9610: out = 1991;
			9611: out = 1994;
			9612: out = 1967;
			9613: out = 1944;
			9614: out = 1931;
			9615: out = 1886;
			9616: out = 1879;
			9617: out = 1842;
			9618: out = 1839;
			9619: out = 1807;
			9620: out = 1792;
			9621: out = 1755;
			9622: out = 1757;
			9623: out = 1720;
			9624: out = 1697;
			9625: out = 1685;
			9626: out = 1677;
			9627: out = 1643;
			9628: out = 1607;
			9629: out = 1602;
			9630: out = 1572;
			9631: out = 1557;
			9632: out = 1549;
			9633: out = 1520;
			9634: out = 1510;
			9635: out = 1484;
			9636: out = 1465;
			9637: out = 1462;
			9638: out = 1433;
			9639: out = 1404;
			9640: out = 1402;
			9641: out = 1379;
			9642: out = 1363;
			9643: out = 1351;
			9644: out = 1312;
			9645: out = 1310;
			9646: out = 1300;
			9647: out = 1284;
			9648: out = 1256;
			9649: out = 1255;
			9650: out = 1240;
			9651: out = 1214;
			9652: out = 1210;
			9653: out = 1186;
			9654: out = 1180;
			9655: out = 1155;
			9656: out = 1135;
			9657: out = 1131;
			9658: out = 1097;
			9659: out = 1097;
			9660: out = 1086;
			9661: out = 1066;
			9662: out = 1049;
			9663: out = 1026;
			9664: out = 1035;
			9665: out = 1008;
			9666: out = 988;
			9667: out = 993;
			9668: out = 974;
			9669: out = 947;
			9670: out = 938;
			9671: out = 933;
			9672: out = 916;
			9673: out = 889;
			9674: out = 891;
			9675: out = 870;
			9676: out = 862;
			9677: out = 846;
			9678: out = 849;
			9679: out = 827;
			9680: out = 817;
			9681: out = 805;
			9682: out = 780;
			9683: out = 779;
			9684: out = 778;
			9685: out = 738;
			9686: out = 739;
			9687: out = 734;
			9688: out = 715;
			9689: out = 711;
			9690: out = 697;
			9691: out = 667;
			9692: out = 646;
			9693: out = 612;
			9694: out = 580;
			9695: out = 559;
			9696: out = 519;
			9697: out = 492;
			9698: out = 469;
			9699: out = 435;
			9700: out = 409;
			9701: out = 386;
			9702: out = 364;
			9703: out = 332;
			9704: out = 318;
			9705: out = 287;
			9706: out = 264;
			9707: out = 226;
			9708: out = 222;
			9709: out = 182;
			9710: out = 161;
			9711: out = 137;
			9712: out = 121;
			9713: out = 91;
			9714: out = 64;
			9715: out = 44;
			9716: out = 16;
			9717: out = 6;
			9718: out = -19;
			9719: out = -42;
			9720: out = -62;
			9721: out = -88;
			9722: out = -112;
			9723: out = -127;
			9724: out = -137;
			9725: out = -178;
			9726: out = -191;
			9727: out = -211;
			9728: out = -237;
			9729: out = -253;
			9730: out = -259;
			9731: out = -288;
			9732: out = -301;
			9733: out = -330;
			9734: out = -347;
			9735: out = -356;
			9736: out = -384;
			9737: out = -401;
			9738: out = -425;
			9739: out = -435;
			9740: out = -456;
			9741: out = -466;
			9742: out = -491;
			9743: out = -502;
			9744: out = -522;
			9745: out = -542;
			9746: out = -554;
			9747: out = -576;
			9748: out = -592;
			9749: out = -617;
			9750: out = -629;
			9751: out = -643;
			9752: out = -664;
			9753: out = -676;
			9754: out = -688;
			9755: out = -723;
			9756: out = -722;
			9757: out = -754;
			9758: out = -759;
			9759: out = -782;
			9760: out = -793;
			9761: out = -820;
			9762: out = -834;
			9763: out = -859;
			9764: out = -859;
			9765: out = -882;
			9766: out = -907;
			9767: out = -920;
			9768: out = -938;
			9769: out = -952;
			9770: out = -962;
			9771: out = -987;
			9772: out = -1018;
			9773: out = -1023;
			9774: out = -1049;
			9775: out = -1070;
			9776: out = -1085;
			9777: out = -1099;
			9778: out = -1121;
			9779: out = -1144;
			9780: out = -1166;
			9781: out = -1182;
			9782: out = -1197;
			9783: out = -1225;
			9784: out = -1234;
			9785: out = -1248;
			9786: out = -1292;
			9787: out = -1295;
			9788: out = -1338;
			9789: out = -1358;
			9790: out = -1392;
			9791: out = -1404;
			9792: out = -1425;
			9793: out = -1466;
			9794: out = -1472;
			9795: out = -1497;
			9796: out = -1525;
			9797: out = -1558;
			9798: out = -1579;
			9799: out = -1610;
			9800: out = -1637;
			9801: out = -1662;
			9802: out = -1694;
			9803: out = -1717;
			9804: out = -1748;
			9805: out = -1779;
			9806: out = -1804;
			9807: out = -1829;
			9808: out = -1872;
			9809: out = -1896;
			9810: out = -1924;
			9811: out = -1960;
			9812: out = -1992;
			9813: out = -2025;
			9814: out = -2057;
			9815: out = -2088;
			9816: out = -2110;
			9817: out = -2171;
			9818: out = -2180;
			9819: out = -2226;
			9820: out = -2258;
			9821: out = -2287;
			9822: out = -2324;
			9823: out = -2353;
			9824: out = -2400;
			9825: out = -2431;
			9826: out = -2468;
			9827: out = -2494;
			9828: out = -2541;
			9829: out = -2555;
			9830: out = -2601;
			9831: out = -2631;
			9832: out = -2658;
			9833: out = -2699;
			9834: out = -2725;
			9835: out = -2758;
			9836: out = -2790;
			9837: out = -2826;
			9838: out = -2854;
			9839: out = -2877;
			9840: out = -2907;
			9841: out = -2942;
			9842: out = -2955;
			9843: out = -2998;
			9844: out = -3016;
			9845: out = -3043;
			9846: out = -3077;
			9847: out = -3097;
			9848: out = -3123;
			9849: out = -3148;
			9850: out = -3165;
			9851: out = -3198;
			9852: out = -3213;
			9853: out = -3236;
			9854: out = -3263;
			9855: out = -3276;
			9856: out = -3298;
			9857: out = -3331;
			9858: out = -3333;
			9859: out = -3358;
			9860: out = -3371;
			9861: out = -3395;
			9862: out = -3421;
			9863: out = -3416;
			9864: out = -3448;
			9865: out = -3470;
			9866: out = -3471;
			9867: out = -3489;
			9868: out = -3495;
			9869: out = -3507;
			9870: out = -3537;
			9871: out = -3536;
			9872: out = -3559;
			9873: out = -3574;
			9874: out = -3587;
			9875: out = -3587;
			9876: out = -3611;
			9877: out = -3606;
			9878: out = -3628;
			9879: out = -3630;
			9880: out = -3640;
			9881: out = -3655;
			9882: out = -3657;
			9883: out = -3665;
			9884: out = -3681;
			9885: out = -3677;
			9886: out = -3695;
			9887: out = -3697;
			9888: out = -3698;
			9889: out = -3706;
			9890: out = -3708;
			9891: out = -3722;
			9892: out = -3719;
			9893: out = -3730;
			9894: out = -3724;
			9895: out = -3732;
			9896: out = -3734;
			9897: out = -3740;
			9898: out = -3741;
			9899: out = -3736;
			9900: out = -3736;
			9901: out = -3747;
			9902: out = -3746;
			9903: out = -3748;
			9904: out = -3747;
			9905: out = -3754;
			9906: out = -3753;
			9907: out = -3742;
			9908: out = -3746;
			9909: out = -3752;
			9910: out = -3747;
			9911: out = -3748;
			9912: out = -3741;
			9913: out = -3749;
			9914: out = -3755;
			9915: out = -3744;
			9916: out = -3746;
			9917: out = -3737;
			9918: out = -3733;
			9919: out = -3744;
			9920: out = -3731;
			9921: out = -3728;
			9922: out = -3735;
			9923: out = -3722;
			9924: out = -3720;
			9925: out = -3711;
			9926: out = -3725;
			9927: out = -3711;
			9928: out = -3707;
			9929: out = -3702;
			9930: out = -3696;
			9931: out = -3690;
			9932: out = -3697;
			9933: out = -3674;
			9934: out = -3686;
			9935: out = -3669;
			9936: out = -3666;
			9937: out = -3671;
			9938: out = -3654;
			9939: out = -3650;
			9940: out = -3652;
			9941: out = -3637;
			9942: out = -3635;
			9943: out = -3623;
			9944: out = -3636;
			9945: out = -3615;
			9946: out = -3606;
			9947: out = -3601;
			9948: out = -3588;
			9949: out = -3599;
			9950: out = -3578;
			9951: out = -3570;
			9952: out = -3568;
			9953: out = -3557;
			9954: out = -3549;
			9955: out = -3540;
			9956: out = -3544;
			9957: out = -3528;
			9958: out = -3517;
			9959: out = -3520;
			9960: out = -3501;
			9961: out = -3500;
			9962: out = -3495;
			9963: out = -3482;
			9964: out = -3477;
			9965: out = -3465;
			9966: out = -3463;
			9967: out = -3433;
			9968: out = -3435;
			9969: out = -3435;
			9970: out = -3413;
			9971: out = -3403;
			9972: out = -3397;
			9973: out = -3394;
			9974: out = -3374;
			9975: out = -3375;
			9976: out = -3352;
			9977: out = -3350;
			9978: out = -3333;
			9979: out = -3331;
			9980: out = -3308;
			9981: out = -3312;
			9982: out = -3288;
			9983: out = -3274;
			9984: out = -3278;
			9985: out = -3247;
			9986: out = -3255;
			9987: out = -3225;
			9988: out = -3223;
			9989: out = -3197;
			9990: out = -3199;
			9991: out = -3187;
			9992: out = -3160;
			9993: out = -3153;
			9994: out = -3132;
			9995: out = -3122;
			9996: out = -3096;
			9997: out = -3094;
			9998: out = -3061;
			9999: out = -3059;
			10000: out = -3030;
			10001: out = -3025;
			10002: out = -3000;
			10003: out = -2988;
			10004: out = -2969;
			10005: out = -2950;
			10006: out = -2921;
			10007: out = -2906;
			10008: out = -2882;
			10009: out = -2864;
			10010: out = -2843;
			10011: out = -2822;
			10012: out = -2795;
			10013: out = -2783;
			10014: out = -2751;
			10015: out = -2730;
			10016: out = -2710;
			10017: out = -2668;
			10018: out = -2668;
			10019: out = -2631;
			10020: out = -2606;
			10021: out = -2577;
			10022: out = -2560;
			10023: out = -2528;
			10024: out = -2507;
			10025: out = -2474;
			10026: out = -2457;
			10027: out = -2434;
			10028: out = -2386;
			10029: out = -2379;
			10030: out = -2355;
			10031: out = -2317;
			10032: out = -2294;
			10033: out = -2271;
			10034: out = -2238;
			10035: out = -2219;
			10036: out = -2193;
			10037: out = -2166;
			10038: out = -2131;
			10039: out = -2121;
			10040: out = -2085;
			10041: out = -2055;
			10042: out = -2040;
			10043: out = -2003;
			10044: out = -1986;
			10045: out = -1965;
			10046: out = -1922;
			10047: out = -1901;
			10048: out = -1874;
			10049: out = -1858;
			10050: out = -1831;
			10051: out = -1809;
			10052: out = -1789;
			10053: out = -1753;
			10054: out = -1740;
			10055: out = -1712;
			10056: out = -1690;
			10057: out = -1674;
			10058: out = -1639;
			10059: out = -1618;
			10060: out = -1604;
			10061: out = -1571;
			10062: out = -1549;
			10063: out = -1534;
			10064: out = -1505;
			10065: out = -1487;
			10066: out = -1465;
			10067: out = -1446;
			10068: out = -1416;
			10069: out = -1409;
			10070: out = -1369;
			10071: out = -1363;
			10072: out = -1344;
			10073: out = -1319;
			10074: out = -1294;
			10075: out = -1268;
			10076: out = -1270;
			10077: out = -1237;
			10078: out = -1219;
			10079: out = -1199;
			10080: out = -1188;
			10081: out = -1163;
			10082: out = -1151;
			10083: out = -1123;
			10084: out = -1107;
			10085: out = -1096;
			10086: out = -1068;
			10087: out = -1059;
			10088: out = -1038;
			10089: out = -1027;
			10090: out = -1006;
			10091: out = -991;
			10092: out = -968;
			10093: out = -954;
			10094: out = -942;
			10095: out = -918;
			10096: out = -917;
			10097: out = -883;
			10098: out = -889;
			10099: out = -860;
			10100: out = -854;
			10101: out = -827;
			10102: out = -822;
			10103: out = -808;
			10104: out = -789;
			10105: out = -775;
			10106: out = -764;
			10107: out = -759;
			10108: out = -735;
			10109: out = -713;
			10110: out = -705;
			10111: out = -706;
			10112: out = -682;
			10113: out = -672;
			10114: out = -654;
			10115: out = -642;
			10116: out = -608;
			10117: out = -601;
			10118: out = -570;
			10119: out = -540;
			10120: out = -531;
			10121: out = -503;
			10122: out = -490;
			10123: out = -459;
			10124: out = -457;
			10125: out = -423;
			10126: out = -411;
			10127: out = -383;
			10128: out = -373;
			10129: out = -349;
			10130: out = -338;
			10131: out = -302;
			10132: out = -303;
			10133: out = -286;
			10134: out = -262;
			10135: out = -240;
			10136: out = -233;
			10137: out = -211;
			10138: out = -192;
			10139: out = -188;
			10140: out = -166;
			10141: out = -135;
			10142: out = -146;
			10143: out = -110;
			10144: out = -104;
			10145: out = -80;
			10146: out = -76;
			10147: out = -60;
			10148: out = -57;
			10149: out = -26;
			10150: out = -14;
			10151: out = 1;
			10152: out = 18;
			10153: out = 20;
			10154: out = 38;
			10155: out = 57;
			10156: out = 72;
			10157: out = 83;
			10158: out = 87;
			10159: out = 112;
			10160: out = 124;
			10161: out = 136;
			10162: out = 141;
			10163: out = 166;
			10164: out = 168;
			10165: out = 185;
			10166: out = 199;
			10167: out = 209;
			10168: out = 217;
			10169: out = 244;
			10170: out = 239;
			10171: out = 263;
			10172: out = 267;
			10173: out = 286;
			10174: out = 301;
			10175: out = 303;
			10176: out = 321;
			10177: out = 336;
			10178: out = 349;
			10179: out = 357;
			10180: out = 371;
			10181: out = 386;
			10182: out = 391;
			10183: out = 406;
			10184: out = 416;
			10185: out = 442;
			10186: out = 432;
			10187: out = 459;
			10188: out = 470;
			10189: out = 480;
			10190: out = 500;
			10191: out = 511;
			10192: out = 531;
			10193: out = 530;
			10194: out = 551;
			10195: out = 560;
			10196: out = 577;
			10197: out = 592;
			10198: out = 594;
			10199: out = 617;
			10200: out = 640;
			10201: out = 641;
			10202: out = 664;
			10203: out = 678;
			10204: out = 692;
			10205: out = 700;
			10206: out = 724;
			10207: out = 738;
			10208: out = 747;
			10209: out = 778;
			10210: out = 775;
			10211: out = 807;
			10212: out = 824;
			10213: out = 839;
			10214: out = 865;
			10215: out = 864;
			10216: out = 904;
			10217: out = 910;
			10218: out = 932;
			10219: out = 945;
			10220: out = 986;
			10221: out = 981;
			10222: out = 1012;
			10223: out = 1037;
			10224: out = 1057;
			10225: out = 1075;
			10226: out = 1098;
			10227: out = 1129;
			10228: out = 1132;
			10229: out = 1174;
			10230: out = 1187;
			10231: out = 1206;
			10232: out = 1241;
			10233: out = 1258;
			10234: out = 1292;
			10235: out = 1300;
			10236: out = 1327;
			10237: out = 1345;
			10238: out = 1386;
			10239: out = 1395;
			10240: out = 1426;
			10241: out = 1444;
			10242: out = 1469;
			10243: out = 1492;
			10244: out = 1503;
			10245: out = 1537;
			10246: out = 1559;
			10247: out = 1581;
			10248: out = 1608;
			10249: out = 1628;
			10250: out = 1664;
			10251: out = 1667;
			10252: out = 1696;
			10253: out = 1720;
			10254: out = 1748;
			10255: out = 1759;
			10256: out = 1794;
			10257: out = 1807;
			10258: out = 1838;
			10259: out = 1844;
			10260: out = 1871;
			10261: out = 1900;
			10262: out = 1915;
			10263: out = 1933;
			10264: out = 1954;
			10265: out = 1984;
			10266: out = 1982;
			10267: out = 2024;
			10268: out = 2030;
			10269: out = 2053;
			10270: out = 2077;
			10271: out = 2084;
			10272: out = 2102;
			10273: out = 2133;
			10274: out = 2150;
			10275: out = 2171;
			10276: out = 2175;
			10277: out = 2203;
			10278: out = 2223;
			10279: out = 2223;
			10280: out = 2257;
			10281: out = 2261;
			10282: out = 2287;
			10283: out = 2300;
			10284: out = 2315;
			10285: out = 2344;
			10286: out = 2349;
			10287: out = 2365;
			10288: out = 2386;
			10289: out = 2400;
			10290: out = 2410;
			10291: out = 2431;
			10292: out = 2446;
			10293: out = 2453;
			10294: out = 2469;
			10295: out = 2481;
			10296: out = 2502;
			10297: out = 2514;
			10298: out = 2539;
			10299: out = 2542;
			10300: out = 2554;
			10301: out = 2569;
			10302: out = 2587;
			10303: out = 2595;
			10304: out = 2614;
			10305: out = 2618;
			10306: out = 2636;
			10307: out = 2658;
			10308: out = 2646;
			10309: out = 2679;
			10310: out = 2689;
			10311: out = 2706;
			10312: out = 2710;
			10313: out = 2720;
			10314: out = 2740;
			10315: out = 2753;
			10316: out = 2750;
			10317: out = 2765;
			10318: out = 2778;
			10319: out = 2785;
			10320: out = 2815;
			10321: out = 2812;
			10322: out = 2832;
			10323: out = 2842;
			10324: out = 2846;
			10325: out = 2877;
			10326: out = 2858;
			10327: out = 2888;
			10328: out = 2892;
			10329: out = 2905;
			10330: out = 2917;
			10331: out = 2919;
			10332: out = 2936;
			10333: out = 2943;
			10334: out = 2953;
			10335: out = 2959;
			10336: out = 2983;
			10337: out = 2979;
			10338: out = 3003;
			10339: out = 3002;
			10340: out = 3009;
			10341: out = 3027;
			10342: out = 3030;
			10343: out = 3049;
			10344: out = 3047;
			10345: out = 3059;
			10346: out = 3062;
			10347: out = 3082;
			10348: out = 3075;
			10349: out = 3090;
			10350: out = 3085;
			10351: out = 3094;
			10352: out = 3095;
			10353: out = 3094;
			10354: out = 3082;
			10355: out = 3073;
			10356: out = 3069;
			10357: out = 3073;
			10358: out = 3074;
			10359: out = 3075;
			10360: out = 3079;
			10361: out = 3072;
			10362: out = 3068;
			10363: out = 3069;
			10364: out = 3054;
			10365: out = 3067;
			10366: out = 3085;
			10367: out = 3063;
			10368: out = 3052;
			10369: out = 3045;
			10370: out = 3031;
			10371: out = 3049;
			10372: out = 3047;
			10373: out = 3038;
			10374: out = 3043;
			10375: out = 3051;
			10376: out = 3038;
			10377: out = 3063;
			10378: out = 3047;
			10379: out = 3049;
			10380: out = 3050;
			10381: out = 3056;
			10382: out = 3057;
			10383: out = 3047;
			10384: out = 3054;
			10385: out = 3048;
			10386: out = 3028;
			10387: out = 3046;
			10388: out = 3044;
			10389: out = 3044;
			10390: out = 3046;
			10391: out = 3031;
			10392: out = 3052;
			10393: out = 3049;
			10394: out = 3047;
			10395: out = 3050;
			10396: out = 3052;
			10397: out = 3021;
			10398: out = 3019;
			10399: out = 3037;
			10400: out = 3013;
			10401: out = 3018;
			10402: out = 3038;
			10403: out = 3007;
			10404: out = 3038;
			10405: out = 3014;
			10406: out = 3014;
			10407: out = 3025;
			10408: out = 3004;
			10409: out = 3014;
			10410: out = 3014;
			10411: out = 3010;
			10412: out = 3026;
			10413: out = 3016;
			10414: out = 2996;
			10415: out = 3006;
			10416: out = 2972;
			10417: out = 2987;
			10418: out = 2983;
			10419: out = 2965;
			10420: out = 2951;
			10421: out = 2966;
			10422: out = 2941;
			10423: out = 2959;
			10424: out = 2938;
			10425: out = 2950;
			10426: out = 2929;
			10427: out = 2941;
			10428: out = 2923;
			10429: out = 2920;
			10430: out = 2900;
			10431: out = 2903;
			10432: out = 2867;
			10433: out = 2858;
			10434: out = 2850;
			10435: out = 2847;
			10436: out = 2823;
			10437: out = 2831;
			10438: out = 2785;
			10439: out = 2803;
			10440: out = 2763;
			10441: out = 2750;
			10442: out = 2751;
			10443: out = 2729;
			10444: out = 2715;
			10445: out = 2715;
			10446: out = 2697;
			10447: out = 2666;
			10448: out = 2660;
			10449: out = 2634;
			10450: out = 2612;
			10451: out = 2600;
			10452: out = 2581;
			10453: out = 2564;
			10454: out = 2557;
			10455: out = 2531;
			10456: out = 2516;
			10457: out = 2489;
			10458: out = 2481;
			10459: out = 2456;
			10460: out = 2430;
			10461: out = 2431;
			10462: out = 2386;
			10463: out = 2383;
			10464: out = 2350;
			10465: out = 2338;
			10466: out = 2312;
			10467: out = 2310;
			10468: out = 2264;
			10469: out = 2254;
			10470: out = 2238;
			10471: out = 2218;
			10472: out = 2198;
			10473: out = 2170;
			10474: out = 2166;
			10475: out = 2142;
			10476: out = 2119;
			10477: out = 2097;
			10478: out = 2080;
			10479: out = 2043;
			10480: out = 2034;
			10481: out = 2016;
			10482: out = 2004;
			10483: out = 1971;
			10484: out = 1960;
			10485: out = 1942;
			10486: out = 1896;
			10487: out = 1896;
			10488: out = 1883;
			10489: out = 1848;
			10490: out = 1833;
			10491: out = 1812;
			10492: out = 1802;
			10493: out = 1774;
			10494: out = 1757;
			10495: out = 1737;
			10496: out = 1722;
			10497: out = 1702;
			10498: out = 1682;
			10499: out = 1660;
			10500: out = 1639;
			10501: out = 1617;
			10502: out = 1610;
			10503: out = 1603;
			10504: out = 1577;
			10505: out = 1558;
			10506: out = 1542;
			10507: out = 1524;
			10508: out = 1493;
			10509: out = 1494;
			10510: out = 1448;
			10511: out = 1448;
			10512: out = 1433;
			10513: out = 1410;
			10514: out = 1403;
			10515: out = 1379;
			10516: out = 1361;
			10517: out = 1348;
			10518: out = 1341;
			10519: out = 1320;
			10520: out = 1294;
			10521: out = 1280;
			10522: out = 1269;
			10523: out = 1258;
			10524: out = 1250;
			10525: out = 1214;
			10526: out = 1206;
			10527: out = 1204;
			10528: out = 1158;
			10529: out = 1168;
			10530: out = 1153;
			10531: out = 1118;
			10532: out = 1115;
			10533: out = 1117;
			10534: out = 1094;
			10535: out = 1081;
			10536: out = 1058;
			10537: out = 1055;
			10538: out = 1027;
			10539: out = 1022;
			10540: out = 1010;
			10541: out = 996;
			10542: out = 983;
			10543: out = 966;
			10544: out = 955;
			10545: out = 953;
			10546: out = 931;
			10547: out = 914;
			10548: out = 904;
			10549: out = 906;
			10550: out = 871;
			10551: out = 867;
			10552: out = 868;
			10553: out = 836;
			10554: out = 834;
			10555: out = 818;
			10556: out = 820;
			10557: out = 790;
			10558: out = 798;
			10559: out = 767;
			10560: out = 771;
			10561: out = 764;
			10562: out = 729;
			10563: out = 738;
			10564: out = 736;
			10565: out = 706;
			10566: out = 707;
			10567: out = 681;
			10568: out = 689;
			10569: out = 669;
			10570: out = 658;
			10571: out = 654;
			10572: out = 642;
			10573: out = 634;
			10574: out = 623;
			10575: out = 624;
			10576: out = 600;
			10577: out = 601;
			10578: out = 577;
			10579: out = 577;
			10580: out = 567;
			10581: out = 553;
			10582: out = 525;
			10583: out = 511;
			10584: out = 480;
			10585: out = 456;
			10586: out = 432;
			10587: out = 412;
			10588: out = 385;
			10589: out = 357;
			10590: out = 345;
			10591: out = 320;
			10592: out = 290;
			10593: out = 280;
			10594: out = 261;
			10595: out = 216;
			10596: out = 220;
			10597: out = 184;
			10598: out = 171;
			10599: out = 148;
			10600: out = 128;
			10601: out = 108;
			10602: out = 84;
			10603: out = 77;
			10604: out = 42;
			10605: out = 17;
			10606: out = 6;
			10607: out = -1;
			10608: out = -43;
			10609: out = -39;
			10610: out = -68;
			10611: out = -78;
			10612: out = -100;
			10613: out = -111;
			10614: out = -122;
			10615: out = -146;
			10616: out = -161;
			10617: out = -171;
			10618: out = -202;
			10619: out = -219;
			10620: out = -227;
			10621: out = -240;
			10622: out = -251;
			10623: out = -274;
			10624: out = -280;
			10625: out = -309;
			10626: out = -304;
			10627: out = -335;
			10628: out = -339;
			10629: out = -357;
			10630: out = -379;
			10631: out = -383;
			10632: out = -399;
			10633: out = -422;
			10634: out = -424;
			10635: out = -448;
			10636: out = -448;
			10637: out = -481;
			10638: out = -480;
			10639: out = -498;
			10640: out = -519;
			10641: out = -525;
			10642: out = -541;
			10643: out = -552;
			10644: out = -578;
			10645: out = -592;
			10646: out = -600;
			10647: out = -623;
			10648: out = -626;
			10649: out = -641;
			10650: out = -660;
			10651: out = -670;
			10652: out = -692;
			10653: out = -692;
			10654: out = -716;
			10655: out = -727;
			10656: out = -741;
			10657: out = -756;
			10658: out = -778;
			10659: out = -779;
			10660: out = -797;
			10661: out = -817;
			10662: out = -818;
			10663: out = -845;
			10664: out = -872;
			10665: out = -853;
			10666: out = -896;
			10667: out = -904;
			10668: out = -927;
			10669: out = -933;
			10670: out = -948;
			10671: out = -968;
			10672: out = -988;
			10673: out = -999;
			10674: out = -1012;
			10675: out = -1044;
			10676: out = -1051;
			10677: out = -1067;
			10678: out = -1087;
			10679: out = -1115;
			10680: out = -1134;
			10681: out = -1135;
			10682: out = -1163;
			10683: out = -1190;
			10684: out = -1197;
			10685: out = -1227;
			10686: out = -1244;
			10687: out = -1269;
			10688: out = -1279;
			10689: out = -1308;
			10690: out = -1321;
			10691: out = -1347;
			10692: out = -1374;
			10693: out = -1397;
			10694: out = -1428;
			10695: out = -1460;
			10696: out = -1466;
			10697: out = -1509;
			10698: out = -1527;
			10699: out = -1544;
			10700: out = -1574;
			10701: out = -1604;
			10702: out = -1612;
			10703: out = -1645;
			10704: out = -1688;
			10705: out = -1702;
			10706: out = -1732;
			10707: out = -1765;
			10708: out = -1799;
			10709: out = -1809;
			10710: out = -1852;
			10711: out = -1865;
			10712: out = -1897;
			10713: out = -1935;
			10714: out = -1953;
			10715: out = -1984;
			10716: out = -2009;
			10717: out = -2048;
			10718: out = -2069;
			10719: out = -2098;
			10720: out = -2125;
			10721: out = -2149;
			10722: out = -2179;
			10723: out = -2197;
			10724: out = -2233;
			10725: out = -2247;
			10726: out = -2282;
			10727: out = -2309;
			10728: out = -2312;
			10729: out = -2368;
			10730: out = -2374;
			10731: out = -2401;
			10732: out = -2419;
			10733: out = -2445;
			10734: out = -2468;
			10735: out = -2482;
			10736: out = -2517;
			10737: out = -2533;
			10738: out = -2553;
			10739: out = -2581;
			10740: out = -2582;
			10741: out = -2621;
			10742: out = -2629;
			10743: out = -2659;
			10744: out = -2661;
			10745: out = -2695;
			10746: out = -2693;
			10747: out = -2720;
			10748: out = -2732;
			10749: out = -2750;
			10750: out = -2763;
			10751: out = -2774;
			10752: out = -2796;
			10753: out = -2798;
			10754: out = -2825;
			10755: out = -2836;
			10756: out = -2849;
			10757: out = -2861;
			10758: out = -2864;
			10759: out = -2894;
			10760: out = -2885;
			10761: out = -2904;
			10762: out = -2903;
			10763: out = -2929;
			10764: out = -2926;
			10765: out = -2943;
			10766: out = -2950;
			10767: out = -2955;
			10768: out = -2969;
			10769: out = -2968;
			10770: out = -2984;
			10771: out = -2980;
			10772: out = -3002;
			10773: out = -2994;
			10774: out = -3006;
			10775: out = -3004;
			10776: out = -3009;
			10777: out = -3034;
			10778: out = -3019;
			10779: out = -3037;
			10780: out = -3028;
			10781: out = -3051;
			10782: out = -3045;
			10783: out = -3056;
			10784: out = -3046;
			10785: out = -3057;
			10786: out = -3063;
			10787: out = -3060;
			10788: out = -3052;
			10789: out = -3074;
			10790: out = -3063;
			10791: out = -3060;
			10792: out = -3072;
			10793: out = -3075;
			10794: out = -3065;
			10795: out = -3068;
			10796: out = -3083;
			10797: out = -3061;
			10798: out = -3072;
			10799: out = -3063;
			10800: out = -3068;
			10801: out = -3075;
			10802: out = -3068;
			10803: out = -3060;
			10804: out = -3066;
			10805: out = -3065;
			10806: out = -3068;
			10807: out = -3054;
			10808: out = -3063;
			10809: out = -3061;
			10810: out = -3050;
			10811: out = -3046;
			10812: out = -3051;
			10813: out = -3043;
			10814: out = -3046;
			10815: out = -3036;
			10816: out = -3033;
			10817: out = -3047;
			10818: out = -3033;
			10819: out = -3021;
			10820: out = -3026;
			10821: out = -3013;
			10822: out = -3023;
			10823: out = -3000;
			10824: out = -3009;
			10825: out = -3008;
			10826: out = -2994;
			10827: out = -2987;
			10828: out = -2999;
			10829: out = -2980;
			10830: out = -2983;
			10831: out = -2968;
			10832: out = -2978;
			10833: out = -2959;
			10834: out = -2952;
			10835: out = -2953;
			10836: out = -2947;
			10837: out = -2939;
			10838: out = -2932;
			10839: out = -2924;
			10840: out = -2923;
			10841: out = -2921;
			10842: out = -2917;
			10843: out = -2890;
			10844: out = -2910;
			10845: out = -2892;
			10846: out = -2880;
			10847: out = -2886;
			10848: out = -2868;
			10849: out = -2864;
			10850: out = -2865;
			10851: out = -2848;
			10852: out = -2843;
			10853: out = -2844;
			10854: out = -2832;
			10855: out = -2820;
			10856: out = -2822;
			10857: out = -2805;
			10858: out = -2805;
			10859: out = -2797;
			10860: out = -2782;
			10861: out = -2785;
			10862: out = -2771;
			10863: out = -2766;
			10864: out = -2760;
			10865: out = -2746;
			10866: out = -2748;
			10867: out = -2725;
			10868: out = -2739;
			10869: out = -2716;
			10870: out = -2706;
			10871: out = -2700;
			10872: out = -2694;
			10873: out = -2669;
			10874: out = -2673;
			10875: out = -2654;
			10876: out = -2653;
			10877: out = -2635;
			10878: out = -2626;
			10879: out = -2619;
			10880: out = -2599;
			10881: out = -2600;
			10882: out = -2585;
			10883: out = -2573;
			10884: out = -2557;
			10885: out = -2545;
			10886: out = -2530;
			10887: out = -2524;
			10888: out = -2506;
			10889: out = -2498;
			10890: out = -2472;
			10891: out = -2466;
			10892: out = -2455;
			10893: out = -2440;
			10894: out = -2415;
			10895: out = -2408;
			10896: out = -2389;
			10897: out = -2367;
			10898: out = -2359;
			10899: out = -2333;
			10900: out = -2329;
			10901: out = -2306;
			10902: out = -2284;
			10903: out = -2268;
			10904: out = -2243;
			10905: out = -2234;
			10906: out = -2208;
			10907: out = -2190;
			10908: out = -2175;
			10909: out = -2152;
			10910: out = -2133;
			10911: out = -2107;
			10912: out = -2089;
			10913: out = -2076;
			10914: out = -2033;
			10915: out = -2034;
			10916: out = -2015;
			10917: out = -1982;
			10918: out = -1966;
			10919: out = -1944;
			10920: out = -1921;
			10921: out = -1900;
			10922: out = -1875;
			10923: out = -1852;
			10924: out = -1840;
			10925: out = -1814;
			10926: out = -1793;
			10927: out = -1769;
			10928: out = -1754;
			10929: out = -1724;
			10930: out = -1714;
			10931: out = -1686;
			10932: out = -1666;
			10933: out = -1642;
			10934: out = -1627;
			10935: out = -1606;
			10936: out = -1575;
			10937: out = -1570;
			10938: out = -1540;
			10939: out = -1521;
			10940: out = -1507;
			10941: out = -1487;
			10942: out = -1457;
			10943: out = -1448;
			10944: out = -1422;
			10945: out = -1401;
			10946: out = -1391;
			10947: out = -1371;
			10948: out = -1350;
			10949: out = -1317;
			10950: out = -1328;
			10951: out = -1296;
			10952: out = -1264;
			10953: out = -1256;
			10954: out = -1234;
			10955: out = -1228;
			10956: out = -1194;
			10957: out = -1189;
			10958: out = -1169;
			10959: out = -1150;
			10960: out = -1146;
			10961: out = -1115;
			10962: out = -1099;
			10963: out = -1094;
			10964: out = -1067;
			10965: out = -1055;
			10966: out = -1039;
			10967: out = -1021;
			10968: out = -1013;
			10969: out = -995;
			10970: out = -974;
			10971: out = -964;
			10972: out = -943;
			10973: out = -928;
			10974: out = -920;
			10975: out = -898;
			10976: out = -892;
			10977: out = -881;
			10978: out = -860;
			10979: out = -845;
			10980: out = -839;
			10981: out = -819;
			10982: out = -810;
			10983: out = -788;
			10984: out = -780;
			10985: out = -772;
			10986: out = -754;
			10987: out = -738;
			10988: out = -734;
			10989: out = -709;
			10990: out = -705;
			10991: out = -706;
			10992: out = -673;
			10993: out = -678;
			10994: out = -658;
			10995: out = -643;
			10996: out = -640;
			10997: out = -619;
			10998: out = -618;
			10999: out = -599;
			11000: out = -589;
			11001: out = -587;
			11002: out = -569;
			11003: out = -562;
			11004: out = -552;
			11005: out = -536;
			11006: out = -521;
			11007: out = -498;
			11008: out = -478;
			11009: out = -466;
			11010: out = -452;
			11011: out = -427;
			11012: out = -408;
			11013: out = -398;
			11014: out = -386;
			11015: out = -362;
			11016: out = -353;
			11017: out = -326;
			11018: out = -327;
			11019: out = -299;
			11020: out = -277;
			11021: out = -278;
			11022: out = -264;
			11023: out = -230;
			11024: out = -230;
			11025: out = -225;
			11026: out = -194;
			11027: out = -183;
			11028: out = -181;
			11029: out = -157;
			11030: out = -143;
			11031: out = -147;
			11032: out = -110;
			11033: out = -111;
			11034: out = -101;
			11035: out = -84;
			11036: out = -79;
			11037: out = -58;
			11038: out = -44;
			11039: out = -44;
			11040: out = -26;
			11041: out = -16;
			11042: out = 6;
			11043: out = 4;
			11044: out = 12;
			11045: out = 37;
			11046: out = 46;
			11047: out = 51;
			11048: out = 56;
			11049: out = 78;
			11050: out = 72;
			11051: out = 112;
			11052: out = 83;
			11053: out = 114;
			11054: out = 117;
			11055: out = 144;
			11056: out = 140;
			11057: out = 148;
			11058: out = 169;
			11059: out = 182;
			11060: out = 188;
			11061: out = 194;
			11062: out = 209;
			11063: out = 220;
			11064: out = 222;
			11065: out = 241;
			11066: out = 240;
			11067: out = 259;
			11068: out = 268;
			11069: out = 274;
			11070: out = 291;
			11071: out = 294;
			11072: out = 309;
			11073: out = 318;
			11074: out = 330;
			11075: out = 342;
			11076: out = 346;
			11077: out = 360;
			11078: out = 359;
			11079: out = 380;
			11080: out = 388;
			11081: out = 398;
			11082: out = 403;
			11083: out = 417;
			11084: out = 436;
			11085: out = 438;
			11086: out = 453;
			11087: out = 459;
			11088: out = 475;
			11089: out = 482;
			11090: out = 496;
			11091: out = 510;
			11092: out = 518;
			11093: out = 537;
			11094: out = 545;
			11095: out = 553;
			11096: out = 566;
			11097: out = 589;
			11098: out = 594;
			11099: out = 610;
			11100: out = 626;
			11101: out = 636;
			11102: out = 657;
			11103: out = 661;
			11104: out = 682;
			11105: out = 689;
			11106: out = 718;
			11107: out = 722;
			11108: out = 744;
			11109: out = 755;
			11110: out = 778;
			11111: out = 789;
			11112: out = 802;
			11113: out = 827;
			11114: out = 838;
			11115: out = 856;
			11116: out = 888;
			11117: out = 895;
			11118: out = 925;
			11119: out = 931;
			11120: out = 948;
			11121: out = 976;
			11122: out = 995;
			11123: out = 993;
			11124: out = 1038;
			11125: out = 1037;
			11126: out = 1073;
			11127: out = 1082;
			11128: out = 1101;
			11129: out = 1122;
			11130: out = 1137;
			11131: out = 1169;
			11132: out = 1182;
			11133: out = 1201;
			11134: out = 1220;
			11135: out = 1244;
			11136: out = 1251;
			11137: out = 1283;
			11138: out = 1303;
			11139: out = 1304;
			11140: out = 1344;
			11141: out = 1353;
			11142: out = 1378;
			11143: out = 1387;
			11144: out = 1401;
			11145: out = 1432;
			11146: out = 1435;
			11147: out = 1457;
			11148: out = 1476;
			11149: out = 1497;
			11150: out = 1515;
			11151: out = 1534;
			11152: out = 1542;
			11153: out = 1566;
			11154: out = 1577;
			11155: out = 1586;
			11156: out = 1611;
			11157: out = 1638;
			11158: out = 1646;
			11159: out = 1662;
			11160: out = 1675;
			11161: out = 1695;
			11162: out = 1712;
			11163: out = 1709;
			11164: out = 1738;
			11165: out = 1747;
			11166: out = 1767;
			11167: out = 1780;
			11168: out = 1802;
			11169: out = 1797;
			11170: out = 1832;
			11171: out = 1837;
			11172: out = 1844;
			11173: out = 1873;
			11174: out = 1875;
			11175: out = 1868;
			11176: out = 1915;
			11177: out = 1914;
			11178: out = 1934;
			11179: out = 1937;
			11180: out = 1955;
			11181: out = 1963;
			11182: out = 1975;
			11183: out = 1996;
			11184: out = 1991;
			11185: out = 2024;
			11186: out = 2014;
			11187: out = 2042;
			11188: out = 2041;
			11189: out = 2058;
			11190: out = 2079;
			11191: out = 2075;
			11192: out = 2089;
			11193: out = 2107;
			11194: out = 2110;
			11195: out = 2134;
			11196: out = 2124;
			11197: out = 2146;
			11198: out = 2156;
			11199: out = 2169;
			11200: out = 2172;
			11201: out = 2193;
			11202: out = 2203;
			11203: out = 2205;
			11204: out = 2216;
			11205: out = 2227;
			11206: out = 2233;
			11207: out = 2244;
			11208: out = 2254;
			11209: out = 2268;
			11210: out = 2271;
			11211: out = 2281;
			11212: out = 2301;
			11213: out = 2302;
			11214: out = 2306;
			11215: out = 2323;
			11216: out = 2333;
			11217: out = 2332;
			11218: out = 2349;
			11219: out = 2353;
			11220: out = 2363;
			11221: out = 2368;
			11222: out = 2383;
			11223: out = 2387;
			11224: out = 2401;
			11225: out = 2404;
			11226: out = 2412;
			11227: out = 2427;
			11228: out = 2420;
			11229: out = 2441;
			11230: out = 2440;
			11231: out = 2448;
			11232: out = 2452;
			11233: out = 2471;
			11234: out = 2467;
			11235: out = 2480;
			11236: out = 2487;
			11237: out = 2488;
			11238: out = 2492;
			11239: out = 2498;
			11240: out = 2492;
			11241: out = 2506;
			11242: out = 2501;
			11243: out = 2495;
			11244: out = 2507;
			11245: out = 2499;
			11246: out = 2497;
			11247: out = 2506;
			11248: out = 2483;
			11249: out = 2495;
			11250: out = 2482;
			11251: out = 2484;
			11252: out = 2491;
			11253: out = 2491;
			11254: out = 2488;
			11255: out = 2490;
			11256: out = 2490;
			11257: out = 2497;
			11258: out = 2491;
			11259: out = 2491;
			11260: out = 2494;
			11261: out = 2478;
			11262: out = 2490;
			11263: out = 2464;
			11264: out = 2469;
			11265: out = 2475;
			11266: out = 2486;
			11267: out = 2464;
			11268: out = 2480;
			11269: out = 2469;
			11270: out = 2478;
			11271: out = 2484;
			11272: out = 2459;
			11273: out = 2476;
			11274: out = 2474;
			11275: out = 2490;
			11276: out = 2480;
			11277: out = 2467;
			11278: out = 2482;
			11279: out = 2480;
			11280: out = 2491;
			11281: out = 2477;
			11282: out = 2483;
			11283: out = 2484;
			11284: out = 2491;
			11285: out = 2471;
			11286: out = 2477;
			11287: out = 2471;
			11288: out = 2477;
			11289: out = 2463;
			11290: out = 2462;
			11291: out = 2470;
			11292: out = 2483;
			11293: out = 2448;
			11294: out = 2455;
			11295: out = 2454;
			11296: out = 2436;
			11297: out = 2442;
			11298: out = 2454;
			11299: out = 2443;
			11300: out = 2430;
			11301: out = 2447;
			11302: out = 2424;
			11303: out = 2420;
			11304: out = 2440;
			11305: out = 2433;
			11306: out = 2415;
			11307: out = 2411;
			11308: out = 2410;
			11309: out = 2415;
			11310: out = 2410;
			11311: out = 2396;
			11312: out = 2400;
			11313: out = 2396;
			11314: out = 2385;
			11315: out = 2389;
			11316: out = 2352;
			11317: out = 2356;
			11318: out = 2344;
			11319: out = 2357;
			11320: out = 2339;
			11321: out = 2325;
			11322: out = 2330;
			11323: out = 2315;
			11324: out = 2314;
			11325: out = 2310;
			11326: out = 2292;
			11327: out = 2285;
			11328: out = 2279;
			11329: out = 2262;
			11330: out = 2240;
			11331: out = 2246;
			11332: out = 2215;
			11333: out = 2217;
			11334: out = 2200;
			11335: out = 2194;
			11336: out = 2175;
			11337: out = 2173;
			11338: out = 2147;
			11339: out = 2146;
			11340: out = 2137;
			11341: out = 2120;
			11342: out = 2108;
			11343: out = 2078;
			11344: out = 2079;
			11345: out = 2053;
			11346: out = 2040;
			11347: out = 2031;
			11348: out = 2005;
			11349: out = 1992;
			11350: out = 1980;
			11351: out = 1971;
			11352: out = 1938;
			11353: out = 1930;
			11354: out = 1924;
			11355: out = 1904;
			11356: out = 1883;
			11357: out = 1871;
			11358: out = 1851;
			11359: out = 1849;
			11360: out = 1819;
			11361: out = 1794;
			11362: out = 1795;
			11363: out = 1777;
			11364: out = 1750;
			11365: out = 1743;
			11366: out = 1718;
			11367: out = 1694;
			11368: out = 1693;
			11369: out = 1670;
			11370: out = 1669;
			11371: out = 1623;
			11372: out = 1625;
			11373: out = 1612;
			11374: out = 1586;
			11375: out = 1571;
			11376: out = 1565;
			11377: out = 1536;
			11378: out = 1537;
			11379: out = 1505;
			11380: out = 1492;
			11381: out = 1482;
			11382: out = 1471;
			11383: out = 1437;
			11384: out = 1422;
			11385: out = 1426;
			11386: out = 1389;
			11387: out = 1385;
			11388: out = 1369;
			11389: out = 1352;
			11390: out = 1346;
			11391: out = 1320;
			11392: out = 1311;
			11393: out = 1297;
			11394: out = 1279;
			11395: out = 1262;
			11396: out = 1248;
			11397: out = 1237;
			11398: out = 1236;
			11399: out = 1211;
			11400: out = 1193;
			11401: out = 1196;
			11402: out = 1177;
			11403: out = 1155;
			11404: out = 1134;
			11405: out = 1128;
			11406: out = 1127;
			11407: out = 1084;
			11408: out = 1083;
			11409: out = 1082;
			11410: out = 1056;
			11411: out = 1048;
			11412: out = 1031;
			11413: out = 1028;
			11414: out = 1006;
			11415: out = 998;
			11416: out = 987;
			11417: out = 965;
			11418: out = 957;
			11419: out = 944;
			11420: out = 936;
			11421: out = 915;
			11422: out = 904;
			11423: out = 902;
			11424: out = 893;
			11425: out = 871;
			11426: out = 868;
			11427: out = 854;
			11428: out = 838;
			11429: out = 821;
			11430: out = 827;
			11431: out = 797;
			11432: out = 797;
			11433: out = 782;
			11434: out = 770;
			11435: out = 767;
			11436: out = 751;
			11437: out = 751;
			11438: out = 726;
			11439: out = 725;
			11440: out = 711;
			11441: out = 703;
			11442: out = 702;
			11443: out = 680;
			11444: out = 671;
			11445: out = 665;
			11446: out = 653;
			11447: out = 645;
			11448: out = 637;
			11449: out = 628;
			11450: out = 609;
			11451: out = 611;
			11452: out = 597;
			11453: out = 592;
			11454: out = 575;
			11455: out = 581;
			11456: out = 567;
			11457: out = 550;
			11458: out = 557;
			11459: out = 535;
			11460: out = 531;
			11461: out = 535;
			11462: out = 498;
			11463: out = 516;
			11464: out = 500;
			11465: out = 489;
			11466: out = 491;
			11467: out = 474;
			11468: out = 466;
			11469: out = 468;
			11470: out = 459;
			11471: out = 445;
			11472: out = 441;
			11473: out = 399;
			11474: out = 384;
			11475: out = 380;
			11476: out = 345;
			11477: out = 329;
			11478: out = 315;
			11479: out = 285;
			11480: out = 273;
			11481: out = 256;
			11482: out = 231;
			11483: out = 218;
			11484: out = 197;
			11485: out = 186;
			11486: out = 162;
			11487: out = 145;
			11488: out = 133;
			11489: out = 110;
			11490: out = 102;
			11491: out = 79;
			11492: out = 67;
			11493: out = 53;
			11494: out = 37;
			11495: out = 22;
			11496: out = 4;
			11497: out = -14;
			11498: out = -18;
			11499: out = -37;
			11500: out = -46;
			11501: out = -77;
			11502: out = -86;
			11503: out = -97;
			11504: out = -116;
			11505: out = -120;
			11506: out = -128;
			11507: out = -151;
			11508: out = -154;
			11509: out = -170;
			11510: out = -184;
			11511: out = -196;
			11512: out = -208;
			11513: out = -230;
			11514: out = -242;
			11515: out = -240;
			11516: out = -262;
			11517: out = -269;
			11518: out = -282;
			11519: out = -301;
			11520: out = -304;
			11521: out = -316;
			11522: out = -340;
			11523: out = -340;
			11524: out = -360;
			11525: out = -367;
			11526: out = -377;
			11527: out = -391;
			11528: out = -401;
			11529: out = -411;
			11530: out = -418;
			11531: out = -440;
			11532: out = -443;
			11533: out = -468;
			11534: out = -464;
			11535: out = -483;
			11536: out = -489;
			11537: out = -506;
			11538: out = -517;
			11539: out = -516;
			11540: out = -548;
			11541: out = -539;
			11542: out = -563;
			11543: out = -580;
			11544: out = -575;
			11545: out = -588;
			11546: out = -607;
			11547: out = -608;
			11548: out = -635;
			11549: out = -634;
			11550: out = -661;
			11551: out = -653;
			11552: out = -672;
			11553: out = -693;
			11554: out = -701;
			11555: out = -707;
			11556: out = -728;
			11557: out = -739;
			11558: out = -744;
			11559: out = -763;
			11560: out = -779;
			11561: out = -782;
			11562: out = -798;
			11563: out = -823;
			11564: out = -825;
			11565: out = -838;
			11566: out = -857;
			11567: out = -865;
			11568: out = -884;
			11569: out = -898;
			11570: out = -908;
			11571: out = -932;
			11572: out = -961;
			11573: out = -952;
			11574: out = -984;
			11575: out = -981;
			11576: out = -1012;
			11577: out = -1027;
			11578: out = -1048;
			11579: out = -1059;
			11580: out = -1073;
			11581: out = -1099;
			11582: out = -1118;
			11583: out = -1127;
			11584: out = -1167;
			11585: out = -1174;
			11586: out = -1186;
			11587: out = -1210;
			11588: out = -1222;
			11589: out = -1258;
			11590: out = -1265;
			11591: out = -1296;
			11592: out = -1316;
			11593: out = -1351;
			11594: out = -1357;
			11595: out = -1387;
			11596: out = -1399;
			11597: out = -1433;
			11598: out = -1441;
			11599: out = -1471;
			11600: out = -1497;
			11601: out = -1518;
			11602: out = -1534;
			11603: out = -1564;
			11604: out = -1582;
			11605: out = -1605;
			11606: out = -1635;
			11607: out = -1645;
			11608: out = -1675;
			11609: out = -1689;
			11610: out = -1723;
			11611: out = -1731;
			11612: out = -1768;
			11613: out = -1783;
			11614: out = -1803;
			11615: out = -1833;
			11616: out = -1843;
			11617: out = -1868;
			11618: out = -1884;
			11619: out = -1898;
			11620: out = -1935;
			11621: out = -1945;
			11622: out = -1961;
			11623: out = -1992;
			11624: out = -2008;
			11625: out = -2019;
			11626: out = -2038;
			11627: out = -2053;
			11628: out = -2076;
			11629: out = -2091;
			11630: out = -2110;
			11631: out = -2120;
			11632: out = -2132;
			11633: out = -2155;
			11634: out = -2163;
			11635: out = -2181;
			11636: out = -2194;
			11637: out = -2208;
			11638: out = -2219;
			11639: out = -2235;
			11640: out = -2245;
			11641: out = -2261;
			11642: out = -2273;
			11643: out = -2270;
			11644: out = -2290;
			11645: out = -2311;
			11646: out = -2309;
			11647: out = -2322;
			11648: out = -2333;
			11649: out = -2344;
			11650: out = -2348;
			11651: out = -2358;
			11652: out = -2372;
			11653: out = -2369;
			11654: out = -2384;
			11655: out = -2389;
			11656: out = -2393;
			11657: out = -2404;
			11658: out = -2416;
			11659: out = -2417;
			11660: out = -2428;
			11661: out = -2433;
			11662: out = -2432;
			11663: out = -2440;
			11664: out = -2442;
			11665: out = -2462;
			11666: out = -2447;
			11667: out = -2459;
			11668: out = -2474;
			11669: out = -2474;
			11670: out = -2470;
			11671: out = -2467;
			11672: out = -2480;
			11673: out = -2479;
			11674: out = -2490;
			11675: out = -2495;
			11676: out = -2482;
			11677: out = -2495;
			11678: out = -2505;
			11679: out = -2492;
			11680: out = -2499;
			11681: out = -2497;
			11682: out = -2509;
			11683: out = -2504;
			11684: out = -2497;
			11685: out = -2509;
			11686: out = -2507;
			11687: out = -2497;
			11688: out = -2511;
			11689: out = -2499;
			11690: out = -2507;
			11691: out = -2504;
			11692: out = -2499;
			11693: out = -2495;
			11694: out = -2510;
			11695: out = -2502;
			11696: out = -2491;
			11697: out = -2503;
			11698: out = -2495;
			11699: out = -2500;
			11700: out = -2486;
			11701: out = -2494;
			11702: out = -2486;
			11703: out = -2492;
			11704: out = -2481;
			11705: out = -2488;
			11706: out = -2481;
			11707: out = -2476;
			11708: out = -2476;
			11709: out = -2471;
			11710: out = -2476;
			11711: out = -2466;
			11712: out = -2464;
			11713: out = -2464;
			11714: out = -2454;
			11715: out = -2459;
			11716: out = -2446;
			11717: out = -2458;
			11718: out = -2447;
			11719: out = -2441;
			11720: out = -2434;
			11721: out = -2432;
			11722: out = -2436;
			11723: out = -2427;
			11724: out = -2419;
			11725: out = -2409;
			11726: out = -2421;
			11727: out = -2409;
			11728: out = -2405;
			11729: out = -2387;
			11730: out = -2404;
			11731: out = -2387;
			11732: out = -2384;
			11733: out = -2372;
			11734: out = -2385;
			11735: out = -2368;
			11736: out = -2359;
			11737: out = -2363;
			11738: out = -2360;
			11739: out = -2342;
			11740: out = -2347;
			11741: out = -2345;
			11742: out = -2323;
			11743: out = -2325;
			11744: out = -2330;
			11745: out = -2310;
			11746: out = -2310;
			11747: out = -2310;
			11748: out = -2293;
			11749: out = -2297;
			11750: out = -2282;
			11751: out = -2282;
			11752: out = -2270;
			11753: out = -2261;
			11754: out = -2256;
			11755: out = -2258;
			11756: out = -2249;
			11757: out = -2230;
			11758: out = -2228;
			11759: out = -2227;
			11760: out = -2218;
			11761: out = -2214;
			11762: out = -2198;
			11763: out = -2198;
			11764: out = -2186;
			11765: out = -2188;
			11766: out = -2168;
			11767: out = -2169;
			11768: out = -2156;
			11769: out = -2142;
			11770: out = -2145;
			11771: out = -2128;
			11772: out = -2115;
			11773: out = -2107;
			11774: out = -2098;
			11775: out = -2090;
			11776: out = -2083;
			11777: out = -2068;
			11778: out = -2048;
			11779: out = -2050;
			11780: out = -2043;
			11781: out = -2017;
			11782: out = -2012;
			11783: out = -2001;
			11784: out = -1984;
			11785: out = -1979;
			11786: out = -1965;
			11787: out = -1951;
			11788: out = -1930;
			11789: out = -1924;
			11790: out = -1900;
			11791: out = -1895;
			11792: out = -1876;
			11793: out = -1856;
			11794: out = -1854;
			11795: out = -1827;
			11796: out = -1816;
			11797: out = -1795;
			11798: out = -1797;
			11799: out = -1757;
			11800: out = -1754;
			11801: out = -1732;
			11802: out = -1714;
			11803: out = -1707;
			11804: out = -1685;
			11805: out = -1658;
			11806: out = -1655;
			11807: out = -1629;
			11808: out = -1618;
			11809: out = -1599;
			11810: out = -1581;
			11811: out = -1561;
			11812: out = -1545;
			11813: out = -1531;
			11814: out = -1511;
			11815: out = -1492;
			11816: out = -1475;
			11817: out = -1466;
			11818: out = -1448;
			11819: out = -1424;
			11820: out = -1404;
			11821: out = -1391;
			11822: out = -1381;
			11823: out = -1354;
			11824: out = -1338;
			11825: out = -1333;
			11826: out = -1296;
			11827: out = -1305;
			11828: out = -1274;
			11829: out = -1253;
			11830: out = -1237;
			11831: out = -1227;
			11832: out = -1210;
			11833: out = -1189;
			11834: out = -1181;
			11835: out = -1156;
			11836: out = -1142;
			11837: out = -1149;
			11838: out = -1104;
			11839: out = -1099;
			11840: out = -1082;
			11841: out = -1063;
			11842: out = -1066;
			11843: out = -1036;
			11844: out = -1025;
			11845: out = -1003;
			11846: out = -993;
			11847: out = -987;
			11848: out = -965;
			11849: out = -942;
			11850: out = -943;
			11851: out = -921;
			11852: out = -910;
			11853: out = -893;
			11854: out = -885;
			11855: out = -868;
			11856: out = -849;
			11857: out = -858;
			11858: out = -826;
			11859: out = -817;
			11860: out = -810;
			11861: out = -788;
			11862: out = -784;
			11863: out = -767;
			11864: out = -761;
			11865: out = -754;
			11866: out = -737;
			11867: out = -716;
			11868: out = -716;
			11869: out = -697;
			11870: out = -688;
			11871: out = -681;
			11872: out = -660;
			11873: out = -667;
			11874: out = -644;
			11875: out = -633;
			11876: out = -630;
			11877: out = -606;
			11878: out = -609;
			11879: out = -590;
			11880: out = -592;
			11881: out = -570;
			11882: out = -569;
			11883: out = -560;
			11884: out = -542;
			11885: out = -539;
			11886: out = -534;
			11887: out = -518;
			11888: out = -510;
			11889: out = -501;
			11890: out = -505;
			11891: out = -480;
			11892: out = -477;
			11893: out = -464;
			11894: out = -466;
			11895: out = -452;
			11896: out = -436;
			11897: out = -428;
			11898: out = -404;
			11899: out = -400;
			11900: out = -380;
			11901: out = -363;
			11902: out = -349;
			11903: out = -347;
			11904: out = -321;
			11905: out = -312;
			11906: out = -308;
			11907: out = -286;
			11908: out = -277;
			11909: out = -253;
			11910: out = -254;
			11911: out = -232;
			11912: out = -226;
			11913: out = -210;
			11914: out = -198;
			11915: out = -192;
			11916: out = -181;
			11917: out = -170;
			11918: out = -155;
			11919: out = -146;
			11920: out = -139;
			11921: out = -124;
			11922: out = -108;
			11923: out = -101;
			11924: out = -102;
			11925: out = -78;
			11926: out = -78;
			11927: out = -49;
			11928: out = -69;
			11929: out = -46;
			11930: out = -36;
			11931: out = -26;
			11932: out = -15;
			11933: out = -6;
			11934: out = 2;
			11935: out = 20;
			11936: out = 15;
			11937: out = 27;
			11938: out = 42;
			11939: out = 46;
			11940: out = 46;
			11941: out = 66;
			11942: out = 77;
			11943: out = 75;
			11944: out = 90;
			11945: out = 102;
			11946: out = 101;
			11947: out = 108;
			11948: out = 129;
			11949: out = 136;
			11950: out = 131;
			11951: out = 149;
			11952: out = 151;
			11953: out = 157;
			11954: out = 180;
			11955: out = 172;
			11956: out = 191;
			11957: out = 200;
			11958: out = 196;
			11959: out = 212;
			11960: out = 223;
			11961: out = 233;
			11962: out = 235;
			11963: out = 243;
			11964: out = 253;
			11965: out = 253;
			11966: out = 274;
			11967: out = 270;
			11968: out = 282;
			11969: out = 292;
			11970: out = 299;
			11971: out = 312;
			11972: out = 318;
			11973: out = 329;
			11974: out = 332;
			11975: out = 349;
			11976: out = 359;
			11977: out = 361;
			11978: out = 369;
			11979: out = 384;
			11980: out = 388;
			11981: out = 389;
			11982: out = 409;
			11983: out = 418;
			11984: out = 429;
			11985: out = 434;
			11986: out = 454;
			11987: out = 459;
			11988: out = 467;
			11989: out = 480;
			11990: out = 487;
			11991: out = 502;
			11992: out = 510;
			11993: out = 524;
			11994: out = 539;
			11995: out = 543;
			11996: out = 562;
			11997: out = 567;
			11998: out = 587;
			11999: out = 589;
			12000: out = 613;
			12001: out = 620;
			12002: out = 640;
			12003: out = 641;
			12004: out = 666;
			12005: out = 675;
			12006: out = 685;
			12007: out = 703;
			12008: out = 724;
			12009: out = 730;
			12010: out = 747;
			12011: out = 767;
			12012: out = 780;
			12013: out = 798;
			12014: out = 803;
			12015: out = 824;
			12016: out = 836;
			12017: out = 859;
			12018: out = 864;
			12019: out = 892;
			12020: out = 901;
			12021: out = 919;
			12022: out = 933;
			12023: out = 951;
			12024: out = 960;
			12025: out = 984;
			12026: out = 996;
			12027: out = 1009;
			12028: out = 1024;
			12029: out = 1044;
			12030: out = 1055;
			12031: out = 1079;
			12032: out = 1081;
			12033: out = 1089;
			12034: out = 1120;
			12035: out = 1133;
			12036: out = 1156;
			12037: out = 1154;
			12038: out = 1176;
			12039: out = 1192;
			12040: out = 1200;
			12041: out = 1209;
			12042: out = 1226;
			12043: out = 1238;
			12044: out = 1261;
			12045: out = 1272;
			12046: out = 1279;
			12047: out = 1296;
			12048: out = 1312;
			12049: out = 1326;
			12050: out = 1334;
			12051: out = 1335;
			12052: out = 1366;
			12053: out = 1375;
			12054: out = 1389;
			12055: out = 1393;
			12056: out = 1405;
			12057: out = 1423;
			12058: out = 1433;
			12059: out = 1444;
			12060: out = 1452;
			12061: out = 1465;
			12062: out = 1476;
			12063: out = 1495;
			12064: out = 1500;
			12065: out = 1511;
			12066: out = 1516;
			12067: out = 1543;
			12068: out = 1527;
			12069: out = 1552;
			12070: out = 1560;
			12071: out = 1576;
			12072: out = 1586;
			12073: out = 1583;
			12074: out = 1608;
			12075: out = 1613;
			12076: out = 1625;
			12077: out = 1619;
			12078: out = 1641;
			12079: out = 1651;
			12080: out = 1661;
			12081: out = 1659;
			12082: out = 1688;
			12083: out = 1684;
			12084: out = 1690;
			12085: out = 1703;
			12086: out = 1719;
			12087: out = 1713;
			12088: out = 1734;
			12089: out = 1742;
			12090: out = 1745;
			12091: out = 1750;
			12092: out = 1768;
			12093: out = 1769;
			12094: out = 1778;
			12095: out = 1796;
			12096: out = 1791;
			12097: out = 1813;
			12098: out = 1803;
			12099: out = 1824;
			12100: out = 1828;
			12101: out = 1836;
			12102: out = 1849;
			12103: out = 1844;
			12104: out = 1856;
			12105: out = 1871;
			12106: out = 1873;
			12107: out = 1872;
			12108: out = 1886;
			12109: out = 1891;
			12110: out = 1902;
			12111: out = 1914;
			12112: out = 1912;
			12113: out = 1916;
			12114: out = 1935;
			12115: out = 1929;
			12116: out = 1937;
			12117: out = 1949;
			12118: out = 1960;
			12119: out = 1953;
			12120: out = 1977;
			12121: out = 1980;
			12122: out = 1981;
			12123: out = 1991;
			12124: out = 1991;
			12125: out = 2000;
			12126: out = 2010;
			12127: out = 2009;
			12128: out = 2007;
			12129: out = 2024;
			12130: out = 2027;
			12131: out = 2034;
			12132: out = 2027;
			12133: out = 2026;
			12134: out = 2036;
			12135: out = 2027;
			12136: out = 2026;
			12137: out = 2026;
			12138: out = 2013;
			12139: out = 2026;
			12140: out = 2022;
			12141: out = 2016;
			12142: out = 2024;
			12143: out = 2028;
			12144: out = 2017;
			12145: out = 2016;
			12146: out = 2012;
			12147: out = 2013;
			12148: out = 2013;
			12149: out = 2007;
			12150: out = 2001;
			12151: out = 2015;
			12152: out = 2008;
			12153: out = 2015;
			12154: out = 2001;
			12155: out = 2008;
			12156: out = 2009;
			12157: out = 2002;
			12158: out = 2009;
			12159: out = 2006;
			12160: out = 2002;
			12161: out = 2003;
			12162: out = 2004;
			12163: out = 1996;
			12164: out = 2009;
			12165: out = 2003;
			12166: out = 2006;
			12167: out = 2012;
			12168: out = 2009;
			12169: out = 2005;
			12170: out = 1998;
			12171: out = 2000;
			12172: out = 2000;
			12173: out = 1991;
			12174: out = 2000;
			12175: out = 1982;
			12176: out = 1985;
			12177: out = 2003;
			12178: out = 1989;
			12179: out = 1997;
			12180: out = 1986;
			12181: out = 1997;
			12182: out = 1983;
			12183: out = 1986;
			12184: out = 1994;
			12185: out = 1983;
			12186: out = 1982;
			12187: out = 1978;
			12188: out = 1980;
			12189: out = 1967;
			12190: out = 1968;
			12191: out = 1986;
			12192: out = 1969;
			12193: out = 1966;
			12194: out = 1970;
			12195: out = 1962;
			12196: out = 1958;
			12197: out = 1969;
			12198: out = 1958;
			12199: out = 1959;
			12200: out = 1942;
			12201: out = 1942;
			12202: out = 1941;
			12203: out = 1934;
			12204: out = 1924;
			12205: out = 1944;
			12206: out = 1925;
			12207: out = 1922;
			12208: out = 1909;
			12209: out = 1903;
			12210: out = 1911;
			12211: out = 1877;
			12212: out = 1890;
			12213: out = 1880;
			12214: out = 1865;
			12215: out = 1858;
			12216: out = 1856;
			12217: out = 1844;
			12218: out = 1845;
			12219: out = 1830;
			12220: out = 1832;
			12221: out = 1823;
			12222: out = 1809;
			12223: out = 1806;
			12224: out = 1800;
			12225: out = 1781;
			12226: out = 1784;
			12227: out = 1766;
			12228: out = 1745;
			12229: out = 1743;
			12230: out = 1740;
			12231: out = 1723;
			12232: out = 1701;
			12233: out = 1691;
			12234: out = 1693;
			12235: out = 1661;
			12236: out = 1664;
			12237: out = 1653;
			12238: out = 1642;
			12239: out = 1615;
			12240: out = 1613;
			12241: out = 1601;
			12242: out = 1595;
			12243: out = 1566;
			12244: out = 1566;
			12245: out = 1551;
			12246: out = 1534;
			12247: out = 1522;
			12248: out = 1513;
			12249: out = 1509;
			12250: out = 1470;
			12251: out = 1465;
			12252: out = 1462;
			12253: out = 1441;
			12254: out = 1433;
			12255: out = 1414;
			12256: out = 1395;
			12257: out = 1393;
			12258: out = 1374;
			12259: out = 1366;
			12260: out = 1353;
			12261: out = 1333;
			12262: out = 1329;
			12263: out = 1300;
			12264: out = 1299;
			12265: out = 1280;
			12266: out = 1267;
			12267: out = 1257;
			12268: out = 1247;
			12269: out = 1224;
			12270: out = 1227;
			12271: out = 1210;
			12272: out = 1184;
			12273: out = 1186;
			12274: out = 1168;
			12275: out = 1157;
			12276: out = 1142;
			12277: out = 1131;
			12278: out = 1108;
			12279: out = 1101;
			12280: out = 1105;
			12281: out = 1074;
			12282: out = 1068;
			12283: out = 1066;
			12284: out = 1048;
			12285: out = 1037;
			12286: out = 1023;
			12287: out = 1011;
			12288: out = 999;
			12289: out = 992;
			12290: out = 983;
			12291: out = 964;
			12292: out = 944;
			12293: out = 951;
			12294: out = 927;
			12295: out = 917;
			12296: out = 909;
			12297: out = 901;
			12298: out = 900;
			12299: out = 885;
			12300: out = 872;
			12301: out = 860;
			12302: out = 844;
			12303: out = 841;
			12304: out = 830;
			12305: out = 810;
			12306: out = 803;
			12307: out = 803;
			12308: out = 784;
			12309: out = 778;
			12310: out = 750;
			12311: out = 771;
			12312: out = 741;
			12313: out = 727;
			12314: out = 729;
			12315: out = 729;
			12316: out = 706;
			12317: out = 702;
			12318: out = 695;
			12319: out = 676;
			12320: out = 672;
			12321: out = 667;
			12322: out = 643;
			12323: out = 649;
			12324: out = 642;
			12325: out = 628;
			12326: out = 619;
			12327: out = 609;
			12328: out = 605;
			12329: out = 590;
			12330: out = 600;
			12331: out = 564;
			12332: out = 572;
			12333: out = 565;
			12334: out = 547;
			12335: out = 550;
			12336: out = 529;
			12337: out = 531;
			12338: out = 522;
			12339: out = 511;
			12340: out = 515;
			12341: out = 501;
			12342: out = 489;
			12343: out = 481;
			12344: out = 481;
			12345: out = 471;
			12346: out = 465;
			12347: out = 448;
			12348: out = 463;
			12349: out = 435;
			12350: out = 436;
			12351: out = 429;
			12352: out = 442;
			12353: out = 411;
			12354: out = 405;
			12355: out = 407;
			12356: out = 393;
			12357: out = 389;
			12358: out = 385;
			12359: out = 376;
			12360: out = 369;
			12361: out = 371;
			12362: out = 360;
			12363: out = 347;
			12364: out = 332;
			12365: out = 311;
			12366: out = 297;
			12367: out = 285;
			12368: out = 262;
			12369: out = 247;
			12370: out = 232;
			12371: out = 223;
			12372: out = 199;
			12373: out = 182;
			12374: out = 180;
			12375: out = 157;
			12376: out = 156;
			12377: out = 117;
			12378: out = 120;
			12379: out = 101;
			12380: out = 89;
			12381: out = 85;
			12382: out = 60;
			12383: out = 54;
			12384: out = 49;
			12385: out = 15;
			12386: out = 18;
			12387: out = 7;
			12388: out = -15;
			12389: out = -22;
			12390: out = -29;
			12391: out = -45;
			12392: out = -52;
			12393: out = -69;
			12394: out = -83;
			12395: out = -96;
			12396: out = -89;
			12397: out = -114;
			12398: out = -128;
			12399: out = -136;
			12400: out = -147;
			12401: out = -158;
			12402: out = -169;
			12403: out = -175;
			12404: out = -192;
			12405: out = -186;
			12406: out = -210;
			12407: out = -216;
			12408: out = -218;
			12409: out = -247;
			12410: out = -244;
			12411: out = -254;
			12412: out = -263;
			12413: out = -278;
			12414: out = -291;
			12415: out = -294;
			12416: out = -299;
			12417: out = -321;
			12418: out = -321;
			12419: out = -337;
			12420: out = -336;
			12421: out = -352;
			12422: out = -360;
			12423: out = -370;
			12424: out = -379;
			12425: out = -392;
			12426: out = -400;
			12427: out = -407;
			12428: out = -417;
			12429: out = -427;
			12430: out = -443;
			12431: out = -439;
			12432: out = -463;
			12433: out = -460;
			12434: out = -465;
			12435: out = -482;
			12436: out = -502;
			12437: out = -490;
			12438: out = -515;
			12439: out = -523;
			12440: out = -526;
			12441: out = -538;
			12442: out = -557;
			12443: out = -551;
			12444: out = -572;
			12445: out = -577;
			12446: out = -584;
			12447: out = -605;
			12448: out = -610;
			12449: out = -622;
			12450: out = -630;
			12451: out = -636;
			12452: out = -655;
			12453: out = -668;
			12454: out = -670;
			12455: out = -688;
			12456: out = -694;
			12457: out = -706;
			12458: out = -725;
			12459: out = -737;
			12460: out = -748;
			12461: out = -759;
			12462: out = -762;
			12463: out = -784;
			12464: out = -795;
			12465: out = -801;
			12466: out = -830;
			12467: out = -834;
			12468: out = -845;
			12469: out = -864;
			12470: out = -881;
			12471: out = -882;
			12472: out = -917;
			12473: out = -912;
			12474: out = -939;
			12475: out = -948;
			12476: out = -978;
			12477: out = -979;
			12478: out = -998;
			12479: out = -1020;
			12480: out = -1033;
			12481: out = -1056;
			12482: out = -1062;
			12483: out = -1085;
			12484: out = -1090;
			12485: out = -1117;
			12486: out = -1130;
			12487: out = -1145;
			12488: out = -1188;
			12489: out = -1184;
			12490: out = -1216;
			12491: out = -1225;
			12492: out = -1252;
			12493: out = -1262;
			12494: out = -1284;
			12495: out = -1296;
			12496: out = -1312;
			12497: out = -1342;
			12498: out = -1350;
			12499: out = -1376;
			12500: out = -1389;
			12501: out = -1415;
			12502: out = -1424;
			12503: out = -1449;
			12504: out = -1459;
			12505: out = -1485;
			12506: out = -1493;
			12507: out = -1512;
			12508: out = -1529;
			12509: out = -1547;
			12510: out = -1564;
			12511: out = -1570;
			12512: out = -1599;
			12513: out = -1607;
			12514: out = -1617;
			12515: out = -1653;
			12516: out = -1654;
			12517: out = -1662;
			12518: out = -1687;
			12519: out = -1697;
			12520: out = -1709;
			12521: out = -1711;
			12522: out = -1732;
			12523: out = -1757;
			12524: out = -1761;
			12525: out = -1764;
			12526: out = -1793;
			12527: out = -1799;
			12528: out = -1802;
			12529: out = -1818;
			12530: out = -1825;
			12531: out = -1840;
			12532: out = -1835;
			12533: out = -1862;
			12534: out = -1865;
			12535: out = -1874;
			12536: out = -1880;
			12537: out = -1885;
			12538: out = -1908;
			12539: out = -1904;
			12540: out = -1910;
			12541: out = -1916;
			12542: out = -1933;
			12543: out = -1932;
			12544: out = -1945;
			12545: out = -1938;
			12546: out = -1961;
			12547: out = -1961;
			12548: out = -1960;
			12549: out = -1974;
			12550: out = -1977;
			12551: out = -1977;
			12552: out = -1994;
			12553: out = -1984;
			12554: out = -1995;
			12555: out = -2002;
			12556: out = -1992;
			12557: out = -2014;
			12558: out = -2009;
			12559: out = -2012;
			12560: out = -2017;
			12561: out = -2020;
			12562: out = -2018;
			12563: out = -2030;
			12564: out = -2022;
			12565: out = -2029;
			12566: out = -2025;
			12567: out = -2041;
			12568: out = -2024;
			12569: out = -2044;
			12570: out = -2022;
			12571: out = -2041;
			12572: out = -2041;
			12573: out = -2032;
			12574: out = -2037;
			12575: out = -2046;
			12576: out = -2040;
			12577: out = -2039;
			12578: out = -2039;
			12579: out = -2049;
			12580: out = -2041;
			12581: out = -2040;
			12582: out = -2038;
			12583: out = -2043;
			12584: out = -2039;
			12585: out = -2039;
			12586: out = -2025;
			12587: out = -2044;
			12588: out = -2031;
			12589: out = -2028;
			12590: out = -2033;
			12591: out = -2028;
			12592: out = -2031;
			12593: out = -2025;
			12594: out = -2029;
			12595: out = -2017;
			12596: out = -2021;
			12597: out = -2015;
			12598: out = -2018;
			12599: out = -2003;
			12600: out = -2025;
			12601: out = -2003;
			12602: out = -2006;
			12603: out = -2006;
			12604: out = -1995;
			12605: out = -2003;
			12606: out = -1996;
			12607: out = -1987;
			12608: out = -1991;
			12609: out = -1974;
			12610: out = -1989;
			12611: out = -1975;
			12612: out = -1983;
			12613: out = -1972;
			12614: out = -1965;
			12615: out = -1968;
			12616: out = -1963;
			12617: out = -1961;
			12618: out = -1949;
			12619: out = -1956;
			12620: out = -1946;
			12621: out = -1941;
			12622: out = -1941;
			12623: out = -1934;
			12624: out = -1936;
			12625: out = -1932;
			12626: out = -1921;
			12627: out = -1923;
			12628: out = -1915;
			12629: out = -1914;
			12630: out = -1909;
			12631: out = -1896;
			12632: out = -1898;
			12633: out = -1900;
			12634: out = -1886;
			12635: out = -1879;
			12636: out = -1885;
			12637: out = -1877;
			12638: out = -1864;
			12639: out = -1873;
			12640: out = -1861;
			12641: out = -1843;
			12642: out = -1862;
			12643: out = -1841;
			12644: out = -1847;
			12645: out = -1825;
			12646: out = -1836;
			12647: out = -1823;
			12648: out = -1819;
			12649: out = -1807;
			12650: out = -1815;
			12651: out = -1793;
			12652: out = -1795;
			12653: out = -1792;
			12654: out = -1778;
			12655: out = -1777;
			12656: out = -1768;
			12657: out = -1766;
			12658: out = -1750;
			12659: out = -1752;
			12660: out = -1748;
			12661: out = -1733;
			12662: out = -1721;
			12663: out = -1723;
			12664: out = -1716;
			12665: out = -1709;
			12666: out = -1693;
			12667: out = -1694;
			12668: out = -1679;
			12669: out = -1678;
			12670: out = -1662;
			12671: out = -1660;
			12672: out = -1642;
			12673: out = -1640;
			12674: out = -1625;
			12675: out = -1614;
			12676: out = -1608;
			12677: out = -1595;
			12678: out = -1587;
			12679: out = -1568;
			12680: out = -1563;
			12681: out = -1549;
			12682: out = -1539;
			12683: out = -1524;
			12684: out = -1513;
			12685: out = -1498;
			12686: out = -1494;
			12687: out = -1473;
			12688: out = -1471;
			12689: out = -1444;
			12690: out = -1434;
			12691: out = -1433;
			12692: out = -1406;
			12693: out = -1399;
			12694: out = -1387;
			12695: out = -1380;
			12696: out = -1351;
			12697: out = -1343;
			12698: out = -1339;
			12699: out = -1317;
			12700: out = -1299;
			12701: out = -1291;
			12702: out = -1275;
			12703: out = -1257;
			12704: out = -1246;
			12705: out = -1225;
			12706: out = -1221;
			12707: out = -1213;
			12708: out = -1187;
			12709: out = -1169;
			12710: out = -1165;
			12711: out = -1150;
			12712: out = -1133;
			12713: out = -1113;
			12714: out = -1109;
			12715: out = -1094;
			12716: out = -1081;
			12717: out = -1063;
			12718: out = -1056;
			12719: out = -1032;
			12720: out = -1021;
			12721: out = -1020;
			12722: out = -989;
			12723: out = -990;
			12724: out = -973;
			12725: out = -964;
			12726: out = -937;
			12727: out = -948;
			12728: out = -917;
			12729: out = -908;
			12730: out = -895;
			12731: out = -877;
			12732: out = -880;
			12733: out = -858;
			12734: out = -856;
			12735: out = -833;
			12736: out = -825;
			12737: out = -817;
			12738: out = -802;
			12739: out = -782;
			12740: out = -784;
			12741: out = -767;
			12742: out = -752;
			12743: out = -743;
			12744: out = -738;
			12745: out = -728;
			12746: out = -708;
			12747: out = -700;
			12748: out = -699;
			12749: out = -679;
			12750: out = -669;
			12751: out = -666;
			12752: out = -656;
			12753: out = -633;
			12754: out = -634;
			12755: out = -621;
			12756: out = -606;
			12757: out = -589;
			12758: out = -604;
			12759: out = -576;
			12760: out = -587;
			12761: out = -552;
			12762: out = -564;
			12763: out = -555;
			12764: out = -534;
			12765: out = -531;
			12766: out = -522;
			12767: out = -521;
			12768: out = -502;
			12769: out = -498;
			12770: out = -484;
			12771: out = -483;
			12772: out = -468;
			12773: out = -472;
			12774: out = -457;
			12775: out = -450;
			12776: out = -440;
			12777: out = -441;
			12778: out = -420;
			12779: out = -424;
			12780: out = -413;
			12781: out = -399;
			12782: out = -405;
			12783: out = -400;
			12784: out = -374;
			12785: out = -381;
			12786: out = -373;
			12787: out = -358;
			12788: out = -349;
			12789: out = -340;
			12790: out = -330;
			12791: out = -300;
			12792: out = -310;
			12793: out = -288;
			12794: out = -277;
			12795: out = -267;
			12796: out = -263;
			12797: out = -246;
			12798: out = -241;
			12799: out = -233;
			12800: out = -221;
			12801: out = -199;
			12802: out = -198;
			12803: out = -191;
			12804: out = -183;
			12805: out = -161;
			12806: out = -163;
			12807: out = -149;
			12808: out = -141;
			12809: out = -138;
			12810: out = -131;
			12811: out = -112;
			12812: out = -110;
			12813: out = -92;
			12814: out = -95;
			12815: out = -84;
			12816: out = -69;
			12817: out = -72;
			12818: out = -53;
			12819: out = -54;
			12820: out = -44;
			12821: out = -41;
			12822: out = -20;
			12823: out = -19;
			12824: out = -15;
			12825: out = -3;
			12826: out = 1;
			12827: out = 3;
			12828: out = 19;
			12829: out = 26;
			12830: out = 31;
			12831: out = 40;
			12832: out = 36;
			12833: out = 62;
			12834: out = 54;
			12835: out = 66;
			12836: out = 76;
			12837: out = 73;
			12838: out = 83;
			12839: out = 99;
			12840: out = 101;
			12841: out = 108;
			12842: out = 114;
			12843: out = 119;
			12844: out = 120;
			12845: out = 138;
			12846: out = 127;
			12847: out = 148;
			12848: out = 148;
			12849: out = 155;
			12850: out = 168;
			12851: out = 168;
			12852: out = 184;
			12853: out = 175;
			12854: out = 198;
			12855: out = 187;
			12856: out = 204;
			12857: out = 204;
			12858: out = 217;
			12859: out = 220;
			12860: out = 239;
			12861: out = 230;
			12862: out = 249;
			12863: out = 249;
			12864: out = 257;
			12865: out = 269;
			12866: out = 273;
			12867: out = 274;
			12868: out = 283;
			12869: out = 304;
			12870: out = 294;
			12871: out = 305;
			12872: out = 316;
			12873: out = 330;
			12874: out = 325;
			12875: out = 341;
			12876: out = 349;
			12877: out = 362;
			12878: out = 368;
			12879: out = 365;
			12880: out = 381;
			12881: out = 391;
			12882: out = 408;
			12883: out = 408;
			12884: out = 408;
			12885: out = 431;
			12886: out = 434;
			12887: out = 456;
			12888: out = 444;
			12889: out = 467;
			12890: out = 480;
			12891: out = 499;
			12892: out = 493;
			12893: out = 515;
			12894: out = 522;
			12895: out = 535;
			12896: out = 538;
			12897: out = 557;
			12898: out = 558;
			12899: out = 585;
			12900: out = 589;
			12901: out = 602;
			12902: out = 618;
			12903: out = 623;
			12904: out = 644;
			12905: out = 645;
			12906: out = 667;
			12907: out = 671;
			12908: out = 684;
			12909: out = 697;
			12910: out = 722;
			12911: out = 726;
			12912: out = 734;
			12913: out = 753;
			12914: out = 764;
			12915: out = 771;
			12916: out = 793;
			12917: out = 798;
			12918: out = 810;
			12919: out = 833;
			12920: out = 831;
			12921: out = 854;
			12922: out = 854;
			12923: out = 878;
			12924: out = 894;
			12925: out = 894;
			12926: out = 909;
			12927: out = 925;
			12928: out = 943;
			12929: out = 940;
			12930: out = 960;
			12931: out = 964;
			12932: out = 993;
			12933: out = 978;
			12934: out = 1007;
			12935: out = 1012;
			12936: out = 1028;
			12937: out = 1033;
			12938: out = 1051;
			12939: out = 1059;
			12940: out = 1071;
			12941: out = 1083;
			12942: out = 1079;
			12943: out = 1108;
			12944: out = 1096;
			12945: out = 1121;
			12946: out = 1120;
			12947: out = 1137;
			12948: out = 1144;
			12949: out = 1146;
			12950: out = 1169;
			12951: out = 1166;
			12952: out = 1188;
			12953: out = 1184;
			12954: out = 1202;
			12955: out = 1210;
			12956: out = 1219;
			12957: out = 1219;
			12958: out = 1236;
			12959: out = 1239;
			12960: out = 1249;
			12961: out = 1257;
			12962: out = 1274;
			12963: out = 1267;
			12964: out = 1284;
			12965: out = 1294;
			12966: out = 1293;
			12967: out = 1314;
			12968: out = 1309;
			12969: out = 1327;
			12970: out = 1326;
			12971: out = 1330;
			12972: out = 1348;
			12973: out = 1352;
			12974: out = 1358;
			12975: out = 1366;
			12976: out = 1376;
			12977: out = 1370;
			12978: out = 1399;
			12979: out = 1391;
			12980: out = 1403;
			12981: out = 1405;
			12982: out = 1416;
			12983: out = 1425;
			12984: out = 1422;
			12985: out = 1441;
			12986: out = 1434;
			12987: out = 1450;
			12988: out = 1449;
			12989: out = 1462;
			12990: out = 1469;
			12991: out = 1464;
			12992: out = 1481;
			12993: out = 1481;
			12994: out = 1492;
			12995: out = 1493;
			12996: out = 1503;
			12997: out = 1505;
			12998: out = 1521;
			12999: out = 1517;
			13000: out = 1520;
			13001: out = 1530;
			13002: out = 1544;
			13003: out = 1539;
			13004: out = 1543;
			13005: out = 1563;
			13006: out = 1555;
			13007: out = 1558;
			13008: out = 1575;
			13009: out = 1570;
			13010: out = 1582;
			13011: out = 1584;
			13012: out = 1591;
			13013: out = 1598;
			13014: out = 1601;
			13015: out = 1599;
			13016: out = 1614;
			13017: out = 1616;
			13018: out = 1623;
			13019: out = 1624;
			13020: out = 1620;
			13021: out = 1628;
			13022: out = 1628;
			13023: out = 1630;
			13024: out = 1628;
			13025: out = 1631;
			13026: out = 1628;
			13027: out = 1626;
			13028: out = 1627;
			13029: out = 1630;
			13030: out = 1628;
			13031: out = 1637;
			13032: out = 1634;
			13033: out = 1623;
			13034: out = 1618;
			13035: out = 1632;
			13036: out = 1604;
			13037: out = 1616;
			13038: out = 1624;
			13039: out = 1617;
			13040: out = 1618;
			13041: out = 1613;
			13042: out = 1612;
			13043: out = 1619;
			13044: out = 1620;
			13045: out = 1611;
			13046: out = 1615;
			13047: out = 1602;
			13048: out = 1622;
			13049: out = 1624;
			13050: out = 1601;
			13051: out = 1622;
			13052: out = 1623;
			13053: out = 1626;
			13054: out = 1603;
			13055: out = 1606;
			13056: out = 1612;
			13057: out = 1612;
			13058: out = 1607;
			13059: out = 1607;
			13060: out = 1618;
			13061: out = 1625;
			13062: out = 1624;
			13063: out = 1615;
			13064: out = 1618;
			13065: out = 1616;
			13066: out = 1589;
			13067: out = 1600;
			13068: out = 1611;
			13069: out = 1598;
			13070: out = 1593;
			13071: out = 1605;
			13072: out = 1607;
			13073: out = 1600;
			13074: out = 1605;
			13075: out = 1610;
			13076: out = 1599;
			13077: out = 1600;
			13078: out = 1601;
			13079: out = 1587;
			13080: out = 1607;
			13081: out = 1588;
			13082: out = 1593;
			13083: out = 1592;
			13084: out = 1576;
			13085: out = 1595;
			13086: out = 1581;
			13087: out = 1586;
			13088: out = 1581;
			13089: out = 1581;
			13090: out = 1576;
			13091: out = 1574;
			13092: out = 1570;
			13093: out = 1567;
			13094: out = 1555;
			13095: out = 1561;
			13096: out = 1566;
			13097: out = 1554;
			13098: out = 1554;
			13099: out = 1540;
			13100: out = 1548;
			13101: out = 1541;
			13102: out = 1523;
			13103: out = 1522;
			13104: out = 1518;
			13105: out = 1515;
			13106: out = 1513;
			13107: out = 1492;
			13108: out = 1500;
			13109: out = 1484;
			13110: out = 1480;
			13111: out = 1480;
			13112: out = 1478;
			13113: out = 1454;
			13114: out = 1458;
			13115: out = 1451;
			13116: out = 1435;
			13117: out = 1435;
			13118: out = 1422;
			13119: out = 1405;
			13120: out = 1410;
			13121: out = 1394;
			13122: out = 1387;
			13123: out = 1385;
			13124: out = 1364;
			13125: out = 1364;
			13126: out = 1344;
			13127: out = 1347;
			13128: out = 1332;
			13129: out = 1320;
			13130: out = 1303;
			13131: out = 1298;
			13132: out = 1294;
			13133: out = 1274;
			13134: out = 1263;
			13135: out = 1264;
			13136: out = 1244;
			13137: out = 1237;
			13138: out = 1224;
			13139: out = 1212;
			13140: out = 1204;
			13141: out = 1189;
			13142: out = 1177;
			13143: out = 1173;
			13144: out = 1157;
			13145: out = 1157;
			13146: out = 1131;
			13147: out = 1118;
			13148: out = 1119;
			13149: out = 1097;
			13150: out = 1094;
			13151: out = 1091;
			13152: out = 1059;
			13153: out = 1067;
			13154: out = 1047;
			13155: out = 1038;
			13156: out = 1023;
			13157: out = 1018;
			13158: out = 1009;
			13159: out = 988;
			13160: out = 989;
			13161: out = 975;
			13162: out = 963;
			13163: out = 953;
			13164: out = 953;
			13165: out = 931;
			13166: out = 921;
			13167: out = 909;
			13168: out = 890;
			13169: out = 897;
			13170: out = 877;
			13171: out = 858;
			13172: out = 862;
			13173: out = 848;
			13174: out = 848;
			13175: out = 818;
			13176: out = 826;
			13177: out = 803;
			13178: out = 805;
			13179: out = 789;
			13180: out = 782;
			13181: out = 774;
			13182: out = 754;
			13183: out = 763;
			13184: out = 738;
			13185: out = 743;
			13186: out = 719;
			13187: out = 730;
			13188: out = 700;
			13189: out = 703;
			13190: out = 692;
			13191: out = 683;
			13192: out = 676;
			13193: out = 666;
			13194: out = 655;
			13195: out = 655;
			13196: out = 634;
			13197: out = 643;
			13198: out = 623;
			13199: out = 617;
			13200: out = 611;
			13201: out = 600;
			13202: out = 587;
			13203: out = 592;
			13204: out = 590;
			13205: out = 567;
			13206: out = 559;
			13207: out = 554;
			13208: out = 552;
			13209: out = 537;
			13210: out = 526;
			13211: out = 523;
			13212: out = 521;
			13213: out = 518;
			13214: out = 496;
			13215: out = 489;
			13216: out = 490;
			13217: out = 476;
			13218: out = 484;
			13219: out = 453;
			13220: out = 458;
			13221: out = 460;
			13222: out = 450;
			13223: out = 441;
			13224: out = 435;
			13225: out = 433;
			13226: out = 422;
			13227: out = 411;
			13228: out = 411;
			13229: out = 403;
			13230: out = 385;
			13231: out = 394;
			13232: out = 392;
			13233: out = 387;
			13234: out = 367;
			13235: out = 374;
			13236: out = 364;
			13237: out = 356;
			13238: out = 356;
			13239: out = 345;
			13240: out = 327;
			13241: out = 348;
			13242: out = 323;
			13243: out = 329;
			13244: out = 309;
			13245: out = 314;
			13246: out = 315;
			13247: out = 296;
			13248: out = 305;
			13249: out = 300;
			13250: out = 288;
			13251: out = 287;
			13252: out = 287;
			13253: out = 265;
			13254: out = 266;
			13255: out = 267;
			13256: out = 226;
			13257: out = 221;
			13258: out = 219;
			13259: out = 196;
			13260: out = 192;
			13261: out = 170;
			13262: out = 162;
			13263: out = 148;
			13264: out = 149;
			13265: out = 114;
			13266: out = 120;
			13267: out = 103;
			13268: out = 87;
			13269: out = 81;
			13270: out = 72;
			13271: out = 52;
			13272: out = 62;
			13273: out = 34;
			13274: out = 33;
			13275: out = 17;
			13276: out = 5;
			13277: out = 4;
			13278: out = -19;
			13279: out = -19;
			13280: out = -28;
			13281: out = -51;
			13282: out = -40;
			13283: out = -64;
			13284: out = -64;
			13285: out = -76;
			13286: out = -90;
			13287: out = -96;
			13288: out = -113;
			13289: out = -113;
			13290: out = -117;
			13291: out = -139;
			13292: out = -138;
			13293: out = -151;
			13294: out = -152;
			13295: out = -167;
			13296: out = -169;
			13297: out = -185;
			13298: out = -186;
			13299: out = -198;
			13300: out = -206;
			13301: out = -206;
			13302: out = -223;
			13303: out = -228;
			13304: out = -239;
			13305: out = -250;
			13306: out = -251;
			13307: out = -259;
			13308: out = -270;
			13309: out = -268;
			13310: out = -287;
			13311: out = -286;
			13312: out = -299;
			13313: out = -308;
			13314: out = -309;
			13315: out = -312;
			13316: out = -330;
			13317: out = -335;
			13318: out = -329;
			13319: out = -348;
			13320: out = -351;
			13321: out = -368;
			13322: out = -371;
			13323: out = -377;
			13324: out = -391;
			13325: out = -391;
			13326: out = -398;
			13327: out = -407;
			13328: out = -415;
			13329: out = -416;
			13330: out = -427;
			13331: out = -432;
			13332: out = -445;
			13333: out = -450;
			13334: out = -468;
			13335: out = -466;
			13336: out = -471;
			13337: out = -492;
			13338: out = -492;
			13339: out = -498;
			13340: out = -506;
			13341: out = -522;
			13342: out = -513;
			13343: out = -530;
			13344: out = -553;
			13345: out = -549;
			13346: out = -559;
			13347: out = -577;
			13348: out = -577;
			13349: out = -597;
			13350: out = -590;
			13351: out = -610;
			13352: out = -618;
			13353: out = -629;
			13354: out = -637;
			13355: out = -647;
			13356: out = -663;
			13357: out = -677;
			13358: out = -681;
			13359: out = -685;
			13360: out = -707;
			13361: out = -717;
			13362: out = -730;
			13363: out = -736;
			13364: out = -755;
			13365: out = -760;
			13366: out = -779;
			13367: out = -788;
			13368: out = -795;
			13369: out = -822;
			13370: out = -827;
			13371: out = -846;
			13372: out = -839;
			13373: out = -881;
			13374: out = -886;
			13375: out = -890;
			13376: out = -910;
			13377: out = -919;
			13378: out = -948;
			13379: out = -950;
			13380: out = -971;
			13381: out = -972;
			13382: out = -1003;
			13383: out = -1010;
			13384: out = -1035;
			13385: out = -1033;
			13386: out = -1058;
			13387: out = -1078;
			13388: out = -1085;
			13389: out = -1102;
			13390: out = -1102;
			13391: out = -1143;
			13392: out = -1134;
			13393: out = -1158;
			13394: out = -1175;
			13395: out = -1189;
			13396: out = -1197;
			13397: out = -1212;
			13398: out = -1238;
			13399: out = -1244;
			13400: out = -1245;
			13401: out = -1279;
			13402: out = -1273;
			13403: out = -1296;
			13404: out = -1306;
			13405: out = -1316;
			13406: out = -1341;
			13407: out = -1324;
			13408: out = -1358;
			13409: out = -1362;
			13410: out = -1377;
			13411: out = -1374;
			13412: out = -1395;
			13413: out = -1410;
			13414: out = -1414;
			13415: out = -1419;
			13416: out = -1438;
			13417: out = -1451;
			13418: out = -1450;
			13419: out = -1465;
			13420: out = -1463;
			13421: out = -1488;
			13422: out = -1478;
			13423: out = -1496;
			13424: out = -1504;
			13425: out = -1505;
			13426: out = -1519;
			13427: out = -1523;
			13428: out = -1532;
			13429: out = -1539;
			13430: out = -1541;
			13431: out = -1554;
			13432: out = -1551;
			13433: out = -1563;
			13434: out = -1571;
			13435: out = -1571;
			13436: out = -1577;
			13437: out = -1580;
			13438: out = -1594;
			13439: out = -1591;
			13440: out = -1592;
			13441: out = -1602;
			13442: out = -1602;
			13443: out = -1612;
			13444: out = -1608;
			13445: out = -1613;
			13446: out = -1626;
			13447: out = -1613;
			13448: out = -1630;
			13449: out = -1627;
			13450: out = -1624;
			13451: out = -1640;
			13452: out = -1638;
			13453: out = -1627;
			13454: out = -1637;
			13455: out = -1645;
			13456: out = -1637;
			13457: out = -1640;
			13458: out = -1650;
			13459: out = -1648;
			13460: out = -1643;
			13461: out = -1654;
			13462: out = -1648;
			13463: out = -1651;
			13464: out = -1654;
			13465: out = -1650;
			13466: out = -1654;
			13467: out = -1652;
			13468: out = -1647;
			13469: out = -1664;
			13470: out = -1651;
			13471: out = -1653;
			13472: out = -1648;
			13473: out = -1648;
			13474: out = -1650;
			13475: out = -1651;
			13476: out = -1653;
			13477: out = -1648;
			13478: out = -1652;
			13479: out = -1657;
			13480: out = -1650;
			13481: out = -1647;
			13482: out = -1642;
			13483: out = -1652;
			13484: out = -1637;
			13485: out = -1645;
			13486: out = -1645;
			13487: out = -1632;
			13488: out = -1638;
			13489: out = -1639;
			13490: out = -1634;
			13491: out = -1636;
			13492: out = -1624;
			13493: out = -1634;
			13494: out = -1632;
			13495: out = -1620;
			13496: out = -1615;
			13497: out = -1625;
			13498: out = -1611;
			13499: out = -1613;
			13500: out = -1618;
			13501: out = -1607;
			13502: out = -1607;
			13503: out = -1619;
			13504: out = -1603;
			13505: out = -1595;
			13506: out = -1592;
			13507: out = -1603;
			13508: out = -1590;
			13509: out = -1583;
			13510: out = -1592;
			13511: out = -1580;
			13512: out = -1574;
			13513: out = -1580;
			13514: out = -1569;
			13515: out = -1571;
			13516: out = -1567;
			13517: out = -1561;
			13518: out = -1558;
			13519: out = -1557;
			13520: out = -1560;
			13521: out = -1537;
			13522: out = -1549;
			13523: out = -1545;
			13524: out = -1535;
			13525: out = -1532;
			13526: out = -1528;
			13527: out = -1539;
			13528: out = -1513;
			13529: out = -1527;
			13530: out = -1513;
			13531: out = -1519;
			13532: out = -1504;
			13533: out = -1503;
			13534: out = -1500;
			13535: out = -1496;
			13536: out = -1486;
			13537: out = -1486;
			13538: out = -1486;
			13539: out = -1482;
			13540: out = -1469;
			13541: out = -1473;
			13542: out = -1462;
			13543: out = -1462;
			13544: out = -1454;
			13545: out = -1447;
			13546: out = -1449;
			13547: out = -1435;
			13548: out = -1437;
			13549: out = -1429;
			13550: out = -1425;
			13551: out = -1413;
			13552: out = -1415;
			13553: out = -1400;
			13554: out = -1400;
			13555: out = -1388;
			13556: out = -1391;
			13557: out = -1374;
			13558: out = -1381;
			13559: out = -1367;
			13560: out = -1354;
			13561: out = -1355;
			13562: out = -1331;
			13563: out = -1341;
			13564: out = -1329;
			13565: out = -1317;
			13566: out = -1315;
			13567: out = -1299;
			13568: out = -1298;
			13569: out = -1285;
			13570: out = -1279;
			13571: out = -1265;
			13572: out = -1263;
			13573: out = -1241;
			13574: out = -1246;
			13575: out = -1238;
			13576: out = -1216;
			13577: out = -1208;
			13578: out = -1208;
			13579: out = -1181;
			13580: out = -1182;
			13581: out = -1174;
			13582: out = -1152;
			13583: out = -1149;
			13584: out = -1143;
			13585: out = -1126;
			13586: out = -1114;
			13587: out = -1097;
			13588: out = -1099;
			13589: out = -1077;
			13590: out = -1071;
			13591: out = -1060;
			13592: out = -1046;
			13593: out = -1037;
			13594: out = -1019;
			13595: out = -1015;
			13596: out = -1003;
			13597: out = -989;
			13598: out = -983;
			13599: out = -965;
			13600: out = -962;
			13601: out = -940;
			13602: out = -933;
			13603: out = -930;
			13604: out = -904;
			13605: out = -903;
			13606: out = -881;
			13607: out = -882;
			13608: out = -868;
			13609: out = -858;
			13610: out = -853;
			13611: out = -833;
			13612: out = -819;
			13613: out = -820;
			13614: out = -810;
			13615: out = -788;
			13616: out = -778;
			13617: out = -771;
			13618: out = -763;
			13619: out = -754;
			13620: out = -743;
			13621: out = -728;
			13622: out = -719;
			13623: out = -714;
			13624: out = -695;
			13625: out = -699;
			13626: out = -677;
			13627: out = -677;
			13628: out = -665;
			13629: out = -655;
			13630: out = -648;
			13631: out = -628;
			13632: out = -634;
			13633: out = -617;
			13634: out = -604;
			13635: out = -604;
			13636: out = -595;
			13637: out = -582;
			13638: out = -574;
			13639: out = -572;
			13640: out = -555;
			13641: out = -545;
			13642: out = -540;
			13643: out = -539;
			13644: out = -517;
			13645: out = -526;
			13646: out = -514;
			13647: out = -495;
			13648: out = -499;
			13649: out = -487;
			13650: out = -480;
			13651: out = -476;
			13652: out = -454;
			13653: out = -458;
			13654: out = -448;
			13655: out = -446;
			13656: out = -438;
			13657: out = -421;
			13658: out = -424;
			13659: out = -415;
			13660: out = -421;
			13661: out = -398;
			13662: out = -400;
			13663: out = -395;
			13664: out = -386;
			13665: out = -377;
			13666: out = -365;
			13667: out = -375;
			13668: out = -351;
			13669: out = -354;
			13670: out = -351;
			13671: out = -342;
			13672: out = -334;
			13673: out = -339;
			13674: out = -318;
			13675: out = -332;
			13676: out = -304;
			13677: out = -317;
			13678: out = -303;
			13679: out = -291;
			13680: out = -281;
			13681: out = -279;
			13682: out = -264;
			13683: out = -249;
			13684: out = -247;
			13685: out = -240;
			13686: out = -231;
			13687: out = -217;
			13688: out = -209;
			13689: out = -208;
			13690: out = -200;
			13691: out = -186;
			13692: out = -178;
			13693: out = -164;
			13694: out = -171;
			13695: out = -147;
			13696: out = -146;
			13697: out = -145;
			13698: out = -134;
			13699: out = -119;
			13700: out = -114;
			13701: out = -112;
			13702: out = -109;
			13703: out = -95;
			13704: out = -89;
			13705: out = -80;
			13706: out = -86;
			13707: out = -69;
			13708: out = -56;
			13709: out = -54;
			13710: out = -52;
			13711: out = -39;
			13712: out = -42;
			13713: out = -32;
			13714: out = -17;
			13715: out = -27;
			13716: out = -10;
			13717: out = -5;
			13718: out = 0;
			13719: out = 7;
			13720: out = -5;
			13721: out = 26;
			13722: out = 24;
			13723: out = 25;
			13724: out = 27;
			13725: out = 49;
			13726: out = 38;
			13727: out = 53;
			13728: out = 57;
			13729: out = 58;
			13730: out = 70;
			13731: out = 72;
			13732: out = 74;
			13733: out = 86;
			13734: out = 89;
			13735: out = 95;
			13736: out = 100;
			13737: out = 99;
			13738: out = 116;
			13739: out = 117;
			13740: out = 113;
			13741: out = 123;
			13742: out = 134;
			13743: out = 136;
			13744: out = 139;
			13745: out = 141;
			13746: out = 170;
			13747: out = 147;
			13748: out = 164;
			13749: out = 172;
			13750: out = 176;
			13751: out = 172;
			13752: out = 194;
			13753: out = 184;
			13754: out = 200;
			13755: out = 195;
			13756: out = 206;
			13757: out = 211;
			13758: out = 218;
			13759: out = 222;
			13760: out = 230;
			13761: out = 239;
			13762: out = 238;
			13763: out = 254;
			13764: out = 257;
			13765: out = 255;
			13766: out = 271;
			13767: out = 279;
			13768: out = 264;
			13769: out = 300;
			13770: out = 288;
			13771: out = 312;
			13772: out = 306;
			13773: out = 314;
			13774: out = 328;
			13775: out = 325;
			13776: out = 348;
			13777: out = 345;
			13778: out = 353;
			13779: out = 367;
			13780: out = 375;
			13781: out = 375;
			13782: out = 389;
			13783: out = 399;
			13784: out = 410;
			13785: out = 410;
			13786: out = 423;
			13787: out = 438;
			13788: out = 442;
			13789: out = 450;
			13790: out = 454;
			13791: out = 479;
			13792: out = 472;
			13793: out = 489;
			13794: out = 504;
			13795: out = 510;
			13796: out = 517;
			13797: out = 529;
			13798: out = 543;
			13799: out = 549;
			13800: out = 557;
			13801: out = 563;
			13802: out = 583;
			13803: out = 589;
			13804: out = 595;
			13805: out = 610;
			13806: out = 620;
			13807: out = 634;
			13808: out = 640;
			13809: out = 643;
			13810: out = 663;
			13811: out = 673;
			13812: out = 680;
			13813: out = 693;
			13814: out = 695;
			13815: out = 707;
			13816: out = 726;
			13817: out = 717;
			13818: out = 744;
			13819: out = 748;
			13820: out = 752;
			13821: out = 770;
			13822: out = 773;
			13823: out = 790;
			13824: out = 786;
			13825: out = 799;
			13826: out = 814;
			13827: out = 820;
			13828: out = 819;
			13829: out = 839;
			13830: out = 847;
			13831: out = 857;
			13832: out = 860;
			13833: out = 862;
			13834: out = 882;
			13835: out = 885;
			13836: out = 890;
			13837: out = 901;
			13838: out = 915;
			13839: out = 905;
			13840: out = 938;
			13841: out = 929;
			13842: out = 938;
			13843: out = 948;
			13844: out = 959;
			13845: out = 953;
			13846: out = 967;
			13847: out = 975;
			13848: out = 976;
			13849: out = 1000;
			13850: out = 990;
			13851: out = 1000;
			13852: out = 1010;
			13853: out = 1023;
			13854: out = 1012;
			13855: out = 1033;
			13856: out = 1035;
			13857: out = 1040;
			13858: out = 1047;
			13859: out = 1056;
			13860: out = 1059;
			13861: out = 1062;
			13862: out = 1082;
			13863: out = 1069;
			13864: out = 1085;
			13865: out = 1090;
			13866: out = 1093;
			13867: out = 1105;
			13868: out = 1101;
			13869: out = 1119;
			13870: out = 1117;
			13871: out = 1121;
			13872: out = 1130;
			13873: out = 1130;
			13874: out = 1135;
			13875: out = 1149;
			13876: out = 1150;
			13877: out = 1151;
			13878: out = 1155;
			13879: out = 1177;
			13880: out = 1168;
			13881: out = 1172;
			13882: out = 1187;
			13883: out = 1179;
			13884: out = 1198;
			13885: out = 1188;
			13886: out = 1208;
			13887: out = 1202;
			13888: out = 1211;
			13889: out = 1211;
			13890: out = 1219;
			13891: out = 1226;
			13892: out = 1225;
			13893: out = 1237;
			13894: out = 1243;
			13895: out = 1237;
			13896: out = 1246;
			13897: out = 1252;
			13898: out = 1256;
			13899: out = 1263;
			13900: out = 1247;
			13901: out = 1271;
			13902: out = 1274;
			13903: out = 1272;
			13904: out = 1286;
			13905: out = 1280;
			13906: out = 1288;
			13907: out = 1298;
			13908: out = 1283;
			13909: out = 1305;
			13910: out = 1296;
			13911: out = 1298;
			13912: out = 1311;
			13913: out = 1300;
			13914: out = 1310;
			13915: out = 1306;
			13916: out = 1315;
			13917: out = 1300;
			13918: out = 1299;
			13919: out = 1308;
			13920: out = 1305;
			13921: out = 1308;
			13922: out = 1295;
			13923: out = 1304;
			13924: out = 1311;
			13925: out = 1300;
			13926: out = 1295;
			13927: out = 1294;
			13928: out = 1308;
			13929: out = 1300;
			13930: out = 1291;
			13931: out = 1287;
			13932: out = 1292;
			13933: out = 1283;
			13934: out = 1286;
			13935: out = 1292;
			13936: out = 1292;
			13937: out = 1280;
			13938: out = 1298;
			13939: out = 1288;
			13940: out = 1297;
			13941: out = 1282;
			13942: out = 1295;
			13943: out = 1293;
			13944: out = 1284;
			13945: out = 1295;
			13946: out = 1290;
			13947: out = 1270;
			13948: out = 1298;
			13949: out = 1279;
			13950: out = 1276;
			13951: out = 1288;
			13952: out = 1279;
			13953: out = 1288;
			13954: out = 1270;
			13955: out = 1283;
			13956: out = 1288;
			13957: out = 1281;
			13958: out = 1277;
			13959: out = 1279;
			13960: out = 1286;
			13961: out = 1281;
			13962: out = 1269;
			13963: out = 1281;
			13964: out = 1285;
			13965: out = 1270;
			13966: out = 1281;
			13967: out = 1282;
			13968: out = 1276;
			13969: out = 1279;
			13970: out = 1264;
			13971: out = 1268;
			13972: out = 1274;
			13973: out = 1272;
			13974: out = 1260;
			13975: out = 1268;
			13976: out = 1249;
			13977: out = 1274;
			13978: out = 1255;
			13979: out = 1260;
			13980: out = 1253;
			13981: out = 1270;
			13982: out = 1261;
			13983: out = 1253;
			13984: out = 1247;
			13985: out = 1255;
			13986: out = 1240;
			13987: out = 1229;
			13988: out = 1243;
			13989: out = 1231;
			13990: out = 1227;
			13991: out = 1228;
			13992: out = 1214;
			13993: out = 1213;
			13994: out = 1215;
			13995: out = 1208;
			13996: out = 1194;
			13997: out = 1206;
			13998: out = 1190;
			13999: out = 1191;
			14000: out = 1190;
			14001: out = 1168;
			14002: out = 1175;
			14003: out = 1167;
			14004: out = 1170;
			14005: out = 1138;
			14006: out = 1161;
			14007: out = 1142;
			14008: out = 1149;
			14009: out = 1128;
			14010: out = 1120;
			14011: out = 1118;
			14012: out = 1117;
			14013: out = 1101;
			14014: out = 1089;
			14015: out = 1085;
			14016: out = 1083;
			14017: out = 1069;
			14018: out = 1060;
			14019: out = 1054;
			14020: out = 1047;
			14021: out = 1035;
			14022: out = 1026;
			14023: out = 1018;
			14024: out = 1021;
			14025: out = 1000;
			14026: out = 998;
			14027: out = 992;
			14028: out = 974;
			14029: out = 978;
			14030: out = 957;
			14031: out = 953;
			14032: out = 945;
			14033: out = 936;
			14034: out = 936;
			14035: out = 915;
			14036: out = 912;
			14037: out = 908;
			14038: out = 901;
			14039: out = 885;
			14040: out = 880;
			14041: out = 868;
			14042: out = 862;
			14043: out = 850;
			14044: out = 838;
			14045: out = 843;
			14046: out = 815;
			14047: out = 817;
			14048: out = 818;
			14049: out = 807;
			14050: out = 789;
			14051: out = 780;
			14052: out = 772;
			14053: out = 766;
			14054: out = 758;
			14055: out = 746;
			14056: out = 728;
			14057: out = 739;
			14058: out = 727;
			14059: out = 723;
			14060: out = 702;
			14061: out = 707;
			14062: out = 701;
			14063: out = 678;
			14064: out = 681;
			14065: out = 677;
			14066: out = 654;
			14067: out = 665;
			14068: out = 642;
			14069: out = 641;
			14070: out = 631;
			14071: out = 623;
			14072: out = 618;
			14073: out = 611;
			14074: out = 598;
			14075: out = 592;
			14076: out = 597;
			14077: out = 575;
			14078: out = 572;
			14079: out = 566;
			14080: out = 560;
			14081: out = 549;
			14082: out = 541;
			14083: out = 541;
			14084: out = 533;
			14085: out = 517;
			14086: out = 518;
			14087: out = 507;
			14088: out = 504;
			14089: out = 499;
			14090: out = 496;
			14091: out = 482;
			14092: out = 479;
			14093: out = 474;
			14094: out = 455;
			14095: out = 464;
			14096: out = 442;
			14097: out = 442;
			14098: out = 444;
			14099: out = 430;
			14100: out = 430;
			14101: out = 434;
			14102: out = 422;
			14103: out = 407;
			14104: out = 410;
			14105: out = 405;
			14106: out = 389;
			14107: out = 391;
			14108: out = 375;
			14109: out = 376;
			14110: out = 373;
			14111: out = 360;
			14112: out = 358;
			14113: out = 357;
			14114: out = 359;
			14115: out = 337;
			14116: out = 340;
			14117: out = 332;
			14118: out = 328;
			14119: out = 323;
			14120: out = 318;
			14121: out = 306;
			14122: out = 309;
			14123: out = 305;
			14124: out = 303;
			14125: out = 296;
			14126: out = 289;
			14127: out = 275;
			14128: out = 287;
			14129: out = 276;
			14130: out = 259;
			14131: out = 267;
			14132: out = 267;
			14133: out = 259;
			14134: out = 252;
			14135: out = 252;
			14136: out = 245;
			14137: out = 244;
			14138: out = 234;
			14139: out = 233;
			14140: out = 228;
			14141: out = 227;
			14142: out = 223;
			14143: out = 219;
			14144: out = 208;
			14145: out = 205;
			14146: out = 191;
			14147: out = 178;
			14148: out = 174;
			14149: out = 160;
			14150: out = 149;
			14151: out = 143;
			14152: out = 128;
			14153: out = 119;
			14154: out = 110;
			14155: out = 102;
			14156: out = 88;
			14157: out = 91;
			14158: out = 65;
			14159: out = 76;
			14160: out = 46;
			14161: out = 53;
			14162: out = 30;
			14163: out = 38;
			14164: out = 17;
			14165: out = 17;
			14166: out = 7;
			14167: out = -2;
			14168: out = -13;
			14169: out = -19;
			14170: out = -24;
			14171: out = -40;
			14172: out = -41;
			14173: out = -51;
			14174: out = -51;
			14175: out = -66;
			14176: out = -72;
			14177: out = -74;
			14178: out = -87;
			14179: out = -95;
			14180: out = -93;
			14181: out = -109;
			14182: out = -115;
			14183: out = -127;
			14184: out = -126;
			14185: out = -136;
			14186: out = -137;
			14187: out = -138;
			14188: out = -166;
			14189: out = -152;
			14190: out = -162;
			14191: out = -172;
			14192: out = -174;
			14193: out = -195;
			14194: out = -192;
			14195: out = -202;
			14196: out = -206;
			14197: out = -206;
			14198: out = -219;
			14199: out = -221;
			14200: out = -227;
			14201: out = -228;
			14202: out = -252;
			14203: out = -249;
			14204: out = -252;
			14205: out = -279;
			14206: out = -259;
			14207: out = -269;
			14208: out = -280;
			14209: out = -276;
			14210: out = -292;
			14211: out = -294;
			14212: out = -304;
			14213: out = -299;
			14214: out = -320;
			14215: out = -308;
			14216: out = -334;
			14217: out = -327;
			14218: out = -327;
			14219: out = -352;
			14220: out = -341;
			14221: out = -353;
			14222: out = -364;
			14223: out = -368;
			14224: out = -373;
			14225: out = -380;
			14226: out = -384;
			14227: out = -388;
			14228: out = -410;
			14229: out = -398;
			14230: out = -418;
			14231: out = -422;
			14232: out = -420;
			14233: out = -443;
			14234: out = -441;
			14235: out = -446;
			14236: out = -453;
			14237: out = -464;
			14238: out = -467;
			14239: out = -480;
			14240: out = -480;
			14241: out = -492;
			14242: out = -507;
			14243: out = -511;
			14244: out = -509;
			14245: out = -528;
			14246: out = -538;
			14247: out = -536;
			14248: out = -552;
			14249: out = -564;
			14250: out = -558;
			14251: out = -585;
			14252: out = -585;
			14253: out = -606;
			14254: out = -602;
			14255: out = -607;
			14256: out = -632;
			14257: out = -643;
			14258: out = -642;
			14259: out = -652;
			14260: out = -671;
			14261: out = -669;
			14262: out = -691;
			14263: out = -695;
			14264: out = -717;
			14265: out = -716;
			14266: out = -728;
			14267: out = -752;
			14268: out = -761;
			14269: out = -763;
			14270: out = -782;
			14271: out = -790;
			14272: out = -814;
			14273: out = -806;
			14274: out = -829;
			14275: out = -834;
			14276: out = -856;
			14277: out = -870;
			14278: out = -871;
			14279: out = -888;
			14280: out = -902;
			14281: out = -910;
			14282: out = -929;
			14283: out = -926;
			14284: out = -952;
			14285: out = -955;
			14286: out = -964;
			14287: out = -976;
			14288: out = -991;
			14289: out = -988;
			14290: out = -1013;
			14291: out = -1014;
			14292: out = -1038;
			14293: out = -1046;
			14294: out = -1054;
			14295: out = -1063;
			14296: out = -1074;
			14297: out = -1081;
			14298: out = -1086;
			14299: out = -1105;
			14300: out = -1105;
			14301: out = -1120;
			14302: out = -1125;
			14303: out = -1135;
			14304: out = -1146;
			14305: out = -1150;
			14306: out = -1156;
			14307: out = -1165;
			14308: out = -1177;
			14309: out = -1184;
			14310: out = -1181;
			14311: out = -1192;
			14312: out = -1197;
			14313: out = -1213;
			14314: out = -1204;
			14315: out = -1221;
			14316: out = -1227;
			14317: out = -1229;
			14318: out = -1236;
			14319: out = -1245;
			14320: out = -1241;
			14321: out = -1256;
			14322: out = -1258;
			14323: out = -1260;
			14324: out = -1261;
			14325: out = -1273;
			14326: out = -1275;
			14327: out = -1280;
			14328: out = -1270;
			14329: out = -1288;
			14330: out = -1293;
			14331: out = -1292;
			14332: out = -1288;
			14333: out = -1298;
			14334: out = -1309;
			14335: out = -1302;
			14336: out = -1304;
			14337: out = -1315;
			14338: out = -1311;
			14339: out = -1315;
			14340: out = -1316;
			14341: out = -1328;
			14342: out = -1307;
			14343: out = -1332;
			14344: out = -1331;
			14345: out = -1320;
			14346: out = -1331;
			14347: out = -1323;
			14348: out = -1341;
			14349: out = -1328;
			14350: out = -1338;
			14351: out = -1330;
			14352: out = -1336;
			14353: out = -1338;
			14354: out = -1331;
			14355: out = -1333;
			14356: out = -1342;
			14357: out = -1335;
			14358: out = -1329;
			14359: out = -1341;
			14360: out = -1343;
			14361: out = -1327;
			14362: out = -1336;
			14363: out = -1345;
			14364: out = -1329;
			14365: out = -1334;
			14366: out = -1340;
			14367: out = -1336;
			14368: out = -1331;
			14369: out = -1329;
			14370: out = -1341;
			14371: out = -1321;
			14372: out = -1327;
			14373: out = -1329;
			14374: out = -1333;
			14375: out = -1329;
			14376: out = -1320;
			14377: out = -1324;
			14378: out = -1322;
			14379: out = -1319;
			14380: out = -1319;
			14381: out = -1323;
			14382: out = -1310;
			14383: out = -1322;
			14384: out = -1321;
			14385: out = -1310;
			14386: out = -1316;
			14387: out = -1312;
			14388: out = -1308;
			14389: out = -1309;
			14390: out = -1299;
			14391: out = -1300;
			14392: out = -1303;
			14393: out = -1297;
			14394: out = -1300;
			14395: out = -1288;
			14396: out = -1294;
			14397: out = -1295;
			14398: out = -1284;
			14399: out = -1291;
			14400: out = -1271;
			14401: out = -1291;
			14402: out = -1277;
			14403: out = -1280;
			14404: out = -1263;
			14405: out = -1272;
			14406: out = -1269;
			14407: out = -1270;
			14408: out = -1255;
			14409: out = -1256;
			14410: out = -1263;
			14411: out = -1256;
			14412: out = -1247;
			14413: out = -1247;
			14414: out = -1259;
			14415: out = -1237;
			14416: out = -1239;
			14417: out = -1250;
			14418: out = -1232;
			14419: out = -1237;
			14420: out = -1226;
			14421: out = -1235;
			14422: out = -1221;
			14423: out = -1216;
			14424: out = -1219;
			14425: out = -1216;
			14426: out = -1208;
			14427: out = -1202;
			14428: out = -1201;
			14429: out = -1196;
			14430: out = -1202;
			14431: out = -1191;
			14432: out = -1179;
			14433: out = -1190;
			14434: out = -1180;
			14435: out = -1168;
			14436: out = -1166;
			14437: out = -1175;
			14438: out = -1164;
			14439: out = -1154;
			14440: out = -1157;
			14441: out = -1154;
			14442: out = -1138;
			14443: out = -1139;
			14444: out = -1137;
			14445: out = -1135;
			14446: out = -1121;
			14447: out = -1122;
			14448: out = -1118;
			14449: out = -1113;
			14450: out = -1108;
			14451: out = -1101;
			14452: out = -1086;
			14453: out = -1097;
			14454: out = -1077;
			14455: out = -1069;
			14456: out = -1074;
			14457: out = -1059;
			14458: out = -1054;
			14459: out = -1049;
			14460: out = -1044;
			14461: out = -1036;
			14462: out = -1025;
			14463: out = -1025;
			14464: out = -1011;
			14465: out = -1004;
			14466: out = -1009;
			14467: out = -985;
			14468: out = -983;
			14469: out = -975;
			14470: out = -959;
			14471: out = -957;
			14472: out = -952;
			14473: out = -936;
			14474: out = -926;
			14475: out = -922;
			14476: out = -919;
			14477: out = -895;
			14478: out = -894;
			14479: out = -882;
			14480: out = -876;
			14481: out = -856;
			14482: out = -861;
			14483: out = -847;
			14484: out = -839;
			14485: out = -834;
			14486: out = -810;
			14487: out = -825;
			14488: out = -802;
			14489: out = -790;
			14490: out = -784;
			14491: out = -771;
			14492: out = -767;
			14493: out = -754;
			14494: out = -742;
			14495: out = -740;
			14496: out = -728;
			14497: out = -722;
			14498: out = -713;
			14499: out = -697;
			14500: out = -704;
			14501: out = -680;
			14502: out = -679;
			14503: out = -663;
			14504: out = -667;
			14505: out = -644;
			14506: out = -648;
			14507: out = -625;
			14508: out = -635;
			14509: out = -611;
			14510: out = -610;
			14511: out = -600;
			14512: out = -598;
			14513: out = -578;
			14514: out = -583;
			14515: out = -576;
			14516: out = -546;
			14517: out = -559;
			14518: out = -550;
			14519: out = -538;
			14520: out = -528;
			14521: out = -528;
			14522: out = -506;
			14523: out = -514;
			14524: out = -504;
			14525: out = -490;
			14526: out = -487;
			14527: out = -480;
			14528: out = -472;
			14529: out = -463;
			14530: out = -456;
			14531: out = -460;
			14532: out = -438;
			14533: out = -433;
			14534: out = -444;
			14535: out = -427;
			14536: out = -412;
			14537: out = -416;
			14538: out = -417;
			14539: out = -392;
			14540: out = -398;
			14541: out = -392;
			14542: out = -382;
			14543: out = -381;
			14544: out = -371;
			14545: out = -362;
			14546: out = -368;
			14547: out = -357;
			14548: out = -342;
			14549: out = -354;
			14550: out = -338;
			14551: out = -323;
			14552: out = -335;
			14553: out = -313;
			14554: out = -325;
			14555: out = -310;
			14556: out = -305;
			14557: out = -308;
			14558: out = -301;
			14559: out = -297;
			14560: out = -281;
			14561: out = -290;
			14562: out = -276;
			14563: out = -277;
			14564: out = -273;
			14565: out = -271;
			14566: out = -254;
			14567: out = -254;
			14568: out = -253;
			14569: out = -247;
			14570: out = -234;
			14571: out = -232;
			14572: out = -223;
			14573: out = -226;
			14574: out = -208;
			14575: out = -195;
			14576: out = -207;
			14577: out = -173;
			14578: out = -191;
			14579: out = -170;
			14580: out = -169;
			14581: out = -160;
			14582: out = -159;
			14583: out = -141;
			14584: out = -144;
			14585: out = -135;
			14586: out = -132;
			14587: out = -124;
			14588: out = -114;
			14589: out = -111;
			14590: out = -101;
			14591: out = -102;
			14592: out = -95;
			14593: out = -84;
			14594: out = -87;
			14595: out = -79;
			14596: out = -69;
			14597: out = -70;
			14598: out = -55;
			14599: out = -57;
			14600: out = -45;
			14601: out = -43;
			14602: out = -45;
			14603: out = -29;
			14604: out = -36;
			14605: out = -20;
			14606: out = -20;
			14607: out = -17;
			14608: out = -10;
			14609: out = -12;
			14610: out = 1;
			14611: out = 7;
			14612: out = -4;
			14613: out = 20;
			14614: out = 9;
			14615: out = 21;
			14616: out = 27;
			14617: out = 27;
			14618: out = 37;
			14619: out = 36;
			14620: out = 38;
			14621: out = 42;
			14622: out = 60;
			14623: out = 52;
			14624: out = 61;
			14625: out = 68;
			14626: out = 67;
			14627: out = 64;
			14628: out = 87;
			14629: out = 76;
			14630: out = 84;
			14631: out = 91;
			14632: out = 85;
			14633: out = 97;
			14634: out = 107;
			14635: out = 100;
			14636: out = 101;
			14637: out = 124;
			14638: out = 110;
			14639: out = 133;
			14640: out = 128;
			14641: out = 114;
			14642: out = 143;
			14643: out = 138;
			14644: out = 147;
			14645: out = 146;
			14646: out = 150;
			14647: out = 154;
			14648: out = 172;
			14649: out = 166;
			14650: out = 158;
			14651: out = 172;
			14652: out = 182;
			14653: out = 188;
			14654: out = 184;
			14655: out = 195;
			14656: out = 194;
			14657: out = 220;
			14658: out = 202;
			14659: out = 220;
			14660: out = 218;
			14661: out = 231;
			14662: out = 222;
			14663: out = 240;
			14664: out = 247;
			14665: out = 242;
			14666: out = 257;
			14667: out = 259;
			14668: out = 264;
			14669: out = 279;
			14670: out = 273;
			14671: out = 286;
			14672: out = 289;
			14673: out = 297;
			14674: out = 308;
			14675: out = 310;
			14676: out = 321;
			14677: out = 325;
			14678: out = 340;
			14679: out = 342;
			14680: out = 346;
			14681: out = 358;
			14682: out = 358;
			14683: out = 367;
			14684: out = 391;
			14685: out = 384;
			14686: out = 393;
			14687: out = 405;
			14688: out = 418;
			14689: out = 419;
			14690: out = 429;
			14691: out = 440;
			14692: out = 440;
			14693: out = 454;
			14694: out = 463;
			14695: out = 466;
			14696: out = 469;
			14697: out = 495;
			14698: out = 487;
			14699: out = 507;
			14700: out = 510;
			14701: out = 519;
			14702: out = 525;
			14703: out = 543;
			14704: out = 536;
			14705: out = 552;
			14706: out = 555;
			14707: out = 566;
			14708: out = 566;
			14709: out = 584;
			14710: out = 584;
			14711: out = 594;
			14712: out = 610;
			14713: out = 604;
			14714: out = 628;
			14715: out = 624;
			14716: out = 625;
			14717: out = 642;
			14718: out = 647;
			14719: out = 655;
			14720: out = 661;
			14721: out = 661;
			14722: out = 677;
			14723: out = 682;
			14724: out = 681;
			14725: out = 691;
			14726: out = 700;
			14727: out = 708;
			14728: out = 716;
			14729: out = 719;
			14730: out = 719;
			14731: out = 730;
			14732: out = 740;
			14733: out = 750;
			14734: out = 739;
			14735: out = 754;
			14736: out = 771;
			14737: out = 771;
			14738: out = 771;
			14739: out = 776;
			14740: out = 787;
			14741: out = 796;
			14742: out = 785;
			14743: out = 801;
			14744: out = 806;
			14745: out = 806;
			14746: out = 818;
			14747: out = 818;
			14748: out = 829;
			14749: out = 822;
			14750: out = 847;
			14751: out = 830;
			14752: out = 849;
			14753: out = 842;
			14754: out = 851;
			14755: out = 862;
			14756: out = 855;
			14757: out = 870;
			14758: out = 866;
			14759: out = 884;
			14760: out = 878;
			14761: out = 890;
			14762: out = 886;
			14763: out = 896;
			14764: out = 897;
			14765: out = 898;
			14766: out = 908;
			14767: out = 910;
			14768: out = 913;
			14769: out = 922;
			14770: out = 918;
			14771: out = 931;
			14772: out = 925;
			14773: out = 942;
			14774: out = 935;
			14775: out = 945;
			14776: out = 944;
			14777: out = 961;
			14778: out = 941;
			14779: out = 966;
			14780: out = 964;
			14781: out = 956;
			14782: out = 968;
			14783: out = 972;
			14784: out = 973;
			14785: out = 978;
			14786: out = 983;
			14787: out = 996;
			14788: out = 984;
			14789: out = 995;
			14790: out = 999;
			14791: out = 1003;
			14792: out = 995;
			14793: out = 1016;
			14794: out = 1013;
			14795: out = 1010;
			14796: out = 1020;
			14797: out = 1030;
			14798: out = 1019;
			14799: out = 1025;
			14800: out = 1039;
			14801: out = 1033;
			14802: out = 1038;
			14803: out = 1036;
			14804: out = 1038;
			14805: out = 1032;
			14806: out = 1051;
			14807: out = 1035;
			14808: out = 1045;
			14809: out = 1035;
			14810: out = 1046;
			14811: out = 1032;
			14812: out = 1038;
			14813: out = 1047;
			14814: out = 1032;
			14815: out = 1036;
			14816: out = 1040;
			14817: out = 1039;
			14818: out = 1028;
			14819: out = 1035;
			14820: out = 1035;
			14821: out = 1024;
			14822: out = 1031;
			14823: out = 1031;
			14824: out = 1035;
			14825: out = 1024;
			14826: out = 1023;
			14827: out = 1027;
			14828: out = 1018;
			14829: out = 1030;
			14830: out = 1021;
			14831: out = 1016;
			14832: out = 1031;
			14833: out = 1035;
			14834: out = 1012;
			14835: out = 1034;
			14836: out = 1019;
			14837: out = 1036;
			14838: out = 1014;
			14839: out = 1022;
			14840: out = 1032;
			14841: out = 1016;
			14842: out = 1020;
			14843: out = 1036;
			14844: out = 1018;
			14845: out = 1025;
			14846: out = 1030;
			14847: out = 1027;
			14848: out = 1023;
			14849: out = 1024;
			14850: out = 1020;
			14851: out = 1019;
			14852: out = 1026;
			14853: out = 1015;
			14854: out = 1007;
			14855: out = 1016;
			14856: out = 1015;
			14857: out = 1010;
			14858: out = 1012;
			14859: out = 1016;
			14860: out = 1022;
			14861: out = 1009;
			14862: out = 1015;
			14863: out = 1016;
			14864: out = 1007;
			14865: out = 1002;
			14866: out = 1006;
			14867: out = 999;
			14868: out = 1002;
			14869: out = 1003;
			14870: out = 1001;
			14871: out = 1011;
			14872: out = 1002;
			14873: out = 1004;
			14874: out = 998;
			14875: out = 999;
			14876: out = 989;
			14877: out = 992;
			14878: out = 978;
			14879: out = 981;
			14880: out = 987;
			14881: out = 978;
			14882: out = 978;
			14883: out = 975;
			14884: out = 979;
			14885: out = 955;
			14886: out = 952;
			14887: out = 971;
			14888: out = 950;
			14889: out = 947;
			14890: out = 948;
			14891: out = 937;
			14892: out = 947;
			14893: out = 926;
			14894: out = 930;
			14895: out = 922;
			14896: out = 927;
			14897: out = 925;
			14898: out = 914;
			14899: out = 906;
			14900: out = 904;
			14901: out = 897;
			14902: out = 874;
			14903: out = 888;
			14904: out = 878;
			14905: out = 860;
			14906: out = 866;
			14907: out = 862;
			14908: out = 850;
			14909: out = 844;
			14910: out = 850;
			14911: out = 824;
			14912: out = 831;
			14913: out = 822;
			14914: out = 800;
			14915: out = 805;
			14916: out = 796;
			14917: out = 786;
			14918: out = 790;
			14919: out = 784;
			14920: out = 774;
			14921: out = 776;
			14922: out = 754;
			14923: out = 756;
			14924: out = 744;
			14925: out = 736;
			14926: out = 735;
			14927: out = 720;
			14928: out = 720;
			14929: out = 715;
			14930: out = 709;
			14931: out = 695;
			14932: out = 699;
			14933: out = 685;
			14934: out = 676;
			14935: out = 665;
			14936: out = 655;
			14937: out = 665;
			14938: out = 634;
			14939: out = 646;
			14940: out = 630;
			14941: out = 634;
			14942: out = 622;
			14943: out = 606;
			14944: out = 614;
			14945: out = 602;
			14946: out = 586;
			14947: out = 592;
			14948: out = 576;
			14949: out = 576;
			14950: out = 575;
			14951: out = 554;
			14952: out = 550;
			14953: out = 558;
			14954: out = 534;
			14955: out = 534;
			14956: out = 537;
			14957: out = 518;
			14958: out = 516;
			14959: out = 514;
			14960: out = 502;
			14961: out = 492;
			14962: out = 492;
			14963: out = 493;
			14964: out = 456;
			14965: out = 488;
			14966: out = 454;
			14967: out = 466;
			14968: out = 459;
			14969: out = 439;
			14970: out = 453;
			14971: out = 436;
			14972: out = 434;
			14973: out = 428;
			14974: out = 422;
			14975: out = 421;
			14976: out = 412;
			14977: out = 389;
			14978: out = 412;
			14979: out = 392;
			14980: out = 379;
			14981: out = 384;
			14982: out = 385;
			14983: out = 371;
			14984: out = 363;
			14985: out = 367;
			14986: out = 357;
			14987: out = 350;
			14988: out = 349;
			14989: out = 332;
			14990: out = 346;
			14991: out = 327;
			14992: out = 330;
			14993: out = 327;
			14994: out = 311;
			14995: out = 313;
			14996: out = 316;
			14997: out = 306;
			14998: out = 306;
			14999: out = 306;
			15000: out = 289;
			15001: out = 292;
			15002: out = 281;
			15003: out = 278;
			15004: out = 269;
			15005: out = 270;
			15006: out = 262;
			15007: out = 264;
			15008: out = 259;
			15009: out = 247;
			15010: out = 259;
			15011: out = 241;
			15012: out = 242;
			15013: out = 233;
			15014: out = 230;
			15015: out = 243;
			15016: out = 219;
			15017: out = 226;
			15018: out = 223;
			15019: out = 222;
			15020: out = 210;
			15021: out = 210;
			15022: out = 216;
			15023: out = 193;
			15024: out = 198;
			15025: out = 196;
			15026: out = 197;
			15027: out = 183;
			15028: out = 186;
			15029: out = 188;
			15030: out = 180;
			15031: out = 182;
			15032: out = 167;
			15033: out = 171;
			15034: out = 169;
			15035: out = 155;
			15036: out = 157;
			15037: out = 154;
			15038: out = 144;
			15039: out = 125;
			15040: out = 128;
			15041: out = 117;
			15042: out = 97;
			15043: out = 102;
			15044: out = 88;
			15045: out = 84;
			15046: out = 64;
			15047: out = 75;
			15048: out = 63;
			15049: out = 39;
			15050: out = 49;
			15051: out = 38;
			15052: out = 38;
			15053: out = 16;
			15054: out = 24;
			15055: out = 1;
			15056: out = 9;
			15057: out = -4;
			15058: out = -7;
			15059: out = -19;
			15060: out = -18;
			15061: out = -20;
			15062: out = -49;
			15063: out = -29;
			15064: out = -57;
			15065: out = -43;
			15066: out = -61;
			15067: out = -60;
			15068: out = -65;
			15069: out = -80;
			15070: out = -76;
			15071: out = -85;
			15072: out = -99;
			15073: out = -97;
			15074: out = -101;
			15075: out = -110;
			15076: out = -115;
			15077: out = -124;
			15078: out = -120;
			15079: out = -125;
			15080: out = -140;
			15081: out = -146;
			15082: out = -140;
			15083: out = -150;
			15084: out = -162;
			15085: out = -159;
			15086: out = -159;
			15087: out = -173;
			15088: out = -174;
			15089: out = -181;
			15090: out = -185;
			15091: out = -193;
			15092: out = -206;
			15093: out = -193;
			15094: out = -207;
			15095: out = -211;
			15096: out = -209;
			15097: out = -222;
			15098: out = -212;
			15099: out = -240;
			15100: out = -238;
			15101: out = -234;
			15102: out = -244;
			15103: out = -253;
			15104: out = -239;
			15105: out = -264;
			15106: out = -259;
			15107: out = -267;
			15108: out = -269;
			15109: out = -277;
			15110: out = -285;
			15111: out = -288;
			15112: out = -291;
			15113: out = -296;
			15114: out = -300;
			15115: out = -314;
			15116: out = -305;
			15117: out = -322;
			15118: out = -316;
			15119: out = -335;
			15120: out = -327;
			15121: out = -350;
			15122: out = -336;
			15123: out = -352;
			15124: out = -356;
			15125: out = -361;
			15126: out = -371;
			15127: out = -372;
			15128: out = -380;
			15129: out = -382;
			15130: out = -388;
			15131: out = -392;
			15132: out = -410;
			15133: out = -403;
			15134: out = -418;
			15135: out = -429;
			15136: out = -424;
			15137: out = -433;
			15138: out = -440;
			15139: out = -452;
			15140: out = -447;
			15141: out = -470;
			15142: out = -468;
			15143: out = -472;
			15144: out = -492;
			15145: out = -494;
			15146: out = -496;
			15147: out = -503;
			15148: out = -516;
			15149: out = -535;
			15150: out = -526;
			15151: out = -548;
			15152: out = -547;
			15153: out = -558;
			15154: out = -573;
			15155: out = -580;
			15156: out = -583;
			15157: out = -596;
			15158: out = -607;
			15159: out = -614;
			15160: out = -621;
			15161: out = -632;
			15162: out = -640;
			15163: out = -648;
			15164: out = -673;
			15165: out = -663;
			15166: out = -680;
			15167: out = -683;
			15168: out = -701;
			15169: out = -705;
			15170: out = -719;
			15171: out = -717;
			15172: out = -752;
			15173: out = -735;
			15174: out = -749;
			15175: out = -771;
			15176: out = -770;
			15177: out = -767;
			15178: out = -791;
			15179: out = -798;
			15180: out = -805;
			15181: out = -814;
			15182: out = -825;
			15183: out = -833;
			15184: out = -838;
			15185: out = -850;
			15186: out = -846;
			15187: out = -867;
			15188: out = -866;
			15189: out = -873;
			15190: out = -889;
			15191: out = -896;
			15192: out = -896;
			15193: out = -906;
			15194: out = -913;
			15195: out = -922;
			15196: out = -927;
			15197: out = -928;
			15198: out = -943;
			15199: out = -943;
			15200: out = -948;
			15201: out = -951;
			15202: out = -966;
			15203: out = -957;
			15204: out = -969;
			15205: out = -981;
			15206: out = -975;
			15207: out = -989;
			15208: out = -995;
			15209: out = -989;
			15210: out = -998;
			15211: out = -998;
			15212: out = -1016;
			15213: out = -1004;
			15214: out = -1015;
			15215: out = -1020;
			15216: out = -1010;
			15217: out = -1036;
			15218: out = -1024;
			15219: out = -1026;
			15220: out = -1044;
			15221: out = -1028;
			15222: out = -1046;
			15223: out = -1040;
			15224: out = -1040;
			15225: out = -1055;
			15226: out = -1046;
			15227: out = -1056;
			15228: out = -1050;
			15229: out = -1055;
			15230: out = -1057;
			15231: out = -1062;
			15232: out = -1056;
			15233: out = -1062;
			15234: out = -1067;
			15235: out = -1060;
			15236: out = -1072;
			15237: out = -1073;
			15238: out = -1063;
			15239: out = -1067;
			15240: out = -1075;
			15241: out = -1067;
			15242: out = -1074;
			15243: out = -1073;
			15244: out = -1075;
			15245: out = -1067;
			15246: out = -1091;
			15247: out = -1066;
			15248: out = -1074;
			15249: out = -1075;
			15250: out = -1071;
			15251: out = -1074;
			15252: out = -1077;
			15253: out = -1075;
			15254: out = -1071;
			15255: out = -1063;
			15256: out = -1072;
			15257: out = -1079;
			15258: out = -1078;
			15259: out = -1066;
			15260: out = -1083;
			15261: out = -1066;
			15262: out = -1073;
			15263: out = -1074;
			15264: out = -1067;
			15265: out = -1070;
			15266: out = -1066;
			15267: out = -1066;
			15268: out = -1066;
			15269: out = -1061;
			15270: out = -1062;
			15271: out = -1061;
			15272: out = -1063;
			15273: out = -1055;
			15274: out = -1063;
			15275: out = -1059;
			15276: out = -1061;
			15277: out = -1058;
			15278: out = -1058;
			15279: out = -1055;
			15280: out = -1044;
			15281: out = -1064;
			15282: out = -1043;
			15283: out = -1052;
			15284: out = -1045;
			15285: out = -1042;
			15286: out = -1049;
			15287: out = -1046;
			15288: out = -1033;
			15289: out = -1044;
			15290: out = -1031;
			15291: out = -1034;
			15292: out = -1032;
			15293: out = -1030;
			15294: out = -1025;
			15295: out = -1022;
			15296: out = -1019;
			15297: out = -1028;
			15298: out = -1016;
			15299: out = -1018;
			15300: out = -1019;
			15301: out = -1012;
			15302: out = -1011;
			15303: out = -1007;
			15304: out = -1013;
			15305: out = -1002;
			15306: out = -1000;
			15307: out = -1008;
			15308: out = -996;
			15309: out = -992;
			15310: out = -995;
			15311: out = -988;
			15312: out = -991;
			15313: out = -987;
			15314: out = -990;
			15315: out = -966;
			15316: out = -979;
			15317: out = -979;
			15318: out = -973;
			15319: out = -962;
			15320: out = -974;
			15321: out = -953;
			15322: out = -964;
			15323: out = -957;
			15324: out = -944;
			15325: out = -959;
			15326: out = -940;
			15327: out = -945;
			15328: out = -945;
			15329: out = -931;
			15330: out = -938;
			15331: out = -929;
			15332: out = -930;
			15333: out = -916;
			15334: out = -929;
			15335: out = -910;
			15336: out = -913;
			15337: out = -904;
			15338: out = -897;
			15339: out = -909;
			15340: out = -898;
			15341: out = -882;
			15342: out = -888;
			15343: out = -881;
			15344: out = -881;
			15345: out = -859;
			15346: out = -866;
			15347: out = -870;
			15348: out = -851;
			15349: out = -858;
			15350: out = -853;
			15351: out = -838;
			15352: out = -836;
			15353: out = -824;
			15354: out = -824;
			15355: out = -821;
			15356: out = -801;
			15357: out = -803;
			15358: out = -803;
			15359: out = -789;
			15360: out = -779;
			15361: out = -783;
			15362: out = -772;
			15363: out = -764;
			15364: out = -763;
			15365: out = -752;
			15366: out = -734;
			15367: out = -752;
			15368: out = -720;
			15369: out = -728;
			15370: out = -714;
			15371: out = -704;
			15372: out = -711;
			15373: out = -694;
			15374: out = -681;
			15375: out = -675;
			15376: out = -675;
			15377: out = -660;
			15378: out = -658;
			15379: out = -651;
			15380: out = -647;
			15381: out = -633;
			15382: out = -635;
			15383: out = -624;
			15384: out = -612;
			15385: out = -610;
			15386: out = -595;
			15387: out = -597;
			15388: out = -588;
			15389: out = -575;
			15390: out = -571;
			15391: out = -567;
			15392: out = -562;
			15393: out = -551;
			15394: out = -548;
			15395: out = -531;
			15396: out = -531;
			15397: out = -529;
			15398: out = -513;
			15399: out = -511;
			15400: out = -499;
			15401: out = -500;
			15402: out = -494;
			15403: out = -483;
			15404: out = -472;
			15405: out = -477;
			15406: out = -463;
			15407: out = -458;
			15408: out = -448;
			15409: out = -455;
			15410: out = -441;
			15411: out = -439;
			15412: out = -434;
			15413: out = -421;
			15414: out = -423;
			15415: out = -411;
			15416: out = -411;
			15417: out = -401;
			15418: out = -397;
			15419: out = -384;
			15420: out = -386;
			15421: out = -392;
			15422: out = -367;
			15423: out = -369;
			15424: out = -357;
			15425: out = -362;
			15426: out = -361;
			15427: out = -347;
			15428: out = -339;
			15429: out = -340;
			15430: out = -338;
			15431: out = -329;
			15432: out = -322;
			15433: out = -317;
			15434: out = -312;
			15435: out = -309;
			15436: out = -298;
			15437: out = -301;
			15438: out = -302;
			15439: out = -289;
			15440: out = -286;
			15441: out = -290;
			15442: out = -282;
			15443: out = -273;
			15444: out = -270;
			15445: out = -271;
			15446: out = -258;
			15447: out = -255;
			15448: out = -257;
			15449: out = -249;
			15450: out = -242;
			15451: out = -256;
			15452: out = -234;
			15453: out = -237;
			15454: out = -238;
			15455: out = -230;
			15456: out = -222;
			15457: out = -220;
			15458: out = -218;
			15459: out = -204;
			15460: out = -209;
			15461: out = -198;
			15462: out = -204;
			15463: out = -176;
			15464: out = -190;
			15465: out = -181;
			15466: out = -167;
			15467: out = -160;
			15468: out = -163;
			15469: out = -148;
			15470: out = -145;
			15471: out = -144;
			15472: out = -131;
			15473: out = -138;
			15474: out = -136;
			15475: out = -119;
			15476: out = -111;
			15477: out = -116;
			15478: out = -110;
			15479: out = -100;
			15480: out = -97;
			15481: out = -97;
			15482: out = -90;
			15483: out = -81;
			15484: out = -85;
			15485: out = -69;
			15486: out = -69;
			15487: out = -60;
			15488: out = -74;
			15489: out = -52;
			15490: out = -54;
			15491: out = -54;
			15492: out = -41;
			15493: out = -43;
			15494: out = -31;
			15495: out = -37;
			15496: out = -20;
			15497: out = -27;
			15498: out = -12;
			15499: out = -19;
			15500: out = -16;
			15501: out = -7;
			15502: out = -5;
			15503: out = -1;
			15504: out = 7;
			15505: out = 4;
			15506: out = 7;
			15507: out = 14;
			15508: out = 20;
			15509: out = 17;
			15510: out = 29;
			15511: out = 21;
			15512: out = 27;
			15513: out = 40;
			15514: out = 36;
			15515: out = 41;
			15516: out = 41;
			15517: out = 46;
			15518: out = 51;
			15519: out = 57;
			15520: out = 54;
			15521: out = 65;
			15522: out = 58;
			15523: out = 80;
			15524: out = 68;
			15525: out = 63;
			15526: out = 83;
			15527: out = 85;
			15528: out = 87;
			15529: out = 83;
			15530: out = 93;
			15531: out = 98;
			15532: out = 103;
			15533: out = 100;
			15534: out = 111;
			15535: out = 109;
			15536: out = 117;
			15537: out = 121;
			15538: out = 123;
			15539: out = 128;
			15540: out = 128;
			15541: out = 132;
			15542: out = 137;
			15543: out = 145;
			15544: out = 136;
			15545: out = 149;
			15546: out = 160;
			15547: out = 145;
			15548: out = 171;
			15549: out = 155;
			15550: out = 171;
			15551: out = 163;
			15552: out = 188;
			15553: out = 174;
			15554: out = 187;
			15555: out = 186;
			15556: out = 208;
			15557: out = 193;
			15558: out = 212;
			15559: out = 211;
			15560: out = 220;
			15561: out = 221;
			15562: out = 222;
			15563: out = 234;
			15564: out = 237;
			15565: out = 237;
			15566: out = 254;
			15567: out = 250;
			15568: out = 261;
			15569: out = 269;
			15570: out = 268;
			15571: out = 280;
			15572: out = 281;
			15573: out = 292;
			15574: out = 297;
			15575: out = 308;
			15576: out = 298;
			15577: out = 326;
			15578: out = 311;
			15579: out = 336;
			15580: out = 332;
			15581: out = 335;
			15582: out = 344;
			15583: out = 353;
			15584: out = 372;
			15585: out = 353;
			15586: out = 381;
			15587: out = 371;
			15588: out = 397;
			15589: out = 388;
			15590: out = 398;
			15591: out = 404;
			15592: out = 420;
			15593: out = 416;
			15594: out = 432;
			15595: out = 430;
			15596: out = 443;
			15597: out = 444;
			15598: out = 445;
			15599: out = 452;
			15600: out = 459;
			15601: out = 472;
			15602: out = 468;
			15603: out = 476;
			15604: out = 490;
			15605: out = 493;
			15606: out = 492;
			15607: out = 496;
			15608: out = 517;
			15609: out = 514;
			15610: out = 518;
			15611: out = 521;
			15612: out = 529;
			15613: out = 535;
			15614: out = 548;
			15615: out = 541;
			15616: out = 545;
			15617: out = 560;
			15618: out = 559;
			15619: out = 577;
			15620: out = 560;
			15621: out = 573;
			15622: out = 582;
			15623: out = 597;
			15624: out = 589;
			15625: out = 593;
			15626: out = 599;
			15627: out = 609;
			15628: out = 609;
			15629: out = 608;
			15630: out = 617;
			15631: out = 620;
			15632: out = 631;
			15633: out = 625;
			15634: out = 636;
			15635: out = 641;
			15636: out = 642;
			15637: out = 645;
			15638: out = 656;
			15639: out = 654;
			15640: out = 655;
			15641: out = 659;
			15642: out = 670;
			15643: out = 672;
			15644: out = 667;
			15645: out = 678;
			15646: out = 683;
			15647: out = 694;
			15648: out = 684;
			15649: out = 695;
			15650: out = 693;
			15651: out = 701;
			15652: out = 712;
			15653: out = 705;
			15654: out = 705;
			15655: out = 713;
			15656: out = 727;
			15657: out = 712;
			15658: out = 731;
			15659: out = 725;
			15660: out = 729;
			15661: out = 735;
			15662: out = 735;
			15663: out = 746;
			15664: out = 744;
			15665: out = 742;
			15666: out = 752;
			15667: out = 752;
			15668: out = 762;
			15669: out = 746;
			15670: out = 765;
			15671: out = 762;
			15672: out = 764;
			15673: out = 776;
			15674: out = 765;
			15675: out = 777;
			15676: out = 778;
			15677: out = 783;
			15678: out = 782;
			15679: out = 783;
			15680: out = 789;
			15681: out = 795;
			15682: out = 796;
			15683: out = 789;
			15684: out = 807;
			15685: out = 800;
			15686: out = 805;
			15687: out = 803;
			15688: out = 813;
			15689: out = 817;
			15690: out = 813;
			15691: out = 814;
			15692: out = 819;
			15693: out = 819;
			15694: out = 822;
			15695: out = 819;
			15696: out = 811;
			15697: out = 824;
			15698: out = 819;
			15699: out = 822;
			15700: out = 810;
			15701: out = 822;
			15702: out = 818;
			15703: out = 819;
			15704: out = 807;
			15705: out = 824;
			15706: out = 812;
			15707: out = 821;
			15708: out = 813;
			15709: out = 797;
			15710: out = 818;
			15711: out = 801;
			15712: out = 818;
			15713: out = 811;
			15714: out = 810;
			15715: out = 813;
			15716: out = 812;
			15717: out = 812;
			15718: out = 822;
			15719: out = 811;
			15720: out = 805;
			15721: out = 813;
			15722: out = 814;
			15723: out = 813;
			15724: out = 801;
			15725: out = 799;
			15726: out = 811;
			15727: out = 791;
			15728: out = 805;
			15729: out = 807;
			15730: out = 793;
			15731: out = 810;
			15732: out = 811;
			15733: out = 800;
			15734: out = 799;
			15735: out = 799;
			15736: out = 801;
			15737: out = 788;
			15738: out = 808;
			15739: out = 796;
			15740: out = 793;
			15741: out = 805;
			15742: out = 799;
			15743: out = 805;
			15744: out = 789;
			15745: out = 798;
			15746: out = 808;
			15747: out = 793;
			15748: out = 797;
			15749: out = 807;
			15750: out = 801;
			15751: out = 796;
			15752: out = 796;
			15753: out = 785;
			15754: out = 806;
			15755: out = 788;
			15756: out = 782;
			15757: out = 786;
			15758: out = 800;
			15759: out = 782;
			15760: out = 778;
			15761: out = 789;
			15762: out = 780;
			15763: out = 778;
			15764: out = 785;
			15765: out = 775;
			15766: out = 784;
			15767: out = 773;
			15768: out = 774;
			15769: out = 777;
			15770: out = 771;
			15771: out = 762;
			15772: out = 770;
			15773: out = 771;
			15774: out = 753;
			15775: out = 766;
			15776: out = 749;
			15777: out = 760;
			15778: out = 741;
			15779: out = 749;
			15780: out = 747;
			15781: out = 740;
			15782: out = 736;
			15783: out = 732;
			15784: out = 734;
			15785: out = 719;
			15786: out = 731;
			15787: out = 707;
			15788: out = 714;
			15789: out = 716;
			15790: out = 707;
			15791: out = 704;
			15792: out = 693;
			15793: out = 702;
			15794: out = 696;
			15795: out = 684;
			15796: out = 679;
			15797: out = 678;
			15798: out = 669;
			15799: out = 667;
			15800: out = 668;
			15801: out = 645;
			15802: out = 656;
			15803: out = 633;
			15804: out = 634;
			15805: out = 637;
			15806: out = 620;
			15807: out = 624;
			15808: out = 617;
			15809: out = 616;
			15810: out = 604;
			15811: out = 607;
			15812: out = 596;
			15813: out = 597;
			15814: out = 582;
			15815: out = 580;
			15816: out = 572;
			15817: out = 565;
			15818: out = 563;
			15819: out = 559;
			15820: out = 542;
			15821: out = 543;
			15822: out = 538;
			15823: out = 538;
			15824: out = 531;
			15825: out = 514;
			15826: out = 526;
			15827: out = 511;
			15828: out = 515;
			15829: out = 498;
			15830: out = 500;
			15831: out = 491;
			15832: out = 490;
			15833: out = 469;
			15834: out = 481;
			15835: out = 472;
			15836: out = 466;
			15837: out = 460;
			15838: out = 454;
			15839: out = 456;
			15840: out = 441;
			15841: out = 436;
			15842: out = 431;
			15843: out = 419;
			15844: out = 430;
			15845: out = 411;
			15846: out = 408;
			15847: out = 415;
			15848: out = 399;
			15849: out = 406;
			15850: out = 386;
			15851: out = 392;
			15852: out = 386;
			15853: out = 373;
			15854: out = 376;
			15855: out = 363;
			15856: out = 363;
			15857: out = 360;
			15858: out = 349;
			15859: out = 349;
			15860: out = 345;
			15861: out = 341;
			15862: out = 328;
			15863: out = 333;
			15864: out = 327;
			15865: out = 324;
			15866: out = 312;
			15867: out = 315;
			15868: out = 306;
			15869: out = 309;
			15870: out = 297;
			15871: out = 304;
			15872: out = 285;
			15873: out = 294;
			15874: out = 286;
			15875: out = 277;
			15876: out = 267;
			15877: out = 276;
			15878: out = 274;
			15879: out = 251;
			15880: out = 257;
			15881: out = 266;
			15882: out = 250;
			15883: out = 242;
			15884: out = 250;
			15885: out = 242;
			15886: out = 232;
			15887: out = 238;
			15888: out = 227;
			15889: out = 217;
			15890: out = 228;
			15891: out = 209;
			15892: out = 208;
			15893: out = 216;
			15894: out = 199;
			15895: out = 204;
			15896: out = 209;
			15897: out = 191;
			15898: out = 199;
			15899: out = 187;
			15900: out = 187;
			15901: out = 188;
			15902: out = 178;
			15903: out = 178;
			15904: out = 180;
			15905: out = 176;
			15906: out = 172;
			15907: out = 169;
			15908: out = 164;
			15909: out = 164;
			15910: out = 158;
			15911: out = 149;
			15912: out = 160;
			15913: out = 139;
			15914: out = 152;
			15915: out = 147;
			15916: out = 133;
			15917: out = 140;
			15918: out = 133;
			15919: out = 141;
			15920: out = 128;
			15921: out = 125;
			15922: out = 123;
			15923: out = 128;
			15924: out = 129;
			15925: out = 108;
			15926: out = 113;
			15927: out = 111;
			15928: out = 104;
			15929: out = 85;
			15930: out = 93;
			15931: out = 78;
			15932: out = 74;
			15933: out = 68;
			15934: out = 65;
			15935: out = 55;
			15936: out = 51;
			15937: out = 43;
			15938: out = 32;
			15939: out = 33;
			15940: out = 30;
			15941: out = 19;
			15942: out = 8;
			15943: out = 12;
			15944: out = 15;
			15945: out = -9;
			15946: out = -1;
			15947: out = -7;
			15948: out = -9;
			15949: out = -25;
			15950: out = -24;
			15951: out = -25;
			15952: out = -32;
			15953: out = -38;
			15954: out = -52;
			15955: out = -49;
			15956: out = -50;
			15957: out = -60;
			15958: out = -63;
			15959: out = -69;
			15960: out = -68;
			15961: out = -79;
			15962: out = -73;
			15963: out = -91;
			15964: out = -81;
			15965: out = -97;
			15966: out = -103;
			15967: out = -108;
			15968: out = -97;
			15969: out = -108;
			15970: out = -117;
			15971: out = -119;
			15972: out = -113;
			15973: out = -131;
			15974: out = -125;
			15975: out = -133;
			15976: out = -140;
			15977: out = -138;
			15978: out = -146;
			15979: out = -144;
			15980: out = -154;
			15981: out = -156;
			15982: out = -157;
			15983: out = -158;
			15984: out = -167;
			15985: out = -171;
			15986: out = -167;
			15987: out = -179;
			15988: out = -179;
			15989: out = -185;
			15990: out = -195;
			15991: out = -191;
			15992: out = -192;
			15993: out = -211;
			15994: out = -195;
			15995: out = -217;
			15996: out = -205;
			15997: out = -217;
			15998: out = -219;
			15999: out = -228;
			16000: out = -221;
			16001: out = -235;
			16002: out = -241;
			16003: out = -238;
			16004: out = -246;
			16005: out = -252;
			16006: out = -257;
			16007: out = -249;
			16008: out = -268;
			16009: out = -258;
			16010: out = -274;
			16011: out = -271;
			16012: out = -278;
			16013: out = -287;
			16014: out = -283;
			16015: out = -286;
			16016: out = -301;
			16017: out = -297;
			16018: out = -304;
			16019: out = -303;
			16020: out = -318;
			16021: out = -312;
			16022: out = -323;
			16023: out = -325;
			16024: out = -336;
			16025: out = -337;
			16026: out = -342;
			16027: out = -350;
			16028: out = -348;
			16029: out = -365;
			16030: out = -369;
			16031: out = -367;
			16032: out = -370;
			16033: out = -384;
			16034: out = -386;
			16035: out = -393;
			16036: out = -405;
			16037: out = -405;
			16038: out = -408;
			16039: out = -421;
			16040: out = -424;
			16041: out = -433;
			16042: out = -431;
			16043: out = -448;
			16044: out = -452;
			16045: out = -463;
			16046: out = -466;
			16047: out = -476;
			16048: out = -481;
			16049: out = -477;
			16050: out = -505;
			16051: out = -502;
			16052: out = -507;
			16053: out = -523;
			16054: out = -525;
			16055: out = -535;
			16056: out = -539;
			16057: out = -542;
			16058: out = -551;
			16059: out = -560;
			16060: out = -581;
			16061: out = -571;
			16062: out = -585;
			16063: out = -586;
			16064: out = -609;
			16065: out = -610;
			16066: out = -614;
			16067: out = -613;
			16068: out = -632;
			16069: out = -637;
			16070: out = -647;
			16071: out = -637;
			16072: out = -660;
			16073: out = -663;
			16074: out = -669;
			16075: out = -672;
			16076: out = -683;
			16077: out = -695;
			16078: out = -692;
			16079: out = -694;
			16080: out = -706;
			16081: out = -720;
			16082: out = -712;
			16083: out = -727;
			16084: out = -723;
			16085: out = -742;
			16086: out = -740;
			16087: out = -747;
			16088: out = -748;
			16089: out = -753;
			16090: out = -760;
			16091: out = -758;
			16092: out = -774;
			16093: out = -766;
			16094: out = -778;
			16095: out = -783;
			16096: out = -786;
			16097: out = -790;
			16098: out = -787;
			16099: out = -795;
			16100: out = -794;
			16101: out = -811;
			16102: out = -794;
			16103: out = -812;
			16104: out = -819;
			16105: out = -806;
			16106: out = -824;
			16107: out = -813;
			16108: out = -826;
			16109: out = -821;
			16110: out = -833;
			16111: out = -823;
			16112: out = -837;
			16113: out = -835;
			16114: out = -834;
			16115: out = -842;
			16116: out = -836;
			16117: out = -843;
			16118: out = -847;
			16119: out = -838;
			16120: out = -857;
			16121: out = -838;
			16122: out = -857;
			16123: out = -850;
			16124: out = -847;
			16125: out = -859;
			16126: out = -853;
			16127: out = -857;
			16128: out = -851;
			16129: out = -865;
			16130: out = -848;
			16131: out = -866;
			16132: out = -855;
			16133: out = -870;
			16134: out = -853;
			16135: out = -864;
			16136: out = -867;
			16137: out = -862;
			16138: out = -858;
			16139: out = -861;
			16140: out = -867;
			16141: out = -867;
			16142: out = -857;
			16143: out = -865;
			16144: out = -867;
			16145: out = -859;
			16146: out = -861;
			16147: out = -865;
			16148: out = -866;
			16149: out = -858;
			16150: out = -873;
			16151: out = -853;
			16152: out = -864;
			16153: out = -865;
			16154: out = -859;
			16155: out = -862;
			16156: out = -843;
			16157: out = -879;
			16158: out = -847;
			16159: out = -859;
			16160: out = -846;
			16161: out = -865;
			16162: out = -846;
			16163: out = -853;
			16164: out = -846;
			16165: out = -847;
			16166: out = -855;
			16167: out = -843;
			16168: out = -846;
			16169: out = -839;
			16170: out = -850;
			16171: out = -848;
			16172: out = -842;
			16173: out = -844;
			16174: out = -830;
			16175: out = -848;
			16176: out = -836;
			16177: out = -839;
			16178: out = -826;
			16179: out = -832;
			16180: out = -841;
			16181: out = -833;
			16182: out = -822;
			16183: out = -823;
			16184: out = -842;
			16185: out = -818;
			16186: out = -823;
			16187: out = -814;
			16188: out = -825;
			16189: out = -821;
			16190: out = -812;
			16191: out = -818;
			16192: out = -812;
			16193: out = -819;
			16194: out = -803;
			16195: out = -812;
			16196: out = -801;
			16197: out = -808;
			16198: out = -801;
			16199: out = -800;
			16200: out = -806;
			16201: out = -794;
			16202: out = -791;
			16203: out = -797;
			16204: out = -794;
			16205: out = -785;
			16206: out = -785;
			16207: out = -790;
			16208: out = -784;
			16209: out = -779;
			16210: out = -775;
			16211: out = -782;
			16212: out = -770;
			16213: out = -773;
			16214: out = -777;
			16215: out = -761;
			16216: out = -765;
			16217: out = -763;
			16218: out = -758;
			16219: out = -758;
			16220: out = -744;
			16221: out = -754;
			16222: out = -758;
			16223: out = -742;
			16224: out = -742;
			16225: out = -741;
			16226: out = -730;
			16227: out = -740;
			16228: out = -725;
			16229: out = -729;
			16230: out = -724;
			16231: out = -716;
			16232: out = -717;
			16233: out = -709;
			16234: out = -708;
			16235: out = -711;
			16236: out = -703;
			16237: out = -694;
			16238: out = -691;
			16239: out = -700;
			16240: out = -683;
			16241: out = -680;
			16242: out = -669;
			16243: out = -681;
			16244: out = -667;
			16245: out = -663;
			16246: out = -660;
			16247: out = -651;
			16248: out = -648;
			16249: out = -645;
			16250: out = -635;
			16251: out = -630;
			16252: out = -640;
			16253: out = -613;
			16254: out = -620;
			16255: out = -613;
			16256: out = -599;
			16257: out = -611;
			16258: out = -590;
			16259: out = -589;
			16260: out = -584;
			16261: out = -570;
			16262: out = -580;
			16263: out = -567;
			16264: out = -557;
			16265: out = -548;
			16266: out = -550;
			16267: out = -549;
			16268: out = -527;
			16269: out = -534;
			16270: out = -518;
			16271: out = -525;
			16272: out = -515;
			16273: out = -500;
			16274: out = -503;
			16275: out = -498;
			16276: out = -483;
			16277: out = -488;
			16278: out = -476;
			16279: out = -474;
			16280: out = -460;
			16281: out = -458;
			16282: out = -458;
			16283: out = -448;
			16284: out = -443;
			16285: out = -441;
			16286: out = -438;
			16287: out = -431;
			16288: out = -418;
			16289: out = -421;
			16290: out = -416;
			16291: out = -404;
			16292: out = -401;
			16293: out = -401;
			16294: out = -391;
			16295: out = -386;
			16296: out = -386;
			16297: out = -376;
			16298: out = -374;
			16299: out = -361;
			16300: out = -365;
			16301: out = -360;
			16302: out = -354;
			16303: out = -339;
			16304: out = -347;
			16305: out = -339;
			16306: out = -327;
			16307: out = -335;
			16308: out = -317;
			16309: out = -330;
			16310: out = -306;
			16311: out = -320;
			16312: out = -302;
			16313: out = -302;
			16314: out = -300;
			16315: out = -288;
			16316: out = -298;
			16317: out = -282;
			16318: out = -278;
			16319: out = -271;
			16320: out = -280;
			16321: out = -262;
			16322: out = -264;
			16323: out = -267;
			16324: out = -255;
			16325: out = -251;
			16326: out = -265;
			16327: out = -239;
			16328: out = -247;
			16329: out = -245;
			16330: out = -242;
			16331: out = -226;
			16332: out = -238;
			16333: out = -231;
			16334: out = -221;
			16335: out = -227;
			16336: out = -210;
			16337: out = -212;
			16338: out = -226;
			16339: out = -207;
			16340: out = -203;
			16341: out = -199;
			16342: out = -193;
			16343: out = -204;
			16344: out = -184;
			16345: out = -190;
			16346: out = -185;
			16347: out = -184;
			16348: out = -181;
			16349: out = -180;
			16350: out = -173;
			16351: out = -172;
			16352: out = -162;
			16353: out = -161;
			16354: out = -154;
			16355: out = -147;
			16356: out = -147;
			16357: out = -139;
			16358: out = -138;
			16359: out = -133;
			16360: out = -133;
			16361: out = -126;
			16362: out = -113;
			16363: out = -114;
			16364: out = -108;
			16365: out = -110;
			16366: out = -98;
			16367: out = -93;
			16368: out = -95;
			16369: out = -101;
			16370: out = -86;
			16371: out = -78;
			16372: out = -74;
			16373: out = -83;
			16374: out = -68;
			16375: out = -64;
			16376: out = -67;
			16377: out = -65;
			16378: out = -56;
			16379: out = -61;
			16380: out = -51;
			16381: out = -49;
			16382: out = -45;
			16383: out = -45;
			16384: out = -38;
			16385: out = -41;
			16386: out = -29;
			16387: out = -34;
			16388: out = -24;
			16389: out = -21;
			16390: out = -17;
			16391: out = -15;
			16392: out = -16;
			16393: out = -8;
			16394: out = -3;
			16395: out = -12;
			16396: out = -4;
			16397: out = 0;
			16398: out = 0;
			16399: out = 7;
			16400: out = 9;
			16401: out = 3;
			16402: out = 20;
			16403: out = 10;
			16404: out = 20;
			16405: out = 16;
			16406: out = 24;
			16407: out = 31;
			16408: out = 32;
			16409: out = 32;
			16410: out = 33;
			16411: out = 45;
			16412: out = 38;
			16413: out = 39;
			16414: out = 45;
			16415: out = 44;
			16416: out = 57;
			16417: out = 50;
			16418: out = 56;
			16419: out = 60;
			16420: out = 70;
			16421: out = 62;
			16422: out = 68;
			16423: out = 72;
			16424: out = 85;
			16425: out = 69;
			16426: out = 77;
			16427: out = 86;
			16428: out = 89;
			16429: out = 79;
			16430: out = 102;
			16431: out = 90;
			16432: out = 101;
			16433: out = 101;
			16434: out = 101;
			16435: out = 113;
			16436: out = 111;
			16437: out = 109;
			16438: out = 119;
			16439: out = 122;
			16440: out = 127;
			16441: out = 116;
			16442: out = 133;
			16443: out = 132;
			16444: out = 131;
			16445: out = 147;
			16446: out = 133;
			16447: out = 154;
			16448: out = 143;
			16449: out = 166;
			16450: out = 157;
			16451: out = 161;
			16452: out = 172;
			16453: out = 180;
			16454: out = 176;
			16455: out = 180;
			16456: out = 190;
			16457: out = 191;
			16458: out = 191;
			16459: out = 196;
			16460: out = 219;
			16461: out = 203;
			16462: out = 212;
			16463: out = 219;
			16464: out = 229;
			16465: out = 225;
			16466: out = 240;
			16467: out = 245;
			16468: out = 242;
			16469: out = 252;
			16470: out = 255;
			16471: out = 259;
			16472: out = 264;
			16473: out = 270;
			16474: out = 280;
			16475: out = 273;
			16476: out = 282;
			16477: out = 293;
			16478: out = 297;
			16479: out = 292;
			16480: out = 309;
			16481: out = 313;
			16482: out = 318;
			16483: out = 320;
			16484: out = 328;
			16485: out = 327;
			16486: out = 344;
			16487: out = 340;
			16488: out = 342;
			16489: out = 353;
			16490: out = 353;
			16491: out = 357;
			16492: out = 367;
			16493: out = 368;
			16494: out = 380;
			16495: out = 374;
			16496: out = 397;
			16497: out = 383;
			16498: out = 383;
			16499: out = 401;
			16500: out = 404;
			16501: out = 407;
			16502: out = 417;
			16503: out = 400;
			16504: out = 432;
			16505: out = 420;
			16506: out = 422;
			16507: out = 444;
			16508: out = 429;
			16509: out = 428;
			16510: out = 452;
			16511: out = 451;
			16512: out = 456;
			16513: out = 446;
			16514: out = 460;
			16515: out = 467;
			16516: out = 457;
			16517: out = 468;
			16518: out = 465;
			16519: out = 484;
			16520: out = 474;
			16521: out = 488;
			16522: out = 483;
			16523: out = 495;
			16524: out = 495;
			16525: out = 492;
			16526: out = 502;
			16527: out = 498;
			16528: out = 507;
			16529: out = 506;
			16530: out = 514;
			16531: out = 514;
			16532: out = 530;
			16533: out = 516;
			16534: out = 521;
			16535: out = 533;
			16536: out = 529;
			16537: out = 529;
			16538: out = 531;
			16539: out = 540;
			16540: out = 547;
			16541: out = 531;
			16542: out = 552;
			16543: out = 546;
			16544: out = 557;
			16545: out = 548;
			16546: out = 561;
			16547: out = 563;
			16548: out = 561;
			16549: out = 564;
			16550: out = 569;
			16551: out = 567;
			16552: out = 572;
			16553: out = 566;
			16554: out = 583;
			16555: out = 575;
			16556: out = 581;
			16557: out = 585;
			16558: out = 592;
			16559: out = 583;
			16560: out = 587;
			16561: out = 598;
			16562: out = 604;
			16563: out = 587;
			16564: out = 605;
			16565: out = 605;
			16566: out = 601;
			16567: out = 613;
			16568: out = 602;
			16569: out = 617;
			16570: out = 611;
			16571: out = 619;
			16572: out = 620;
			16573: out = 625;
			16574: out = 620;
			16575: out = 630;
			16576: out = 620;
			16577: out = 637;
			16578: out = 621;
			16579: out = 626;
			16580: out = 633;
			16581: out = 630;
			16582: out = 647;
			16583: out = 625;
			16584: out = 646;
			16585: out = 633;
			16586: out = 646;
			16587: out = 635;
			16588: out = 646;
			16589: out = 640;
			16590: out = 649;
			16591: out = 632;
			16592: out = 640;
			16593: out = 638;
			16594: out = 641;
			16595: out = 622;
			16596: out = 634;
			16597: out = 630;
			16598: out = 625;
			16599: out = 644;
			16600: out = 623;
			16601: out = 637;
			16602: out = 631;
			16603: out = 638;
			16604: out = 632;
			16605: out = 626;
			16606: out = 638;
			16607: out = 628;
			16608: out = 634;
			16609: out = 623;
			16610: out = 642;
			16611: out = 631;
			16612: out = 638;
			16613: out = 622;
			16614: out = 638;
			16615: out = 634;
			16616: out = 625;
			16617: out = 628;
			16618: out = 625;
			16619: out = 632;
			16620: out = 633;
			16621: out = 621;
			16622: out = 632;
			16623: out = 622;
			16624: out = 623;
			16625: out = 622;
			16626: out = 626;
			16627: out = 622;
			16628: out = 623;
			16629: out = 628;
			16630: out = 619;
			16631: out = 619;
			16632: out = 631;
			16633: out = 618;
			16634: out = 614;
			16635: out = 629;
			16636: out = 614;
			16637: out = 635;
			16638: out = 616;
			16639: out = 620;
			16640: out = 614;
			16641: out = 636;
			16642: out = 611;
			16643: out = 619;
			16644: out = 619;
			16645: out = 628;
			16646: out = 605;
			16647: out = 622;
			16648: out = 610;
			16649: out = 618;
			16650: out = 616;
			16651: out = 607;
			16652: out = 619;
			16653: out = 611;
			16654: out = 614;
			16655: out = 601;
			16656: out = 610;
			16657: out = 607;
			16658: out = 600;
			16659: out = 596;
			16660: out = 602;
			16661: out = 602;
			16662: out = 593;
			16663: out = 592;
			16664: out = 598;
			16665: out = 596;
			16666: out = 590;
			16667: out = 575;
			16668: out = 598;
			16669: out = 581;
			16670: out = 580;
			16671: out = 573;
			16672: out = 583;
			16673: out = 567;
			16674: out = 569;
			16675: out = 565;
			16676: out = 558;
			16677: out = 573;
			16678: out = 545;
			16679: out = 557;
			16680: out = 549;
			16681: out = 553;
			16682: out = 547;
			16683: out = 524;
			16684: out = 543;
			16685: out = 533;
			16686: out = 533;
			16687: out = 522;
			16688: out = 526;
			16689: out = 517;
			16690: out = 517;
			16691: out = 512;
			16692: out = 505;
			16693: out = 499;
			16694: out = 504;
			16695: out = 492;
			16696: out = 477;
			16697: out = 493;
			16698: out = 477;
			16699: out = 466;
			16700: out = 477;
			16701: out = 468;
			16702: out = 459;
			16703: out = 459;
			16704: out = 454;
			16705: out = 451;
			16706: out = 439;
			16707: out = 442;
			16708: out = 445;
			16709: out = 424;
			16710: out = 431;
			16711: out = 422;
			16712: out = 425;
			16713: out = 412;
			16714: out = 407;
			16715: out = 408;
			16716: out = 404;
			16717: out = 401;
			16718: out = 395;
			16719: out = 389;
			16720: out = 392;
			16721: out = 371;
			16722: out = 377;
			16723: out = 379;
			16724: out = 363;
			16725: out = 358;
			16726: out = 360;
			16727: out = 354;
			16728: out = 347;
			16729: out = 349;
			16730: out = 339;
			16731: out = 345;
			16732: out = 333;
			16733: out = 329;
			16734: out = 327;
			16735: out = 324;
			16736: out = 312;
			16737: out = 310;
			16738: out = 311;
			16739: out = 299;
			16740: out = 314;
			16741: out = 292;
			16742: out = 293;
			16743: out = 289;
			16744: out = 296;
			16745: out = 282;
			16746: out = 276;
			16747: out = 280;
			16748: out = 267;
			16749: out = 262;
			16750: out = 264;
			16751: out = 266;
			16752: out = 255;
			16753: out = 261;
			16754: out = 245;
			16755: out = 251;
			16756: out = 245;
			16757: out = 238;
			16758: out = 231;
			16759: out = 228;
			16760: out = 231;
			16761: out = 230;
			16762: out = 220;
			16763: out = 222;
			16764: out = 220;
			16765: out = 207;
			16766: out = 218;
			16767: out = 202;
			16768: out = 202;
			16769: out = 203;
			16770: out = 191;
			16771: out = 202;
			16772: out = 185;
			16773: out = 191;
			16774: out = 185;
			16775: out = 186;
			16776: out = 176;
			16777: out = 175;
			16778: out = 174;
			16779: out = 168;
			16780: out = 173;
			16781: out = 160;
			16782: out = 159;
			16783: out = 161;
			16784: out = 161;
			16785: out = 152;
			16786: out = 148;
			16787: out = 149;
			16788: out = 160;
			16789: out = 136;
			16790: out = 145;
			16791: out = 146;
			16792: out = 134;
			16793: out = 124;
			16794: out = 137;
			16795: out = 133;
			16796: out = 124;
			16797: out = 123;
			16798: out = 129;
			16799: out = 119;
			16800: out = 121;
			16801: out = 112;
			16802: out = 114;
			16803: out = 112;
			16804: out = 110;
			16805: out = 114;
			16806: out = 102;
			16807: out = 111;
			16808: out = 92;
			16809: out = 111;
			16810: out = 97;
			16811: out = 99;
			16812: out = 97;
			16813: out = 96;
			16814: out = 85;
			16815: out = 96;
			16816: out = 88;
			16817: out = 64;
			16818: out = 86;
			16819: out = 64;
			16820: out = 67;
			16821: out = 60;
			16822: out = 54;
			16823: out = 48;
			16824: out = 50;
			16825: out = 41;
			16826: out = 33;
			16827: out = 30;
			16828: out = 31;
			16829: out = 10;
			16830: out = 13;
			16831: out = 15;
			16832: out = 3;
			16833: out = 5;
			16834: out = -7;
			16835: out = -4;
			16836: out = -7;
			16837: out = -16;
			16838: out = -18;
			16839: out = -32;
			16840: out = -16;
			16841: out = -37;
			16842: out = -31;
			16843: out = -42;
			16844: out = -38;
			16845: out = -55;
			16846: out = -40;
			16847: out = -61;
			16848: out = -53;
			16849: out = -62;
			16850: out = -65;
			16851: out = -63;
			16852: out = -75;
			16853: out = -74;
			16854: out = -73;
			16855: out = -85;
			16856: out = -85;
			16857: out = -87;
			16858: out = -90;
			16859: out = -96;
			16860: out = -102;
			16861: out = -97;
			16862: out = -111;
			16863: out = -105;
			16864: out = -123;
			16865: out = -103;
			16866: out = -123;
			16867: out = -120;
			16868: out = -127;
			16869: out = -125;
			16870: out = -125;
			16871: out = -138;
			16872: out = -132;
			16873: out = -141;
			16874: out = -144;
			16875: out = -145;
			16876: out = -148;
			16877: out = -160;
			16878: out = -156;
			16879: out = -149;
			16880: out = -173;
			16881: out = -164;
			16882: out = -170;
			16883: out = -161;
			16884: out = -181;
			16885: out = -176;
			16886: out = -178;
			16887: out = -183;
			16888: out = -181;
			16889: out = -193;
			16890: out = -186;
			16891: out = -191;
			16892: out = -199;
			16893: out = -191;
			16894: out = -212;
			16895: out = -208;
			16896: out = -205;
			16897: out = -217;
			16898: out = -211;
			16899: out = -229;
			16900: out = -210;
			16901: out = -227;
			16902: out = -225;
			16903: out = -235;
			16904: out = -235;
			16905: out = -234;
			16906: out = -243;
			16907: out = -243;
			16908: out = -249;
			16909: out = -249;
			16910: out = -261;
			16911: out = -266;
			16912: out = -261;
			16913: out = -270;
			16914: out = -275;
			16915: out = -275;
			16916: out = -283;
			16917: out = -280;
			16918: out = -286;
			16919: out = -305;
			16920: out = -292;
			16921: out = -298;
			16922: out = -312;
			16923: out = -302;
			16924: out = -320;
			16925: out = -316;
			16926: out = -326;
			16927: out = -323;
			16928: out = -337;
			16929: out = -340;
			16930: out = -339;
			16931: out = -349;
			16932: out = -359;
			16933: out = -354;
			16934: out = -357;
			16935: out = -373;
			16936: out = -379;
			16937: out = -368;
			16938: out = -391;
			16939: out = -389;
			16940: out = -396;
			16941: out = -412;
			16942: out = -407;
			16943: out = -412;
			16944: out = -415;
			16945: out = -435;
			16946: out = -430;
			16947: out = -438;
			16948: out = -440;
			16949: out = -457;
			16950: out = -454;
			16951: out = -460;
			16952: out = -458;
			16953: out = -467;
			16954: out = -481;
			16955: out = -483;
			16956: out = -484;
			16957: out = -494;
			16958: out = -504;
			16959: out = -506;
			16960: out = -518;
			16961: out = -505;
			16962: out = -525;
			16963: out = -527;
			16964: out = -527;
			16965: out = -542;
			16966: out = -531;
			16967: out = -553;
			16968: out = -554;
			16969: out = -560;
			16970: out = -560;
			16971: out = -567;
			16972: out = -559;
			16973: out = -577;
			16974: out = -575;
			16975: out = -581;
			16976: out = -590;
			16977: out = -595;
			16978: out = -590;
			16979: out = -602;
			16980: out = -605;
			16981: out = -598;
			16982: out = -621;
			16983: out = -602;
			16984: out = -618;
			16985: out = -625;
			16986: out = -624;
			16987: out = -623;
			16988: out = -629;
			16989: out = -632;
			16990: out = -633;
			16991: out = -636;
			16992: out = -642;
			16993: out = -641;
			16994: out = -652;
			16995: out = -642;
			16996: out = -645;
			16997: out = -659;
			16998: out = -646;
			16999: out = -654;
			17000: out = -658;
			17001: out = -651;
			17002: out = -667;
			17003: out = -656;
			17004: out = -665;
			17005: out = -660;
			17006: out = -668;
			17007: out = -666;
			17008: out = -675;
			17009: out = -676;
			17010: out = -664;
			17011: out = -672;
			17012: out = -677;
			17013: out = -667;
			17014: out = -685;
			17015: out = -669;
			17016: out = -681;
			17017: out = -687;
			17018: out = -679;
			17019: out = -680;
			17020: out = -681;
			17021: out = -678;
			17022: out = -689;
			17023: out = -671;
			17024: out = -688;
			17025: out = -683;
			17026: out = -687;
			17027: out = -683;
			17028: out = -690;
			17029: out = -683;
			17030: out = -691;
			17031: out = -681;
			17032: out = -688;
			17033: out = -691;
			17034: out = -682;
			17035: out = -689;
			17036: out = -687;
			17037: out = -687;
			17038: out = -685;
			17039: out = -685;
			17040: out = -684;
			17041: out = -695;
			17042: out = -679;
			17043: out = -684;
			17044: out = -684;
			17045: out = -683;
			17046: out = -682;
			17047: out = -680;
			17048: out = -681;
			17049: out = -684;
			17050: out = -678;
			17051: out = -691;
			17052: out = -679;
			17053: out = -671;
			17054: out = -687;
			17055: out = -677;
			17056: out = -679;
			17057: out = -672;
			17058: out = -679;
			17059: out = -679;
			17060: out = -663;
			17061: out = -683;
			17062: out = -664;
			17063: out = -678;
			17064: out = -670;
			17065: out = -672;
			17066: out = -659;
			17067: out = -673;
			17068: out = -666;
			17069: out = -660;
			17070: out = -669;
			17071: out = -652;
			17072: out = -668;
			17073: out = -659;
			17074: out = -656;
			17075: out = -665;
			17076: out = -656;
			17077: out = -654;
			17078: out = -657;
			17079: out = -652;
			17080: out = -656;
			17081: out = -646;
			17082: out = -643;
			17083: out = -649;
			17084: out = -645;
			17085: out = -643;
			17086: out = -641;
			17087: out = -642;
			17088: out = -646;
			17089: out = -638;
			17090: out = -641;
			17091: out = -641;
			17092: out = -633;
			17093: out = -636;
			17094: out = -633;
			17095: out = -629;
			17096: out = -629;
			17097: out = -629;
			17098: out = -623;
			17099: out = -631;
			17100: out = -610;
			17101: out = -630;
			17102: out = -622;
			17103: out = -610;
			17104: out = -617;
			17105: out = -613;
			17106: out = -605;
			17107: out = -610;
			17108: out = -610;
			17109: out = -599;
			17110: out = -604;
			17111: out = -595;
			17112: out = -602;
			17113: out = -594;
			17114: out = -588;
			17115: out = -597;
			17116: out = -583;
			17117: out = -587;
			17118: out = -589;
			17119: out = -582;
			17120: out = -576;
			17121: out = -576;
			17122: out = -573;
			17123: out = -576;
			17124: out = -560;
			17125: out = -567;
			17126: out = -564;
			17127: out = -557;
			17128: out = -548;
			17129: out = -552;
			17130: out = -546;
			17131: out = -549;
			17132: out = -540;
			17133: out = -533;
			17134: out = -535;
			17135: out = -547;
			17136: out = -516;
			17137: out = -530;
			17138: out = -513;
			17139: out = -524;
			17140: out = -509;
			17141: out = -510;
			17142: out = -502;
			17143: out = -500;
			17144: out = -494;
			17145: out = -490;
			17146: out = -489;
			17147: out = -479;
			17148: out = -476;
			17149: out = -468;
			17150: out = -480;
			17151: out = -460;
			17152: out = -463;
			17153: out = -455;
			17154: out = -450;
			17155: out = -453;
			17156: out = -438;
			17157: out = -436;
			17158: out = -428;
			17159: out = -429;
			17160: out = -432;
			17161: out = -404;
			17162: out = -420;
			17163: out = -416;
			17164: out = -397;
			17165: out = -397;
			17166: out = -395;
			17167: out = -395;
			17168: out = -381;
			17169: out = -381;
			17170: out = -379;
			17171: out = -374;
			17172: out = -369;
			17173: out = -367;
			17174: out = -356;
			17175: out = -357;
			17176: out = -356;
			17177: out = -345;
			17178: out = -340;
			17179: out = -350;
			17180: out = -330;
			17181: out = -344;
			17182: out = -326;
			17183: out = -322;
			17184: out = -327;
			17185: out = -311;
			17186: out = -320;
			17187: out = -305;
			17188: out = -308;
			17189: out = -294;
			17190: out = -303;
			17191: out = -286;
			17192: out = -294;
			17193: out = -280;
			17194: out = -277;
			17195: out = -282;
			17196: out = -276;
			17197: out = -265;
			17198: out = -269;
			17199: out = -266;
			17200: out = -262;
			17201: out = -258;
			17202: out = -250;
			17203: out = -265;
			17204: out = -232;
			17205: out = -254;
			17206: out = -235;
			17207: out = -234;
			17208: out = -239;
			17209: out = -232;
			17210: out = -230;
			17211: out = -219;
			17212: out = -219;
			17213: out = -221;
			17214: out = -214;
			17215: out = -217;
			17216: out = -208;
			17217: out = -206;
			17218: out = -205;
			17219: out = -208;
			17220: out = -193;
			17221: out = -196;
			17222: out = -195;
			17223: out = -193;
			17224: out = -180;
			17225: out = -199;
			17226: out = -178;
			17227: out = -180;
			17228: out = -184;
			17229: out = -170;
			17230: out = -181;
			17231: out = -172;
			17232: out = -170;
			17233: out = -164;
			17234: out = -160;
			17235: out = -171;
			17236: out = -154;
			17237: out = -154;
			17238: out = -164;
			17239: out = -152;
			17240: out = -147;
			17241: out = -148;
			17242: out = -145;
			17243: out = -138;
			17244: out = -131;
			17245: out = -128;
			17246: out = -129;
			17247: out = -111;
			17248: out = -128;
			17249: out = -115;
			17250: out = -104;
			17251: out = -115;
			17252: out = -105;
			17253: out = -100;
			17254: out = -98;
			17255: out = -95;
			17256: out = -95;
			17257: out = -89;
			17258: out = -89;
			17259: out = -77;
			17260: out = -76;
			17261: out = -83;
			17262: out = -76;
			17263: out = -58;
			17264: out = -78;
			17265: out = -61;
			17266: out = -67;
			17267: out = -50;
			17268: out = -53;
			17269: out = -54;
			17270: out = -52;
			17271: out = -44;
			17272: out = -40;
			17273: out = -44;
			17274: out = -40;
			17275: out = -40;
			17276: out = -41;
			17277: out = -24;
			17278: out = -33;
			17279: out = -36;
			17280: out = -21;
			17281: out = -21;
			17282: out = -15;
			17283: out = -16;
			17284: out = -22;
			17285: out = -15;
			17286: out = -9;
			17287: out = -8;
			17288: out = -8;
			17289: out = -5;
			17290: out = -5;
			17291: out = 6;
			17292: out = -6;
			17293: out = 4;
			17294: out = 6;
			17295: out = 17;
			17296: out = 13;
			17297: out = 2;
			17298: out = 20;
			17299: out = 21;
			17300: out = 21;
			17301: out = 21;
			17302: out = 20;
			17303: out = 26;
			17304: out = 34;
			17305: out = 28;
			17306: out = 34;
			17307: out = 36;
			17308: out = 38;
			17309: out = 45;
			17310: out = 41;
			17311: out = 41;
			17312: out = 54;
			17313: out = 43;
			17314: out = 45;
			17315: out = 53;
			17316: out = 56;
			17317: out = 52;
			17318: out = 62;
			17319: out = 58;
			17320: out = 67;
			17321: out = 54;
			17322: out = 75;
			17323: out = 67;
			17324: out = 67;
			17325: out = 83;
			17326: out = 64;
			17327: out = 85;
			17328: out = 79;
			17329: out = 85;
			17330: out = 93;
			17331: out = 87;
			17332: out = 96;
			17333: out = 101;
			17334: out = 103;
			17335: out = 102;
			17336: out = 103;
			17337: out = 107;
			17338: out = 121;
			17339: out = 110;
			17340: out = 113;
			17341: out = 122;
			17342: out = 133;
			17343: out = 126;
			17344: out = 125;
			17345: out = 144;
			17346: out = 138;
			17347: out = 143;
			17348: out = 134;
			17349: out = 155;
			17350: out = 147;
			17351: out = 152;
			17352: out = 158;
			17353: out = 161;
			17354: out = 170;
			17355: out = 167;
			17356: out = 176;
			17357: out = 179;
			17358: out = 176;
			17359: out = 183;
			17360: out = 194;
			17361: out = 185;
			17362: out = 206;
			17363: out = 199;
			17364: out = 202;
			17365: out = 216;
			17366: out = 210;
			17367: out = 212;
			17368: out = 221;
			17369: out = 233;
			17370: out = 234;
			17371: out = 238;
			17372: out = 228;
			17373: out = 254;
			17374: out = 245;
			17375: out = 251;
			17376: out = 255;
			17377: out = 257;
			17378: out = 262;
			17379: out = 266;
			17380: out = 276;
			17381: out = 269;
			17382: out = 285;
			17383: out = 279;
			17384: out = 278;
			17385: out = 296;
			17386: out = 291;
			17387: out = 287;
			17388: out = 306;
			17389: out = 297;
			17390: out = 313;
			17391: out = 309;
			17392: out = 315;
			17393: out = 316;
			17394: out = 329;
			17395: out = 315;
			17396: out = 326;
			17397: out = 334;
			17398: out = 329;
			17399: out = 341;
			17400: out = 333;
			17401: out = 340;
			17402: out = 340;
			17403: out = 350;
			17404: out = 340;
			17405: out = 358;
			17406: out = 352;
			17407: out = 361;
			17408: out = 364;
			17409: out = 364;
			17410: out = 375;
			17411: out = 372;
			17412: out = 373;
			17413: out = 374;
			17414: out = 383;
			17415: out = 380;
			17416: out = 384;
			17417: out = 381;
			17418: out = 397;
			17419: out = 393;
			17420: out = 386;
			17421: out = 401;
			17422: out = 403;
			17423: out = 403;
			17424: out = 400;
			17425: out = 399;
			17426: out = 413;
			17427: out = 417;
			17428: out = 413;
			17429: out = 409;
			17430: out = 420;
			17431: out = 430;
			17432: out = 418;
			17433: out = 422;
			17434: out = 430;
			17435: out = 438;
			17436: out = 422;
			17437: out = 432;
			17438: out = 439;
			17439: out = 428;
			17440: out = 444;
			17441: out = 441;
			17442: out = 444;
			17443: out = 441;
			17444: out = 450;
			17445: out = 456;
			17446: out = 442;
			17447: out = 456;
			17448: out = 450;
			17449: out = 455;
			17450: out = 465;
			17451: out = 456;
			17452: out = 474;
			17453: out = 455;
			17454: out = 468;
			17455: out = 465;
			17456: out = 467;
			17457: out = 477;
			17458: out = 469;
			17459: out = 470;
			17460: out = 486;
			17461: out = 469;
			17462: out = 488;
			17463: out = 478;
			17464: out = 483;
			17465: out = 486;
			17466: out = 489;
			17467: out = 488;
			17468: out = 489;
			17469: out = 488;
			17470: out = 487;
			17471: out = 490;
			17472: out = 489;
			17473: out = 491;
			17474: out = 492;
			17475: out = 495;
			17476: out = 482;
			17477: out = 500;
			17478: out = 491;
			17479: out = 489;
			17480: out = 493;
			17481: out = 494;
			17482: out = 489;
			17483: out = 492;
			17484: out = 500;
			17485: out = 480;
			17486: out = 500;
			17487: out = 478;
			17488: out = 501;
			17489: out = 481;
			17490: out = 487;
			17491: out = 500;
			17492: out = 493;
			17493: out = 489;
			17494: out = 493;
			17495: out = 498;
			17496: out = 486;
			17497: out = 493;
			17498: out = 484;
			17499: out = 482;
			17500: out = 490;
			17501: out = 487;
			17502: out = 474;
			17503: out = 489;
			17504: out = 482;
			17505: out = 480;
			17506: out = 481;
			17507: out = 483;
			17508: out = 482;
			17509: out = 483;
			17510: out = 480;
			17511: out = 490;
			17512: out = 475;
			17513: out = 484;
			17514: out = 487;
			17515: out = 487;
			17516: out = 476;
			17517: out = 488;
			17518: out = 479;
			17519: out = 487;
			17520: out = 470;
			17521: out = 480;
			17522: out = 474;
			17523: out = 482;
			17524: out = 468;
			17525: out = 483;
			17526: out = 480;
			17527: out = 477;
			17528: out = 479;
			17529: out = 470;
			17530: out = 484;
			17531: out = 474;
			17532: out = 462;
			17533: out = 483;
			17534: out = 472;
			17535: out = 470;
			17536: out = 482;
			17537: out = 471;
			17538: out = 477;
			17539: out = 474;
			17540: out = 472;
			17541: out = 467;
			17542: out = 468;
			17543: out = 471;
			17544: out = 465;
			17545: out = 462;
			17546: out = 470;
			17547: out = 464;
			17548: out = 463;
			17549: out = 469;
			17550: out = 456;
			17551: out = 467;
			17552: out = 458;
			17553: out = 463;
			17554: out = 458;
			17555: out = 451;
			17556: out = 447;
			17557: out = 455;
			17558: out = 444;
			17559: out = 435;
			17560: out = 444;
			17561: out = 440;
			17562: out = 442;
			17563: out = 431;
			17564: out = 436;
			17565: out = 429;
			17566: out = 434;
			17567: out = 430;
			17568: out = 417;
			17569: out = 423;
			17570: out = 417;
			17571: out = 428;
			17572: out = 411;
			17573: out = 408;
			17574: out = 411;
			17575: out = 417;
			17576: out = 405;
			17577: out = 403;
			17578: out = 394;
			17579: out = 405;
			17580: out = 391;
			17581: out = 389;
			17582: out = 396;
			17583: out = 379;
			17584: out = 377;
			17585: out = 387;
			17586: out = 364;
			17587: out = 372;
			17588: out = 362;
			17589: out = 370;
			17590: out = 350;
			17591: out = 359;
			17592: out = 352;
			17593: out = 349;
			17594: out = 341;
			17595: out = 340;
			17596: out = 341;
			17597: out = 333;
			17598: out = 333;
			17599: out = 328;
			17600: out = 327;
			17601: out = 320;
			17602: out = 317;
			17603: out = 324;
			17604: out = 305;
			17605: out = 304;
			17606: out = 309;
			17607: out = 305;
			17608: out = 289;
			17609: out = 291;
			17610: out = 294;
			17611: out = 286;
			17612: out = 286;
			17613: out = 283;
			17614: out = 279;
			17615: out = 270;
			17616: out = 277;
			17617: out = 258;
			17618: out = 267;
			17619: out = 258;
			17620: out = 253;
			17621: out = 262;
			17622: out = 243;
			17623: out = 256;
			17624: out = 241;
			17625: out = 238;
			17626: out = 245;
			17627: out = 237;
			17628: out = 223;
			17629: out = 234;
			17630: out = 230;
			17631: out = 215;
			17632: out = 220;
			17633: out = 214;
			17634: out = 216;
			17635: out = 211;
			17636: out = 197;
			17637: out = 208;
			17638: out = 203;
			17639: out = 196;
			17640: out = 193;
			17641: out = 192;
			17642: out = 185;
			17643: out = 184;
			17644: out = 186;
			17645: out = 179;
			17646: out = 171;
			17647: out = 176;
			17648: out = 170;
			17649: out = 169;
			17650: out = 171;
			17651: out = 164;
			17652: out = 161;
			17653: out = 164;
			17654: out = 156;
			17655: out = 155;
			17656: out = 149;
			17657: out = 150;
			17658: out = 148;
			17659: out = 147;
			17660: out = 139;
			17661: out = 135;
			17662: out = 144;
			17663: out = 138;
			17664: out = 120;
			17665: out = 139;
			17666: out = 119;
			17667: out = 128;
			17668: out = 124;
			17669: out = 125;
			17670: out = 122;
			17671: out = 111;
			17672: out = 119;
			17673: out = 113;
			17674: out = 115;
			17675: out = 111;
			17676: out = 93;
			17677: out = 104;
			17678: out = 112;
			17679: out = 98;
			17680: out = 98;
			17681: out = 91;
			17682: out = 101;
			17683: out = 96;
			17684: out = 88;
			17685: out = 92;
			17686: out = 88;
			17687: out = 81;
			17688: out = 80;
			17689: out = 84;
			17690: out = 74;
			17691: out = 81;
			17692: out = 74;
			17693: out = 77;
			17694: out = 73;
			17695: out = 73;
			17696: out = 65;
			17697: out = 66;
			17698: out = 77;
			17699: out = 55;
			17700: out = 53;
			17701: out = 68;
			17702: out = 64;
			17703: out = 56;
			17704: out = 51;
			17705: out = 61;
			17706: out = 54;
			17707: out = 50;
			17708: out = 44;
			17709: out = 50;
			17710: out = 31;
			17711: out = 39;
			17712: out = 36;
			17713: out = 22;
			17714: out = 25;
			17715: out = 22;
			17716: out = 14;
			17717: out = 17;
			17718: out = 5;
			17719: out = 4;
			17720: out = 5;
			17721: out = -3;
			17722: out = -6;
			17723: out = -13;
			17724: out = -5;
			17725: out = -22;
			17726: out = -6;
			17727: out = -30;
			17728: out = -21;
			17729: out = -26;
			17730: out = -29;
			17731: out = -38;
			17732: out = -32;
			17733: out = -42;
			17734: out = -32;
			17735: out = -49;
			17736: out = -48;
			17737: out = -44;
			17738: out = -57;
			17739: out = -57;
			17740: out = -60;
			17741: out = -57;
			17742: out = -64;
			17743: out = -69;
			17744: out = -63;
			17745: out = -72;
			17746: out = -83;
			17747: out = -73;
			17748: out = -76;
			17749: out = -74;
			17750: out = -93;
			17751: out = -91;
			17752: out = -81;
			17753: out = -95;
			17754: out = -97;
			17755: out = -97;
			17756: out = -97;
			17757: out = -102;
			17758: out = -103;
			17759: out = -108;
			17760: out = -104;
			17761: out = -110;
			17762: out = -112;
			17763: out = -124;
			17764: out = -111;
			17765: out = -114;
			17766: out = -136;
			17767: out = -123;
			17768: out = -131;
			17769: out = -122;
			17770: out = -139;
			17771: out = -137;
			17772: out = -133;
			17773: out = -146;
			17774: out = -135;
			17775: out = -145;
			17776: out = -155;
			17777: out = -141;
			17778: out = -150;
			17779: out = -151;
			17780: out = -156;
			17781: out = -152;
			17782: out = -170;
			17783: out = -154;
			17784: out = -169;
			17785: out = -169;
			17786: out = -159;
			17787: out = -184;
			17788: out = -182;
			17789: out = -168;
			17790: out = -179;
			17791: out = -183;
			17792: out = -183;
			17793: out = -193;
			17794: out = -183;
			17795: out = -195;
			17796: out = -196;
			17797: out = -209;
			17798: out = -194;
			17799: out = -205;
			17800: out = -206;
			17801: out = -204;
			17802: out = -211;
			17803: out = -216;
			17804: out = -214;
			17805: out = -218;
			17806: out = -221;
			17807: out = -232;
			17808: out = -229;
			17809: out = -235;
			17810: out = -235;
			17811: out = -238;
			17812: out = -247;
			17813: out = -245;
			17814: out = -246;
			17815: out = -254;
			17816: out = -255;
			17817: out = -253;
			17818: out = -275;
			17819: out = -271;
			17820: out = -261;
			17821: out = -282;
			17822: out = -277;
			17823: out = -279;
			17824: out = -298;
			17825: out = -297;
			17826: out = -294;
			17827: out = -297;
			17828: out = -310;
			17829: out = -311;
			17830: out = -310;
			17831: out = -318;
			17832: out = -314;
			17833: out = -339;
			17834: out = -338;
			17835: out = -325;
			17836: out = -348;
			17837: out = -342;
			17838: out = -350;
			17839: out = -348;
			17840: out = -365;
			17841: out = -361;
			17842: out = -362;
			17843: out = -373;
			17844: out = -379;
			17845: out = -382;
			17846: out = -391;
			17847: out = -391;
			17848: out = -391;
			17849: out = -400;
			17850: out = -410;
			17851: out = -405;
			17852: out = -410;
			17853: out = -415;
			17854: out = -411;
			17855: out = -439;
			17856: out = -424;
			17857: out = -428;
			17858: out = -434;
			17859: out = -434;
			17860: out = -445;
			17861: out = -451;
			17862: out = -451;
			17863: out = -442;
			17864: out = -468;
			17865: out = -462;
			17866: out = -464;
			17867: out = -462;
			17868: out = -462;
			17869: out = -484;
			17870: out = -467;
			17871: out = -477;
			17872: out = -472;
			17873: out = -491;
			17874: out = -488;
			17875: out = -483;
			17876: out = -483;
			17877: out = -501;
			17878: out = -490;
			17879: out = -493;
			17880: out = -503;
			17881: out = -496;
			17882: out = -506;
			17883: out = -507;
			17884: out = -505;
			17885: out = -516;
			17886: out = -510;
			17887: out = -511;
			17888: out = -518;
			17889: out = -522;
			17890: out = -513;
			17891: out = -522;
			17892: out = -526;
			17893: out = -521;
			17894: out = -518;
			17895: out = -535;
			17896: out = -526;
			17897: out = -529;
			17898: out = -530;
			17899: out = -533;
			17900: out = -540;
			17901: out = -519;
			17902: out = -531;
			17903: out = -534;
			17904: out = -531;
			17905: out = -525;
			17906: out = -535;
			17907: out = -537;
			17908: out = -538;
			17909: out = -537;
			17910: out = -533;
			17911: out = -542;
			17912: out = -540;
			17913: out = -531;
			17914: out = -539;
			17915: out = -539;
			17916: out = -543;
			17917: out = -531;
			17918: out = -541;
			17919: out = -542;
			17920: out = -533;
			17921: out = -546;
			17922: out = -551;
			17923: out = -525;
			17924: out = -553;
			17925: out = -534;
			17926: out = -547;
			17927: out = -540;
			17928: out = -539;
			17929: out = -546;
			17930: out = -534;
			17931: out = -540;
			17932: out = -540;
			17933: out = -537;
			17934: out = -537;
			17935: out = -539;
			17936: out = -545;
			17937: out = -537;
			17938: out = -537;
			17939: out = -547;
			17940: out = -537;
			17941: out = -542;
			17942: out = -528;
			17943: out = -546;
			17944: out = -538;
			17945: out = -535;
			17946: out = -539;
			17947: out = -531;
			17948: out = -534;
			17949: out = -548;
			17950: out = -528;
			17951: out = -529;
			17952: out = -531;
			17953: out = -537;
			17954: out = -530;
			17955: out = -528;
			17956: out = -528;
			17957: out = -530;
			17958: out = -528;
			17959: out = -525;
			17960: out = -519;
			17961: out = -522;
			17962: out = -536;
			17963: out = -516;
			17964: out = -518;
			17965: out = -525;
			17966: out = -531;
			17967: out = -507;
			17968: out = -527;
			17969: out = -510;
			17970: out = -524;
			17971: out = -510;
			17972: out = -516;
			17973: out = -514;
			17974: out = -510;
			17975: out = -513;
			17976: out = -507;
			17977: out = -517;
			17978: out = -506;
			17979: out = -503;
			17980: out = -515;
			17981: out = -502;
			17982: out = -511;
			17983: out = -495;
			17984: out = -519;
			17985: out = -490;
			17986: out = -504;
			17987: out = -498;
			17988: out = -501;
			17989: out = -498;
			17990: out = -488;
			17991: out = -493;
			17992: out = -496;
			17993: out = -488;
			17994: out = -479;
			17995: out = -491;
			17996: out = -487;
			17997: out = -478;
			17998: out = -492;
			17999: out = -476;
			18000: out = -486;
			18001: out = -477;
			18002: out = -480;
			18003: out = -476;
			18004: out = -470;
			18005: out = -480;
			18006: out = -469;
			18007: out = -468;
			18008: out = -467;
			18009: out = -470;
			18010: out = -455;
			18011: out = -468;
			18012: out = -460;
			18013: out = -454;
			18014: out = -458;
			18015: out = -454;
			18016: out = -454;
			18017: out = -441;
			18018: out = -444;
			18019: out = -444;
			18020: out = -433;
			18021: out = -438;
			18022: out = -438;
			18023: out = -427;
			18024: out = -432;
			18025: out = -419;
			18026: out = -432;
			18027: out = -424;
			18028: out = -413;
			18029: out = -416;
			18030: out = -405;
			18031: out = -407;
			18032: out = -397;
			18033: out = -408;
			18034: out = -399;
			18035: out = -384;
			18036: out = -399;
			18037: out = -388;
			18038: out = -373;
			18039: out = -387;
			18040: out = -369;
			18041: out = -377;
			18042: out = -365;
			18043: out = -363;
			18044: out = -369;
			18045: out = -359;
			18046: out = -353;
			18047: out = -354;
			18048: out = -350;
			18049: out = -338;
			18050: out = -347;
			18051: out = -339;
			18052: out = -332;
			18053: out = -335;
			18054: out = -336;
			18055: out = -322;
			18056: out = -329;
			18057: out = -314;
			18058: out = -313;
			18059: out = -318;
			18060: out = -298;
			18061: out = -304;
			18062: out = -304;
			18063: out = -291;
			18064: out = -297;
			18065: out = -288;
			18066: out = -282;
			18067: out = -282;
			18068: out = -275;
			18069: out = -278;
			18070: out = -268;
			18071: out = -266;
			18072: out = -269;
			18073: out = -267;
			18074: out = -257;
			18075: out = -249;
			18076: out = -247;
			18077: out = -259;
			18078: out = -243;
			18079: out = -238;
			18080: out = -241;
			18081: out = -244;
			18082: out = -225;
			18083: out = -244;
			18084: out = -220;
			18085: out = -234;
			18086: out = -216;
			18087: out = -228;
			18088: out = -214;
			18089: out = -217;
			18090: out = -216;
			18091: out = -207;
			18092: out = -217;
			18093: out = -204;
			18094: out = -197;
			18095: out = -207;
			18096: out = -195;
			18097: out = -199;
			18098: out = -185;
			18099: out = -202;
			18100: out = -183;
			18101: out = -186;
			18102: out = -191;
			18103: out = -178;
			18104: out = -183;
			18105: out = -174;
			18106: out = -171;
			18107: out = -179;
			18108: out = -162;
			18109: out = -171;
			18110: out = -163;
			18111: out = -168;
			18112: out = -150;
			18113: out = -170;
			18114: out = -152;
			18115: out = -157;
			18116: out = -150;
			18117: out = -147;
			18118: out = -156;
			18119: out = -145;
			18120: out = -143;
			18121: out = -143;
			18122: out = -140;
			18123: out = -138;
			18124: out = -137;
			18125: out = -135;
			18126: out = -135;
			18127: out = -135;
			18128: out = -134;
			18129: out = -131;
			18130: out = -128;
			18131: out = -120;
			18132: out = -120;
			18133: out = -126;
			18134: out = -115;
			18135: out = -108;
			18136: out = -120;
			18137: out = -102;
			18138: out = -105;
			18139: out = -96;
			18140: out = -95;
			18141: out = -103;
			18142: out = -96;
			18143: out = -79;
			18144: out = -98;
			18145: out = -76;
			18146: out = -85;
			18147: out = -72;
			18148: out = -75;
			18149: out = -81;
			18150: out = -67;
			18151: out = -67;
			18152: out = -73;
			18153: out = -56;
			18154: out = -65;
			18155: out = -64;
			18156: out = -52;
			18157: out = -62;
			18158: out = -44;
			18159: out = -67;
			18160: out = -44;
			18161: out = -49;
			18162: out = -49;
			18163: out = -49;
			18164: out = -36;
			18165: out = -45;
			18166: out = -42;
			18167: out = -30;
			18168: out = -36;
			18169: out = -36;
			18170: out = -30;
			18171: out = -29;
			18172: out = -24;
			18173: out = -28;
			18174: out = -18;
			18175: out = -16;
			18176: out = -25;
			18177: out = -18;
			18178: out = -17;
			18179: out = -10;
			18180: out = -15;
			18181: out = -12;
			18182: out = -8;
			18183: out = -4;
			18184: out = -1;
			18185: out = -6;
			18186: out = 1;
			18187: out = -4;
			18188: out = 2;
			18189: out = 6;
			18190: out = 9;
			18191: out = 9;
			18192: out = 4;
			18193: out = 17;
			18194: out = 5;
			18195: out = 17;
			18196: out = 21;
			18197: out = 2;
			18198: out = 30;
			18199: out = 25;
			18200: out = 19;
			18201: out = 30;
			18202: out = 22;
			18203: out = 37;
			18204: out = 32;
			18205: out = 19;
			18206: out = 41;
			18207: out = 34;
			18208: out = 36;
			18209: out = 45;
			18210: out = 37;
			18211: out = 49;
			18212: out = 42;
			18213: out = 48;
			18214: out = 44;
			18215: out = 56;
			18216: out = 43;
			18217: out = 53;
			18218: out = 51;
			18219: out = 65;
			18220: out = 51;
			18221: out = 66;
			18222: out = 63;
			18223: out = 68;
			18224: out = 62;
			18225: out = 72;
			18226: out = 74;
			18227: out = 72;
			18228: out = 79;
			18229: out = 80;
			18230: out = 74;
			18231: out = 90;
			18232: out = 86;
			18233: out = 81;
			18234: out = 99;
			18235: out = 84;
			18236: out = 111;
			18237: out = 91;
			18238: out = 103;
			18239: out = 102;
			18240: out = 116;
			18241: out = 109;
			18242: out = 115;
			18243: out = 119;
			18244: out = 128;
			18245: out = 126;
			18246: out = 115;
			18247: out = 136;
			18248: out = 136;
			18249: out = 129;
			18250: out = 139;
			18251: out = 144;
			18252: out = 143;
			18253: out = 145;
			18254: out = 160;
			18255: out = 150;
			18256: out = 155;
			18257: out = 167;
			18258: out = 168;
			18259: out = 168;
			18260: out = 174;
			18261: out = 160;
			18262: out = 175;
			18263: out = 186;
			18264: out = 179;
			18265: out = 187;
			18266: out = 193;
			18267: out = 191;
			18268: out = 203;
			18269: out = 193;
			18270: out = 206;
			18271: out = 207;
			18272: out = 211;
			18273: out = 206;
			18274: out = 214;
			18275: out = 209;
			18276: out = 218;
			18277: out = 222;
			18278: out = 214;
			18279: out = 223;
			18280: out = 232;
			18281: out = 230;
			18282: out = 231;
			18283: out = 238;
			18284: out = 241;
			18285: out = 241;
			18286: out = 246;
			18287: out = 243;
			18288: out = 253;
			18289: out = 251;
			18290: out = 256;
			18291: out = 251;
			18292: out = 262;
			18293: out = 265;
			18294: out = 270;
			18295: out = 262;
			18296: out = 277;
			18297: out = 274;
			18298: out = 267;
			18299: out = 278;
			18300: out = 283;
			18301: out = 265;
			18302: out = 282;
			18303: out = 283;
			18304: out = 283;
			18305: out = 282;
			18306: out = 288;
			18307: out = 293;
			18308: out = 294;
			18309: out = 291;
			18310: out = 298;
			18311: out = 294;
			18312: out = 291;
			18313: out = 312;
			18314: out = 303;
			18315: out = 302;
			18316: out = 306;
			18317: out = 313;
			18318: out = 309;
			18319: out = 315;
			18320: out = 312;
			18321: out = 306;
			18322: out = 318;
			18323: out = 322;
			18324: out = 322;
			18325: out = 314;
			18326: out = 336;
			18327: out = 320;
			18328: out = 322;
			18329: out = 327;
			18330: out = 335;
			18331: out = 330;
			18332: out = 327;
			18333: out = 330;
			18334: out = 342;
			18335: out = 334;
			18336: out = 340;
			18337: out = 335;
			18338: out = 344;
			18339: out = 346;
			18340: out = 338;
			18341: out = 347;
			18342: out = 357;
			18343: out = 339;
			18344: out = 347;
			18345: out = 357;
			18346: out = 346;
			18347: out = 356;
			18348: out = 348;
			18349: out = 360;
			18350: out = 352;
			18351: out = 349;
			18352: out = 361;
			18353: out = 364;
			18354: out = 362;
			18355: out = 352;
			18356: out = 367;
			18357: out = 367;
			18358: out = 369;
			18359: out = 364;
			18360: out = 369;
			18361: out = 371;
			18362: out = 367;
			18363: out = 373;
			18364: out = 380;
			18365: out = 361;
			18366: out = 374;
			18367: out = 372;
			18368: out = 380;
			18369: out = 368;
			18370: out = 374;
			18371: out = 376;
			18372: out = 364;
			18373: out = 369;
			18374: out = 373;
			18375: out = 375;
			18376: out = 367;
			18377: out = 367;
			18378: out = 367;
			18379: out = 375;
			18380: out = 363;
			18381: out = 361;
			18382: out = 368;
			18383: out = 367;
			18384: out = 374;
			18385: out = 363;
			18386: out = 361;
			18387: out = 376;
			18388: out = 372;
			18389: out = 363;
			18390: out = 367;
			18391: out = 363;
			18392: out = 374;
			18393: out = 357;
			18394: out = 363;
			18395: out = 364;
			18396: out = 373;
			18397: out = 359;
			18398: out = 351;
			18399: out = 376;
			18400: out = 348;
			18401: out = 369;
			18402: out = 361;
			18403: out = 358;
			18404: out = 358;
			18405: out = 373;
			18406: out = 360;
			18407: out = 362;
			18408: out = 359;
			18409: out = 364;
			18410: out = 356;
			18411: out = 357;
			18412: out = 364;
			18413: out = 353;
			18414: out = 365;
			18415: out = 360;
			18416: out = 363;
			18417: out = 354;
			18418: out = 367;
			18419: out = 358;
			18420: out = 352;
			18421: out = 360;
			18422: out = 351;
			18423: out = 354;
			18424: out = 361;
			18425: out = 351;
			18426: out = 357;
			18427: out = 350;
			18428: out = 361;
			18429: out = 354;
			18430: out = 356;
			18431: out = 357;
			18432: out = 351;
			18433: out = 357;
			18434: out = 356;
			18435: out = 344;
			18436: out = 357;
			18437: out = 339;
			18438: out = 345;
			18439: out = 351;
			18440: out = 342;
			18441: out = 348;
			18442: out = 346;
			18443: out = 342;
			18444: out = 341;
			18445: out = 344;
			18446: out = 335;
			18447: out = 329;
			18448: out = 330;
			18449: out = 345;
			18450: out = 318;
			18451: out = 329;
			18452: out = 333;
			18453: out = 321;
			18454: out = 329;
			18455: out = 325;
			18456: out = 317;
			18457: out = 320;
			18458: out = 317;
			18459: out = 324;
			18460: out = 311;
			18461: out = 304;
			18462: out = 315;
			18463: out = 309;
			18464: out = 308;
			18465: out = 302;
			18466: out = 309;
			18467: out = 304;
			18468: out = 306;
			18469: out = 291;
			18470: out = 302;
			18471: out = 292;
			18472: out = 281;
			18473: out = 290;
			18474: out = 287;
			18475: out = 265;
			18476: out = 288;
			18477: out = 271;
			18478: out = 276;
			18479: out = 263;
			18480: out = 269;
			18481: out = 267;
			18482: out = 258;
			18483: out = 265;
			18484: out = 256;
			18485: out = 257;
			18486: out = 246;
			18487: out = 261;
			18488: out = 235;
			18489: out = 255;
			18490: out = 239;
			18491: out = 243;
			18492: out = 232;
			18493: out = 237;
			18494: out = 234;
			18495: out = 230;
			18496: out = 219;
			18497: out = 225;
			18498: out = 221;
			18499: out = 220;
			18500: out = 210;
			18501: out = 214;
			18502: out = 210;
			18503: out = 215;
			18504: out = 202;
			18505: out = 207;
			18506: out = 197;
			18507: out = 202;
			18508: out = 187;
			18509: out = 195;
			18510: out = 175;
			18511: out = 199;
			18512: out = 171;
			18513: out = 187;
			18514: out = 181;
			18515: out = 172;
			18516: out = 178;
			18517: out = 172;
			18518: out = 172;
			18519: out = 168;
			18520: out = 167;
			18521: out = 161;
			18522: out = 167;
			18523: out = 160;
			18524: out = 150;
			18525: out = 146;
			18526: out = 154;
			18527: out = 148;
			18528: out = 143;
			18529: out = 141;
			18530: out = 146;
			18531: out = 139;
			18532: out = 133;
			18533: out = 140;
			18534: out = 137;
			18535: out = 126;
			18536: out = 131;
			18537: out = 127;
			18538: out = 122;
			18539: out = 124;
			18540: out = 112;
			18541: out = 122;
			18542: out = 119;
			18543: out = 114;
			18544: out = 119;
			18545: out = 110;
			18546: out = 116;
			18547: out = 102;
			18548: out = 100;
			18549: out = 108;
			18550: out = 103;
			18551: out = 98;
			18552: out = 97;
			18553: out = 103;
			18554: out = 88;
			18555: out = 100;
			18556: out = 85;
			18557: out = 90;
			18558: out = 89;
			18559: out = 87;
			18560: out = 83;
			18561: out = 73;
			18562: out = 88;
			18563: out = 74;
			18564: out = 81;
			18565: out = 67;
			18566: out = 80;
			18567: out = 68;
			18568: out = 80;
			18569: out = 63;
			18570: out = 76;
			18571: out = 67;
			18572: out = 68;
			18573: out = 62;
			18574: out = 64;
			18575: out = 57;
			18576: out = 63;
			18577: out = 50;
			18578: out = 61;
			18579: out = 50;
			18580: out = 52;
			18581: out = 52;
			18582: out = 50;
			18583: out = 48;
			18584: out = 48;
			18585: out = 46;
			18586: out = 46;
			18587: out = 44;
			18588: out = 48;
			18589: out = 37;
			18590: out = 38;
			18591: out = 43;
			18592: out = 36;
			18593: out = 34;
			18594: out = 34;
			18595: out = 36;
			18596: out = 36;
			18597: out = 32;
			18598: out = 29;
			18599: out = 28;
			18600: out = 30;
			18601: out = 20;
			18602: out = 17;
			18603: out = 14;
			18604: out = 6;
			18605: out = 14;
			18606: out = -1;
			18607: out = 2;
			18608: out = 2;
			18609: out = -4;
			18610: out = -10;
			18611: out = -9;
			18612: out = -5;
			18613: out = -29;
			18614: out = -10;
			18615: out = -19;
			18616: out = -16;
			18617: out = -31;
			18618: out = -24;
			18619: out = -31;
			18620: out = -24;
			18621: out = -39;
			18622: out = -27;
			18623: out = -38;
			18624: out = -42;
			18625: out = -43;
			18626: out = -49;
			18627: out = -45;
			18628: out = -54;
			18629: out = -54;
			18630: out = -54;
			18631: out = -55;
			18632: out = -55;
			18633: out = -61;
			18634: out = -60;
			18635: out = -64;
			18636: out = -67;
			18637: out = -68;
			18638: out = -69;
			18639: out = -74;
			18640: out = -83;
			18641: out = -76;
			18642: out = -74;
			18643: out = -84;
			18644: out = -83;
			18645: out = -87;
			18646: out = -80;
			18647: out = -85;
			18648: out = -86;
			18649: out = -95;
			18650: out = -89;
			18651: out = -88;
			18652: out = -109;
			18653: out = -102;
			18654: out = -91;
			18655: out = -107;
			18656: out = -109;
			18657: out = -100;
			18658: out = -104;
			18659: out = -109;
			18660: out = -116;
			18661: out = -103;
			18662: out = -122;
			18663: out = -120;
			18664: out = -110;
			18665: out = -132;
			18666: out = -116;
			18667: out = -124;
			18668: out = -128;
			18669: out = -124;
			18670: out = -129;
			18671: out = -132;
			18672: out = -134;
			18673: out = -132;
			18674: out = -134;
			18675: out = -135;
			18676: out = -151;
			18677: out = -133;
			18678: out = -141;
			18679: out = -158;
			18680: out = -144;
			18681: out = -148;
			18682: out = -150;
			18683: out = -152;
			18684: out = -159;
			18685: out = -148;
			18686: out = -163;
			18687: out = -157;
			18688: out = -166;
			18689: out = -168;
			18690: out = -164;
			18691: out = -171;
			18692: out = -166;
			18693: out = -174;
			18694: out = -176;
			18695: out = -172;
			18696: out = -183;
			18697: out = -182;
			18698: out = -179;
			18699: out = -186;
			18700: out = -192;
			18701: out = -190;
			18702: out = -190;
			18703: out = -197;
			18704: out = -196;
			18705: out = -208;
			18706: out = -204;
			18707: out = -217;
			18708: out = -203;
			18709: out = -221;
			18710: out = -203;
			18711: out = -230;
			18712: out = -217;
			18713: out = -225;
			18714: out = -229;
			18715: out = -232;
			18716: out = -234;
			18717: out = -242;
			18718: out = -237;
			18719: out = -242;
			18720: out = -249;
			18721: out = -246;
			18722: out = -254;
			18723: out = -256;
			18724: out = -256;
			18725: out = -266;
			18726: out = -258;
			18727: out = -278;
			18728: out = -273;
			18729: out = -273;
			18730: out = -288;
			18731: out = -290;
			18732: out = -289;
			18733: out = -286;
			18734: out = -293;
			18735: out = -300;
			18736: out = -299;
			18737: out = -301;
			18738: out = -306;
			18739: out = -308;
			18740: out = -313;
			18741: out = -321;
			18742: out = -310;
			18743: out = -327;
			18744: out = -336;
			18745: out = -323;
			18746: out = -333;
			18747: out = -334;
			18748: out = -342;
			18749: out = -339;
			18750: out = -348;
			18751: out = -340;
			18752: out = -360;
			18753: out = -348;
			18754: out = -358;
			18755: out = -362;
			18756: out = -359;
			18757: out = -361;
			18758: out = -367;
			18759: out = -370;
			18760: out = -367;
			18761: out = -374;
			18762: out = -373;
			18763: out = -374;
			18764: out = -380;
			18765: out = -384;
			18766: out = -377;
			18767: out = -381;
			18768: out = -386;
			18769: out = -386;
			18770: out = -388;
			18771: out = -392;
			18772: out = -396;
			18773: out = -382;
			18774: out = -409;
			18775: out = -386;
			18776: out = -407;
			18777: out = -385;
			18778: out = -401;
			18779: out = -408;
			18780: out = -394;
			18781: out = -404;
			18782: out = -410;
			18783: out = -406;
			18784: out = -403;
			18785: out = -408;
			18786: out = -408;
			18787: out = -417;
			18788: out = -407;
			18789: out = -413;
			18790: out = -416;
			18791: out = -408;
			18792: out = -422;
			18793: out = -420;
			18794: out = -418;
			18795: out = -419;
			18796: out = -417;
			18797: out = -425;
			18798: out = -419;
			18799: out = -422;
			18800: out = -415;
			18801: out = -428;
			18802: out = -429;
			18803: out = -419;
			18804: out = -427;
			18805: out = -421;
			18806: out = -432;
			18807: out = -420;
			18808: out = -425;
			18809: out = -420;
			18810: out = -427;
			18811: out = -418;
			18812: out = -423;
			18813: out = -420;
			18814: out = -422;
			18815: out = -429;
			18816: out = -411;
			18817: out = -430;
			18818: out = -430;
			18819: out = -423;
			18820: out = -420;
			18821: out = -423;
			18822: out = -439;
			18823: out = -417;
			18824: out = -428;
			18825: out = -422;
			18826: out = -430;
			18827: out = -418;
			18828: out = -427;
			18829: out = -419;
			18830: out = -424;
			18831: out = -422;
			18832: out = -419;
			18833: out = -417;
			18834: out = -436;
			18835: out = -418;
			18836: out = -416;
			18837: out = -425;
			18838: out = -420;
			18839: out = -423;
			18840: out = -421;
			18841: out = -419;
			18842: out = -419;
			18843: out = -413;
			18844: out = -422;
			18845: out = -413;
			18846: out = -413;
			18847: out = -425;
			18848: out = -415;
			18849: out = -420;
			18850: out = -404;
			18851: out = -418;
			18852: out = -419;
			18853: out = -407;
			18854: out = -405;
			18855: out = -417;
			18856: out = -408;
			18857: out = -405;
			18858: out = -411;
			18859: out = -400;
			18860: out = -411;
			18861: out = -406;
			18862: out = -400;
			18863: out = -404;
			18864: out = -407;
			18865: out = -407;
			18866: out = -392;
			18867: out = -411;
			18868: out = -397;
			18869: out = -400;
			18870: out = -397;
			18871: out = -398;
			18872: out = -400;
			18873: out = -393;
			18874: out = -395;
			18875: out = -391;
			18876: out = -399;
			18877: out = -401;
			18878: out = -381;
			18879: out = -401;
			18880: out = -382;
			18881: out = -393;
			18882: out = -393;
			18883: out = -380;
			18884: out = -388;
			18885: out = -379;
			18886: out = -384;
			18887: out = -376;
			18888: out = -381;
			18889: out = -373;
			18890: out = -381;
			18891: out = -380;
			18892: out = -377;
			18893: out = -371;
			18894: out = -382;
			18895: out = -371;
			18896: out = -377;
			18897: out = -369;
			18898: out = -361;
			18899: out = -370;
			18900: out = -365;
			18901: out = -364;
			18902: out = -354;
			18903: out = -362;
			18904: out = -363;
			18905: out = -360;
			18906: out = -353;
			18907: out = -353;
			18908: out = -356;
			18909: out = -351;
			18910: out = -341;
			18911: out = -338;
			18912: out = -356;
			18913: out = -337;
			18914: out = -335;
			18915: out = -345;
			18916: out = -332;
			18917: out = -327;
			18918: out = -341;
			18919: out = -330;
			18920: out = -322;
			18921: out = -320;
			18922: out = -330;
			18923: out = -316;
			18924: out = -316;
			18925: out = -318;
			18926: out = -300;
			18927: out = -324;
			18928: out = -304;
			18929: out = -302;
			18930: out = -302;
			18931: out = -296;
			18932: out = -293;
			18933: out = -293;
			18934: out = -289;
			18935: out = -293;
			18936: out = -278;
			18937: out = -277;
			18938: out = -291;
			18939: out = -271;
			18940: out = -275;
			18941: out = -265;
			18942: out = -273;
			18943: out = -269;
			18944: out = -256;
			18945: out = -265;
			18946: out = -262;
			18947: out = -252;
			18948: out = -252;
			18949: out = -258;
			18950: out = -241;
			18951: out = -249;
			18952: out = -250;
			18953: out = -238;
			18954: out = -235;
			18955: out = -244;
			18956: out = -232;
			18957: out = -225;
			18958: out = -235;
			18959: out = -220;
			18960: out = -219;
			18961: out = -218;
			18962: out = -227;
			18963: out = -208;
			18964: out = -210;
			18965: out = -208;
			18966: out = -200;
			18967: out = -216;
			18968: out = -200;
			18969: out = -203;
			18970: out = -194;
			18971: out = -196;
			18972: out = -205;
			18973: out = -181;
			18974: out = -188;
			18975: out = -180;
			18976: out = -191;
			18977: out = -178;
			18978: out = -174;
			18979: out = -175;
			18980: out = -176;
			18981: out = -171;
			18982: out = -168;
			18983: out = -163;
			18984: out = -179;
			18985: out = -159;
			18986: out = -161;
			18987: out = -161;
			18988: out = -172;
			18989: out = -143;
			18990: out = -171;
			18991: out = -146;
			18992: out = -159;
			18993: out = -148;
			18994: out = -150;
			18995: out = -154;
			18996: out = -144;
			18997: out = -154;
			18998: out = -132;
			18999: out = -148;
			19000: out = -141;
			19001: out = -136;
			19002: out = -135;
			19003: out = -136;
			19004: out = -132;
			19005: out = -131;
			19006: out = -127;
			19007: out = -128;
			19008: out = -119;
			19009: out = -122;
			19010: out = -127;
			19011: out = -121;
			19012: out = -110;
			19013: out = -126;
			19014: out = -115;
			19015: out = -115;
			19016: out = -120;
			19017: out = -109;
			19018: out = -112;
			19019: out = -107;
			19020: out = -113;
			19021: out = -99;
			19022: out = -108;
			19023: out = -97;
			19024: out = -102;
			19025: out = -91;
			19026: out = -102;
			19027: out = -85;
			19028: out = -88;
			19029: out = -87;
			19030: out = -88;
			19031: out = -75;
			19032: out = -90;
			19033: out = -81;
			19034: out = -74;
			19035: out = -85;
			19036: out = -66;
			19037: out = -76;
			19038: out = -74;
			19039: out = -67;
			19040: out = -63;
			19041: out = -62;
			19042: out = -68;
			19043: out = -56;
			19044: out = -51;
			19045: out = -63;
			19046: out = -58;
			19047: out = -48;
			19048: out = -51;
			19049: out = -50;
			19050: out = -40;
			19051: out = -55;
			19052: out = -39;
			19053: out = -46;
			19054: out = -37;
			19055: out = -39;
			19056: out = -46;
			19057: out = -33;
			19058: out = -30;
			19059: out = -38;
			19060: out = -25;
			19061: out = -33;
			19062: out = -19;
			19063: out = -24;
			19064: out = -27;
			19065: out = -22;
			19066: out = -25;
			19067: out = -26;
			19068: out = -18;
			19069: out = -17;
			19070: out = -27;
			19071: out = -6;
			19072: out = -19;
			19073: out = -12;
			19074: out = -16;
			19075: out = -16;
			19076: out = -8;
			19077: out = -14;
			19078: out = -8;
			19079: out = -10;
			19080: out = 1;
			19081: out = -7;
			19082: out = -1;
			19083: out = 3;
			19084: out = -2;
			19085: out = 0;
			19086: out = 1;
			19087: out = 7;
			19088: out = 2;
			19089: out = 7;
			19090: out = 9;
			19091: out = 12;
			19092: out = 16;
			19093: out = 3;
			19094: out = 15;
			19095: out = 17;
			19096: out = 22;
			19097: out = 13;
			19098: out = 22;
			19099: out = 14;
			19100: out = 33;
			19101: out = 16;
			19102: out = 26;
			19103: out = 26;
			19104: out = 27;
			19105: out = 24;
			19106: out = 27;
			19107: out = 39;
			19108: out = 21;
			19109: out = 39;
			19110: out = 36;
			19111: out = 28;
			19112: out = 44;
			19113: out = 34;
			19114: out = 38;
			19115: out = 46;
			19116: out = 38;
			19117: out = 49;
			19118: out = 46;
			19119: out = 51;
			19120: out = 52;
			19121: out = 46;
			19122: out = 58;
			19123: out = 69;
			19124: out = 49;
			19125: out = 66;
			19126: out = 68;
			19127: out = 65;
			19128: out = 72;
			19129: out = 68;
			19130: out = 76;
			19131: out = 72;
			19132: out = 79;
			19133: out = 75;
			19134: out = 85;
			19135: out = 89;
			19136: out = 80;
			19137: out = 98;
			19138: out = 91;
			19139: out = 100;
			19140: out = 96;
			19141: out = 91;
			19142: out = 112;
			19143: out = 97;
			19144: out = 105;
			19145: out = 103;
			19146: out = 119;
			19147: out = 115;
			19148: out = 112;
			19149: out = 121;
			19150: out = 127;
			19151: out = 123;
			19152: out = 124;
			19153: out = 128;
			19154: out = 132;
			19155: out = 136;
			19156: out = 127;
			19157: out = 137;
			19158: out = 138;
			19159: out = 146;
			19160: out = 135;
			19161: out = 156;
			19162: out = 145;
			19163: out = 145;
			19164: out = 154;
			19165: out = 163;
			19166: out = 160;
			19167: out = 154;
			19168: out = 163;
			19169: out = 166;
			19170: out = 174;
			19171: out = 166;
			19172: out = 170;
			19173: out = 168;
			19174: out = 185;
			19175: out = 176;
			19176: out = 172;
			19177: out = 186;
			19178: out = 181;
			19179: out = 184;
			19180: out = 186;
			19181: out = 185;
			19182: out = 188;
			19183: out = 199;
			19184: out = 190;
			19185: out = 200;
			19186: out = 193;
			19187: out = 197;
			19188: out = 200;
			19189: out = 203;
			19190: out = 200;
			19191: out = 205;
			19192: out = 203;
			19193: out = 206;
			19194: out = 215;
			19195: out = 219;
			19196: out = 208;
			19197: out = 210;
			19198: out = 222;
			19199: out = 217;
			19200: out = 220;
			19201: out = 219;
			19202: out = 222;
			19203: out = 225;
			19204: out = 227;
			19205: out = 226;
			19206: out = 229;
			19207: out = 239;
			19208: out = 216;
			19209: out = 230;
			19210: out = 242;
			19211: out = 230;
			19212: out = 240;
			19213: out = 234;
			19214: out = 233;
			19215: out = 243;
			19216: out = 247;
			19217: out = 234;
			19218: out = 251;
			19219: out = 239;
			19220: out = 255;
			19221: out = 245;
			19222: out = 243;
			19223: out = 245;
			19224: out = 256;
			19225: out = 255;
			19226: out = 244;
			19227: out = 255;
			19228: out = 255;
			19229: out = 263;
			19230: out = 244;
			19231: out = 261;
			19232: out = 252;
			19233: out = 258;
			19234: out = 265;
			19235: out = 252;
			19236: out = 269;
			19237: out = 258;
			19238: out = 264;
			19239: out = 262;
			19240: out = 263;
			19241: out = 274;
			19242: out = 257;
			19243: out = 268;
			19244: out = 273;
			19245: out = 267;
			19246: out = 276;
			19247: out = 265;
			19248: out = 273;
			19249: out = 275;
			19250: out = 277;
			19251: out = 270;
			19252: out = 270;
			19253: out = 281;
			19254: out = 268;
			19255: out = 275;
			19256: out = 275;
			19257: out = 268;
			19258: out = 287;
			19259: out = 262;
			19260: out = 282;
			19261: out = 270;
			19262: out = 276;
			19263: out = 269;
			19264: out = 278;
			19265: out = 273;
			19266: out = 285;
			19267: out = 271;
			19268: out = 275;
			19269: out = 271;
			19270: out = 268;
			19271: out = 282;
			19272: out = 255;
			19273: out = 266;
			19274: out = 271;
			19275: out = 271;
			19276: out = 267;
			19277: out = 259;
			19278: out = 276;
			19279: out = 266;
			19280: out = 267;
			19281: out = 273;
			19282: out = 262;
			19283: out = 269;
			19284: out = 274;
			19285: out = 265;
			19286: out = 273;
			19287: out = 266;
			19288: out = 262;
			19289: out = 266;
			19290: out = 271;
			19291: out = 257;
			19292: out = 261;
			19293: out = 267;
			19294: out = 263;
			19295: out = 271;
			19296: out = 254;
			19297: out = 275;
			19298: out = 258;
			19299: out = 266;
			19300: out = 267;
			19301: out = 259;
			19302: out = 267;
			19303: out = 269;
			19304: out = 256;
			19305: out = 274;
			19306: out = 258;
			19307: out = 264;
			19308: out = 268;
			19309: out = 255;
			19310: out = 264;
			19311: out = 267;
			19312: out = 253;
			19313: out = 269;
			19314: out = 254;
			19315: out = 259;
			19316: out = 261;
			19317: out = 254;
			19318: out = 255;
			19319: out = 261;
			19320: out = 251;
			19321: out = 254;
			19322: out = 258;
			19323: out = 246;
			19324: out = 265;
			19325: out = 239;
			19326: out = 255;
			19327: out = 252;
			19328: out = 250;
			19329: out = 249;
			19330: out = 255;
			19331: out = 249;
			19332: out = 246;
			19333: out = 255;
			19334: out = 240;
			19335: out = 242;
			19336: out = 252;
			19337: out = 239;
			19338: out = 242;
			19339: out = 245;
			19340: out = 237;
			19341: out = 245;
			19342: out = 239;
			19343: out = 233;
			19344: out = 240;
			19345: out = 239;
			19346: out = 235;
			19347: out = 234;
			19348: out = 238;
			19349: out = 225;
			19350: out = 241;
			19351: out = 216;
			19352: out = 222;
			19353: out = 228;
			19354: out = 223;
			19355: out = 218;
			19356: out = 223;
			19357: out = 214;
			19358: out = 218;
			19359: out = 218;
			19360: out = 203;
			19361: out = 209;
			19362: out = 200;
			19363: out = 212;
			19364: out = 194;
			19365: out = 212;
			19366: out = 197;
			19367: out = 190;
			19368: out = 207;
			19369: out = 190;
			19370: out = 195;
			19371: out = 190;
			19372: out = 183;
			19373: out = 200;
			19374: out = 182;
			19375: out = 181;
			19376: out = 184;
			19377: out = 183;
			19378: out = 169;
			19379: out = 181;
			19380: out = 175;
			19381: out = 170;
			19382: out = 168;
			19383: out = 167;
			19384: out = 161;
			19385: out = 166;
			19386: out = 158;
			19387: out = 158;
			19388: out = 157;
			19389: out = 157;
			19390: out = 158;
			19391: out = 143;
			19392: out = 158;
			19393: out = 144;
			19394: out = 143;
			19395: out = 144;
			19396: out = 136;
			19397: out = 147;
			19398: out = 136;
			19399: out = 129;
			19400: out = 139;
			19401: out = 132;
			19402: out = 123;
			19403: out = 126;
			19404: out = 128;
			19405: out = 114;
			19406: out = 127;
			19407: out = 119;
			19408: out = 116;
			19409: out = 119;
			19410: out = 115;
			19411: out = 101;
			19412: out = 115;
			19413: out = 104;
			19414: out = 103;
			19415: out = 104;
			19416: out = 107;
			19417: out = 91;
			19418: out = 103;
			19419: out = 99;
			19420: out = 89;
			19421: out = 100;
			19422: out = 88;
			19423: out = 96;
			19424: out = 86;
			19425: out = 95;
			19426: out = 89;
			19427: out = 89;
			19428: out = 79;
			19429: out = 85;
			19430: out = 79;
			19431: out = 83;
			19432: out = 68;
			19433: out = 78;
			19434: out = 73;
			19435: out = 74;
			19436: out = 84;
			19437: out = 53;
			19438: out = 67;
			19439: out = 62;
			19440: out = 73;
			19441: out = 57;
			19442: out = 57;
			19443: out = 61;
			19444: out = 60;
			19445: out = 51;
			19446: out = 58;
			19447: out = 53;
			19448: out = 49;
			19449: out = 51;
			19450: out = 50;
			19451: out = 56;
			19452: out = 41;
			19453: out = 49;
			19454: out = 49;
			19455: out = 46;
			19456: out = 42;
			19457: out = 41;
			19458: out = 40;
			19459: out = 39;
			19460: out = 37;
			19461: out = 37;
			19462: out = 43;
			19463: out = 29;
			19464: out = 41;
			19465: out = 31;
			19466: out = 25;
			19467: out = 37;
			19468: out = 37;
			19469: out = 21;
			19470: out = 30;
			19471: out = 22;
			19472: out = 29;
			19473: out = 24;
			19474: out = 25;
			19475: out = 21;
			19476: out = 16;
			19477: out = 28;
			19478: out = 20;
			19479: out = 17;
			19480: out = 25;
			19481: out = 13;
			19482: out = 15;
			19483: out = 8;
			19484: out = 25;
			19485: out = 9;
			19486: out = 12;
			19487: out = 5;
			19488: out = 9;
			19489: out = 10;
			19490: out = 6;
			19491: out = 4;
			19492: out = 2;
			19493: out = 8;
			19494: out = -9;
			19495: out = -4;
			19496: out = 1;
			19497: out = -18;
			19498: out = -7;
			19499: out = -15;
			19500: out = -16;
			19501: out = -13;
			19502: out = -26;
			19503: out = -17;
			19504: out = -30;
			19505: out = -21;
			19506: out = -32;
			19507: out = -20;
			19508: out = -41;
			19509: out = -25;
			19510: out = -40;
			19511: out = -29;
			19512: out = -38;
			19513: out = -41;
			19514: out = -46;
			19515: out = -43;
			19516: out = -29;
			19517: out = -61;
			19518: out = -43;
			19519: out = -48;
			19520: out = -49;
			19521: out = -52;
			19522: out = -56;
			19523: out = -55;
			19524: out = -53;
			19525: out = -55;
			19526: out = -49;
			19527: out = -68;
			19528: out = -57;
			19529: out = -55;
			19530: out = -63;
			19531: out = -70;
			19532: out = -61;
			19533: out = -68;
			19534: out = -72;
			19535: out = -74;
			19536: out = -77;
			19537: out = -67;
			19538: out = -83;
			19539: out = -75;
			19540: out = -72;
			19541: out = -79;
			19542: out = -84;
			19543: out = -79;
			19544: out = -80;
			19545: out = -86;
			19546: out = -89;
			19547: out = -92;
			19548: out = -96;
			19549: out = -87;
			19550: out = -95;
			19551: out = -88;
			19552: out = -105;
			19553: out = -86;
			19554: out = -100;
			19555: out = -95;
			19556: out = -104;
			19557: out = -98;
			19558: out = -100;
			19559: out = -104;
			19560: out = -113;
			19561: out = -100;
			19562: out = -112;
			19563: out = -108;
			19564: out = -122;
			19565: out = -105;
			19566: out = -120;
			19567: out = -116;
			19568: out = -117;
			19569: out = -113;
			19570: out = -131;
			19571: out = -112;
			19572: out = -127;
			19573: out = -113;
			19574: out = -127;
			19575: out = -134;
			19576: out = -120;
			19577: out = -131;
			19578: out = -134;
			19579: out = -132;
			19580: out = -132;
			19581: out = -137;
			19582: out = -138;
			19583: out = -137;
			19584: out = -137;
			19585: out = -140;
			19586: out = -145;
			19587: out = -145;
			19588: out = -143;
			19589: out = -150;
			19590: out = -152;
			19591: out = -152;
			19592: out = -156;
			19593: out = -156;
			19594: out = -161;
			19595: out = -157;
			19596: out = -163;
			19597: out = -168;
			19598: out = -166;
			19599: out = -169;
			19600: out = -175;
			19601: out = -173;
			19602: out = -175;
			19603: out = -171;
			19604: out = -174;
			19605: out = -191;
			19606: out = -182;
			19607: out = -180;
			19608: out = -193;
			19609: out = -187;
			19610: out = -190;
			19611: out = -207;
			19612: out = -187;
			19613: out = -205;
			19614: out = -200;
			19615: out = -205;
			19616: out = -215;
			19617: out = -200;
			19618: out = -225;
			19619: out = -211;
			19620: out = -226;
			19621: out = -214;
			19622: out = -227;
			19623: out = -219;
			19624: out = -239;
			19625: out = -220;
			19626: out = -239;
			19627: out = -238;
			19628: out = -243;
			19629: out = -235;
			19630: out = -244;
			19631: out = -245;
			19632: out = -250;
			19633: out = -250;
			19634: out = -251;
			19635: out = -267;
			19636: out = -254;
			19637: out = -273;
			19638: out = -263;
			19639: out = -265;
			19640: out = -271;
			19641: out = -261;
			19642: out = -282;
			19643: out = -263;
			19644: out = -282;
			19645: out = -271;
			19646: out = -276;
			19647: out = -290;
			19648: out = -279;
			19649: out = -280;
			19650: out = -288;
			19651: out = -286;
			19652: out = -279;
			19653: out = -296;
			19654: out = -291;
			19655: out = -292;
			19656: out = -286;
			19657: out = -304;
			19658: out = -297;
			19659: out = -298;
			19660: out = -300;
			19661: out = -300;
			19662: out = -306;
			19663: out = -302;
			19664: out = -305;
			19665: out = -305;
			19666: out = -310;
			19667: out = -304;
			19668: out = -312;
			19669: out = -314;
			19670: out = -313;
			19671: out = -300;
			19672: out = -316;
			19673: out = -314;
			19674: out = -308;
			19675: out = -316;
			19676: out = -324;
			19677: out = -310;
			19678: out = -318;
			19679: out = -321;
			19680: out = -313;
			19681: out = -323;
			19682: out = -321;
			19683: out = -317;
			19684: out = -322;
			19685: out = -317;
			19686: out = -315;
			19687: out = -329;
			19688: out = -322;
			19689: out = -323;
			19690: out = -324;
			19691: out = -317;
			19692: out = -333;
			19693: out = -323;
			19694: out = -320;
			19695: out = -325;
			19696: out = -323;
			19697: out = -328;
			19698: out = -320;
			19699: out = -323;
			19700: out = -333;
			19701: out = -321;
			19702: out = -324;
			19703: out = -328;
			19704: out = -328;
			19705: out = -329;
			19706: out = -327;
			19707: out = -334;
			19708: out = -326;
			19709: out = -330;
			19710: out = -332;
			19711: out = -328;
			19712: out = -323;
			19713: out = -332;
			19714: out = -332;
			19715: out = -329;
			19716: out = -318;
			19717: out = -329;
			19718: out = -335;
			19719: out = -321;
			19720: out = -327;
			19721: out = -320;
			19722: out = -337;
			19723: out = -329;
			19724: out = -313;
			19725: out = -333;
			19726: out = -329;
			19727: out = -320;
			19728: out = -321;
			19729: out = -333;
			19730: out = -323;
			19731: out = -320;
			19732: out = -330;
			19733: out = -326;
			19734: out = -322;
			19735: out = -330;
			19736: out = -320;
			19737: out = -328;
			19738: out = -320;
			19739: out = -324;
			19740: out = -328;
			19741: out = -314;
			19742: out = -321;
			19743: out = -318;
			19744: out = -321;
			19745: out = -322;
			19746: out = -324;
			19747: out = -317;
			19748: out = -321;
			19749: out = -326;
			19750: out = -309;
			19751: out = -327;
			19752: out = -309;
			19753: out = -318;
			19754: out = -314;
			19755: out = -313;
			19756: out = -316;
			19757: out = -310;
			19758: out = -305;
			19759: out = -326;
			19760: out = -309;
			19761: out = -301;
			19762: out = -321;
			19763: out = -313;
			19764: out = -305;
			19765: out = -313;
			19766: out = -310;
			19767: out = -306;
			19768: out = -310;
			19769: out = -305;
			19770: out = -298;
			19771: out = -320;
			19772: out = -309;
			19773: out = -299;
			19774: out = -311;
			19775: out = -288;
			19776: out = -316;
			19777: out = -298;
			19778: out = -297;
			19779: out = -300;
			19780: out = -299;
			19781: out = -297;
			19782: out = -300;
			19783: out = -287;
			19784: out = -298;
			19785: out = -300;
			19786: out = -288;
			19787: out = -288;
			19788: out = -296;
			19789: out = -291;
			19790: out = -286;
			19791: out = -286;
			19792: out = -293;
			19793: out = -283;
			19794: out = -286;
			19795: out = -283;
			19796: out = -285;
			19797: out = -277;
			19798: out = -273;
			19799: out = -275;
			19800: out = -283;
			19801: out = -269;
			19802: out = -279;
			19803: out = -273;
			19804: out = -266;
			19805: out = -276;
			19806: out = -273;
			19807: out = -258;
			19808: out = -262;
			19809: out = -266;
			19810: out = -261;
			19811: out = -249;
			19812: out = -268;
			19813: out = -256;
			19814: out = -245;
			19815: out = -261;
			19816: out = -250;
			19817: out = -250;
			19818: out = -247;
			19819: out = -244;
			19820: out = -241;
			19821: out = -241;
			19822: out = -238;
			19823: out = -242;
			19824: out = -219;
			19825: out = -234;
			19826: out = -239;
			19827: out = -221;
			19828: out = -227;
			19829: out = -219;
			19830: out = -225;
			19831: out = -216;
			19832: out = -212;
			19833: out = -215;
			19834: out = -214;
			19835: out = -210;
			19836: out = -207;
			19837: out = -204;
			19838: out = -203;
			19839: out = -199;
			19840: out = -203;
			19841: out = -193;
			19842: out = -197;
			19843: out = -195;
			19844: out = -190;
			19845: out = -197;
			19846: out = -181;
			19847: out = -194;
			19848: out = -179;
			19849: out = -183;
			19850: out = -183;
			19851: out = -178;
			19852: out = -175;
			19853: out = -175;
			19854: out = -172;
			19855: out = -167;
			19856: out = -171;
			19857: out = -163;
			19858: out = -169;
			19859: out = -164;
			19860: out = -150;
			19861: out = -169;
			19862: out = -168;
			19863: out = -143;
			19864: out = -162;
			19865: out = -151;
			19866: out = -152;
			19867: out = -144;
			19868: out = -156;
			19869: out = -143;
			19870: out = -143;
			19871: out = -140;
			19872: out = -135;
			19873: out = -148;
			19874: out = -145;
			19875: out = -124;
			19876: out = -146;
			19877: out = -125;
			19878: out = -131;
			19879: out = -132;
			19880: out = -131;
			19881: out = -121;
			19882: out = -124;
			19883: out = -136;
			19884: out = -119;
			19885: out = -121;
			19886: out = -117;
			19887: out = -123;
			19888: out = -121;
			19889: out = -119;
			19890: out = -103;
			19891: out = -120;
			19892: out = -116;
			19893: out = -109;
			19894: out = -111;
			19895: out = -112;
			19896: out = -103;
			19897: out = -112;
			19898: out = -105;
			19899: out = -99;
			19900: out = -104;
			19901: out = -101;
			19902: out = -92;
			19903: out = -103;
			19904: out = -105;
			19905: out = -95;
			19906: out = -90;
			19907: out = -95;
			19908: out = -104;
			19909: out = -85;
			19910: out = -100;
			19911: out = -81;
			19912: out = -88;
			19913: out = -89;
			19914: out = -88;
			19915: out = -84;
			19916: out = -85;
			19917: out = -80;
			19918: out = -78;
			19919: out = -85;
			19920: out = -79;
			19921: out = -67;
			19922: out = -76;
			19923: out = -73;
			19924: out = -70;
			19925: out = -68;
			19926: out = -74;
			19927: out = -68;
			19928: out = -61;
			19929: out = -68;
			19930: out = -57;
			19931: out = -65;
			19932: out = -48;
			19933: out = -61;
			19934: out = -58;
			19935: out = -52;
			19936: out = -46;
			19937: out = -45;
			19938: out = -54;
			19939: out = -45;
			19940: out = -49;
			19941: out = -37;
			19942: out = -44;
			19943: out = -56;
			19944: out = -36;
			19945: out = -38;
			19946: out = -37;
			19947: out = -37;
			19948: out = -37;
			19949: out = -31;
			19950: out = -38;
			19951: out = -32;
			19952: out = -31;
			19953: out = -34;
			19954: out = -24;
			19955: out = -42;
			19956: out = -21;
			19957: out = -24;
			19958: out = -30;
			19959: out = -22;
			19960: out = -25;
			19961: out = -24;
			19962: out = -20;
			19963: out = -17;
			19964: out = -20;
			19965: out = -22;
			19966: out = -14;
			19967: out = -16;
			19968: out = -18;
			19969: out = -17;
			19970: out = -18;
			19971: out = -4;
			19972: out = -20;
			19973: out = -15;
			19974: out = -5;
			19975: out = -5;
			19976: out = -9;
			19977: out = -5;
			19978: out = 0;
			19979: out = 6;
			19980: out = -13;
			19981: out = 4;
			19982: out = 5;
			19983: out = -10;
			19984: out = 1;
			19985: out = -4;
			19986: out = 14;
			19987: out = -3;
			19988: out = 3;
			19989: out = 14;
			19990: out = 0;
			19991: out = 8;
			19992: out = 14;
			19993: out = 10;
			19994: out = 15;
			19995: out = 15;
			19996: out = 14;
			19997: out = 12;
			19998: out = 25;
			19999: out = 7;
			20000: out = 13;
			20001: out = 33;
			20002: out = 13;
			20003: out = 18;
			20004: out = 28;
			20005: out = 29;
			20006: out = 22;
			20007: out = 29;
			20008: out = 28;
			20009: out = 24;
			20010: out = 33;
			20011: out = 36;
			20012: out = 30;
			20013: out = 38;
			20014: out = 37;
			20015: out = 40;
			20016: out = 43;
			20017: out = 46;
			20018: out = 43;
			20019: out = 45;
			20020: out = 50;
			20021: out = 51;
			20022: out = 41;
			20023: out = 55;
			20024: out = 53;
			20025: out = 55;
			20026: out = 55;
			20027: out = 58;
			20028: out = 66;
			20029: out = 56;
			20030: out = 68;
			20031: out = 64;
			20032: out = 69;
			20033: out = 62;
			20034: out = 78;
			20035: out = 64;
			20036: out = 77;
			20037: out = 74;
			20038: out = 85;
			20039: out = 80;
			20040: out = 83;
			20041: out = 87;
			20042: out = 87;
			20043: out = 93;
			20044: out = 86;
			20045: out = 92;
			20046: out = 87;
			20047: out = 100;
			20048: out = 95;
			20049: out = 105;
			20050: out = 96;
			20051: out = 109;
			20052: out = 100;
			20053: out = 108;
			20054: out = 112;
			20055: out = 110;
			20056: out = 98;
			20057: out = 122;
			20058: out = 111;
			20059: out = 122;
			20060: out = 113;
			20061: out = 115;
			20062: out = 126;
			20063: out = 121;
			20064: out = 122;
			20065: out = 128;
			20066: out = 131;
			20067: out = 120;
			20068: out = 136;
			20069: out = 129;
			20070: out = 128;
			20071: out = 132;
			20072: out = 139;
			20073: out = 124;
			20074: out = 141;
			20075: out = 141;
			20076: out = 134;
			20077: out = 144;
			20078: out = 127;
			20079: out = 150;
			20080: out = 143;
			20081: out = 145;
			20082: out = 140;
			20083: out = 156;
			20084: out = 146;
			20085: out = 155;
			20086: out = 154;
			20087: out = 146;
			20088: out = 157;
			20089: out = 161;
			20090: out = 143;
			20091: out = 157;
			20092: out = 156;
			20093: out = 157;
			20094: out = 171;
			20095: out = 159;
			20096: out = 155;
			20097: out = 167;
			20098: out = 166;
			20099: out = 167;
			20100: out = 166;
			20101: out = 161;
			20102: out = 166;
			20103: out = 173;
			20104: out = 167;
			20105: out = 170;
			20106: out = 174;
			20107: out = 170;
			20108: out = 174;
			20109: out = 171;
			20110: out = 176;
			20111: out = 164;
			20112: out = 182;
			20113: out = 171;
			20114: out = 176;
			20115: out = 183;
			20116: out = 164;
			20117: out = 178;
			20118: out = 182;
			20119: out = 185;
			20120: out = 182;
			20121: out = 180;
			20122: out = 185;
			20123: out = 180;
			20124: out = 179;
			20125: out = 196;
			20126: out = 172;
			20127: out = 186;
			20128: out = 188;
			20129: out = 188;
			20130: out = 193;
			20131: out = 185;
			20132: out = 191;
			20133: out = 188;
			20134: out = 188;
			20135: out = 194;
			20136: out = 194;
			20137: out = 191;
			20138: out = 196;
			20139: out = 184;
			20140: out = 198;
			20141: out = 192;
			20142: out = 196;
			20143: out = 186;
			20144: out = 199;
			20145: out = 195;
			20146: out = 188;
			20147: out = 195;
			20148: out = 199;
			20149: out = 190;
			20150: out = 204;
			20151: out = 194;
			20152: out = 188;
			20153: out = 202;
			20154: out = 185;
			20155: out = 209;
			20156: out = 183;
			20157: out = 192;
			20158: out = 202;
			20159: out = 196;
			20160: out = 190;
			20161: out = 198;
			20162: out = 196;
			20163: out = 194;
			20164: out = 199;
			20165: out = 188;
			20166: out = 188;
			20167: out = 193;
			20168: out = 194;
			20169: out = 183;
			20170: out = 195;
			20171: out = 192;
			20172: out = 179;
			20173: out = 199;
			20174: out = 190;
			20175: out = 181;
			20176: out = 198;
			20177: out = 181;
			20178: out = 194;
			20179: out = 192;
			20180: out = 179;
			20181: out = 192;
			20182: out = 191;
			20183: out = 183;
			20184: out = 192;
			20185: out = 190;
			20186: out = 181;
			20187: out = 192;
			20188: out = 183;
			20189: out = 188;
			20190: out = 179;
			20191: out = 183;
			20192: out = 187;
			20193: out = 188;
			20194: out = 188;
			20195: out = 174;
			20196: out = 195;
			20197: out = 182;
			20198: out = 183;
			20199: out = 192;
			20200: out = 173;
			20201: out = 179;
			20202: out = 190;
			20203: out = 179;
			20204: out = 185;
			20205: out = 181;
			20206: out = 183;
			20207: out = 181;
			20208: out = 183;
			20209: out = 187;
			20210: out = 185;
			20211: out = 170;
			20212: out = 185;
			20213: out = 183;
			20214: out = 175;
			20215: out = 170;
			20216: out = 183;
			20217: out = 181;
			20218: out = 167;
			20219: out = 178;
			20220: out = 176;
			20221: out = 174;
			20222: out = 173;
			20223: out = 170;
			20224: out = 162;
			20225: out = 169;
			20226: out = 172;
			20227: out = 167;
			20228: out = 164;
			20229: out = 164;
			20230: out = 171;
			20231: out = 168;
			20232: out = 164;
			20233: out = 161;
			20234: out = 167;
			20235: out = 158;
			20236: out = 172;
			20237: out = 158;
			20238: out = 161;
			20239: out = 161;
			20240: out = 149;
			20241: out = 166;
			20242: out = 151;
			20243: out = 157;
			20244: out = 154;
			20245: out = 156;
			20246: out = 158;
			20247: out = 146;
			20248: out = 148;
			20249: out = 152;
			20250: out = 141;
			20251: out = 150;
			20252: out = 143;
			20253: out = 140;
			20254: out = 144;
			20255: out = 139;
			20256: out = 139;
			20257: out = 136;
			20258: out = 138;
			20259: out = 124;
			20260: out = 140;
			20261: out = 123;
			20262: out = 139;
			20263: out = 116;
			20264: out = 119;
			20265: out = 125;
			20266: out = 125;
			20267: out = 115;
			20268: out = 116;
			20269: out = 124;
			20270: out = 110;
			20271: out = 116;
			20272: out = 114;
			20273: out = 102;
			20274: out = 105;
			20275: out = 114;
			20276: out = 102;
			20277: out = 104;
			20278: out = 110;
			20279: out = 99;
			20280: out = 107;
			20281: out = 97;
			20282: out = 105;
			20283: out = 97;
			20284: out = 98;
			20285: out = 92;
			20286: out = 93;
			20287: out = 86;
			20288: out = 98;
			20289: out = 90;
			20290: out = 79;
			20291: out = 87;
			20292: out = 91;
			20293: out = 78;
			20294: out = 84;
			20295: out = 75;
			20296: out = 76;
			20297: out = 78;
			20298: out = 76;
			20299: out = 67;
			20300: out = 75;
			20301: out = 69;
			20302: out = 69;
			20303: out = 77;
			20304: out = 63;
			20305: out = 74;
			20306: out = 54;
			20307: out = 66;
			20308: out = 70;
			20309: out = 57;
			20310: out = 54;
			20311: out = 65;
			20312: out = 62;
			20313: out = 69;
			20314: out = 48;
			20315: out = 57;
			20316: out = 62;
			20317: out = 54;
			20318: out = 46;
			20319: out = 53;
			20320: out = 50;
			20321: out = 52;
			20322: out = 36;
			20323: out = 52;
			20324: out = 38;
			20325: out = 46;
			20326: out = 32;
			20327: out = 49;
			20328: out = 33;
			20329: out = 34;
			20330: out = 40;
			20331: out = 34;
			20332: out = 44;
			20333: out = 22;
			20334: out = 37;
			20335: out = 29;
			20336: out = 40;
			20337: out = 34;
			20338: out = 15;
			20339: out = 39;
			20340: out = 24;
			20341: out = 40;
			20342: out = 14;
			20343: out = 28;
			20344: out = 26;
			20345: out = 32;
			20346: out = 18;
			20347: out = 25;
			20348: out = 28;
			20349: out = 28;
			20350: out = 14;
			20351: out = 17;
			20352: out = 15;
			20353: out = 26;
			20354: out = 3;
			20355: out = 22;
			20356: out = 12;
			20357: out = 7;
			20358: out = 10;
			20359: out = 7;
			20360: out = 12;
			20361: out = 1;
			20362: out = 9;
			20363: out = 7;
			20364: out = 8;
			20365: out = 9;
			20366: out = -5;
			20367: out = 6;
			20368: out = 6;
			20369: out = 4;
			20370: out = 0;
			20371: out = -3;
			20372: out = 8;
			20373: out = -2;
			20374: out = 7;
			20375: out = -9;
			20376: out = 10;
			20377: out = -3;
			20378: out = 1;
			20379: out = 4;
			20380: out = -14;
			20381: out = -1;
			20382: out = -5;
			20383: out = -6;
			20384: out = -8;
			20385: out = -13;
			20386: out = -8;
			20387: out = -24;
			20388: out = -4;
			20389: out = -24;
			20390: out = -13;
			20391: out = -22;
			20392: out = -21;
			20393: out = -31;
			20394: out = -27;
			20395: out = -28;
			20396: out = -27;
			20397: out = -36;
			20398: out = -29;
			20399: out = -34;
			20400: out = -37;
			20401: out = -33;
			20402: out = -39;
			20403: out = -45;
			20404: out = -45;
			20405: out = -38;
			20406: out = -37;
			20407: out = -55;
			20408: out = -42;
			20409: out = -49;
			20410: out = -42;
			20411: out = -48;
			20412: out = -54;
			20413: out = -45;
			20414: out = -53;
			20415: out = -57;
			20416: out = -49;
			20417: out = -53;
			20418: out = -54;
			20419: out = -64;
			20420: out = -43;
			20421: out = -67;
			20422: out = -58;
			20423: out = -56;
			20424: out = -69;
			20425: out = -62;
			20426: out = -63;
			20427: out = -63;
			20428: out = -64;
			20429: out = -69;
			20430: out = -65;
			20431: out = -67;
			20432: out = -77;
			20433: out = -73;
			20434: out = -67;
			20435: out = -72;
			20436: out = -78;
			20437: out = -74;
			20438: out = -77;
			20439: out = -85;
			20440: out = -74;
			20441: out = -85;
			20442: out = -79;
			20443: out = -85;
			20444: out = -75;
			20445: out = -81;
			20446: out = -92;
			20447: out = -76;
			20448: out = -86;
			20449: out = -102;
			20450: out = -78;
			20451: out = -92;
			20452: out = -83;
			20453: out = -100;
			20454: out = -91;
			20455: out = -84;
			20456: out = -100;
			20457: out = -96;
			20458: out = -87;
			20459: out = -93;
			20460: out = -101;
			20461: out = -98;
			20462: out = -99;
			20463: out = -95;
			20464: out = -101;
			20465: out = -111;
			20466: out = -104;
			20467: out = -103;
			20468: out = -104;
			20469: out = -115;
			20470: out = -103;
			20471: out = -112;
			20472: out = -103;
			20473: out = -122;
			20474: out = -105;
			20475: out = -114;
			20476: out = -112;
			20477: out = -115;
			20478: out = -126;
			20479: out = -110;
			20480: out = -122;
			20481: out = -114;
			20482: out = -121;
			20483: out = -132;
			20484: out = -120;
			20485: out = -119;
			20486: out = -132;
			20487: out = -127;
			20488: out = -132;
			20489: out = -131;
			20490: out = -125;
			20491: out = -141;
			20492: out = -139;
			20493: out = -128;
			20494: out = -136;
			20495: out = -148;
			20496: out = -137;
			20497: out = -145;
			20498: out = -143;
			20499: out = -146;
			20500: out = -160;
			20501: out = -145;
			20502: out = -148;
			20503: out = -157;
			20504: out = -152;
			20505: out = -161;
			20506: out = -154;
			20507: out = -167;
			20508: out = -159;
			20509: out = -174;
			20510: out = -171;
			20511: out = -167;
			20512: out = -167;
			20513: out = -184;
			20514: out = -172;
			20515: out = -173;
			20516: out = -173;
			20517: out = -185;
			20518: out = -179;
			20519: out = -188;
			20520: out = -185;
			20521: out = -183;
			20522: out = -195;
			20523: out = -187;
			20524: out = -197;
			20525: out = -193;
			20526: out = -204;
			20527: out = -202;
			20528: out = -200;
			20529: out = -198;
			20530: out = -204;
			20531: out = -206;
			20532: out = -207;
			20533: out = -202;
			20534: out = -218;
			20535: out = -206;
			20536: out = -207;
			20537: out = -211;
			20538: out = -223;
			20539: out = -204;
			20540: out = -222;
			20541: out = -225;
			20542: out = -214;
			20543: out = -227;
			20544: out = -222;
			20545: out = -222;
			20546: out = -230;
			20547: out = -226;
			20548: out = -225;
			20549: out = -232;
			20550: out = -229;
			20551: out = -233;
			20552: out = -233;
			20553: out = -240;
			20554: out = -225;
			20555: out = -243;
			20556: out = -233;
			20557: out = -237;
			20558: out = -237;
			20559: out = -230;
			20560: out = -235;
			20561: out = -240;
			20562: out = -242;
			20563: out = -243;
			20564: out = -233;
			20565: out = -244;
			20566: out = -254;
			20567: out = -233;
			20568: out = -241;
			20569: out = -243;
			20570: out = -253;
			20571: out = -234;
			20572: out = -250;
			20573: out = -246;
			20574: out = -249;
			20575: out = -249;
			20576: out = -253;
			20577: out = -247;
			20578: out = -250;
			20579: out = -247;
			20580: out = -245;
			20581: out = -257;
			20582: out = -252;
			20583: out = -250;
			20584: out = -245;
			20585: out = -247;
			20586: out = -263;
			20587: out = -245;
			20588: out = -254;
			20589: out = -258;
			20590: out = -247;
			20591: out = -261;
			20592: out = -252;
			20593: out = -256;
			20594: out = -245;
			20595: out = -255;
			20596: out = -251;
			20597: out = -257;
			20598: out = -241;
			20599: out = -259;
			20600: out = -261;
			20601: out = -251;
			20602: out = -246;
			20603: out = -256;
			20604: out = -253;
			20605: out = -246;
			20606: out = -251;
			20607: out = -245;
			20608: out = -257;
			20609: out = -251;
			20610: out = -251;
			20611: out = -252;
			20612: out = -250;
			20613: out = -253;
			20614: out = -254;
			20615: out = -250;
			20616: out = -251;
			20617: out = -255;
			20618: out = -252;
			20619: out = -249;
			20620: out = -253;
			20621: out = -252;
			20622: out = -254;
			20623: out = -253;
			20624: out = -255;
			20625: out = -244;
			20626: out = -259;
			20627: out = -241;
			20628: out = -255;
			20629: out = -239;
			20630: out = -254;
			20631: out = -247;
			20632: out = -243;
			20633: out = -251;
			20634: out = -253;
			20635: out = -237;
			20636: out = -256;
			20637: out = -251;
			20638: out = -245;
			20639: out = -238;
			20640: out = -252;
			20641: out = -244;
			20642: out = -235;
			20643: out = -245;
			20644: out = -245;
			20645: out = -244;
			20646: out = -242;
			20647: out = -243;
			20648: out = -240;
			20649: out = -237;
			20650: out = -240;
			20651: out = -241;
			20652: out = -238;
			20653: out = -244;
			20654: out = -230;
			20655: out = -238;
			20656: out = -241;
			20657: out = -234;
			20658: out = -237;
			20659: out = -234;
			20660: out = -242;
			20661: out = -226;
			20662: out = -249;
			20663: out = -233;
			20664: out = -233;
			20665: out = -234;
			20666: out = -230;
			20667: out = -237;
			20668: out = -233;
			20669: out = -229;
			20670: out = -223;
			20671: out = -239;
			20672: out = -223;
			20673: out = -229;
			20674: out = -242;
			20675: out = -216;
			20676: out = -230;
			20677: out = -230;
			20678: out = -222;
			20679: out = -229;
			20680: out = -210;
			20681: out = -234;
			20682: out = -221;
			20683: out = -220;
			20684: out = -214;
			20685: out = -232;
			20686: out = -209;
			20687: out = -226;
			20688: out = -207;
			20689: out = -220;
			20690: out = -222;
			20691: out = -218;
			20692: out = -214;
			20693: out = -210;
			20694: out = -212;
			20695: out = -211;
			20696: out = -209;
			20697: out = -204;
			20698: out = -206;
			20699: out = -210;
			20700: out = -196;
			20701: out = -209;
			20702: out = -197;
			20703: out = -210;
			20704: out = -184;
			20705: out = -198;
			20706: out = -199;
			20707: out = -191;
			20708: out = -194;
			20709: out = -192;
			20710: out = -188;
			20711: out = -190;
			20712: out = -186;
			20713: out = -180;
			20714: out = -192;
			20715: out = -182;
			20716: out = -180;
			20717: out = -184;
			20718: out = -186;
			20719: out = -174;
			20720: out = -176;
			20721: out = -182;
			20722: out = -173;
			20723: out = -172;
			20724: out = -176;
			20725: out = -166;
			20726: out = -171;
			20727: out = -168;
			20728: out = -161;
			20729: out = -161;
			20730: out = -158;
			20731: out = -160;
			20732: out = -164;
			20733: out = -151;
			20734: out = -154;
			20735: out = -157;
			20736: out = -143;
			20737: out = -152;
			20738: out = -148;
			20739: out = -149;
			20740: out = -136;
			20741: out = -148;
			20742: out = -139;
			20743: out = -140;
			20744: out = -129;
			20745: out = -144;
			20746: out = -133;
			20747: out = -133;
			20748: out = -137;
			20749: out = -132;
			20750: out = -123;
			20751: out = -139;
			20752: out = -117;
			20753: out = -141;
			20754: out = -122;
			20755: out = -125;
			20756: out = -133;
			20757: out = -115;
			20758: out = -126;
			20759: out = -117;
			20760: out = -121;
			20761: out = -112;
			20762: out = -119;
			20763: out = -115;
			20764: out = -115;
			20765: out = -120;
			20766: out = -119;
			20767: out = -101;
			20768: out = -119;
			20769: out = -105;
			20770: out = -110;
			20771: out = -102;
			20772: out = -111;
			20773: out = -99;
			20774: out = -102;
			20775: out = -105;
			20776: out = -101;
			20777: out = -96;
			20778: out = -101;
			20779: out = -93;
			20780: out = -97;
			20781: out = -105;
			20782: out = -93;
			20783: out = -100;
			20784: out = -85;
			20785: out = -98;
			20786: out = -96;
			20787: out = -90;
			20788: out = -83;
			20789: out = -83;
			20790: out = -92;
			20791: out = -85;
			20792: out = -81;
			20793: out = -89;
			20794: out = -86;
			20795: out = -81;
			20796: out = -80;
			20797: out = -86;
			20798: out = -83;
			20799: out = -72;
			20800: out = -80;
			20801: out = -75;
			20802: out = -77;
			20803: out = -69;
			20804: out = -77;
			20805: out = -66;
			20806: out = -69;
			20807: out = -75;
			20808: out = -66;
			20809: out = -69;
			20810: out = -72;
			20811: out = -75;
			20812: out = -56;
			20813: out = -67;
			20814: out = -58;
			20815: out = -66;
			20816: out = -52;
			20817: out = -62;
			20818: out = -51;
			20819: out = -61;
			20820: out = -60;
			20821: out = -57;
			20822: out = -43;
			20823: out = -53;
			20824: out = -51;
			20825: out = -50;
			20826: out = -45;
			20827: out = -50;
			20828: out = -52;
			20829: out = -42;
			20830: out = -48;
			20831: out = -40;
			20832: out = -45;
			20833: out = -38;
			20834: out = -34;
			20835: out = -41;
			20836: out = -42;
			20837: out = -40;
			20838: out = -39;
			20839: out = -33;
			20840: out = -31;
			20841: out = -38;
			20842: out = -37;
			20843: out = -27;
			20844: out = -30;
			20845: out = -27;
			20846: out = -33;
			20847: out = -34;
			20848: out = -28;
			20849: out = -20;
			20850: out = -31;
			20851: out = -28;
			20852: out = -21;
			20853: out = -21;
			20854: out = -25;
			20855: out = -18;
			20856: out = -26;
			20857: out = -26;
			20858: out = -20;
			20859: out = -19;
			20860: out = -19;
			20861: out = -21;
			20862: out = -22;
			20863: out = -12;
			20864: out = -21;
			20865: out = -17;
			20866: out = -16;
			20867: out = -8;
			20868: out = -9;
			20869: out = -25;
			20870: out = -8;
			20871: out = -6;
			20872: out = -10;
			20873: out = -13;
			20874: out = -7;
			20875: out = -10;
			20876: out = -9;
			20877: out = 0;
			20878: out = -15;
			20879: out = -1;
			20880: out = -8;
			20881: out = 2;
			20882: out = -5;
			20883: out = -8;
			20884: out = 0;
			20885: out = 0;
			20886: out = -1;
			20887: out = -7;
			20888: out = 2;
			20889: out = 7;
			20890: out = -6;
			20891: out = 4;
			20892: out = 10;
			20893: out = -9;
			20894: out = 19;
			20895: out = 1;
			20896: out = 7;
			20897: out = 5;
			20898: out = 7;
			20899: out = 18;
			20900: out = 6;
			20901: out = 17;
			20902: out = 6;
			20903: out = 24;
			20904: out = 12;
			20905: out = 21;
			20906: out = 21;
			20907: out = 19;
			20908: out = 22;
			20909: out = 20;
			20910: out = 22;
			20911: out = 25;
			20912: out = 26;
			20913: out = 22;
			20914: out = 28;
			20915: out = 28;
			20916: out = 29;
			20917: out = 24;
			20918: out = 32;
			20919: out = 36;
			20920: out = 37;
			20921: out = 36;
			20922: out = 31;
			20923: out = 41;
			20924: out = 38;
			20925: out = 40;
			20926: out = 45;
			20927: out = 38;
			20928: out = 49;
			20929: out = 55;
			20930: out = 45;
			20931: out = 46;
			20932: out = 54;
			20933: out = 63;
			20934: out = 52;
			20935: out = 57;
			20936: out = 64;
			20937: out = 58;
			20938: out = 51;
			20939: out = 74;
			20940: out = 58;
			20941: out = 62;
			20942: out = 65;
			20943: out = 73;
			20944: out = 64;
			20945: out = 70;
			20946: out = 68;
			20947: out = 74;
			20948: out = 68;
			20949: out = 76;
			20950: out = 70;
			20951: out = 84;
			20952: out = 74;
			20953: out = 69;
			20954: out = 89;
			20955: out = 70;
			20956: out = 81;
			20957: out = 84;
			20958: out = 87;
			20959: out = 77;
			20960: out = 85;
			20961: out = 95;
			20962: out = 86;
			20963: out = 89;
			20964: out = 90;
			20965: out = 89;
			20966: out = 95;
			20967: out = 100;
			20968: out = 90;
			20969: out = 97;
			20970: out = 97;
			20971: out = 102;
			20972: out = 102;
			20973: out = 91;
			20974: out = 104;
			20975: out = 105;
			20976: out = 97;
			20977: out = 103;
			20978: out = 101;
			20979: out = 110;
			20980: out = 107;
			20981: out = 101;
			20982: out = 113;
			20983: out = 107;
			20984: out = 108;
			20985: out = 105;
			20986: out = 116;
			20987: out = 108;
			20988: out = 108;
			20989: out = 116;
			20990: out = 109;
			20991: out = 114;
			20992: out = 115;
			20993: out = 115;
			20994: out = 104;
			20995: out = 122;
			20996: out = 113;
			20997: out = 113;
			20998: out = 117;
			20999: out = 117;
			21000: out = 123;
			21001: out = 111;
			21002: out = 125;
			21003: out = 116;
			21004: out = 121;
			21005: out = 120;
			21006: out = 125;
			21007: out = 128;
			21008: out = 117;
			21009: out = 125;
			21010: out = 125;
			21011: out = 125;
			21012: out = 116;
			21013: out = 128;
			21014: out = 119;
			21015: out = 127;
			21016: out = 128;
			21017: out = 117;
			21018: out = 128;
			21019: out = 123;
			21020: out = 133;
			21021: out = 122;
			21022: out = 131;
			21023: out = 127;
			21024: out = 133;
			21025: out = 135;
			21026: out = 121;
			21027: out = 131;
			21028: out = 128;
			21029: out = 141;
			21030: out = 119;
			21031: out = 131;
			21032: out = 133;
			21033: out = 128;
			21034: out = 139;
			21035: out = 121;
			21036: out = 134;
			21037: out = 129;
			21038: out = 144;
			21039: out = 122;
			21040: out = 132;
			21041: out = 134;
			21042: out = 128;
			21043: out = 120;
			21044: out = 141;
			21045: out = 127;
			21046: out = 127;
			21047: out = 135;
			21048: out = 127;
			21049: out = 133;
			21050: out = 128;
			21051: out = 129;
			21052: out = 127;
			21053: out = 117;
			21054: out = 140;
			21055: out = 123;
			21056: out = 121;
			21057: out = 133;
			21058: out = 128;
			21059: out = 125;
			21060: out = 125;
			21061: out = 126;
			21062: out = 125;
			21063: out = 121;
			21064: out = 135;
			21065: out = 124;
			21066: out = 123;
			21067: out = 123;
			21068: out = 132;
			21069: out = 121;
			21070: out = 124;
			21071: out = 116;
			21072: out = 128;
			21073: out = 129;
			21074: out = 121;
			21075: out = 123;
			21076: out = 132;
			21077: out = 128;
			21078: out = 115;
			21079: out = 129;
			21080: out = 124;
			21081: out = 113;
			21082: out = 127;
			21083: out = 115;
			21084: out = 124;
			21085: out = 119;
			21086: out = 122;
			21087: out = 125;
			21088: out = 117;
			21089: out = 124;
			21090: out = 117;
			21091: out = 123;
			21092: out = 122;
			21093: out = 110;
			21094: out = 120;
			21095: out = 117;
			21096: out = 122;
			21097: out = 116;
			21098: out = 122;
			21099: out = 112;
			21100: out = 121;
			21101: out = 120;
			21102: out = 117;
			21103: out = 115;
			21104: out = 122;
			21105: out = 109;
			21106: out = 127;
			21107: out = 111;
			21108: out = 121;
			21109: out = 115;
			21110: out = 113;
			21111: out = 116;
			21112: out = 117;
			21113: out = 110;
			21114: out = 113;
			21115: out = 116;
			21116: out = 112;
			21117: out = 107;
			21118: out = 114;
			21119: out = 112;
			21120: out = 105;
			21121: out = 113;
			21122: out = 108;
			21123: out = 104;
			21124: out = 109;
			21125: out = 110;
			21126: out = 101;
			21127: out = 100;
			21128: out = 98;
			21129: out = 101;
			21130: out = 109;
			21131: out = 98;
			21132: out = 103;
			21133: out = 101;
			21134: out = 98;
			21135: out = 108;
			21136: out = 87;
			21137: out = 95;
			21138: out = 104;
			21139: out = 96;
			21140: out = 99;
			21141: out = 89;
			21142: out = 98;
			21143: out = 95;
			21144: out = 97;
			21145: out = 86;
			21146: out = 88;
			21147: out = 91;
			21148: out = 97;
			21149: out = 80;
			21150: out = 88;
			21151: out = 80;
			21152: out = 92;
			21153: out = 83;
			21154: out = 81;
			21155: out = 80;
			21156: out = 79;
			21157: out = 78;
			21158: out = 75;
			21159: out = 78;
			21160: out = 72;
			21161: out = 77;
			21162: out = 67;
			21163: out = 68;
			21164: out = 65;
			21165: out = 77;
			21166: out = 55;
			21167: out = 64;
			21168: out = 66;
			21169: out = 61;
			21170: out = 61;
			21171: out = 63;
			21172: out = 51;
			21173: out = 57;
			21174: out = 61;
			21175: out = 52;
			21176: out = 48;
			21177: out = 60;
			21178: out = 49;
			21179: out = 50;
			21180: out = 49;
			21181: out = 50;
			21182: out = 55;
			21183: out = 50;
			21184: out = 36;
			21185: out = 50;
			21186: out = 48;
			21187: out = 48;
			21188: out = 49;
			21189: out = 38;
			21190: out = 46;
			21191: out = 42;
			21192: out = 37;
			21193: out = 38;
			21194: out = 33;
			21195: out = 42;
			21196: out = 36;
			21197: out = 40;
			21198: out = 27;
			21199: out = 46;
			21200: out = 28;
			21201: out = 31;
			21202: out = 38;
			21203: out = 21;
			21204: out = 15;
			21205: out = 37;
			21206: out = 22;
			21207: out = 24;
			21208: out = 20;
			21209: out = 27;
			21210: out = 26;
			21211: out = 9;
			21212: out = 24;
			21213: out = 17;
			21214: out = 22;
			21215: out = 13;
			21216: out = 15;
			21217: out = 24;
			21218: out = 14;
			21219: out = 6;
			21220: out = 19;
			21221: out = 8;
			21222: out = 17;
			21223: out = 12;
			21224: out = 5;
			21225: out = 21;
			21226: out = 2;
			21227: out = 6;
			21228: out = 13;
			21229: out = 9;
			21230: out = -3;
			21231: out = 14;
			21232: out = 4;
			21233: out = 8;
			21234: out = -1;
			21235: out = 3;
			21236: out = 5;
			21237: out = 0;
			21238: out = -3;
			21239: out = 5;
			21240: out = 2;
			21241: out = -6;
			21242: out = -1;
			21243: out = 5;
			21244: out = -12;
			21245: out = 3;
			21246: out = -8;
			21247: out = -4;
			21248: out = 0;
			21249: out = -9;
			21250: out = -4;
			21251: out = -8;
			21252: out = -6;
			21253: out = -1;
			21254: out = -13;
			21255: out = -3;
			21256: out = -10;
			21257: out = -9;
			21258: out = -4;
			21259: out = -9;
			21260: out = -19;
			21261: out = -7;
			21262: out = -9;
			21263: out = -14;
			21264: out = -12;
			21265: out = -16;
			21266: out = -10;
			21267: out = -20;
			21268: out = -14;
			21269: out = -12;
			21270: out = -16;
			21271: out = -22;
			21272: out = -21;
			21273: out = -18;
			21274: out = -16;
			21275: out = -36;
			21276: out = -24;
			21277: out = -22;
			21278: out = -34;
			21279: out = -27;
			21280: out = -24;
			21281: out = -32;
			21282: out = -36;
			21283: out = -33;
			21284: out = -27;
			21285: out = -36;
			21286: out = -33;
			21287: out = -38;
			21288: out = -37;
			21289: out = -34;
			21290: out = -33;
			21291: out = -39;
			21292: out = -38;
			21293: out = -33;
			21294: out = -46;
			21295: out = -31;
			21296: out = -40;
			21297: out = -57;
			21298: out = -33;
			21299: out = -48;
			21300: out = -44;
			21301: out = -46;
			21302: out = -48;
			21303: out = -41;
			21304: out = -58;
			21305: out = -44;
			21306: out = -50;
			21307: out = -49;
			21308: out = -58;
			21309: out = -43;
			21310: out = -56;
			21311: out = -50;
			21312: out = -56;
			21313: out = -53;
			21314: out = -57;
			21315: out = -61;
			21316: out = -54;
			21317: out = -62;
			21318: out = -64;
			21319: out = -67;
			21320: out = -58;
			21321: out = -65;
			21322: out = -67;
			21323: out = -63;
			21324: out = -66;
			21325: out = -63;
			21326: out = -73;
			21327: out = -49;
			21328: out = -79;
			21329: out = -73;
			21330: out = -64;
			21331: out = -73;
			21332: out = -72;
			21333: out = -70;
			21334: out = -65;
			21335: out = -67;
			21336: out = -75;
			21337: out = -72;
			21338: out = -64;
			21339: out = -85;
			21340: out = -67;
			21341: out = -75;
			21342: out = -77;
			21343: out = -73;
			21344: out = -76;
			21345: out = -80;
			21346: out = -73;
			21347: out = -80;
			21348: out = -77;
			21349: out = -83;
			21350: out = -76;
			21351: out = -84;
			21352: out = -83;
			21353: out = -78;
			21354: out = -83;
			21355: out = -89;
			21356: out = -79;
			21357: out = -88;
			21358: out = -98;
			21359: out = -93;
			21360: out = -86;
			21361: out = -90;
			21362: out = -90;
			21363: out = -98;
			21364: out = -91;
			21365: out = -97;
			21366: out = -91;
			21367: out = -87;
			21368: out = -95;
			21369: out = -105;
			21370: out = -89;
			21371: out = -95;
			21372: out = -100;
			21373: out = -100;
			21374: out = -96;
			21375: out = -105;
			21376: out = -99;
			21377: out = -107;
			21378: out = -105;
			21379: out = -107;
			21380: out = -107;
			21381: out = -102;
			21382: out = -114;
			21383: out = -105;
			21384: out = -110;
			21385: out = -111;
			21386: out = -114;
			21387: out = -116;
			21388: out = -115;
			21389: out = -119;
			21390: out = -113;
			21391: out = -117;
			21392: out = -119;
			21393: out = -124;
			21394: out = -120;
			21395: out = -123;
			21396: out = -128;
			21397: out = -133;
			21398: out = -120;
			21399: out = -135;
			21400: out = -128;
			21401: out = -131;
			21402: out = -134;
			21403: out = -127;
			21404: out = -140;
			21405: out = -139;
			21406: out = -138;
			21407: out = -137;
			21408: out = -139;
			21409: out = -152;
			21410: out = -145;
			21411: out = -138;
			21412: out = -148;
			21413: out = -146;
			21414: out = -149;
			21415: out = -144;
			21416: out = -149;
			21417: out = -157;
			21418: out = -145;
			21419: out = -148;
			21420: out = -164;
			21421: out = -152;
			21422: out = -158;
			21423: out = -158;
			21424: out = -160;
			21425: out = -163;
			21426: out = -152;
			21427: out = -164;
			21428: out = -167;
			21429: out = -156;
			21430: out = -166;
			21431: out = -169;
			21432: out = -166;
			21433: out = -168;
			21434: out = -174;
			21435: out = -162;
			21436: out = -174;
			21437: out = -170;
			21438: out = -174;
			21439: out = -176;
			21440: out = -166;
			21441: out = -172;
			21442: out = -186;
			21443: out = -172;
			21444: out = -172;
			21445: out = -171;
			21446: out = -179;
			21447: out = -170;
			21448: out = -184;
			21449: out = -174;
			21450: out = -172;
			21451: out = -191;
			21452: out = -163;
			21453: out = -185;
			21454: out = -184;
			21455: out = -172;
			21456: out = -181;
			21457: out = -185;
			21458: out = -176;
			21459: out = -179;
			21460: out = -181;
			21461: out = -192;
			21462: out = -178;
			21463: out = -186;
			21464: out = -181;
			21465: out = -191;
			21466: out = -182;
			21467: out = -180;
			21468: out = -191;
			21469: out = -183;
			21470: out = -186;
			21471: out = -184;
			21472: out = -190;
			21473: out = -190;
			21474: out = -183;
			21475: out = -184;
			21476: out = -192;
			21477: out = -183;
			21478: out = -185;
			21479: out = -190;
			21480: out = -190;
			21481: out = -193;
			21482: out = -185;
			21483: out = -196;
			21484: out = -191;
			21485: out = -183;
			21486: out = -198;
			21487: out = -185;
			21488: out = -187;
			21489: out = -193;
			21490: out = -185;
			21491: out = -199;
			21492: out = -186;
			21493: out = -184;
			21494: out = -202;
			21495: out = -185;
			21496: out = -184;
			21497: out = -193;
			21498: out = -188;
			21499: out = -188;
			21500: out = -182;
			21501: out = -184;
			21502: out = -199;
			21503: out = -187;
			21504: out = -190;
			21505: out = -191;
			21506: out = -188;
			21507: out = -194;
			21508: out = -185;
			21509: out = -186;
			21510: out = -180;
			21511: out = -198;
			21512: out = -180;
			21513: out = -191;
			21514: out = -196;
			21515: out = -192;
			21516: out = -179;
			21517: out = -188;
			21518: out = -192;
			21519: out = -186;
			21520: out = -182;
			21521: out = -187;
			21522: out = -184;
			21523: out = -188;
			21524: out = -191;
			21525: out = -179;
			21526: out = -191;
			21527: out = -186;
			21528: out = -191;
			21529: out = -190;
			21530: out = -196;
			21531: out = -176;
			21532: out = -194;
			21533: out = -188;
			21534: out = -178;
			21535: out = -192;
			21536: out = -182;
			21537: out = -185;
			21538: out = -187;
			21539: out = -179;
			21540: out = -187;
			21541: out = -182;
			21542: out = -176;
			21543: out = -186;
			21544: out = -181;
			21545: out = -180;
			21546: out = -181;
			21547: out = -181;
			21548: out = -184;
			21549: out = -179;
			21550: out = -182;
			21551: out = -167;
			21552: out = -194;
			21553: out = -178;
			21554: out = -179;
			21555: out = -178;
			21556: out = -178;
			21557: out = -181;
			21558: out = -176;
			21559: out = -174;
			21560: out = -184;
			21561: out = -170;
			21562: out = -181;
			21563: out = -176;
			21564: out = -178;
			21565: out = -173;
			21566: out = -179;
			21567: out = -181;
			21568: out = -163;
			21569: out = -184;
			21570: out = -170;
			21571: out = -175;
			21572: out = -179;
			21573: out = -163;
			21574: out = -181;
			21575: out = -159;
			21576: out = -175;
			21577: out = -171;
			21578: out = -169;
			21579: out = -160;
			21580: out = -164;
			21581: out = -159;
			21582: out = -174;
			21583: out = -159;
			21584: out = -159;
			21585: out = -167;
			21586: out = -161;
			21587: out = -161;
			21588: out = -167;
			21589: out = -152;
			21590: out = -160;
			21591: out = -158;
			21592: out = -161;
			21593: out = -152;
			21594: out = -156;
			21595: out = -158;
			21596: out = -155;
			21597: out = -151;
			21598: out = -154;
			21599: out = -144;
			21600: out = -158;
			21601: out = -148;
			21602: out = -146;
			21603: out = -141;
			21604: out = -150;
			21605: out = -146;
			21606: out = -136;
			21607: out = -135;
			21608: out = -143;
			21609: out = -139;
			21610: out = -133;
			21611: out = -137;
			21612: out = -137;
			21613: out = -131;
			21614: out = -138;
			21615: out = -123;
			21616: out = -132;
			21617: out = -135;
			21618: out = -124;
			21619: out = -138;
			21620: out = -124;
			21621: out = -119;
			21622: out = -133;
			21623: out = -122;
			21624: out = -127;
			21625: out = -111;
			21626: out = -133;
			21627: out = -117;
			21628: out = -116;
			21629: out = -116;
			21630: out = -113;
			21631: out = -123;
			21632: out = -105;
			21633: out = -111;
			21634: out = -112;
			21635: out = -112;
			21636: out = -101;
			21637: out = -107;
			21638: out = -110;
			21639: out = -103;
			21640: out = -108;
			21641: out = -107;
			21642: out = -101;
			21643: out = -111;
			21644: out = -100;
			21645: out = -102;
			21646: out = -103;
			21647: out = -104;
			21648: out = -95;
			21649: out = -109;
			21650: out = -100;
			21651: out = -95;
			21652: out = -98;
			21653: out = -92;
			21654: out = -86;
			21655: out = -102;
			21656: out = -85;
			21657: out = -97;
			21658: out = -84;
			21659: out = -89;
			21660: out = -96;
			21661: out = -93;
			21662: out = -81;
			21663: out = -85;
			21664: out = -86;
			21665: out = -88;
			21666: out = -77;
			21667: out = -79;
			21668: out = -87;
			21669: out = -78;
			21670: out = -83;
			21671: out = -81;
			21672: out = -76;
			21673: out = -79;
			21674: out = -85;
			21675: out = -64;
			21676: out = -81;
			21677: out = -83;
			21678: out = -70;
			21679: out = -73;
			21680: out = -77;
			21681: out = -77;
			21682: out = -77;
			21683: out = -69;
			21684: out = -79;
			21685: out = -70;
			21686: out = -79;
			21687: out = -68;
			21688: out = -68;
			21689: out = -75;
			21690: out = -61;
			21691: out = -67;
			21692: out = -77;
			21693: out = -61;
			21694: out = -64;
			21695: out = -69;
			21696: out = -66;
			21697: out = -65;
			21698: out = -61;
			21699: out = -61;
			21700: out = -63;
			21701: out = -61;
			21702: out = -57;
			21703: out = -60;
			21704: out = -60;
			21705: out = -56;
			21706: out = -60;
			21707: out = -53;
			21708: out = -46;
			21709: out = -56;
			21710: out = -58;
			21711: out = -45;
			21712: out = -49;
			21713: out = -49;
			21714: out = -51;
			21715: out = -48;
			21716: out = -42;
			21717: out = -45;
			21718: out = -52;
			21719: out = -41;
			21720: out = -43;
			21721: out = -54;
			21722: out = -40;
			21723: out = -37;
			21724: out = -54;
			21725: out = -40;
			21726: out = -38;
			21727: out = -43;
			21728: out = -37;
			21729: out = -42;
			21730: out = -30;
			21731: out = -46;
			21732: out = -33;
			21733: out = -40;
			21734: out = -33;
			21735: out = -32;
			21736: out = -37;
			21737: out = -28;
			21738: out = -45;
			21739: out = -25;
			21740: out = -38;
			21741: out = -32;
			21742: out = -30;
			21743: out = -27;
			21744: out = -28;
			21745: out = -28;
			21746: out = -24;
			21747: out = -27;
			21748: out = -27;
			21749: out = -24;
			21750: out = -26;
			21751: out = -24;
			21752: out = -24;
			21753: out = -25;
			21754: out = -27;
			21755: out = -20;
			21756: out = -20;
			21757: out = -32;
			21758: out = -26;
			21759: out = -18;
			21760: out = -22;
			21761: out = -28;
			21762: out = -9;
			21763: out = -26;
			21764: out = -24;
			21765: out = -14;
			21766: out = -19;
			21767: out = -14;
			21768: out = -17;
			21769: out = -22;
			21770: out = -9;
			21771: out = -13;
			21772: out = -14;
			21773: out = -15;
			21774: out = -13;
			21775: out = -7;
			21776: out = -2;
			21777: out = -21;
			21778: out = -9;
			21779: out = -2;
			21780: out = -6;
			21781: out = -9;
			21782: out = -4;
			21783: out = -5;
			21784: out = -12;
			21785: out = 0;
			default: out = 0;
		endcase
	end
endmodule
