module ride_lookup(index, out);
	input logic unsigned [15:0] index;
	output logic signed [15:0] out;
	always_comb begin
		case(index)
			0: out = 16'(0);
			1: out = 16'(0);
			2: out = 16'(18);
			3: out = 16'(-93);
			4: out = 16'(16);
			5: out = 16'(-97);
			6: out = 16'(38);
			7: out = 16'(-126);
			8: out = 16'(71);
			9: out = 16'(-169);
			10: out = 16'(69);
			11: out = 16'(-585);
			12: out = 16'(21);
			13: out = 16'(-2506);
			14: out = 16'(-3841);
			15: out = 16'(-8349);
			16: out = 16'(8299);
			17: out = 16'(9420);
			18: out = 16'(-22012);
			19: out = 16'(-26602);
			20: out = 16'(-26790);
			21: out = 16'(23837);
			22: out = 16'(620);
			23: out = 16'(-27834);
			24: out = 16'(-624);
			25: out = 16'(-2956);
			26: out = 16'(-3601);
			27: out = 16'(38);
			28: out = 16'(3163);
			29: out = 16'(764);
			30: out = 16'(6420);
			31: out = 16'(1912);
			32: out = 16'(-5883);
			33: out = 16'(1596);
			34: out = 16'(1327);
			35: out = 16'(-32767);
			36: out = 16'(5972);
			37: out = 16'(27312);
			38: out = 16'(20281);
			39: out = 16'(-7778);
			40: out = 16'(-31196);
			41: out = 16'(-22403);
			42: out = 16'(-351);
			43: out = 16'(26805);
			44: out = 16'(21790);
			45: out = 16'(24563);
			46: out = 16'(22227);
			47: out = 16'(-13671);
			48: out = 16'(-25864);
			49: out = 16'(-8746);
			50: out = 16'(-6210);
			51: out = 16'(3771);
			52: out = 16'(2007);
			53: out = 16'(13635);
			54: out = 16'(11822);
			55: out = 16'(3428);
			56: out = 16'(-13956);
			57: out = 16'(-24412);
			58: out = 16'(-705);
			59: out = 16'(2608);
			60: out = 16'(4175);
			61: out = 16'(21207);
			62: out = 16'(9747);
			63: out = 16'(-15861);
			64: out = 16'(9642);
			65: out = 16'(13815);
			66: out = 16'(19235);
			67: out = 16'(-13223);
			68: out = 16'(-26317);
			69: out = 16'(-19990);
			70: out = 16'(-8521);
			71: out = 16'(6276);
			72: out = 16'(19007);
			73: out = 16'(18222);
			74: out = 16'(6635);
			75: out = 16'(-26092);
			76: out = 16'(-29177);
			77: out = 16'(-27222);
			78: out = 16'(8717);
			79: out = 16'(21553);
			80: out = 16'(22250);
			81: out = 16'(6043);
			82: out = 16'(-170);
			83: out = 16'(1745);
			84: out = 16'(-2054);
			85: out = 16'(-334);
			86: out = 16'(4263);
			87: out = 16'(-2026);
			88: out = 16'(-4989);
			89: out = 16'(1419);
			90: out = 16'(-411);
			91: out = 16'(-1800);
			92: out = 16'(-15057);
			93: out = 16'(-5068);
			94: out = 16'(4243);
			95: out = 16'(-21759);
			96: out = 16'(-17665);
			97: out = 16'(-5652);
			98: out = 16'(-1118);
			99: out = 16'(-4358);
			100: out = 16'(-20738);
			101: out = 16'(10830);
			102: out = 16'(21237);
			103: out = 16'(27651);
			104: out = 16'(8190);
			105: out = 16'(-8997);
			106: out = 16'(-32767);
			107: out = 16'(-7546);
			108: out = 16'(17093);
			109: out = 16'(24529);
			110: out = 16'(819);
			111: out = 16'(-25338);
			112: out = 16'(-18636);
			113: out = 16'(-10472);
			114: out = 16'(7773);
			115: out = 16'(5367);
			116: out = 16'(13564);
			117: out = 16'(16501);
			118: out = 16'(10631);
			119: out = 16'(4451);
			120: out = 16'(2697);
			121: out = 16'(-4913);
			122: out = 16'(-1127);
			123: out = 16'(17694);
			124: out = 16'(8495);
			125: out = 16'(1810);
			126: out = 16'(-7909);
			127: out = 16'(-8111);
			128: out = 16'(-5795);
			129: out = 16'(19902);
			130: out = 16'(-5662);
			131: out = 16'(-32563);
			132: out = 16'(-2613);
			133: out = 16'(12995);
			134: out = 16'(24813);
			135: out = 16'(-11509);
			136: out = 16'(-23140);
			137: out = 16'(-22691);
			138: out = 16'(-2470);
			139: out = 16'(7998);
			140: out = 16'(-5300);
			141: out = 16'(14954);
			142: out = 16'(17109);
			143: out = 16'(11750);
			144: out = 16'(-680);
			145: out = 16'(-7461);
			146: out = 16'(-25301);
			147: out = 16'(1464);
			148: out = 16'(26018);
			149: out = 16'(20224);
			150: out = 16'(-3547);
			151: out = 16'(-32767);
			152: out = 16'(-23367);
			153: out = 16'(-13458);
			154: out = 16'(8344);
			155: out = 16'(2345);
			156: out = 16'(8175);
			157: out = 16'(11919);
			158: out = 16'(18874);
			159: out = 16'(12375);
			160: out = 16'(-16412);
			161: out = 16'(-7615);
			162: out = 16'(1465);
			163: out = 16'(9474);
			164: out = 16'(6340);
			165: out = 16'(-2568);
			166: out = 16'(-26034);
			167: out = 16'(-23504);
			168: out = 16'(-7810);
			169: out = 16'(-15231);
			170: out = 16'(-1568);
			171: out = 16'(17224);
			172: out = 16'(5297);
			173: out = 16'(1778);
			174: out = 16'(-648);
			175: out = 16'(5986);
			176: out = 16'(7519);
			177: out = 16'(1903);
			178: out = 16'(-3267);
			179: out = 16'(-4557);
			180: out = 16'(20595);
			181: out = 16'(-11448);
			182: out = 16'(-30296);
			183: out = 16'(13958);
			184: out = 16'(16147);
			185: out = 16'(7125);
			186: out = 16'(10447);
			187: out = 16'(-1981);
			188: out = 16'(-14115);
			189: out = 16'(-19825);
			190: out = 16'(-6676);
			191: out = 16'(20965);
			192: out = 16'(22248);
			193: out = 16'(12566);
			194: out = 16'(-31181);
			195: out = 16'(-4231);
			196: out = 16'(6750);
			197: out = 16'(1486);
			198: out = 16'(-5121);
			199: out = 16'(-4549);
			200: out = 16'(25234);
			201: out = 16'(19127);
			202: out = 16'(7952);
			203: out = 16'(2041);
			204: out = 16'(-17694);
			205: out = 16'(-30328);
			206: out = 16'(-20597);
			207: out = 16'(1151);
			208: out = 16'(24999);
			209: out = 16'(13369);
			210: out = 16'(4788);
			211: out = 16'(-11443);
			212: out = 16'(3398);
			213: out = 16'(7365);
			214: out = 16'(-10848);
			215: out = 16'(12002);
			216: out = 16'(22641);
			217: out = 16'(8398);
			218: out = 16'(1450);
			219: out = 16'(-7561);
			220: out = 16'(6667);
			221: out = 16'(-1804);
			222: out = 16'(-11759);
			223: out = 16'(-28149);
			224: out = 16'(-22748);
			225: out = 16'(-2129);
			226: out = 16'(-2554);
			227: out = 16'(4834);
			228: out = 16'(14724);
			229: out = 16'(14333);
			230: out = 16'(9180);
			231: out = 16'(-12049);
			232: out = 16'(10078);
			233: out = 16'(18884);
			234: out = 16'(941);
			235: out = 16'(4290);
			236: out = 16'(2614);
			237: out = 16'(-4493);
			238: out = 16'(-16282);
			239: out = 16'(-26478);
			240: out = 16'(-1320);
			241: out = 16'(12547);
			242: out = 16'(28419);
			243: out = 16'(-7770);
			244: out = 16'(-4799);
			245: out = 16'(13219);
			246: out = 16'(13318);
			247: out = 16'(11835);
			248: out = 16'(13238);
			249: out = 16'(-13888);
			250: out = 16'(-22345);
			251: out = 16'(2674);
			252: out = 16'(16612);
			253: out = 16'(21851);
			254: out = 16'(-12057);
			255: out = 16'(-21987);
			256: out = 16'(-28277);
			257: out = 16'(9003);
			258: out = 16'(13531);
			259: out = 16'(9760);
			260: out = 16'(8771);
			261: out = 16'(401);
			262: out = 16'(-10591);
			263: out = 16'(-8484);
			264: out = 16'(-10863);
			265: out = 16'(-23166);
			266: out = 16'(1612);
			267: out = 16'(10006);
			268: out = 16'(1468);
			269: out = 16'(-1785);
			270: out = 16'(-5614);
			271: out = 16'(-14457);
			272: out = 16'(-1343);
			273: out = 16'(12527);
			274: out = 16'(24050);
			275: out = 16'(14933);
			276: out = 16'(-2697);
			277: out = 16'(-24163);
			278: out = 16'(-28210);
			279: out = 16'(-17560);
			280: out = 16'(-2719);
			281: out = 16'(4941);
			282: out = 16'(1358);
			283: out = 16'(3912);
			284: out = 16'(1543);
			285: out = 16'(-10);
			286: out = 16'(1190);
			287: out = 16'(4327);
			288: out = 16'(7963);
			289: out = 16'(2815);
			290: out = 16'(-2901);
			291: out = 16'(6199);
			292: out = 16'(408);
			293: out = 16'(-6091);
			294: out = 16'(-28146);
			295: out = 16'(-18216);
			296: out = 16'(8816);
			297: out = 16'(-4682);
			298: out = 16'(1678);
			299: out = 16'(12830);
			300: out = 16'(10841);
			301: out = 16'(6644);
			302: out = 16'(-2121);
			303: out = 16'(1785);
			304: out = 16'(7575);
			305: out = 16'(16988);
			306: out = 16'(19500);
			307: out = 16'(12267);
			308: out = 16'(-27354);
			309: out = 16'(-23791);
			310: out = 16'(-9872);
			311: out = 16'(15107);
			312: out = 16'(20557);
			313: out = 16'(18242);
			314: out = 16'(734);
			315: out = 16'(-13817);
			316: out = 16'(-29317);
			317: out = 16'(1735);
			318: out = 16'(12870);
			319: out = 16'(4985);
			320: out = 16'(-3562);
			321: out = 16'(-9398);
			322: out = 16'(14072);
			323: out = 16'(-14394);
			324: out = 16'(-26384);
			325: out = 16'(-13485);
			326: out = 16'(119);
			327: out = 16'(10241);
			328: out = 16'(17278);
			329: out = 16'(5597);
			330: out = 16'(-10305);
			331: out = 16'(-10627);
			332: out = 16'(-11522);
			333: out = 16'(-10749);
			334: out = 16'(17492);
			335: out = 16'(14271);
			336: out = 16'(-15799);
			337: out = 16'(-23882);
			338: out = 16'(-25840);
			339: out = 16'(6372);
			340: out = 16'(-7166);
			341: out = 16'(-5773);
			342: out = 16'(10625);
			343: out = 16'(18911);
			344: out = 16'(20210);
			345: out = 16'(17154);
			346: out = 16'(-5720);
			347: out = 16'(-30190);
			348: out = 16'(38);
			349: out = 16'(7554);
			350: out = 16'(14591);
			351: out = 16'(-14823);
			352: out = 16'(-14457);
			353: out = 16'(3902);
			354: out = 16'(1288);
			355: out = 16'(5050);
			356: out = 16'(11991);
			357: out = 16'(3819);
			358: out = 16'(368);
			359: out = 16'(6395);
			360: out = 16'(10189);
			361: out = 16'(13236);
			362: out = 16'(4070);
			363: out = 16'(282);
			364: out = 16'(-5812);
			365: out = 16'(14899);
			366: out = 16'(521);
			367: out = 16'(-18293);
			368: out = 16'(-6526);
			369: out = 16'(5544);
			370: out = 16'(21714);
			371: out = 16'(6149);
			372: out = 16'(379);
			373: out = 16'(-2404);
			374: out = 16'(601);
			375: out = 16'(2042);
			376: out = 16'(-5247);
			377: out = 16'(7972);
			378: out = 16'(14002);
			379: out = 16'(10421);
			380: out = 16'(3098);
			381: out = 16'(-5042);
			382: out = 16'(-11707);
			383: out = 16'(-8887);
			384: out = 16'(-1144);
			385: out = 16'(1982);
			386: out = 16'(7603);
			387: out = 16'(12458);
			388: out = 16'(-6261);
			389: out = 16'(-10063);
			390: out = 16'(-3560);
			391: out = 16'(1500);
			392: out = 16'(-2194);
			393: out = 16'(-30850);
			394: out = 16'(-2568);
			395: out = 16'(10125);
			396: out = 16'(-11106);
			397: out = 16'(-6452);
			398: out = 16'(-1522);
			399: out = 16'(29322);
			400: out = 16'(10982);
			401: out = 16'(-9851);
			402: out = 16'(-5866);
			403: out = 16'(-11577);
			404: out = 16'(-16645);
			405: out = 16'(5100);
			406: out = 16'(16224);
			407: out = 16'(26747);
			408: out = 16'(-16832);
			409: out = 16'(-29416);
			410: out = 16'(-21099);
			411: out = 16'(1146);
			412: out = 16'(13351);
			413: out = 16'(7819);
			414: out = 16'(7613);
			415: out = 16'(5133);
			416: out = 16'(2838);
			417: out = 16'(5341);
			418: out = 16'(8018);
			419: out = 16'(25071);
			420: out = 16'(4317);
			421: out = 16'(-23907);
			422: out = 16'(-4490);
			423: out = 16'(-912);
			424: out = 16'(1395);
			425: out = 16'(11037);
			426: out = 16'(8389);
			427: out = 16'(-5029);
			428: out = 16'(-1717);
			429: out = 16'(-2709);
			430: out = 16'(-13644);
			431: out = 16'(11964);
			432: out = 16'(21583);
			433: out = 16'(2250);
			434: out = 16'(-9199);
			435: out = 16'(-19526);
			436: out = 16'(3234);
			437: out = 16'(6895);
			438: out = 16'(11913);
			439: out = 16'(-5050);
			440: out = 16'(-425);
			441: out = 16'(8218);
			442: out = 16'(-5572);
			443: out = 16'(-338);
			444: out = 16'(19207);
			445: out = 16'(713);
			446: out = 16'(-4504);
			447: out = 16'(-10504);
			448: out = 16'(5406);
			449: out = 16'(9913);
			450: out = 16'(2095);
			451: out = 16'(-13619);
			452: out = 16'(-22000);
			453: out = 16'(15985);
			454: out = 16'(13860);
			455: out = 16'(11811);
			456: out = 16'(-24067);
			457: out = 16'(-11813);
			458: out = 16'(13177);
			459: out = 16'(4072);
			460: out = 16'(6810);
			461: out = 16'(6434);
			462: out = 16'(1952);
			463: out = 16'(-8750);
			464: out = 16'(-24610);
			465: out = 16'(-19798);
			466: out = 16'(-7878);
			467: out = 16'(15450);
			468: out = 16'(13427);
			469: out = 16'(8305);
			470: out = 16'(-9725);
			471: out = 16'(-7255);
			472: out = 16'(-1911);
			473: out = 16'(12334);
			474: out = 16'(309);
			475: out = 16'(-18925);
			476: out = 16'(9847);
			477: out = 16'(9562);
			478: out = 16'(8041);
			479: out = 16'(-14229);
			480: out = 16'(-18364);
			481: out = 16'(-13374);
			482: out = 16'(5910);
			483: out = 16'(16695);
			484: out = 16'(23047);
			485: out = 16'(-6092);
			486: out = 16'(-22347);
			487: out = 16'(10225);
			488: out = 16'(2101);
			489: out = 16'(645);
			490: out = 16'(-22172);
			491: out = 16'(2002);
			492: out = 16'(26178);
			493: out = 16'(4966);
			494: out = 16'(-422);
			495: out = 16'(-10362);
			496: out = 16'(3243);
			497: out = 16'(-1051);
			498: out = 16'(-10150);
			499: out = 16'(-2859);
			500: out = 16'(3066);
			501: out = 16'(1084);
			502: out = 16'(15320);
			503: out = 16'(14111);
			504: out = 16'(-1511);
			505: out = 16'(-12139);
			506: out = 16'(-16637);
			507: out = 16'(-10392);
			508: out = 16'(5066);
			509: out = 16'(17651);
			510: out = 16'(11698);
			511: out = 16'(11073);
			512: out = 16'(10461);
			513: out = 16'(-16858);
			514: out = 16'(-18635);
			515: out = 16'(-9505);
			516: out = 16'(14004);
			517: out = 16'(17370);
			518: out = 16'(5598);
			519: out = 16'(-11303);
			520: out = 16'(-15568);
			521: out = 16'(13401);
			522: out = 16'(-154);
			523: out = 16'(-4761);
			524: out = 16'(8341);
			525: out = 16'(3828);
			526: out = 16'(952);
			527: out = 16'(-23279);
			528: out = 16'(-5789);
			529: out = 16'(16394);
			530: out = 16'(21962);
			531: out = 16'(5783);
			532: out = 16'(-26587);
			533: out = 16'(-23658);
			534: out = 16'(-18069);
			535: out = 16'(2964);
			536: out = 16'(8926);
			537: out = 16'(12727);
			538: out = 16'(975);
			539: out = 16'(1996);
			540: out = 16'(-2664);
			541: out = 16'(1004);
			542: out = 16'(-10221);
			543: out = 16'(-12946);
			544: out = 16'(5126);
			545: out = 16'(13542);
			546: out = 16'(17122);
			547: out = 16'(-13316);
			548: out = 16'(-15759);
			549: out = 16'(-8437);
			550: out = 16'(-241);
			551: out = 16'(4874);
			552: out = 16'(3539);
			553: out = 16'(10361);
			554: out = 16'(7873);
			555: out = 16'(848);
			556: out = 16'(-5895);
			557: out = 16'(-6873);
			558: out = 16'(4511);
			559: out = 16'(4537);
			560: out = 16'(5436);
			561: out = 16'(659);
			562: out = 16'(2349);
			563: out = 16'(2801);
			564: out = 16'(15857);
			565: out = 16'(-3902);
			566: out = 16'(-31062);
			567: out = 16'(-759);
			568: out = 16'(10115);
			569: out = 16'(21601);
			570: out = 16'(-6115);
			571: out = 16'(-13456);
			572: out = 16'(-16394);
			573: out = 16'(4856);
			574: out = 16'(10495);
			575: out = 16'(766);
			576: out = 16'(-4470);
			577: out = 16'(-5488);
			578: out = 16'(1148);
			579: out = 16'(10464);
			580: out = 16'(15123);
			581: out = 16'(16550);
			582: out = 16'(794);
			583: out = 16'(-15509);
			584: out = 16'(-16935);
			585: out = 16'(456);
			586: out = 16'(27296);
			587: out = 16'(9978);
			588: out = 16'(1738);
			589: out = 16'(-11799);
			590: out = 16'(-8576);
			591: out = 16'(-5266);
			592: out = 16'(592);
			593: out = 16'(9541);
			594: out = 16'(14833);
			595: out = 16'(17012);
			596: out = 16'(8633);
			597: out = 16'(-812);
			598: out = 16'(-22930);
			599: out = 16'(-15244);
			600: out = 16'(-934);
			601: out = 16'(21520);
			602: out = 16'(12527);
			603: out = 16'(-7449);
			604: out = 16'(-6663);
			605: out = 16'(-5047);
			606: out = 16'(4299);
			607: out = 16'(7142);
			608: out = 16'(2574);
			609: out = 16'(-19820);
			610: out = 16'(-11725);
			611: out = 16'(-5758);
			612: out = 16'(11477);
			613: out = 16'(-5957);
			614: out = 16'(-13518);
			615: out = 16'(16912);
			616: out = 16'(6832);
			617: out = 16'(-2035);
			618: out = 16'(-23155);
			619: out = 16'(-14093);
			620: out = 16'(3368);
			621: out = 16'(1105);
			622: out = 16'(9119);
			623: out = 16'(20397);
			624: out = 16'(-17527);
			625: out = 16'(-17389);
			626: out = 16'(16012);
			627: out = 16'(3330);
			628: out = 16'(1880);
			629: out = 16'(-1788);
			630: out = 16'(380);
			631: out = 16'(1269);
			632: out = 16'(8037);
			633: out = 16'(8836);
			634: out = 16'(6835);
			635: out = 16'(-27146);
			636: out = 16'(-16673);
			637: out = 16'(1868);
			638: out = 16'(4867);
			639: out = 16'(6254);
			640: out = 16'(1525);
			641: out = 16'(12638);
			642: out = 16'(3310);
			643: out = 16'(-19227);
			644: out = 16'(-9438);
			645: out = 16'(-3607);
			646: out = 16'(9663);
			647: out = 16'(-6311);
			648: out = 16'(-8661);
			649: out = 16'(7962);
			650: out = 16'(15800);
			651: out = 16'(17348);
			652: out = 16'(-9745);
			653: out = 16'(-9746);
			654: out = 16'(-7357);
			655: out = 16'(12921);
			656: out = 16'(3644);
			657: out = 16'(-13566);
			658: out = 16'(10478);
			659: out = 16'(12964);
			660: out = 16'(15444);
			661: out = 16'(-14257);
			662: out = 16'(-15969);
			663: out = 16'(6733);
			664: out = 16'(15004);
			665: out = 16'(14268);
			666: out = 16'(-22628);
			667: out = 16'(3478);
			668: out = 16'(15153);
			669: out = 16'(9979);
			670: out = 16'(4393);
			671: out = 16'(-678);
			672: out = 16'(-1898);
			673: out = 16'(2181);
			674: out = 16'(7001);
			675: out = 16'(-2390);
			676: out = 16'(-3315);
			677: out = 16'(-1493);
			678: out = 16'(-701);
			679: out = 16'(-319);
			680: out = 16'(-4293);
			681: out = 16'(-277);
			682: out = 16'(282);
			683: out = 16'(9035);
			684: out = 16'(-14807);
			685: out = 16'(-23661);
			686: out = 16'(-8154);
			687: out = 16'(-879);
			688: out = 16'(5719);
			689: out = 16'(17627);
			690: out = 16'(3903);
			691: out = 16'(-11216);
			692: out = 16'(-12136);
			693: out = 16'(-6560);
			694: out = 16'(3689);
			695: out = 16'(12403);
			696: out = 16'(6608);
			697: out = 16'(-10808);
			698: out = 16'(-13911);
			699: out = 16'(-11606);
			700: out = 16'(5395);
			701: out = 16'(-69);
			702: out = 16'(499);
			703: out = 16'(7537);
			704: out = 16'(-10127);
			705: out = 16'(-18434);
			706: out = 16'(14538);
			707: out = 16'(14589);
			708: out = 16'(13928);
			709: out = 16'(-25131);
			710: out = 16'(-15820);
			711: out = 16'(2772);
			712: out = 16'(2518);
			713: out = 16'(-7094);
			714: out = 16'(-30415);
			715: out = 16'(10219);
			716: out = 16'(15536);
			717: out = 16'(3469);
			718: out = 16'(-3684);
			719: out = 16'(-8955);
			720: out = 16'(-3612);
			721: out = 16'(-8711);
			722: out = 16'(-5574);
			723: out = 16'(11108);
			724: out = 16'(9514);
			725: out = 16'(6362);
			726: out = 16'(4036);
			727: out = 16'(-1581);
			728: out = 16'(-6249);
			729: out = 16'(7250);
			730: out = 16'(8896);
			731: out = 16'(9717);
			732: out = 16'(-4763);
			733: out = 16'(2335);
			734: out = 16'(25563);
			735: out = 16'(5234);
			736: out = 16'(-1265);
			737: out = 16'(-8175);
			738: out = 16'(11418);
			739: out = 16'(19916);
			740: out = 16'(9949);
			741: out = 16'(6100);
			742: out = 16'(836);
			743: out = 16'(16534);
			744: out = 16'(7851);
			745: out = 16'(2777);
			746: out = 16'(-21733);
			747: out = 16'(-6055);
			748: out = 16'(18575);
			749: out = 16'(14775);
			750: out = 16'(4887);
			751: out = 16'(-19662);
			752: out = 16'(-7106);
			753: out = 16'(-3639);
			754: out = 16'(3570);
			755: out = 16'(861);
			756: out = 16'(-2613);
			757: out = 16'(-23647);
			758: out = 16'(-7386);
			759: out = 16'(3845);
			760: out = 16'(13732);
			761: out = 16'(-2146);
			762: out = 16'(-16283);
			763: out = 16'(11177);
			764: out = 16'(9462);
			765: out = 16'(6552);
			766: out = 16'(1955);
			767: out = 16'(-3300);
			768: out = 16'(-12435);
			769: out = 16'(3557);
			770: out = 16'(-2245);
			771: out = 16'(-26542);
			772: out = 16'(-10320);
			773: out = 16'(-802);
			774: out = 16'(6224);
			775: out = 16'(3929);
			776: out = 16'(942);
			777: out = 16'(-2370);
			778: out = 16'(-3080);
			779: out = 16'(-2467);
			780: out = 16'(-4916);
			781: out = 16'(6145);
			782: out = 16'(17463);
			783: out = 16'(-5354);
			784: out = 16'(-11603);
			785: out = 16'(-20572);
			786: out = 16'(4483);
			787: out = 16'(3624);
			788: out = 16'(-5399);
			789: out = 16'(-21117);
			790: out = 16'(-19724);
			791: out = 16'(5600);
			792: out = 16'(7638);
			793: out = 16'(9576);
			794: out = 16'(4213);
			795: out = 16'(-635);
			796: out = 16'(-7220);
			797: out = 16'(-14467);
			798: out = 16'(-7931);
			799: out = 16'(4494);
			800: out = 16'(13479);
			801: out = 16'(11262);
			802: out = 16'(-604);
			803: out = 16'(13097);
			804: out = 16'(10165);
			805: out = 16'(10019);
			806: out = 16'(-1308);
			807: out = 16'(-1782);
			808: out = 16'(-4084);
			809: out = 16'(15923);
			810: out = 16'(21242);
			811: out = 16'(23722);
			812: out = 16'(-9470);
			813: out = 16'(-28702);
			814: out = 16'(-8980);
			815: out = 16'(5368);
			816: out = 16'(17842);
			817: out = 16'(9493);
			818: out = 16'(1448);
			819: out = 16'(-11181);
			820: out = 16'(213);
			821: out = 16'(5539);
			822: out = 16'(15225);
			823: out = 16'(7124);
			824: out = 16'(4766);
			825: out = 16'(-1998);
			826: out = 16'(331);
			827: out = 16'(-1549);
			828: out = 16'(100);
			829: out = 16'(-8593);
			830: out = 16'(-10787);
			831: out = 16'(-7356);
			832: out = 16'(4089);
			833: out = 16'(11133);
			834: out = 16'(-8602);
			835: out = 16'(3090);
			836: out = 16'(14373);
			837: out = 16'(118);
			838: out = 16'(-4563);
			839: out = 16'(-12018);
			840: out = 16'(15055);
			841: out = 16'(10898);
			842: out = 16'(-5163);
			843: out = 16'(-7101);
			844: out = 16'(-8000);
			845: out = 16'(-5085);
			846: out = 16'(5505);
			847: out = 16'(9390);
			848: out = 16'(-1741);
			849: out = 16'(4267);
			850: out = 16'(5248);
			851: out = 16'(-3821);
			852: out = 16'(-2928);
			853: out = 16'(-1787);
			854: out = 16'(9396);
			855: out = 16'(-4503);
			856: out = 16'(-23796);
			857: out = 16'(-4189);
			858: out = 16'(-175);
			859: out = 16'(3361);
			860: out = 16'(-3763);
			861: out = 16'(-1783);
			862: out = 16'(7902);
			863: out = 16'(-10336);
			864: out = 16'(-11123);
			865: out = 16'(16578);
			866: out = 16'(-1439);
			867: out = 16'(-8149);
			868: out = 16'(-8922);
			869: out = 16'(10552);
			870: out = 16'(19840);
			871: out = 16'(-27525);
			872: out = 16'(-17469);
			873: out = 16'(-298);
			874: out = 16'(11610);
			875: out = 16'(7188);
			876: out = 16'(-6098);
			877: out = 16'(6469);
			878: out = 16'(6472);
			879: out = 16'(7632);
			880: out = 16'(-4962);
			881: out = 16'(-5885);
			882: out = 16'(1925);
			883: out = 16'(700);
			884: out = 16'(-438);
			885: out = 16'(-1324);
			886: out = 16'(-2124);
			887: out = 16'(-2276);
			888: out = 16'(-13367);
			889: out = 16'(-1686);
			890: out = 16'(8699);
			891: out = 16'(10730);
			892: out = 16'(6107);
			893: out = 16'(-894);
			894: out = 16'(-9536);
			895: out = 16'(-5440);
			896: out = 16'(7171);
			897: out = 16'(1923);
			898: out = 16'(3400);
			899: out = 16'(9157);
			900: out = 16'(-13454);
			901: out = 16'(-13760);
			902: out = 16'(25891);
			903: out = 16'(7911);
			904: out = 16'(-3973);
			905: out = 16'(-30971);
			906: out = 16'(-10879);
			907: out = 16'(9769);
			908: out = 16'(864);
			909: out = 16'(7641);
			910: out = 16'(11623);
			911: out = 16'(1736);
			912: out = 16'(-7920);
			913: out = 16'(-22308);
			914: out = 16'(11444);
			915: out = 16'(11994);
			916: out = 16'(-862);
			917: out = 16'(-14260);
			918: out = 16'(-14360);
			919: out = 16'(9157);
			920: out = 16'(11608);
			921: out = 16'(8426);
			922: out = 16'(-31483);
			923: out = 16'(-9318);
			924: out = 16'(7396);
			925: out = 16'(11200);
			926: out = 16'(9051);
			927: out = 16'(5818);
			928: out = 16'(-20754);
			929: out = 16'(-14802);
			930: out = 16'(-515);
			931: out = 16'(15181);
			932: out = 16'(1958);
			933: out = 16'(-32767);
			934: out = 16'(1867);
			935: out = 16'(14035);
			936: out = 16'(11791);
			937: out = 16'(11217);
			938: out = 16'(6325);
			939: out = 16'(5055);
			940: out = 16'(-10101);
			941: out = 16'(-16552);
			942: out = 16'(-8372);
			943: out = 16'(6552);
			944: out = 16'(17616);
			945: out = 16'(6965);
			946: out = 16'(-1015);
			947: out = 16'(-11513);
			948: out = 16'(-6445);
			949: out = 16'(4640);
			950: out = 16'(24650);
			951: out = 16'(-8128);
			952: out = 16'(-10599);
			953: out = 16'(1729);
			954: out = 16'(4889);
			955: out = 16'(8472);
			956: out = 16'(6415);
			957: out = 16'(7947);
			958: out = 16'(6073);
			959: out = 16'(7862);
			960: out = 16'(4301);
			961: out = 16'(2376);
			962: out = 16'(-25187);
			963: out = 16'(-4600);
			964: out = 16'(19293);
			965: out = 16'(17944);
			966: out = 16'(11931);
			967: out = 16'(-1672);
			968: out = 16'(-11795);
			969: out = 16'(-6082);
			970: out = 16'(21353);
			971: out = 16'(311);
			972: out = 16'(-5051);
			973: out = 16'(-20990);
			974: out = 16'(5043);
			975: out = 16'(14800);
			976: out = 16'(19978);
			977: out = 16'(-7180);
			978: out = 16'(-24402);
			979: out = 16'(-1015);
			980: out = 16'(-797);
			981: out = 16'(1239);
			982: out = 16'(16181);
			983: out = 16'(7399);
			984: out = 16'(-7121);
			985: out = 16'(2000);
			986: out = 16'(-1929);
			987: out = 16'(-11386);
			988: out = 16'(5121);
			989: out = 16'(1899);
			990: out = 16'(-13700);
			991: out = 16'(-15057);
			992: out = 16'(-10038);
			993: out = 16'(5222);
			994: out = 16'(7844);
			995: out = 16'(7405);
			996: out = 16'(12218);
			997: out = 16'(-8899);
			998: out = 16'(-25583);
			999: out = 16'(-25912);
			1000: out = 16'(-4155);
			1001: out = 16'(22429);
			1002: out = 16'(4552);
			1003: out = 16'(5678);
			1004: out = 16'(4287);
			1005: out = 16'(-21362);
			1006: out = 16'(-25570);
			1007: out = 16'(-6529);
			1008: out = 16'(-3429);
			1009: out = 16'(3894);
			1010: out = 16'(56);
			1011: out = 16'(16068);
			1012: out = 16'(14223);
			1013: out = 16'(-11416);
			1014: out = 16'(-14490);
			1015: out = 16'(-13799);
			1016: out = 16'(-1789);
			1017: out = 16'(3820);
			1018: out = 16'(8312);
			1019: out = 16'(-2068);
			1020: out = 16'(1775);
			1021: out = 16'(6628);
			1022: out = 16'(3164);
			1023: out = 16'(-1993);
			1024: out = 16'(-8838);
			1025: out = 16'(-2143);
			1026: out = 16'(5391);
			1027: out = 16'(15048);
			1028: out = 16'(9355);
			1029: out = 16'(1937);
			1030: out = 16'(-9935);
			1031: out = 16'(-11216);
			1032: out = 16'(-7934);
			1033: out = 16'(720);
			1034: out = 16'(7836);
			1035: out = 16'(10512);
			1036: out = 16'(3395);
			1037: out = 16'(-8406);
			1038: out = 16'(-20954);
			1039: out = 16'(5195);
			1040: out = 16'(14954);
			1041: out = 16'(22853);
			1042: out = 16'(-2855);
			1043: out = 16'(-11374);
			1044: out = 16'(-11827);
			1045: out = 16'(-2095);
			1046: out = 16'(1001);
			1047: out = 16'(-13723);
			1048: out = 16'(7552);
			1049: out = 16'(15406);
			1050: out = 16'(5088);
			1051: out = 16'(-6716);
			1052: out = 16'(-15894);
			1053: out = 16'(23052);
			1054: out = 16'(-299);
			1055: out = 16'(-23575);
			1056: out = 16'(1968);
			1057: out = 16'(14137);
			1058: out = 16'(25723);
			1059: out = 16'(1650);
			1060: out = 16'(-8344);
			1061: out = 16'(-18199);
			1062: out = 16'(-7904);
			1063: out = 16'(1804);
			1064: out = 16'(18115);
			1065: out = 16'(3955);
			1066: out = 16'(-3787);
			1067: out = 16'(-12903);
			1068: out = 16'(1903);
			1069: out = 16'(13392);
			1070: out = 16'(17861);
			1071: out = 16'(-2123);
			1072: out = 16'(-25387);
			1073: out = 16'(9944);
			1074: out = 16'(4452);
			1075: out = 16'(2085);
			1076: out = 16'(-26572);
			1077: out = 16'(-13309);
			1078: out = 16'(16928);
			1079: out = 16'(14574);
			1080: out = 16'(9608);
			1081: out = 16'(-3646);
			1082: out = 16'(-8285);
			1083: out = 16'(-11446);
			1084: out = 16'(-14714);
			1085: out = 16'(11879);
			1086: out = 16'(23998);
			1087: out = 16'(-4052);
			1088: out = 16'(-6426);
			1089: out = 16'(-12365);
			1090: out = 16'(15103);
			1091: out = 16'(-5668);
			1092: out = 16'(-26374);
			1093: out = 16'(1376);
			1094: out = 16'(7723);
			1095: out = 16'(8594);
			1096: out = 16'(3319);
			1097: out = 16'(5477);
			1098: out = 16'(18541);
			1099: out = 16'(-7168);
			1100: out = 16'(-16895);
			1101: out = 16'(-25396);
			1102: out = 16'(2569);
			1103: out = 16'(14667);
			1104: out = 16'(-2066);
			1105: out = 16'(1499);
			1106: out = 16'(-631);
			1107: out = 16'(-20275);
			1108: out = 16'(-9452);
			1109: out = 16'(4897);
			1110: out = 16'(-271);
			1111: out = 16'(8822);
			1112: out = 16'(18652);
			1113: out = 16'(-15746);
			1114: out = 16'(-13130);
			1115: out = 16'(5735);
			1116: out = 16'(10183);
			1117: out = 16'(3518);
			1118: out = 16'(-24239);
			1119: out = 16'(-18278);
			1120: out = 16'(-10286);
			1121: out = 16'(15922);
			1122: out = 16'(8407);
			1123: out = 16'(3963);
			1124: out = 16'(-9852);
			1125: out = 16'(-2408);
			1126: out = 16'(4844);
			1127: out = 16'(15611);
			1128: out = 16'(-483);
			1129: out = 16'(-23988);
			1130: out = 16'(13388);
			1131: out = 16'(10348);
			1132: out = 16'(4106);
			1133: out = 16'(-21638);
			1134: out = 16'(-20322);
			1135: out = 16'(1627);
			1136: out = 16'(9405);
			1137: out = 16'(13936);
			1138: out = 16'(8971);
			1139: out = 16'(3951);
			1140: out = 16'(-2773);
			1141: out = 16'(-3730);
			1142: out = 16'(-13220);
			1143: out = 16'(-14329);
			1144: out = 16'(22000);
			1145: out = 16'(15607);
			1146: out = 16'(6872);
			1147: out = 16'(-23688);
			1148: out = 16'(-15447);
			1149: out = 16'(7386);
			1150: out = 16'(5699);
			1151: out = 16'(6139);
			1152: out = 16'(829);
			1153: out = 16'(-5762);
			1154: out = 16'(-2384);
			1155: out = 16'(18459);
			1156: out = 16'(12452);
			1157: out = 16'(5406);
			1158: out = 16'(-28733);
			1159: out = 16'(-9416);
			1160: out = 16'(3841);
			1161: out = 16'(6677);
			1162: out = 16'(7733);
			1163: out = 16'(7080);
			1164: out = 16'(-12384);
			1165: out = 16'(-2399);
			1166: out = 16'(12826);
			1167: out = 16'(13112);
			1168: out = 16'(9983);
			1169: out = 16'(-458);
			1170: out = 16'(6372);
			1171: out = 16'(4153);
			1172: out = 16'(429);
			1173: out = 16'(2471);
			1174: out = 16'(3027);
			1175: out = 16'(-1886);
			1176: out = 16'(1236);
			1177: out = 16'(59);
			1178: out = 16'(-4998);
			1179: out = 16'(-9801);
			1180: out = 16'(-8672);
			1181: out = 16'(16472);
			1182: out = 16'(17257);
			1183: out = 16'(13630);
			1184: out = 16'(-3202);
			1185: out = 16'(-6544);
			1186: out = 16'(-3470);
			1187: out = 16'(4759);
			1188: out = 16'(3180);
			1189: out = 16'(-12925);
			1190: out = 16'(11055);
			1191: out = 16'(11396);
			1192: out = 16'(487);
			1193: out = 16'(-20657);
			1194: out = 16'(-25260);
			1195: out = 16'(8612);
			1196: out = 16'(13238);
			1197: out = 16'(15881);
			1198: out = 16'(-64);
			1199: out = 16'(3275);
			1200: out = 16'(2931);
			1201: out = 16'(-4025);
			1202: out = 16'(-12556);
			1203: out = 16'(-18716);
			1204: out = 16'(726);
			1205: out = 16'(4607);
			1206: out = 16'(-2686);
			1207: out = 16'(8207);
			1208: out = 16'(7078);
			1209: out = 16'(8964);
			1210: out = 16'(-17172);
			1211: out = 16'(-18670);
			1212: out = 16'(19172);
			1213: out = 16'(13734);
			1214: out = 16'(9009);
			1215: out = 16'(-8805);
			1216: out = 16'(-6171);
			1217: out = 16'(-3854);
			1218: out = 16'(-23335);
			1219: out = 16'(-14796);
			1220: out = 16'(311);
			1221: out = 16'(8133);
			1222: out = 16'(9165);
			1223: out = 16'(2676);
			1224: out = 16'(10211);
			1225: out = 16'(3355);
			1226: out = 16'(-15178);
			1227: out = 16'(3808);
			1228: out = 16'(6824);
			1229: out = 16'(-2458);
			1230: out = 16'(-19154);
			1231: out = 16'(-23146);
			1232: out = 16'(22907);
			1233: out = 16'(3322);
			1234: out = 16'(-10999);
			1235: out = 16'(-22935);
			1236: out = 16'(-8337);
			1237: out = 16'(13058);
			1238: out = 16'(862);
			1239: out = 16'(9661);
			1240: out = 16'(14548);
			1241: out = 16'(13623);
			1242: out = 16'(5139);
			1243: out = 16'(-3698);
			1244: out = 16'(-11988);
			1245: out = 16'(-11813);
			1246: out = 16'(-9473);
			1247: out = 16'(13651);
			1248: out = 16'(19937);
			1249: out = 16'(5230);
			1250: out = 16'(-10767);
			1251: out = 16'(-22338);
			1252: out = 16'(2006);
			1253: out = 16'(11126);
			1254: out = 16'(21601);
			1255: out = 16'(-7184);
			1256: out = 16'(-2294);
			1257: out = 16'(476);
			1258: out = 16'(19542);
			1259: out = 16'(5299);
			1260: out = 16'(-21186);
			1261: out = 16'(-19295);
			1262: out = 16'(-17345);
			1263: out = 16'(-13415);
			1264: out = 16'(8355);
			1265: out = 16'(18360);
			1266: out = 16'(17237);
			1267: out = 16'(-2474);
			1268: out = 16'(-15239);
			1269: out = 16'(9946);
			1270: out = 16'(-1012);
			1271: out = 16'(-5190);
			1272: out = 16'(-7797);
			1273: out = 16'(-1670);
			1274: out = 16'(2774);
			1275: out = 16'(1812);
			1276: out = 16'(71);
			1277: out = 16'(-566);
			1278: out = 16'(-11600);
			1279: out = 16'(-8075);
			1280: out = 16'(5813);
			1281: out = 16'(9022);
			1282: out = 16'(14406);
			1283: out = 16'(16581);
			1284: out = 16'(9924);
			1285: out = 16'(645);
			1286: out = 16'(-7946);
			1287: out = 16'(-4041);
			1288: out = 16'(1432);
			1289: out = 16'(-24636);
			1290: out = 16'(-4405);
			1291: out = 16'(11238);
			1292: out = 16'(7952);
			1293: out = 16'(-4666);
			1294: out = 16'(-19577);
			1295: out = 16'(-13758);
			1296: out = 16'(-1327);
			1297: out = 16'(15498);
			1298: out = 16'(19594);
			1299: out = 16'(12519);
			1300: out = 16'(-8255);
			1301: out = 16'(-22422);
			1302: out = 16'(-25187);
			1303: out = 16'(3880);
			1304: out = 16'(1994);
			1305: out = 16'(2976);
			1306: out = 16'(-7109);
			1307: out = 16'(-2331);
			1308: out = 16'(1910);
			1309: out = 16'(18389);
			1310: out = 16'(15441);
			1311: out = 16'(10457);
			1312: out = 16'(4175);
			1313: out = 16'(-11034);
			1314: out = 16'(-32106);
			1315: out = 16'(10143);
			1316: out = 16'(19753);
			1317: out = 16'(14455);
			1318: out = 16'(-10748);
			1319: out = 16'(-17832);
			1320: out = 16'(6695);
			1321: out = 16'(250);
			1322: out = 16'(2990);
			1323: out = 16'(-1156);
			1324: out = 16'(16644);
			1325: out = 16'(23274);
			1326: out = 16'(9764);
			1327: out = 16'(-4752);
			1328: out = 16'(-20723);
			1329: out = 16'(5899);
			1330: out = 16'(-486);
			1331: out = 16'(-7396);
			1332: out = 16'(-18481);
			1333: out = 16'(-9963);
			1334: out = 16'(7942);
			1335: out = 16'(7786);
			1336: out = 16'(5426);
			1337: out = 16'(-735);
			1338: out = 16'(-11172);
			1339: out = 16'(-11772);
			1340: out = 16'(6100);
			1341: out = 16'(6829);
			1342: out = 16'(7455);
			1343: out = 16'(1096);
			1344: out = 16'(1203);
			1345: out = 16'(-410);
			1346: out = 16'(-15968);
			1347: out = 16'(-9788);
			1348: out = 16'(1599);
			1349: out = 16'(7983);
			1350: out = 16'(6020);
			1351: out = 16'(-3163);
			1352: out = 16'(644);
			1353: out = 16'(6556);
			1354: out = 16'(22827);
			1355: out = 16'(-1698);
			1356: out = 16'(-10383);
			1357: out = 16'(-11981);
			1358: out = 16'(319);
			1359: out = 16'(5186);
			1360: out = 16'(-14369);
			1361: out = 16'(-3665);
			1362: out = 16'(3223);
			1363: out = 16'(4545);
			1364: out = 16'(-2462);
			1365: out = 16'(-9201);
			1366: out = 16'(10204);
			1367: out = 16'(11525);
			1368: out = 16'(10091);
			1369: out = 16'(6385);
			1370: out = 16'(1040);
			1371: out = 16'(-8032);
			1372: out = 16'(-4111);
			1373: out = 16'(-2616);
			1374: out = 16'(5354);
			1375: out = 16'(-14654);
			1376: out = 16'(-20100);
			1377: out = 16'(-3217);
			1378: out = 16'(7173);
			1379: out = 16'(13433);
			1380: out = 16'(-10525);
			1381: out = 16'(580);
			1382: out = 16'(9976);
			1383: out = 16'(19188);
			1384: out = 16'(9599);
			1385: out = 16'(-5807);
			1386: out = 16'(9317);
			1387: out = 16'(-1855);
			1388: out = 16'(-22061);
			1389: out = 16'(-10085);
			1390: out = 16'(-87);
			1391: out = 16'(16583);
			1392: out = 16'(4942);
			1393: out = 16'(1499);
			1394: out = 16'(-1605);
			1395: out = 16'(8182);
			1396: out = 16'(13672);
			1397: out = 16'(19559);
			1398: out = 16'(2338);
			1399: out = 16'(-12830);
			1400: out = 16'(-7404);
			1401: out = 16'(1990);
			1402: out = 16'(15435);
			1403: out = 16'(-10557);
			1404: out = 16'(-15913);
			1405: out = 16'(-24963);
			1406: out = 16'(11996);
			1407: out = 16'(19520);
			1408: out = 16'(23318);
			1409: out = 16'(-12081);
			1410: out = 16'(-22104);
			1411: out = 16'(-10226);
			1412: out = 16'(6640);
			1413: out = 16'(13910);
			1414: out = 16'(2018);
			1415: out = 16'(-8566);
			1416: out = 16'(-18560);
			1417: out = 16'(-13683);
			1418: out = 16'(-1877);
			1419: out = 16'(12523);
			1420: out = 16'(1756);
			1421: out = 16'(-520);
			1422: out = 16'(-7538);
			1423: out = 16'(14142);
			1424: out = 16'(10927);
			1425: out = 16'(0);
			1426: out = 16'(5471);
			1427: out = 16'(6512);
			1428: out = 16'(9011);
			1429: out = 16'(-18285);
			1430: out = 16'(-25238);
			1431: out = 16'(13550);
			1432: out = 16'(-3473);
			1433: out = 16'(-9819);
			1434: out = 16'(-10039);
			1435: out = 16'(7487);
			1436: out = 16'(19700);
			1437: out = 16'(5657);
			1438: out = 16'(1675);
			1439: out = 16'(-3369);
			1440: out = 16'(-3979);
			1441: out = 16'(118);
			1442: out = 16'(8435);
			1443: out = 16'(6595);
			1444: out = 16'(-3137);
			1445: out = 16'(-30989);
			1446: out = 16'(-5141);
			1447: out = 16'(3787);
			1448: out = 16'(6288);
			1449: out = 16'(-13415);
			1450: out = 16'(-21149);
			1451: out = 16'(3463);
			1452: out = 16'(8843);
			1453: out = 16'(13482);
			1454: out = 16'(-13592);
			1455: out = 16'(-1088);
			1456: out = 16'(10369);
			1457: out = 16'(8546);
			1458: out = 16'(4265);
			1459: out = 16'(-1376);
			1460: out = 16'(-9938);
			1461: out = 16'(-8789);
			1462: out = 16'(-1064);
			1463: out = 16'(11364);
			1464: out = 16'(11808);
			1465: out = 16'(-5425);
			1466: out = 16'(1264);
			1467: out = 16'(5085);
			1468: out = 16'(22725);
			1469: out = 16'(1125);
			1470: out = 16'(-12402);
			1471: out = 16'(-11579);
			1472: out = 16'(-8998);
			1473: out = 16'(-3415);
			1474: out = 16'(6971);
			1475: out = 16'(3426);
			1476: out = 16'(-4456);
			1477: out = 16'(4609);
			1478: out = 16'(7285);
			1479: out = 16'(12066);
			1480: out = 16'(4462);
			1481: out = 16'(4155);
			1482: out = 16'(4397);
			1483: out = 16'(10592);
			1484: out = 16'(9595);
			1485: out = 16'(1025);
			1486: out = 16'(-4290);
			1487: out = 16'(-9264);
			1488: out = 16'(-10354);
			1489: out = 16'(-6258);
			1490: out = 16'(-463);
			1491: out = 16'(-10032);
			1492: out = 16'(-816);
			1493: out = 16'(7487);
			1494: out = 16'(13971);
			1495: out = 16'(11559);
			1496: out = 16'(6469);
			1497: out = 16'(2349);
			1498: out = 16'(99);
			1499: out = 16'(-2195);
			1500: out = 16'(5488);
			1501: out = 16'(3772);
			1502: out = 16'(-4727);
			1503: out = 16'(-15132);
			1504: out = 16'(-15375);
			1505: out = 16'(10513);
			1506: out = 16'(7581);
			1507: out = 16'(6495);
			1508: out = 16'(356);
			1509: out = 16'(-4851);
			1510: out = 16'(-10984);
			1511: out = 16'(8171);
			1512: out = 16'(4082);
			1513: out = 16'(-110);
			1514: out = 16'(-17465);
			1515: out = 16'(-10597);
			1516: out = 16'(9221);
			1517: out = 16'(-321);
			1518: out = 16'(-501);
			1519: out = 16'(1684);
			1520: out = 16'(2850);
			1521: out = 16'(88);
			1522: out = 16'(-19264);
			1523: out = 16'(10975);
			1524: out = 16'(23304);
			1525: out = 16'(-3372);
			1526: out = 16'(-17257);
			1527: out = 16'(-29633);
			1528: out = 16'(15399);
			1529: out = 16'(8476);
			1530: out = 16'(-1346);
			1531: out = 16'(-25996);
			1532: out = 16'(-15062);
			1533: out = 16'(12395);
			1534: out = 16'(8948);
			1535: out = 16'(10681);
			1536: out = 16'(6733);
			1537: out = 16'(906);
			1538: out = 16'(-2558);
			1539: out = 16'(4951);
			1540: out = 16'(5822);
			1541: out = 16'(7225);
			1542: out = 16'(-14680);
			1543: out = 16'(7434);
			1544: out = 16'(17050);
			1545: out = 16'(11392);
			1546: out = 16'(-11874);
			1547: out = 16'(-31002);
			1548: out = 16'(-15988);
			1549: out = 16'(3522);
			1550: out = 16'(24964);
			1551: out = 16'(8249);
			1552: out = 16'(7047);
			1553: out = 16'(3502);
			1554: out = 16'(1879);
			1555: out = 16'(-1435);
			1556: out = 16'(875);
			1557: out = 16'(-771);
			1558: out = 16'(-1884);
			1559: out = 16'(-21902);
			1560: out = 16'(5381);
			1561: out = 16'(16682);
			1562: out = 16'(2241);
			1563: out = 16'(-11545);
			1564: out = 16'(-21712);
			1565: out = 16'(13042);
			1566: out = 16'(8895);
			1567: out = 16'(1205);
			1568: out = 16'(17929);
			1569: out = 16'(11202);
			1570: out = 16'(-1408);
			1571: out = 16'(-9792);
			1572: out = 16'(-12730);
			1573: out = 16'(-8809);
			1574: out = 16'(1546);
			1575: out = 16'(4438);
			1576: out = 16'(-9079);
			1577: out = 16'(5454);
			1578: out = 16'(9782);
			1579: out = 16'(-2153);
			1580: out = 16'(641);
			1581: out = 16'(2747);
			1582: out = 16'(21349);
			1583: out = 16'(-4329);
			1584: out = 16'(-30798);
			1585: out = 16'(-4497);
			1586: out = 16'(6332);
			1587: out = 16'(18655);
			1588: out = 16'(-14805);
			1589: out = 16'(-12483);
			1590: out = 16'(6448);
			1591: out = 16'(459);
			1592: out = 16'(1387);
			1593: out = 16'(976);
			1594: out = 16'(6019);
			1595: out = 16'(5302);
			1596: out = 16'(-1355);
			1597: out = 16'(-5297);
			1598: out = 16'(-6664);
			1599: out = 16'(1842);
			1600: out = 16'(1610);
			1601: out = 16'(1093);
			1602: out = 16'(-821);
			1603: out = 16'(-8792);
			1604: out = 16'(-18833);
			1605: out = 16'(15809);
			1606: out = 16'(13990);
			1607: out = 16'(3583);
			1608: out = 16'(-5325);
			1609: out = 16'(-839);
			1610: out = 16'(19065);
			1611: out = 16'(6998);
			1612: out = 16'(-463);
			1613: out = 16'(-18576);
			1614: out = 16'(-10838);
			1615: out = 16'(-4328);
			1616: out = 16'(11268);
			1617: out = 16'(6438);
			1618: out = 16'(3416);
			1619: out = 16'(-12983);
			1620: out = 16'(4708);
			1621: out = 16'(21089);
			1622: out = 16'(-824);
			1623: out = 16'(-9806);
			1624: out = 16'(-19594);
			1625: out = 16'(-3874);
			1626: out = 16'(7170);
			1627: out = 16'(18842);
			1628: out = 16'(12449);
			1629: out = 16'(4250);
			1630: out = 16'(-13301);
			1631: out = 16'(-11391);
			1632: out = 16'(-7167);
			1633: out = 16'(10059);
			1634: out = 16'(7945);
			1635: out = 16'(6776);
			1636: out = 16'(-10177);
			1637: out = 16'(2817);
			1638: out = 16'(12744);
			1639: out = 16'(6681);
			1640: out = 16'(-10382);
			1641: out = 16'(-31492);
			1642: out = 16'(-5168);
			1643: out = 16'(7809);
			1644: out = 16'(20044);
			1645: out = 16'(2881);
			1646: out = 16'(-1039);
			1647: out = 16'(-4103);
			1648: out = 16'(6817);
			1649: out = 16'(5313);
			1650: out = 16'(-7145);
			1651: out = 16'(-22282);
			1652: out = 16'(-22538);
			1653: out = 16'(24817);
			1654: out = 16'(22156);
			1655: out = 16'(14888);
			1656: out = 16'(-22101);
			1657: out = 16'(-29067);
			1658: out = 16'(-27750);
			1659: out = 16'(-3290);
			1660: out = 16'(2897);
			1661: out = 16'(-1358);
			1662: out = 16'(15924);
			1663: out = 16'(12769);
			1664: out = 16'(-245);
			1665: out = 16'(-5624);
			1666: out = 16'(-5442);
			1667: out = 16'(14684);
			1668: out = 16'(-16608);
			1669: out = 16'(-25524);
			1670: out = 16'(7490);
			1671: out = 16'(11092);
			1672: out = 16'(11247);
			1673: out = 16'(-18034);
			1674: out = 16'(-3862);
			1675: out = 16'(12342);
			1676: out = 16'(-13641);
			1677: out = 16'(-8060);
			1678: out = 16'(2980);
			1679: out = 16'(16740);
			1680: out = 16'(9033);
			1681: out = 16'(-19822);
			1682: out = 16'(8217);
			1683: out = 16'(9005);
			1684: out = 16'(1748);
			1685: out = 16'(-13163);
			1686: out = 16'(-13871);
			1687: out = 16'(7823);
			1688: out = 16'(15412);
			1689: out = 16'(16460);
			1690: out = 16'(-7957);
			1691: out = 16'(-9463);
			1692: out = 16'(-8702);
			1693: out = 16'(3602);
			1694: out = 16'(10212);
			1695: out = 16'(15313);
			1696: out = 16'(-1481);
			1697: out = 16'(-7395);
			1698: out = 16'(-12228);
			1699: out = 16'(-697);
			1700: out = 16'(-730);
			1701: out = 16'(-10953);
			1702: out = 16'(-1083);
			1703: out = 16'(6538);
			1704: out = 16'(21765);
			1705: out = 16'(4093);
			1706: out = 16'(-5905);
			1707: out = 16'(-7169);
			1708: out = 16'(218);
			1709: out = 16'(6046);
			1710: out = 16'(-5291);
			1711: out = 16'(-6949);
			1712: out = 16'(-8273);
			1713: out = 16'(799);
			1714: out = 16'(3587);
			1715: out = 16'(5384);
			1716: out = 16'(8303);
			1717: out = 16'(6729);
			1718: out = 16'(1467);
			1719: out = 16'(-2448);
			1720: out = 16'(-1095);
			1721: out = 16'(13889);
			1722: out = 16'(-4639);
			1723: out = 16'(-6085);
			1724: out = 16'(16990);
			1725: out = 16'(11187);
			1726: out = 16'(3652);
			1727: out = 16'(-23034);
			1728: out = 16'(-16108);
			1729: out = 16'(-2199);
			1730: out = 16'(4280);
			1731: out = 16'(15673);
			1732: out = 16'(20580);
			1733: out = 16'(6807);
			1734: out = 16'(-8828);
			1735: out = 16'(-28599);
			1736: out = 16'(-6309);
			1737: out = 16'(1908);
			1738: out = 16'(-899);
			1739: out = 16'(7340);
			1740: out = 16'(6341);
			1741: out = 16'(429);
			1742: out = 16'(-5004);
			1743: out = 16'(-8031);
			1744: out = 16'(-10621);
			1745: out = 16'(-5971);
			1746: out = 16'(629);
			1747: out = 16'(20651);
			1748: out = 16'(15980);
			1749: out = 16'(7726);
			1750: out = 16'(-23998);
			1751: out = 16'(-18493);
			1752: out = 16'(4616);
			1753: out = 16'(2923);
			1754: out = 16'(5657);
			1755: out = 16'(2494);
			1756: out = 16'(3196);
			1757: out = 16'(-325);
			1758: out = 16'(-5849);
			1759: out = 16'(7848);
			1760: out = 16'(12762);
			1761: out = 16'(-6097);
			1762: out = 16'(4416);
			1763: out = 16'(7690);
			1764: out = 16'(4864);
			1765: out = 16'(2379);
			1766: out = 16'(1185);
			1767: out = 16'(-2998);
			1768: out = 16'(-7383);
			1769: out = 16'(-14517);
			1770: out = 16'(11594);
			1771: out = 16'(10412);
			1772: out = 16'(5483);
			1773: out = 16'(-21278);
			1774: out = 16'(-18622);
			1775: out = 16'(11686);
			1776: out = 16'(17524);
			1777: out = 16'(11993);
			1778: out = 16'(-31129);
			1779: out = 16'(-12275);
			1780: out = 16'(914);
			1781: out = 16'(17147);
			1782: out = 16'(4616);
			1783: out = 16'(-7253);
			1784: out = 16'(-21651);
			1785: out = 16'(-11413);
			1786: out = 16'(6543);
			1787: out = 16'(-566);
			1788: out = 16'(2565);
			1789: out = 16'(5);
			1790: out = 16'(15581);
			1791: out = 16'(13650);
			1792: out = 16'(11365);
			1793: out = 16'(-18331);
			1794: out = 16'(-21321);
			1795: out = 16'(7712);
			1796: out = 16'(9486);
			1797: out = 16'(8624);
			1798: out = 16'(-16397);
			1799: out = 16'(-9862);
			1800: out = 16'(-4675);
			1801: out = 16'(13776);
			1802: out = 16'(4875);
			1803: out = 16'(-2856);
			1804: out = 16'(3047);
			1805: out = 16'(3699);
			1806: out = 16'(2785);
			1807: out = 16'(-1299);
			1808: out = 16'(-2099);
			1809: out = 16'(2965);
			1810: out = 16'(-17520);
			1811: out = 16'(-22027);
			1812: out = 16'(-18384);
			1813: out = 16'(-1732);
			1814: out = 16'(9542);
			1815: out = 16'(16191);
			1816: out = 16'(6909);
			1817: out = 16'(-3045);
			1818: out = 16'(-19648);
			1819: out = 16'(-8109);
			1820: out = 16'(5053);
			1821: out = 16'(5475);
			1822: out = 16'(-6715);
			1823: out = 16'(-25790);
			1824: out = 16'(9189);
			1825: out = 16'(10572);
			1826: out = 16'(8553);
			1827: out = 16'(2293);
			1828: out = 16'(-314);
			1829: out = 16'(-5501);
			1830: out = 16'(6387);
			1831: out = 16'(9622);
			1832: out = 16'(9463);
			1833: out = 16'(7181);
			1834: out = 16'(3665);
			1835: out = 16'(-16220);
			1836: out = 16'(4399);
			1837: out = 16'(17257);
			1838: out = 16'(6790);
			1839: out = 16'(-4558);
			1840: out = 16'(-17743);
			1841: out = 16'(801);
			1842: out = 16'(4146);
			1843: out = 16'(8469);
			1844: out = 16'(5998);
			1845: out = 16'(3965);
			1846: out = 16'(-3699);
			1847: out = 16'(5989);
			1848: out = 16'(7373);
			1849: out = 16'(10696);
			1850: out = 16'(-10496);
			1851: out = 16'(-15146);
			1852: out = 16'(12385);
			1853: out = 16'(4206);
			1854: out = 16'(-1111);
			1855: out = 16'(-22777);
			1856: out = 16'(-9601);
			1857: out = 16'(5270);
			1858: out = 16'(12217);
			1859: out = 16'(7889);
			1860: out = 16'(-2934);
			1861: out = 16'(3217);
			1862: out = 16'(-2149);
			1863: out = 16'(-6701);
			1864: out = 16'(-1816);
			1865: out = 16'(7077);
			1866: out = 16'(19641);
			1867: out = 16'(-1131);
			1868: out = 16'(-6713);
			1869: out = 16'(15637);
			1870: out = 16'(-151);
			1871: out = 16'(-7414);
			1872: out = 16'(-31592);
			1873: out = 16'(-766);
			1874: out = 16'(22362);
			1875: out = 16'(17826);
			1876: out = 16'(1913);
			1877: out = 16'(-18493);
			1878: out = 16'(-20157);
			1879: out = 16'(-8712);
			1880: out = 16'(15132);
			1881: out = 16'(-491);
			1882: out = 16'(-563);
			1883: out = 16'(-1784);
			1884: out = 16'(-6562);
			1885: out = 16'(-4431);
			1886: out = 16'(15669);
			1887: out = 16'(-3723);
			1888: out = 16'(-8799);
			1889: out = 16'(733);
			1890: out = 16'(7691);
			1891: out = 16'(9514);
			1892: out = 16'(-22498);
			1893: out = 16'(-5185);
			1894: out = 16'(12079);
			1895: out = 16'(-10500);
			1896: out = 16'(-13891);
			1897: out = 16'(-17847);
			1898: out = 16'(15525);
			1899: out = 16'(8346);
			1900: out = 16'(-18650);
			1901: out = 16'(13989);
			1902: out = 16'(16562);
			1903: out = 16'(4107);
			1904: out = 16'(1420);
			1905: out = 16'(1244);
			1906: out = 16'(17508);
			1907: out = 16'(-3684);
			1908: out = 16'(-12668);
			1909: out = 16'(3637);
			1910: out = 16'(4549);
			1911: out = 16'(5694);
			1912: out = 16'(-4103);
			1913: out = 16'(75);
			1914: out = 16'(4717);
			1915: out = 16'(-6142);
			1916: out = 16'(-5713);
			1917: out = 16'(-1903);
			1918: out = 16'(7860);
			1919: out = 16'(3897);
			1920: out = 16'(-15720);
			1921: out = 16'(-1765);
			1922: out = 16'(4291);
			1923: out = 16'(19863);
			1924: out = 16'(-5340);
			1925: out = 16'(-16906);
			1926: out = 16'(-19550);
			1927: out = 16'(-2916);
			1928: out = 16'(10055);
			1929: out = 16'(12317);
			1930: out = 16'(6367);
			1931: out = 16'(-1078);
			1932: out = 16'(-12640);
			1933: out = 16'(-5524);
			1934: out = 16'(6272);
			1935: out = 16'(12266);
			1936: out = 16'(91);
			1937: out = 16'(-27263);
			1938: out = 16'(-15065);
			1939: out = 16'(-2339);
			1940: out = 16'(19498);
			1941: out = 16'(13071);
			1942: out = 16'(10635);
			1943: out = 16'(11890);
			1944: out = 16'(-2298);
			1945: out = 16'(-12005);
			1946: out = 16'(-13384);
			1947: out = 16'(-6286);
			1948: out = 16'(3609);
			1949: out = 16'(15540);
			1950: out = 16'(15407);
			1951: out = 16'(10998);
			1952: out = 16'(-18464);
			1953: out = 16'(-23930);
			1954: out = 16'(-19009);
			1955: out = 16'(7980);
			1956: out = 16'(16123);
			1957: out = 16'(12934);
			1958: out = 16'(-4351);
			1959: out = 16'(-12258);
			1960: out = 16'(-6193);
			1961: out = 16'(6183);
			1962: out = 16'(14524);
			1963: out = 16'(6626);
			1964: out = 16'(4307);
			1965: out = 16'(-1948);
			1966: out = 16'(-8007);
			1967: out = 16'(-451);
			1968: out = 16'(11468);
			1969: out = 16'(-4583);
			1970: out = 16'(1566);
			1971: out = 16'(6824);
			1972: out = 16'(-267);
			1973: out = 16'(-7250);
			1974: out = 16'(-13082);
			1975: out = 16'(1503);
			1976: out = 16'(12505);
			1977: out = 16'(16198);
			1978: out = 16'(19852);
			1979: out = 16'(8994);
			1980: out = 16'(-22211);
			1981: out = 16'(-23397);
			1982: out = 16'(-16524);
			1983: out = 16'(1553);
			1984: out = 16'(6954);
			1985: out = 16'(7783);
			1986: out = 16'(23452);
			1987: out = 16'(2467);
			1988: out = 16'(-23619);
			1989: out = 16'(-19289);
			1990: out = 16'(-8169);
			1991: out = 16'(15010);
			1992: out = 16'(-9827);
			1993: out = 16'(-7519);
			1994: out = 16'(9010);
			1995: out = 16'(2107);
			1996: out = 16'(-2817);
			1997: out = 16'(-20093);
			1998: out = 16'(5721);
			1999: out = 16'(16247);
			2000: out = 16'(932);
			2001: out = 16'(-6377);
			2002: out = 16'(-12607);
			2003: out = 16'(6492);
			2004: out = 16'(4156);
			2005: out = 16'(1871);
			2006: out = 16'(-2045);
			2007: out = 16'(2970);
			2008: out = 16'(11225);
			2009: out = 16'(-23968);
			2010: out = 16'(-22321);
			2011: out = 16'(1288);
			2012: out = 16'(12055);
			2013: out = 16'(13379);
			2014: out = 16'(-3934);
			2015: out = 16'(6336);
			2016: out = 16'(5360);
			2017: out = 16'(-3098);
			2018: out = 16'(-5992);
			2019: out = 16'(-4431);
			2020: out = 16'(8666);
			2021: out = 16'(7385);
			2022: out = 16'(4279);
			2023: out = 16'(3131);
			2024: out = 16'(-6108);
			2025: out = 16'(-17273);
			2026: out = 16'(1574);
			2027: out = 16'(8134);
			2028: out = 16'(16460);
			2029: out = 16'(-21563);
			2030: out = 16'(-23085);
			2031: out = 16'(1964);
			2032: out = 16'(19950);
			2033: out = 16'(18885);
			2034: out = 16'(-22874);
			2035: out = 16'(-664);
			2036: out = 16'(7450);
			2037: out = 16'(-107);
			2038: out = 16'(-9233);
			2039: out = 16'(-13399);
			2040: out = 16'(24082);
			2041: out = 16'(15329);
			2042: out = 16'(4164);
			2043: out = 16'(-13803);
			2044: out = 16'(-13752);
			2045: out = 16'(-5129);
			2046: out = 16'(3706);
			2047: out = 16'(11252);
			2048: out = 16'(19656);
			2049: out = 16'(-17172);
			2050: out = 16'(-20949);
			2051: out = 16'(18984);
			2052: out = 16'(9456);
			2053: out = 16'(5234);
			2054: out = 16'(-24442);
			2055: out = 16'(-743);
			2056: out = 16'(11341);
			2057: out = 16'(1995);
			2058: out = 16'(-7892);
			2059: out = 16'(-14893);
			2060: out = 16'(12773);
			2061: out = 16'(14041);
			2062: out = 16'(9985);
			2063: out = 16'(3360);
			2064: out = 16'(-1073);
			2065: out = 16'(-73);
			2066: out = 16'(-11973);
			2067: out = 16'(-7414);
			2068: out = 16'(6840);
			2069: out = 16'(11989);
			2070: out = 16'(9608);
			2071: out = 16'(-5663);
			2072: out = 16'(-3053);
			2073: out = 16'(-98);
			2074: out = 16'(-4119);
			2075: out = 16'(13050);
			2076: out = 16'(21417);
			2077: out = 16'(2610);
			2078: out = 16'(-13570);
			2079: out = 16'(-29494);
			2080: out = 16'(-3949);
			2081: out = 16'(5764);
			2082: out = 16'(11301);
			2083: out = 16'(10715);
			2084: out = 16'(4004);
			2085: out = 16'(-9645);
			2086: out = 16'(-5217);
			2087: out = 16'(-3049);
			2088: out = 16'(-1219);
			2089: out = 16'(1374);
			2090: out = 16'(3658);
			2091: out = 16'(13174);
			2092: out = 16'(-1996);
			2093: out = 16'(-14185);
			2094: out = 16'(-20257);
			2095: out = 16'(-7706);
			2096: out = 16'(9105);
			2097: out = 16'(1505);
			2098: out = 16'(3156);
			2099: out = 16'(42);
			2100: out = 16'(3187);
			2101: out = 16'(-1669);
			2102: out = 16'(-6510);
			2103: out = 16'(-7426);
			2104: out = 16'(-653);
			2105: out = 16'(16077);
			2106: out = 16'(-523);
			2107: out = 16'(-4607);
			2108: out = 16'(12759);
			2109: out = 16'(1169);
			2110: out = 16'(-4289);
			2111: out = 16'(-6001);
			2112: out = 16'(7951);
			2113: out = 16'(16419);
			2114: out = 16'(-27691);
			2115: out = 16'(-16090);
			2116: out = 16'(6346);
			2117: out = 16'(5772);
			2118: out = 16'(862);
			2119: out = 16'(-14588);
			2120: out = 16'(16607);
			2121: out = 16'(8401);
			2122: out = 16'(-29099);
			2123: out = 16'(-11734);
			2124: out = 16'(639);
			2125: out = 16'(25015);
			2126: out = 16'(-815);
			2127: out = 16'(-13480);
			2128: out = 16'(-4467);
			2129: out = 16'(-1770);
			2130: out = 16'(2522);
			2131: out = 16'(6574);
			2132: out = 16'(5699);
			2133: out = 16'(3912);
			2134: out = 16'(-324);
			2135: out = 16'(2176);
			2136: out = 16'(5772);
			2137: out = 16'(18429);
			2138: out = 16'(6853);
			2139: out = 16'(-26050);
			2140: out = 16'(-5589);
			2141: out = 16'(2215);
			2142: out = 16'(9756);
			2143: out = 16'(1962);
			2144: out = 16'(253);
			2145: out = 16'(8158);
			2146: out = 16'(479);
			2147: out = 16'(-2243);
			2148: out = 16'(15591);
			2149: out = 16'(13637);
			2150: out = 16'(10702);
			2151: out = 16'(-20614);
			2152: out = 16'(-10365);
			2153: out = 16'(10892);
			2154: out = 16'(-1131);
			2155: out = 16'(-6115);
			2156: out = 16'(-20685);
			2157: out = 16'(13312);
			2158: out = 16'(14700);
			2159: out = 16'(929);
			2160: out = 16'(-11674);
			2161: out = 16'(-12755);
			2162: out = 16'(12685);
			2163: out = 16'(5891);
			2164: out = 16'(3338);
			2165: out = 16'(-9662);
			2166: out = 16'(-3210);
			2167: out = 16'(621);
			2168: out = 16'(5253);
			2169: out = 16'(1921);
			2170: out = 16'(-306);
			2171: out = 16'(-19648);
			2172: out = 16'(-6163);
			2173: out = 16'(19367);
			2174: out = 16'(5534);
			2175: out = 16'(4320);
			2176: out = 16'(813);
			2177: out = 16'(5442);
			2178: out = 16'(4284);
			2179: out = 16'(319);
			2180: out = 16'(-2781);
			2181: out = 16'(-3774);
			2182: out = 16'(4103);
			2183: out = 16'(-5431);
			2184: out = 16'(-9373);
			2185: out = 16'(2887);
			2186: out = 16'(3525);
			2187: out = 16'(2818);
			2188: out = 16'(727);
			2189: out = 16'(-323);
			2190: out = 16'(1104);
			2191: out = 16'(-3476);
			2192: out = 16'(2321);
			2193: out = 16'(9621);
			2194: out = 16'(8114);
			2195: out = 16'(3981);
			2196: out = 16'(182);
			2197: out = 16'(-8371);
			2198: out = 16'(-12344);
			2199: out = 16'(-22685);
			2200: out = 16'(3881);
			2201: out = 16'(18442);
			2202: out = 16'(19004);
			2203: out = 16'(-3733);
			2204: out = 16'(-25128);
			2205: out = 16'(-7303);
			2206: out = 16'(-2522);
			2207: out = 16'(7155);
			2208: out = 16'(9157);
			2209: out = 16'(8562);
			2210: out = 16'(-228);
			2211: out = 16'(854);
			2212: out = 16'(-5851);
			2213: out = 16'(-9708);
			2214: out = 16'(-14254);
			2215: out = 16'(-7106);
			2216: out = 16'(10475);
			2217: out = 16'(11511);
			2218: out = 16'(9360);
			2219: out = 16'(-6603);
			2220: out = 16'(3987);
			2221: out = 16'(9425);
			2222: out = 16'(3514);
			2223: out = 16'(-5892);
			2224: out = 16'(-17033);
			2225: out = 16'(-3793);
			2226: out = 16'(-6611);
			2227: out = 16'(-6457);
			2228: out = 16'(-24525);
			2229: out = 16'(-8402);
			2230: out = 16'(24781);
			2231: out = 16'(8839);
			2232: out = 16'(-2721);
			2233: out = 16'(-32145);
			2234: out = 16'(4065);
			2235: out = 16'(19164);
			2236: out = 16'(15281);
			2237: out = 16'(6251);
			2238: out = 16'(-6759);
			2239: out = 16'(-26853);
			2240: out = 16'(-19814);
			2241: out = 16'(-5518);
			2242: out = 16'(2233);
			2243: out = 16'(4692);
			2244: out = 16'(635);
			2245: out = 16'(12091);
			2246: out = 16'(11570);
			2247: out = 16'(13683);
			2248: out = 16'(-25361);
			2249: out = 16'(-16321);
			2250: out = 16'(24893);
			2251: out = 16'(15343);
			2252: out = 16'(1949);
			2253: out = 16'(-30834);
			2254: out = 16'(-15335);
			2255: out = 16'(-1574);
			2256: out = 16'(9158);
			2257: out = 16'(8762);
			2258: out = 16'(6394);
			2259: out = 16'(9402);
			2260: out = 16'(-3412);
			2261: out = 16'(-13408);
			2262: out = 16'(18037);
			2263: out = 16'(12455);
			2264: out = 16'(-882);
			2265: out = 16'(1187);
			2266: out = 16'(-3761);
			2267: out = 16'(-4008);
			2268: out = 16'(-14287);
			2269: out = 16'(-6011);
			2270: out = 16'(14426);
			2271: out = 16'(18280);
			2272: out = 16'(13223);
			2273: out = 16'(-8387);
			2274: out = 16'(-12870);
			2275: out = 16'(-11302);
			2276: out = 16'(10600);
			2277: out = 16'(15716);
			2278: out = 16'(17317);
			2279: out = 16'(112);
			2280: out = 16'(-4030);
			2281: out = 16'(-7730);
			2282: out = 16'(-2547);
			2283: out = 16'(-7600);
			2284: out = 16'(-16992);
			2285: out = 16'(8102);
			2286: out = 16'(15314);
			2287: out = 16'(15194);
			2288: out = 16'(5781);
			2289: out = 16'(647);
			2290: out = 16'(194);
			2291: out = 16'(7585);
			2292: out = 16'(10848);
			2293: out = 16'(-688);
			2294: out = 16'(2489);
			2295: out = 16'(725);
			2296: out = 16'(-9213);
			2297: out = 16'(-15488);
			2298: out = 16'(-17876);
			2299: out = 16'(-2039);
			2300: out = 16'(7443);
			2301: out = 16'(15991);
			2302: out = 16'(3555);
			2303: out = 16'(96);
			2304: out = 16'(-5009);
			2305: out = 16'(14405);
			2306: out = 16'(17743);
			2307: out = 16'(14889);
			2308: out = 16'(-12760);
			2309: out = 16'(-24851);
			2310: out = 16'(3783);
			2311: out = 16'(-4922);
			2312: out = 16'(-5841);
			2313: out = 16'(-17461);
			2314: out = 16'(3654);
			2315: out = 16'(18752);
			2316: out = 16'(2473);
			2317: out = 16'(-5118);
			2318: out = 16'(-14435);
			2319: out = 16'(-146);
			2320: out = 16'(9815);
			2321: out = 16'(24899);
			2322: out = 16'(-12275);
			2323: out = 16'(-25748);
			2324: out = 16'(-31086);
			2325: out = 16'(-2344);
			2326: out = 16'(14627);
			2327: out = 16'(2955);
			2328: out = 16'(4347);
			2329: out = 16'(-71);
			2330: out = 16'(11259);
			2331: out = 16'(-14487);
			2332: out = 16'(-27819);
			2333: out = 16'(9353);
			2334: out = 16'(12507);
			2335: out = 16'(8290);
			2336: out = 16'(-2405);
			2337: out = 16'(-10655);
			2338: out = 16'(-16512);
			2339: out = 16'(-4425);
			2340: out = 16'(-8684);
			2341: out = 16'(-31167);
			2342: out = 16'(9355);
			2343: out = 16'(21554);
			2344: out = 16'(17069);
			2345: out = 16'(6817);
			2346: out = 16'(375);
			2347: out = 16'(2538);
			2348: out = 16'(1729);
			2349: out = 16'(1225);
			2350: out = 16'(9178);
			2351: out = 16'(-9078);
			2352: out = 16'(-26619);
			2353: out = 16'(-17419);
			2354: out = 16'(-2703);
			2355: out = 16'(17593);
			2356: out = 16'(-10043);
			2357: out = 16'(-7412);
			2358: out = 16'(2906);
			2359: out = 16'(3462);
			2360: out = 16'(6829);
			2361: out = 16'(9291);
			2362: out = 16'(16046);
			2363: out = 16'(11063);
			2364: out = 16'(-13657);
			2365: out = 16'(-11655);
			2366: out = 16'(-9600);
			2367: out = 16'(1302);
			2368: out = 16'(1830);
			2369: out = 16'(3166);
			2370: out = 16'(-7005);
			2371: out = 16'(6810);
			2372: out = 16'(20733);
			2373: out = 16'(888);
			2374: out = 16'(-3);
			2375: out = 16'(615);
			2376: out = 16'(935);
			2377: out = 16'(1027);
			2378: out = 16'(3126);
			2379: out = 16'(4834);
			2380: out = 16'(6686);
			2381: out = 16'(2425);
			2382: out = 16'(8247);
			2383: out = 16'(6114);
			2384: out = 16'(3815);
			2385: out = 16'(-16572);
			2386: out = 16'(-23945);
			2387: out = 16'(17323);
			2388: out = 16'(13057);
			2389: out = 16'(6267);
			2390: out = 16'(12707);
			2391: out = 16'(6239);
			2392: out = 16'(-15);
			2393: out = 16'(-25177);
			2394: out = 16'(-20652);
			2395: out = 16'(869);
			2396: out = 16'(8363);
			2397: out = 16'(4137);
			2398: out = 16'(-22188);
			2399: out = 16'(-1408);
			2400: out = 16'(6563);
			2401: out = 16'(4389);
			2402: out = 16'(13577);
			2403: out = 16'(17348);
			2404: out = 16'(15483);
			2405: out = 16'(-77);
			2406: out = 16'(-15189);
			2407: out = 16'(5694);
			2408: out = 16'(-7020);
			2409: out = 16'(-19229);
			2410: out = 16'(-12884);
			2411: out = 16'(-5952);
			2412: out = 16'(3840);
			2413: out = 16'(3732);
			2414: out = 16'(8148);
			2415: out = 16'(11949);
			2416: out = 16'(14787);
			2417: out = 16'(12025);
			2418: out = 16'(2403);
			2419: out = 16'(7422);
			2420: out = 16'(6430);
			2421: out = 16'(-8154);
			2422: out = 16'(-6481);
			2423: out = 16'(-5645);
			2424: out = 16'(1805);
			2425: out = 16'(2761);
			2426: out = 16'(4438);
			2427: out = 16'(-27921);
			2428: out = 16'(-11154);
			2429: out = 16'(16742);
			2430: out = 16'(15445);
			2431: out = 16'(7002);
			2432: out = 16'(-14473);
			2433: out = 16'(-9892);
			2434: out = 16'(-6979);
			2435: out = 16'(7706);
			2436: out = 16'(-7581);
			2437: out = 16'(-9728);
			2438: out = 16'(605);
			2439: out = 16'(1018);
			2440: out = 16'(2069);
			2441: out = 16'(496);
			2442: out = 16'(1650);
			2443: out = 16'(2925);
			2444: out = 16'(17230);
			2445: out = 16'(8275);
			2446: out = 16'(-2909);
			2447: out = 16'(560);
			2448: out = 16'(-6297);
			2449: out = 16'(-18037);
			2450: out = 16'(4811);
			2451: out = 16'(5914);
			2452: out = 16'(-304);
			2453: out = 16'(-23905);
			2454: out = 16'(-23649);
			2455: out = 16'(9299);
			2456: out = 16'(17644);
			2457: out = 16'(21698);
			2458: out = 16'(14660);
			2459: out = 16'(3712);
			2460: out = 16'(-8767);
			2461: out = 16'(-4049);
			2462: out = 16'(-10299);
			2463: out = 16'(-10959);
			2464: out = 16'(-11502);
			2465: out = 16'(-4086);
			2466: out = 16'(2225);
			2467: out = 16'(5261);
			2468: out = 16'(-476);
			2469: out = 16'(-12217);
			2470: out = 16'(-3998);
			2471: out = 16'(-799);
			2472: out = 16'(2632);
			2473: out = 16'(-7568);
			2474: out = 16'(-4023);
			2475: out = 16'(29736);
			2476: out = 16'(8411);
			2477: out = 16'(-6707);
			2478: out = 16'(-31979);
			2479: out = 16'(-5426);
			2480: out = 16'(21261);
			2481: out = 16'(2702);
			2482: out = 16'(-12212);
			2483: out = 16'(-30970);
			2484: out = 16'(13600);
			2485: out = 16'(20419);
			2486: out = 16'(18015);
			2487: out = 16'(5607);
			2488: out = 16'(-2350);
			2489: out = 16'(-10108);
			2490: out = 16'(5740);
			2491: out = 16'(9319);
			2492: out = 16'(-3907);
			2493: out = 16'(-1344);
			2494: out = 16'(-915);
			2495: out = 16'(17735);
			2496: out = 16'(-6399);
			2497: out = 16'(-19806);
			2498: out = 16'(-5478);
			2499: out = 16'(9362);
			2500: out = 16'(21894);
			2501: out = 16'(12277);
			2502: out = 16'(5302);
			2503: out = 16'(-6073);
			2504: out = 16'(-896);
			2505: out = 16'(-5487);
			2506: out = 16'(-12299);
			2507: out = 16'(-9763);
			2508: out = 16'(-1865);
			2509: out = 16'(19623);
			2510: out = 16'(-6219);
			2511: out = 16'(-15344);
			2512: out = 16'(-13861);
			2513: out = 16'(9137);
			2514: out = 16'(24280);
			2515: out = 16'(20843);
			2516: out = 16'(11500);
			2517: out = 16'(-2645);
			2518: out = 16'(-7689);
			2519: out = 16'(-18202);
			2520: out = 16'(-24005);
			2521: out = 16'(3606);
			2522: out = 16'(12901);
			2523: out = 16'(16835);
			2524: out = 16'(-8360);
			2525: out = 16'(-17836);
			2526: out = 16'(-19927);
			2527: out = 16'(7066);
			2528: out = 16'(19535);
			2529: out = 16'(13867);
			2530: out = 16'(7335);
			2531: out = 16'(-231);
			2532: out = 16'(5894);
			2533: out = 16'(-3969);
			2534: out = 16'(-8577);
			2535: out = 16'(1140);
			2536: out = 16'(-882);
			2537: out = 16'(-3510);
			2538: out = 16'(-16126);
			2539: out = 16'(-4342);
			2540: out = 16'(17910);
			2541: out = 16'(5436);
			2542: out = 16'(8711);
			2543: out = 16'(10534);
			2544: out = 16'(7267);
			2545: out = 16'(-3207);
			2546: out = 16'(-20738);
			2547: out = 16'(-14727);
			2548: out = 16'(-7870);
			2549: out = 16'(-8690);
			2550: out = 16'(9510);
			2551: out = 16'(18028);
			2552: out = 16'(8727);
			2553: out = 16'(-3192);
			2554: out = 16'(-15812);
			2555: out = 16'(9125);
			2556: out = 16'(5724);
			2557: out = 16'(3427);
			2558: out = 16'(-7339);
			2559: out = 16'(3191);
			2560: out = 16'(21220);
			2561: out = 16'(4289);
			2562: out = 16'(-8562);
			2563: out = 16'(-27947);
			2564: out = 16'(-16089);
			2565: out = 16'(-6111);
			2566: out = 16'(-631);
			2567: out = 16'(13837);
			2568: out = 16'(17518);
			2569: out = 16'(-3000);
			2570: out = 16'(-1461);
			2571: out = 16'(-920);
			2572: out = 16'(10187);
			2573: out = 16'(-6106);
			2574: out = 16'(-26081);
			2575: out = 16'(11292);
			2576: out = 16'(9575);
			2577: out = 16'(2413);
			2578: out = 16'(-22352);
			2579: out = 16'(-20820);
			2580: out = 16'(4508);
			2581: out = 16'(133);
			2582: out = 16'(-77);
			2583: out = 16'(-12939);
			2584: out = 16'(12807);
			2585: out = 16'(18473);
			2586: out = 16'(-10718);
			2587: out = 16'(-3621);
			2588: out = 16'(382);
			2589: out = 16'(13400);
			2590: out = 16'(-7316);
			2591: out = 16'(-29421);
			2592: out = 16'(-8005);
			2593: out = 16'(-814);
			2594: out = 16'(9874);
			2595: out = 16'(-5798);
			2596: out = 16'(9);
			2597: out = 16'(9387);
			2598: out = 16'(9738);
			2599: out = 16'(8092);
			2600: out = 16'(9930);
			2601: out = 16'(-3924);
			2602: out = 16'(-10349);
			2603: out = 16'(-21546);
			2604: out = 16'(4844);
			2605: out = 16'(17581);
			2606: out = 16'(4522);
			2607: out = 16'(-13067);
			2608: out = 16'(-28756);
			2609: out = 16'(892);
			2610: out = 16'(2314);
			2611: out = 16'(2696);
			2612: out = 16'(15781);
			2613: out = 16'(12345);
			2614: out = 16'(2569);
			2615: out = 16'(-9354);
			2616: out = 16'(-5473);
			2617: out = 16'(19914);
			2618: out = 16'(-11659);
			2619: out = 16'(-15991);
			2620: out = 16'(3994);
			2621: out = 16'(1218);
			2622: out = 16'(-359);
			2623: out = 16'(-17192);
			2624: out = 16'(2675);
			2625: out = 16'(17487);
			2626: out = 16'(15947);
			2627: out = 16'(16714);
			2628: out = 16'(12760);
			2629: out = 16'(-9965);
			2630: out = 16'(-14271);
			2631: out = 16'(-12080);
			2632: out = 16'(6779);
			2633: out = 16'(3675);
			2634: out = 16'(-14872);
			2635: out = 16'(-3916);
			2636: out = 16'(2798);
			2637: out = 16'(18511);
			2638: out = 16'(3347);
			2639: out = 16'(-740);
			2640: out = 16'(-48);
			2641: out = 16'(8189);
			2642: out = 16'(10449);
			2643: out = 16'(-2444);
			2644: out = 16'(-1970);
			2645: out = 16'(-761);
			2646: out = 16'(1167);
			2647: out = 16'(1310);
			2648: out = 16'(176);
			2649: out = 16'(11594);
			2650: out = 16'(1339);
			2651: out = 16'(-18460);
			2652: out = 16'(836);
			2653: out = 16'(9468);
			2654: out = 16'(19398);
			2655: out = 16'(2579);
			2656: out = 16'(-7536);
			2657: out = 16'(-19273);
			2658: out = 16'(-6600);
			2659: out = 16'(4301);
			2660: out = 16'(12546);
			2661: out = 16'(4346);
			2662: out = 16'(-3378);
			2663: out = 16'(8887);
			2664: out = 16'(7557);
			2665: out = 16'(8049);
			2666: out = 16'(-24899);
			2667: out = 16'(-15330);
			2668: out = 16'(5992);
			2669: out = 16'(15527);
			2670: out = 16'(9967);
			2671: out = 16'(-13323);
			2672: out = 16'(-2236);
			2673: out = 16'(4010);
			2674: out = 16'(27179);
			2675: out = 16'(-9695);
			2676: out = 16'(-26132);
			2677: out = 16'(-30469);
			2678: out = 16'(-13415);
			2679: out = 16'(4961);
			2680: out = 16'(24747);
			2681: out = 16'(9381);
			2682: out = 16'(-7126);
			2683: out = 16'(-15404);
			2684: out = 16'(-8887);
			2685: out = 16'(4921);
			2686: out = 16'(11341);
			2687: out = 16'(10019);
			2688: out = 16'(457);
			2689: out = 16'(-1434);
			2690: out = 16'(-11324);
			2691: out = 16'(-29288);
			2692: out = 16'(1523);
			2693: out = 16'(15074);
			2694: out = 16'(14325);
			2695: out = 16'(-5691);
			2696: out = 16'(-18409);
			2697: out = 16'(1030);
			2698: out = 16'(-1253);
			2699: out = 16'(3172);
			2700: out = 16'(4916);
			2701: out = 16'(10630);
			2702: out = 16'(9876);
			2703: out = 16'(-10873);
			2704: out = 16'(-13429);
			2705: out = 16'(-4339);
			2706: out = 16'(-14005);
			2707: out = 16'(-2229);
			2708: out = 16'(14324);
			2709: out = 16'(20011);
			2710: out = 16'(10700);
			2711: out = 16'(-19415);
			2712: out = 16'(-13322);
			2713: out = 16'(-6598);
			2714: out = 16'(12073);
			2715: out = 16'(5636);
			2716: out = 16'(88);
			2717: out = 16'(-12478);
			2718: out = 16'(-4104);
			2719: out = 16'(5284);
			2720: out = 16'(-1945);
			2721: out = 16'(-4862);
			2722: out = 16'(-11126);
			2723: out = 16'(9676);
			2724: out = 16'(13420);
			2725: out = 16'(17937);
			2726: out = 16'(-22513);
			2727: out = 16'(-24110);
			2728: out = 16'(-1776);
			2729: out = 16'(21130);
			2730: out = 16'(22671);
			2731: out = 16'(1618);
			2732: out = 16'(-19325);
			2733: out = 16'(-28609);
			2734: out = 16'(1242);
			2735: out = 16'(8677);
			2736: out = 16'(14136);
			2737: out = 16'(15683);
			2738: out = 16'(12591);
			2739: out = 16'(6372);
			2740: out = 16'(-22242);
			2741: out = 16'(-17121);
			2742: out = 16'(5807);
			2743: out = 16'(6257);
			2744: out = 16'(8204);
			2745: out = 16'(-2763);
			2746: out = 16'(9774);
			2747: out = 16'(4709);
			2748: out = 16'(-7696);
			2749: out = 16'(-8075);
			2750: out = 16'(-3698);
			2751: out = 16'(908);
			2752: out = 16'(12698);
			2753: out = 16'(16488);
			2754: out = 16'(10066);
			2755: out = 16'(-11213);
			2756: out = 16'(-30438);
			2757: out = 16'(-1205);
			2758: out = 16'(12456);
			2759: out = 16'(26124);
			2760: out = 16'(-21775);
			2761: out = 16'(-21242);
			2762: out = 16'(-3555);
			2763: out = 16'(19582);
			2764: out = 16'(17142);
			2765: out = 16'(-10475);
			2766: out = 16'(-7109);
			2767: out = 16'(-5647);
			2768: out = 16'(10560);
			2769: out = 16'(1819);
			2770: out = 16'(-1008);
			2771: out = 16'(-7702);
			2772: out = 16'(8288);
			2773: out = 16'(19146);
			2774: out = 16'(690);
			2775: out = 16'(215);
			2776: out = 16'(-1150);
			2777: out = 16'(10126);
			2778: out = 16'(8211);
			2779: out = 16'(5511);
			2780: out = 16'(-9332);
			2781: out = 16'(-6790);
			2782: out = 16'(8234);
			2783: out = 16'(2501);
			2784: out = 16'(2659);
			2785: out = 16'(7546);
			2786: out = 16'(-8091);
			2787: out = 16'(-12657);
			2788: out = 16'(11664);
			2789: out = 16'(3482);
			2790: out = 16'(-1866);
			2791: out = 16'(-15144);
			2792: out = 16'(-8517);
			2793: out = 16'(166);
			2794: out = 16'(-585);
			2795: out = 16'(2669);
			2796: out = 16'(4886);
			2797: out = 16'(5696);
			2798: out = 16'(5789);
			2799: out = 16'(5446);
			2800: out = 16'(-4142);
			2801: out = 16'(-6707);
			2802: out = 16'(1408);
			2803: out = 16'(-9388);
			2804: out = 16'(-7677);
			2805: out = 16'(8612);
			2806: out = 16'(6951);
			2807: out = 16'(4314);
			2808: out = 16'(-2436);
			2809: out = 16'(1397);
			2810: out = 16'(5607);
			2811: out = 16'(-10296);
			2812: out = 16'(-6758);
			2813: out = 16'(-3826);
			2814: out = 16'(11358);
			2815: out = 16'(4050);
			2816: out = 16'(-7659);
			2817: out = 16'(-14543);
			2818: out = 16'(-7427);
			2819: out = 16'(9272);
			2820: out = 16'(17795);
			2821: out = 16'(12249);
			2822: out = 16'(-14184);
			2823: out = 16'(-16904);
			2824: out = 16'(-15387);
			2825: out = 16'(2142);
			2826: out = 16'(2499);
			2827: out = 16'(1261);
			2828: out = 16'(1760);
			2829: out = 16'(-6055);
			2830: out = 16'(-11545);
			2831: out = 16'(-20311);
			2832: out = 16'(-6013);
			2833: out = 16'(13531);
			2834: out = 16'(17616);
			2835: out = 16'(7420);
			2836: out = 16'(-16355);
			2837: out = 16'(-19576);
			2838: out = 16'(-13547);
			2839: out = 16'(14079);
			2840: out = 16'(9837);
			2841: out = 16'(8501);
			2842: out = 16'(-7526);
			2843: out = 16'(-460);
			2844: out = 16'(2222);
			2845: out = 16'(9970);
			2846: out = 16'(2706);
			2847: out = 16'(-2184);
			2848: out = 16'(-2496);
			2849: out = 16'(5303);
			2850: out = 16'(13957);
			2851: out = 16'(721);
			2852: out = 16'(-3902);
			2853: out = 16'(-10303);
			2854: out = 16'(2886);
			2855: out = 16'(5845);
			2856: out = 16'(8232);
			2857: out = 16'(-6826);
			2858: out = 16'(-7261);
			2859: out = 16'(11057);
			2860: out = 16'(7048);
			2861: out = 16'(5221);
			2862: out = 16'(443);
			2863: out = 16'(-2809);
			2864: out = 16'(-5463);
			2865: out = 16'(504);
			2866: out = 16'(404);
			2867: out = 16'(1235);
			2868: out = 16'(1717);
			2869: out = 16'(-2358);
			2870: out = 16'(-10456);
			2871: out = 16'(9565);
			2872: out = 16'(10839);
			2873: out = 16'(8425);
			2874: out = 16'(-2500);
			2875: out = 16'(-6703);
			2876: out = 16'(-9128);
			2877: out = 16'(8287);
			2878: out = 16'(14844);
			2879: out = 16'(6459);
			2880: out = 16'(1482);
			2881: out = 16'(-3572);
			2882: out = 16'(1659);
			2883: out = 16'(4270);
			2884: out = 16'(8684);
			2885: out = 16'(2198);
			2886: out = 16'(5071);
			2887: out = 16'(6006);
			2888: out = 16'(5829);
			2889: out = 16'(2442);
			2890: out = 16'(-863);
			2891: out = 16'(-3226);
			2892: out = 16'(-3130);
			2893: out = 16'(-2146);
			2894: out = 16'(1383);
			2895: out = 16'(2327);
			2896: out = 16'(1104);
			2897: out = 16'(-895);
			2898: out = 16'(-2325);
			2899: out = 16'(-2038);
			2900: out = 16'(-1264);
			2901: out = 16'(-356);
			2902: out = 16'(1415);
			2903: out = 16'(-3047);
			2904: out = 16'(-7981);
			2905: out = 16'(2074);
			2906: out = 16'(1526);
			2907: out = 16'(-56);
			2908: out = 16'(-1860);
			2909: out = 16'(2640);
			2910: out = 16'(13077);
			2911: out = 16'(-7878);
			2912: out = 16'(-15574);
			2913: out = 16'(-13225);
			2914: out = 16'(-7675);
			2915: out = 16'(2198);
			2916: out = 16'(12805);
			2917: out = 16'(18186);
			2918: out = 16'(15043);
			2919: out = 16'(-6168);
			2920: out = 16'(-19872);
			2921: out = 16'(-28261);
			2922: out = 16'(10347);
			2923: out = 16'(13426);
			2924: out = 16'(11417);
			2925: out = 16'(-19199);
			2926: out = 16'(-13234);
			2927: out = 16'(12183);
			2928: out = 16'(3170);
			2929: out = 16'(-1664);
			2930: out = 16'(-21007);
			2931: out = 16'(2134);
			2932: out = 16'(8008);
			2933: out = 16'(4966);
			2934: out = 16'(-5977);
			2935: out = 16'(-11455);
			2936: out = 16'(-2589);
			2937: out = 16'(3474);
			2938: out = 16'(7175);
			2939: out = 16'(-17621);
			2940: out = 16'(-13677);
			2941: out = 16'(-6134);
			2942: out = 16'(13413);
			2943: out = 16'(9808);
			2944: out = 16'(-2446);
			2945: out = 16'(2156);
			2946: out = 16'(3739);
			2947: out = 16'(10766);
			2948: out = 16'(1147);
			2949: out = 16'(-7081);
			2950: out = 16'(-30087);
			2951: out = 16'(-1907);
			2952: out = 16'(13682);
			2953: out = 16'(18525);
			2954: out = 16'(8500);
			2955: out = 16'(-1458);
			2956: out = 16'(-14708);
			2957: out = 16'(-2673);
			2958: out = 16'(12464);
			2959: out = 16'(12576);
			2960: out = 16'(13185);
			2961: out = 16'(8130);
			2962: out = 16'(-7684);
			2963: out = 16'(-16642);
			2964: out = 16'(-19884);
			2965: out = 16'(-3880);
			2966: out = 16'(7974);
			2967: out = 16'(16022);
			2968: out = 16'(6577);
			2969: out = 16'(-4122);
			2970: out = 16'(-22620);
			2971: out = 16'(-8702);
			2972: out = 16'(4097);
			2973: out = 16'(10040);
			2974: out = 16'(5851);
			2975: out = 16'(-1826);
			2976: out = 16'(-4046);
			2977: out = 16'(-6411);
			2978: out = 16'(-3959);
			2979: out = 16'(-183);
			2980: out = 16'(8538);
			2981: out = 16'(16173);
			2982: out = 16'(2223);
			2983: out = 16'(-5316);
			2984: out = 16'(-11811);
			2985: out = 16'(-4236);
			2986: out = 16'(2135);
			2987: out = 16'(8562);
			2988: out = 16'(3541);
			2989: out = 16'(-1398);
			2990: out = 16'(-6600);
			2991: out = 16'(-6581);
			2992: out = 16'(-2718);
			2993: out = 16'(12546);
			2994: out = 16'(7075);
			2995: out = 16'(-812);
			2996: out = 16'(-1971);
			2997: out = 16'(4292);
			2998: out = 16'(17343);
			2999: out = 16'(-15139);
			3000: out = 16'(-12155);
			3001: out = 16'(1384);
			3002: out = 16'(15135);
			3003: out = 16'(8838);
			3004: out = 16'(-22547);
			3005: out = 16'(-12627);
			3006: out = 16'(-7890);
			3007: out = 16'(930);
			3008: out = 16'(412);
			3009: out = 16'(2035);
			3010: out = 16'(4643);
			3011: out = 16'(1564);
			3012: out = 16'(-2281);
			3013: out = 16'(12437);
			3014: out = 16'(3498);
			3015: out = 16'(-6499);
			3016: out = 16'(-9750);
			3017: out = 16'(-1985);
			3018: out = 16'(13770);
			3019: out = 16'(6196);
			3020: out = 16'(1857);
			3021: out = 16'(-13796);
			3022: out = 16'(6423);
			3023: out = 16'(8308);
			3024: out = 16'(2877);
			3025: out = 16'(-14110);
			3026: out = 16'(-18784);
			3027: out = 16'(6182);
			3028: out = 16'(6734);
			3029: out = 16'(6890);
			3030: out = 16'(2511);
			3031: out = 16'(1531);
			3032: out = 16'(1311);
			3033: out = 16'(-11479);
			3034: out = 16'(929);
			3035: out = 16'(20447);
			3036: out = 16'(3804);
			3037: out = 16'(-1524);
			3038: out = 16'(-9657);
			3039: out = 16'(2786);
			3040: out = 16'(3975);
			3041: out = 16'(-5177);
			3042: out = 16'(3206);
			3043: out = 16'(5677);
			3044: out = 16'(6078);
			3045: out = 16'(-2386);
			3046: out = 16'(-7698);
			3047: out = 16'(-2884);
			3048: out = 16'(-2869);
			3049: out = 16'(-1813);
			3050: out = 16'(9995);
			3051: out = 16'(6216);
			3052: out = 16'(542);
			3053: out = 16'(-8121);
			3054: out = 16'(-1424);
			3055: out = 16'(14082);
			3056: out = 16'(8188);
			3057: out = 16'(5738);
			3058: out = 16'(-1430);
			3059: out = 16'(1583);
			3060: out = 16'(-3945);
			3061: out = 16'(-24678);
			3062: out = 16'(-10297);
			3063: out = 16'(3219);
			3064: out = 16'(16399);
			3065: out = 16'(8759);
			3066: out = 16'(-531);
			3067: out = 16'(-696);
			3068: out = 16'(-2570);
			3069: out = 16'(-1308);
			3070: out = 16'(-2217);
			3071: out = 16'(-777);
			3072: out = 16'(-8);
			3073: out = 16'(-5189);
			3074: out = 16'(-1452);
			3075: out = 16'(11694);
			3076: out = 16'(-5271);
			3077: out = 16'(-7816);
			3078: out = 16'(-1515);
			3079: out = 16'(6608);
			3080: out = 16'(6581);
			3081: out = 16'(-18234);
			3082: out = 16'(-10092);
			3083: out = 16'(-2629);
			3084: out = 16'(18639);
			3085: out = 16'(3198);
			3086: out = 16'(-12185);
			3087: out = 16'(-8973);
			3088: out = 16'(110);
			3089: out = 16'(14306);
			3090: out = 16'(-4223);
			3091: out = 16'(-6885);
			3092: out = 16'(-10731);
			3093: out = 16'(8832);
			3094: out = 16'(11844);
			3095: out = 16'(6376);
			3096: out = 16'(1512);
			3097: out = 16'(-5798);
			3098: out = 16'(-19035);
			3099: out = 16'(-10955);
			3100: out = 16'(-2217);
			3101: out = 16'(8286);
			3102: out = 16'(2032);
			3103: out = 16'(-3666);
			3104: out = 16'(12305);
			3105: out = 16'(3416);
			3106: out = 16'(-6814);
			3107: out = 16'(-906);
			3108: out = 16'(-3451);
			3109: out = 16'(-5102);
			3110: out = 16'(-5352);
			3111: out = 16'(4467);
			3112: out = 16'(20794);
			3113: out = 16'(10280);
			3114: out = 16'(-1011);
			3115: out = 16'(-26630);
			3116: out = 16'(-13428);
			3117: out = 16'(-2744);
			3118: out = 16'(9841);
			3119: out = 16'(7610);
			3120: out = 16'(3941);
			3121: out = 16'(-11556);
			3122: out = 16'(-3165);
			3123: out = 16'(6619);
			3124: out = 16'(11381);
			3125: out = 16'(3717);
			3126: out = 16'(-10355);
			3127: out = 16'(5282);
			3128: out = 16'(3324);
			3129: out = 16'(788);
			3130: out = 16'(-7481);
			3131: out = 16'(-4940);
			3132: out = 16'(5173);
			3133: out = 16'(7594);
			3134: out = 16'(2527);
			3135: out = 16'(-24664);
			3136: out = 16'(-7381);
			3137: out = 16'(5685);
			3138: out = 16'(14897);
			3139: out = 16'(7706);
			3140: out = 16'(-1780);
			3141: out = 16'(-4045);
			3142: out = 16'(-6763);
			3143: out = 16'(-4327);
			3144: out = 16'(-5443);
			3145: out = 16'(1714);
			3146: out = 16'(7320);
			3147: out = 16'(9229);
			3148: out = 16'(3036);
			3149: out = 16'(-7427);
			3150: out = 16'(-4285);
			3151: out = 16'(968);
			3152: out = 16'(8215);
			3153: out = 16'(9751);
			3154: out = 16'(7149);
			3155: out = 16'(967);
			3156: out = 16'(-2249);
			3157: out = 16'(-3626);
			3158: out = 16'(-14436);
			3159: out = 16'(-3492);
			3160: out = 16'(6606);
			3161: out = 16'(20347);
			3162: out = 16'(10347);
			3163: out = 16'(-3174);
			3164: out = 16'(-15644);
			3165: out = 16'(-5332);
			3166: out = 16'(19037);
			3167: out = 16'(13834);
			3168: out = 16'(5349);
			3169: out = 16'(-18804);
			3170: out = 16'(-17961);
			3171: out = 16'(-11880);
			3172: out = 16'(18737);
			3173: out = 16'(5948);
			3174: out = 16'(-1189);
			3175: out = 16'(-20912);
			3176: out = 16'(-1954);
			3177: out = 16'(14175);
			3178: out = 16'(-801);
			3179: out = 16'(2636);
			3180: out = 16'(3137);
			3181: out = 16'(19872);
			3182: out = 16'(7702);
			3183: out = 16'(-12422);
			3184: out = 16'(-10146);
			3185: out = 16'(-7513);
			3186: out = 16'(1274);
			3187: out = 16'(5437);
			3188: out = 16'(6782);
			3189: out = 16'(-3022);
			3190: out = 16'(6588);
			3191: out = 16'(6373);
			3192: out = 16'(-4234);
			3193: out = 16'(-7564);
			3194: out = 16'(-7500);
			3195: out = 16'(3255);
			3196: out = 16'(11698);
			3197: out = 16'(17394);
			3198: out = 16'(-19573);
			3199: out = 16'(-16133);
			3200: out = 16'(-4046);
			3201: out = 16'(11802);
			3202: out = 16'(5246);
			3203: out = 16'(-19433);
			3204: out = 16'(5096);
			3205: out = 16'(7413);
			3206: out = 16'(3106);
			3207: out = 16'(-15099);
			3208: out = 16'(-18663);
			3209: out = 16'(14381);
			3210: out = 16'(-5367);
			3211: out = 16'(-14223);
			3212: out = 16'(-22796);
			3213: out = 16'(-4457);
			3214: out = 16'(11186);
			3215: out = 16'(15232);
			3216: out = 16'(4791);
			3217: out = 16'(-10441);
			3218: out = 16'(-14544);
			3219: out = 16'(-10588);
			3220: out = 16'(3112);
			3221: out = 16'(7362);
			3222: out = 16'(10627);
			3223: out = 16'(6372);
			3224: out = 16'(1426);
			3225: out = 16'(-3523);
			3226: out = 16'(427);
			3227: out = 16'(-3606);
			3228: out = 16'(-4161);
			3229: out = 16'(-13670);
			3230: out = 16'(-4928);
			3231: out = 16'(1183);
			3232: out = 16'(12876);
			3233: out = 16'(1397);
			3234: out = 16'(-9631);
			3235: out = 16'(942);
			3236: out = 16'(7274);
			3237: out = 16'(13392);
			3238: out = 16'(7825);
			3239: out = 16'(-2308);
			3240: out = 16'(-21087);
			3241: out = 16'(-8084);
			3242: out = 16'(-1912);
			3243: out = 16'(6069);
			3244: out = 16'(-6188);
			3245: out = 16'(-8083);
			3246: out = 16'(8743);
			3247: out = 16'(8581);
			3248: out = 16'(7343);
			3249: out = 16'(-21775);
			3250: out = 16'(-8588);
			3251: out = 16'(4049);
			3252: out = 16'(18198);
			3253: out = 16'(12518);
			3254: out = 16'(4775);
			3255: out = 16'(-20794);
			3256: out = 16'(-14689);
			3257: out = 16'(6469);
			3258: out = 16'(17779);
			3259: out = 16'(13253);
			3260: out = 16'(-11827);
			3261: out = 16'(-3283);
			3262: out = 16'(184);
			3263: out = 16'(9261);
			3264: out = 16'(11883);
			3265: out = 16'(12944);
			3266: out = 16'(4302);
			3267: out = 16'(-2281);
			3268: out = 16'(-9856);
			3269: out = 16'(-1751);
			3270: out = 16'(-3098);
			3271: out = 16'(574);
			3272: out = 16'(14);
			3273: out = 16'(9957);
			3274: out = 16'(17246);
			3275: out = 16'(7100);
			3276: out = 16'(350);
			3277: out = 16'(-2513);
			3278: out = 16'(-10994);
			3279: out = 16'(-7952);
			3280: out = 16'(1514);
			3281: out = 16'(11356);
			3282: out = 16'(11675);
			3283: out = 16'(89);
			3284: out = 16'(-12387);
			3285: out = 16'(-19221);
			3286: out = 16'(1405);
			3287: out = 16'(2475);
			3288: out = 16'(6565);
			3289: out = 16'(16997);
			3290: out = 16'(11943);
			3291: out = 16'(728);
			3292: out = 16'(10592);
			3293: out = 16'(3606);
			3294: out = 16'(-3805);
			3295: out = 16'(-15217);
			3296: out = 16'(-11363);
			3297: out = 16'(6723);
			3298: out = 16'(5279);
			3299: out = 16'(3813);
			3300: out = 16'(-12398);
			3301: out = 16'(79);
			3302: out = 16'(4970);
			3303: out = 16'(14938);
			3304: out = 16'(-9010);
			3305: out = 16'(-25600);
			3306: out = 16'(-4137);
			3307: out = 16'(4981);
			3308: out = 16'(14204);
			3309: out = 16'(583);
			3310: out = 16'(-225);
			3311: out = 16'(-2573);
			3312: out = 16'(-6073);
			3313: out = 16'(-5621);
			3314: out = 16'(2611);
			3315: out = 16'(-952);
			3316: out = 16'(-930);
			3317: out = 16'(-10700);
			3318: out = 16'(9735);
			3319: out = 16'(13532);
			3320: out = 16'(4576);
			3321: out = 16'(-3235);
			3322: out = 16'(-9680);
			3323: out = 16'(-23561);
			3324: out = 16'(-11768);
			3325: out = 16'(1647);
			3326: out = 16'(13036);
			3327: out = 16'(8478);
			3328: out = 16'(278);
			3329: out = 16'(-21518);
			3330: out = 16'(-14331);
			3331: out = 16'(10256);
			3332: out = 16'(13324);
			3333: out = 16'(12707);
			3334: out = 16'(-1884);
			3335: out = 16'(-5671);
			3336: out = 16'(-10946);
			3337: out = 16'(-1912);
			3338: out = 16'(-14371);
			3339: out = 16'(-14195);
			3340: out = 16'(4601);
			3341: out = 16'(3406);
			3342: out = 16'(-461);
			3343: out = 16'(-6704);
			3344: out = 16'(-9211);
			3345: out = 16'(-7462);
			3346: out = 16'(4259);
			3347: out = 16'(10446);
			3348: out = 16'(12825);
			3349: out = 16'(2291);
			3350: out = 16'(-2695);
			3351: out = 16'(-2945);
			3352: out = 16'(-7540);
			3353: out = 16'(-6109);
			3354: out = 16'(-1994);
			3355: out = 16'(1592);
			3356: out = 16'(3594);
			3357: out = 16'(8563);
			3358: out = 16'(-2171);
			3359: out = 16'(-5395);
			3360: out = 16'(14877);
			3361: out = 16'(17732);
			3362: out = 16'(17743);
			3363: out = 16'(-2197);
			3364: out = 16'(-6946);
			3365: out = 16'(-9917);
			3366: out = 16'(4442);
			3367: out = 16'(-1336);
			3368: out = 16'(-17800);
			3369: out = 16'(3270);
			3370: out = 16'(8079);
			3371: out = 16'(8587);
			3372: out = 16'(2632);
			3373: out = 16'(-680);
			3374: out = 16'(-6122);
			3375: out = 16'(4597);
			3376: out = 16'(9316);
			3377: out = 16'(4311);
			3378: out = 16'(3724);
			3379: out = 16'(310);
			3380: out = 16'(-23480);
			3381: out = 16'(-19935);
			3382: out = 16'(-9827);
			3383: out = 16'(14099);
			3384: out = 16'(16086);
			3385: out = 16'(11626);
			3386: out = 16'(-12789);
			3387: out = 16'(-11997);
			3388: out = 16'(8345);
			3389: out = 16'(6731);
			3390: out = 16'(6128);
			3391: out = 16'(-6997);
			3392: out = 16'(-2453);
			3393: out = 16'(-1213);
			3394: out = 16'(11183);
			3395: out = 16'(-4953);
			3396: out = 16'(-11408);
			3397: out = 16'(6575);
			3398: out = 16'(12175);
			3399: out = 16'(15970);
			3400: out = 16'(-6372);
			3401: out = 16'(-1490);
			3402: out = 16'(6286);
			3403: out = 16'(8557);
			3404: out = 16'(6307);
			3405: out = 16'(651);
			3406: out = 16'(736);
			3407: out = 16'(-3893);
			3408: out = 16'(-14610);
			3409: out = 16'(-8932);
			3410: out = 16'(-2918);
			3411: out = 16'(18078);
			3412: out = 16'(-12158);
			3413: out = 16'(-25221);
			3414: out = 16'(-3099);
			3415: out = 16'(8524);
			3416: out = 16'(17428);
			3417: out = 16'(5583);
			3418: out = 16'(1524);
			3419: out = 16'(-5110);
			3420: out = 16'(5415);
			3421: out = 16'(2916);
			3422: out = 16'(-255);
			3423: out = 16'(266);
			3424: out = 16'(-266);
			3425: out = 16'(-1662);
			3426: out = 16'(-2403);
			3427: out = 16'(-4522);
			3428: out = 16'(-10534);
			3429: out = 16'(3066);
			3430: out = 16'(12259);
			3431: out = 16'(17141);
			3432: out = 16'(9850);
			3433: out = 16'(864);
			3434: out = 16'(-6423);
			3435: out = 16'(-4420);
			3436: out = 16'(1968);
			3437: out = 16'(-10139);
			3438: out = 16'(1577);
			3439: out = 16'(13401);
			3440: out = 16'(2503);
			3441: out = 16'(-9959);
			3442: out = 16'(-29254);
			3443: out = 16'(-5301);
			3444: out = 16'(8851);
			3445: out = 16'(21371);
			3446: out = 16'(4470);
			3447: out = 16'(-10890);
			3448: out = 16'(-30402);
			3449: out = 16'(-12545);
			3450: out = 16'(4963);
			3451: out = 16'(-1030);
			3452: out = 16'(3471);
			3453: out = 16'(615);
			3454: out = 16'(5947);
			3455: out = 16'(-14580);
			3456: out = 16'(-30113);
			3457: out = 16'(-8667);
			3458: out = 16'(12455);
			3459: out = 16'(27746);
			3460: out = 16'(11943);
			3461: out = 16'(-1814);
			3462: out = 16'(-20161);
			3463: out = 16'(-13763);
			3464: out = 16'(-7762);
			3465: out = 16'(-2076);
			3466: out = 16'(-1977);
			3467: out = 16'(-442);
			3468: out = 16'(20133);
			3469: out = 16'(-4611);
			3470: out = 16'(-17230);
			3471: out = 16'(7593);
			3472: out = 16'(14270);
			3473: out = 16'(16631);
			3474: out = 16'(12783);
			3475: out = 16'(1685);
			3476: out = 16'(-9025);
			3477: out = 16'(-25856);
			3478: out = 16'(-15148);
			3479: out = 16'(13464);
			3480: out = 16'(13611);
			3481: out = 16'(6769);
			3482: out = 16'(-18993);
			3483: out = 16'(-16045);
			3484: out = 16'(-12015);
			3485: out = 16'(3248);
			3486: out = 16'(8135);
			3487: out = 16'(12471);
			3488: out = 16'(13600);
			3489: out = 16'(4133);
			3490: out = 16'(-7355);
			3491: out = 16'(-12792);
			3492: out = 16'(-6615);
			3493: out = 16'(7827);
			3494: out = 16'(-5496);
			3495: out = 16'(4156);
			3496: out = 16'(15809);
			3497: out = 16'(10935);
			3498: out = 16'(-1094);
			3499: out = 16'(-27564);
			3500: out = 16'(-5295);
			3501: out = 16'(8280);
			3502: out = 16'(20489);
			3503: out = 16'(6672);
			3504: out = 16'(-3080);
			3505: out = 16'(-6096);
			3506: out = 16'(-623);
			3507: out = 16'(6112);
			3508: out = 16'(1168);
			3509: out = 16'(3327);
			3510: out = 16'(3149);
			3511: out = 16'(2027);
			3512: out = 16'(6081);
			3513: out = 16'(14842);
			3514: out = 16'(-2287);
			3515: out = 16'(-2959);
			3516: out = 16'(-1770);
			3517: out = 16'(11845);
			3518: out = 16'(10229);
			3519: out = 16'(-3603);
			3520: out = 16'(-8810);
			3521: out = 16'(-12253);
			3522: out = 16'(-8326);
			3523: out = 16'(-8996);
			3524: out = 16'(-5294);
			3525: out = 16'(13972);
			3526: out = 16'(6599);
			3527: out = 16'(-1002);
			3528: out = 16'(-6957);
			3529: out = 16'(4057);
			3530: out = 16'(19533);
			3531: out = 16'(10393);
			3532: out = 16'(4062);
			3533: out = 16'(-11146);
			3534: out = 16'(2997);
			3535: out = 16'(2403);
			3536: out = 16'(1926);
			3537: out = 16'(-9258);
			3538: out = 16'(-10233);
			3539: out = 16'(-4862);
			3540: out = 16'(7139);
			3541: out = 16'(12051);
			3542: out = 16'(5631);
			3543: out = 16'(-2643);
			3544: out = 16'(-7839);
			3545: out = 16'(11633);
			3546: out = 16'(13908);
			3547: out = 16'(14636);
			3548: out = 16'(-12493);
			3549: out = 16'(-14659);
			3550: out = 16'(-9762);
			3551: out = 16'(-2002);
			3552: out = 16'(-2091);
			3553: out = 16'(-11399);
			3554: out = 16'(6096);
			3555: out = 16'(10961);
			3556: out = 16'(11178);
			3557: out = 16'(2624);
			3558: out = 16'(-6476);
			3559: out = 16'(-23586);
			3560: out = 16'(-13500);
			3561: out = 16'(-1262);
			3562: out = 16'(14034);
			3563: out = 16'(8330);
			3564: out = 16'(-1793);
			3565: out = 16'(-17689);
			3566: out = 16'(-14723);
			3567: out = 16'(-960);
			3568: out = 16'(-546);
			3569: out = 16'(6488);
			3570: out = 16'(7439);
			3571: out = 16'(16271);
			3572: out = 16'(7874);
			3573: out = 16'(-9132);
			3574: out = 16'(-14870);
			3575: out = 16'(-11538);
			3576: out = 16'(9381);
			3577: out = 16'(3714);
			3578: out = 16'(-41);
			3579: out = 16'(-8450);
			3580: out = 16'(-4419);
			3581: out = 16'(757);
			3582: out = 16'(6418);
			3583: out = 16'(7677);
			3584: out = 16'(6531);
			3585: out = 16'(6402);
			3586: out = 16'(3442);
			3587: out = 16'(1082);
			3588: out = 16'(-8697);
			3589: out = 16'(-5816);
			3590: out = 16'(5427);
			3591: out = 16'(1259);
			3592: out = 16'(-3734);
			3593: out = 16'(-19514);
			3594: out = 16'(-5313);
			3595: out = 16'(2618);
			3596: out = 16'(7568);
			3597: out = 16'(-2802);
			3598: out = 16'(-8138);
			3599: out = 16'(13355);
			3600: out = 16'(11477);
			3601: out = 16'(9881);
			3602: out = 16'(-18348);
			3603: out = 16'(-13880);
			3604: out = 16'(-3713);
			3605: out = 16'(9874);
			3606: out = 16'(8532);
			3607: out = 16'(1253);
			3608: out = 16'(-12466);
			3609: out = 16'(-12979);
			3610: out = 16'(543);
			3611: out = 16'(9688);
			3612: out = 16'(11389);
			3613: out = 16'(-8539);
			3614: out = 16'(1153);
			3615: out = 16'(4153);
			3616: out = 16'(10415);
			3617: out = 16'(3020);
			3618: out = 16'(-1680);
			3619: out = 16'(-2609);
			3620: out = 16'(-2341);
			3621: out = 16'(-2082);
			3622: out = 16'(8862);
			3623: out = 16'(5573);
			3624: out = 16'(-548);
			3625: out = 16'(-9892);
			3626: out = 16'(-4634);
			3627: out = 16'(13452);
			3628: out = 16'(9016);
			3629: out = 16'(4798);
			3630: out = 16'(-15402);
			3631: out = 16'(-3954);
			3632: out = 16'(271);
			3633: out = 16'(13450);
			3634: out = 16'(-4424);
			3635: out = 16'(-14729);
			3636: out = 16'(-25927);
			3637: out = 16'(-1593);
			3638: out = 16'(21582);
			3639: out = 16'(16722);
			3640: out = 16'(5547);
			3641: out = 16'(-13896);
			3642: out = 16'(-1907);
			3643: out = 16'(5739);
			3644: out = 16'(22104);
			3645: out = 16'(-3907);
			3646: out = 16'(-9250);
			3647: out = 16'(-8997);
			3648: out = 16'(-1985);
			3649: out = 16'(973);
			3650: out = 16'(473);
			3651: out = 16'(2248);
			3652: out = 16'(2205);
			3653: out = 16'(-7413);
			3654: out = 16'(-518);
			3655: out = 16'(6684);
			3656: out = 16'(17699);
			3657: out = 16'(8771);
			3658: out = 16'(-5173);
			3659: out = 16'(1950);
			3660: out = 16'(-7);
			3661: out = 16'(2115);
			3662: out = 16'(-15746);
			3663: out = 16'(-15407);
			3664: out = 16'(-6544);
			3665: out = 16'(7452);
			3666: out = 16'(13831);
			3667: out = 16'(11801);
			3668: out = 16'(5002);
			3669: out = 16'(-3755);
			3670: out = 16'(-14650);
			3671: out = 16'(-6658);
			3672: out = 16'(3720);
			3673: out = 16'(1562);
			3674: out = 16'(2969);
			3675: out = 16'(-996);
			3676: out = 16'(12381);
			3677: out = 16'(1576);
			3678: out = 16'(-9415);
			3679: out = 16'(-18190);
			3680: out = 16'(-7358);
			3681: out = 16'(15517);
			3682: out = 16'(6775);
			3683: out = 16'(4599);
			3684: out = 16'(3073);
			3685: out = 16'(-6253);
			3686: out = 16'(-9870);
			3687: out = 16'(-3991);
			3688: out = 16'(953);
			3689: out = 16'(4881);
			3690: out = 16'(1136);
			3691: out = 16'(1082);
			3692: out = 16'(114);
			3693: out = 16'(-1549);
			3694: out = 16'(2341);
			3695: out = 16'(6882);
			3696: out = 16'(1120);
			3697: out = 16'(-2742);
			3698: out = 16'(-7596);
			3699: out = 16'(-1582);
			3700: out = 16'(982);
			3701: out = 16'(1446);
			3702: out = 16'(2025);
			3703: out = 16'(1960);
			3704: out = 16'(6330);
			3705: out = 16'(-3308);
			3706: out = 16'(-10344);
			3707: out = 16'(-27737);
			3708: out = 16'(-5451);
			3709: out = 16'(14289);
			3710: out = 16'(13482);
			3711: out = 16'(11953);
			3712: out = 16'(4205);
			3713: out = 16'(-4634);
			3714: out = 16'(-9698);
			3715: out = 16'(-8818);
			3716: out = 16'(3494);
			3717: out = 16'(8249);
			3718: out = 16'(5659);
			3719: out = 16'(-377);
			3720: out = 16'(-7885);
			3721: out = 16'(-10590);
			3722: out = 16'(-14095);
			3723: out = 16'(-7638);
			3724: out = 16'(7799);
			3725: out = 16'(15265);
			3726: out = 16'(14443);
			3727: out = 16'(-7617);
			3728: out = 16'(-12044);
			3729: out = 16'(-13267);
			3730: out = 16'(7143);
			3731: out = 16'(7376);
			3732: out = 16'(5066);
			3733: out = 16'(-9246);
			3734: out = 16'(-7822);
			3735: out = 16'(1720);
			3736: out = 16'(-364);
			3737: out = 16'(1626);
			3738: out = 16'(1869);
			3739: out = 16'(210);
			3740: out = 16'(908);
			3741: out = 16'(11933);
			3742: out = 16'(1131);
			3743: out = 16'(-3706);
			3744: out = 16'(-10784);
			3745: out = 16'(1873);
			3746: out = 16'(10037);
			3747: out = 16'(7652);
			3748: out = 16'(-3511);
			3749: out = 16'(-15486);
			3750: out = 16'(-1213);
			3751: out = 16'(8250);
			3752: out = 16'(20504);
			3753: out = 16'(951);
			3754: out = 16'(-3170);
			3755: out = 16'(-7940);
			3756: out = 16'(7778);
			3757: out = 16'(10484);
			3758: out = 16'(6314);
			3759: out = 16'(2291);
			3760: out = 16'(-2457);
			3761: out = 16'(-10484);
			3762: out = 16'(-9614);
			3763: out = 16'(-6044);
			3764: out = 16'(12645);
			3765: out = 16'(7382);
			3766: out = 16'(2820);
			3767: out = 16'(-16744);
			3768: out = 16'(-364);
			3769: out = 16'(21092);
			3770: out = 16'(13793);
			3771: out = 16'(-790);
			3772: out = 16'(-30979);
			3773: out = 16'(-4914);
			3774: out = 16'(3513);
			3775: out = 16'(13798);
			3776: out = 16'(177);
			3777: out = 16'(-6712);
			3778: out = 16'(-25406);
			3779: out = 16'(5808);
			3780: out = 16'(19182);
			3781: out = 16'(8028);
			3782: out = 16'(-8920);
			3783: out = 16'(-22337);
			3784: out = 16'(14795);
			3785: out = 16'(8409);
			3786: out = 16'(3348);
			3787: out = 16'(-12527);
			3788: out = 16'(-5918);
			3789: out = 16'(6848);
			3790: out = 16'(1809);
			3791: out = 16'(-317);
			3792: out = 16'(-6613);
			3793: out = 16'(266);
			3794: out = 16'(1114);
			3795: out = 16'(1789);
			3796: out = 16'(-2075);
			3797: out = 16'(-1722);
			3798: out = 16'(880);
			3799: out = 16'(4445);
			3800: out = 16'(5511);
			3801: out = 16'(8642);
			3802: out = 16'(141);
			3803: out = 16'(-7463);
			3804: out = 16'(-16378);
			3805: out = 16'(-9024);
			3806: out = 16'(2981);
			3807: out = 16'(-1629);
			3808: out = 16'(1598);
			3809: out = 16'(6206);
			3810: out = 16'(-4996);
			3811: out = 16'(-4934);
			3812: out = 16'(288);
			3813: out = 16'(13173);
			3814: out = 16'(10868);
			3815: out = 16'(-14279);
			3816: out = 16'(-17302);
			3817: out = 16'(-15130);
			3818: out = 16'(18421);
			3819: out = 16'(8054);
			3820: out = 16'(2276);
			3821: out = 16'(-8844);
			3822: out = 16'(-427);
			3823: out = 16'(8312);
			3824: out = 16'(13202);
			3825: out = 16'(10202);
			3826: out = 16'(4559);
			3827: out = 16'(-1513);
			3828: out = 16'(-4267);
			3829: out = 16'(-6194);
			3830: out = 16'(6051);
			3831: out = 16'(6897);
			3832: out = 16'(-567);
			3833: out = 16'(-7297);
			3834: out = 16'(-8974);
			3835: out = 16'(379);
			3836: out = 16'(4840);
			3837: out = 16'(7351);
			3838: out = 16'(-50);
			3839: out = 16'(-4679);
			3840: out = 16'(-8932);
			3841: out = 16'(650);
			3842: out = 16'(3577);
			3843: out = 16'(6944);
			3844: out = 16'(-860);
			3845: out = 16'(-729);
			3846: out = 16'(1060);
			3847: out = 16'(-6935);
			3848: out = 16'(-7838);
			3849: out = 16'(-2066);
			3850: out = 16'(853);
			3851: out = 16'(3573);
			3852: out = 16'(-583);
			3853: out = 16'(3725);
			3854: out = 16'(4581);
			3855: out = 16'(11126);
			3856: out = 16'(1132);
			3857: out = 16'(-6020);
			3858: out = 16'(-15391);
			3859: out = 16'(-5827);
			3860: out = 16'(6148);
			3861: out = 16'(8325);
			3862: out = 16'(6268);
			3863: out = 16'(27);
			3864: out = 16'(-5794);
			3865: out = 16'(-4764);
			3866: out = 16'(3998);
			3867: out = 16'(4245);
			3868: out = 16'(3920);
			3869: out = 16'(-3991);
			3870: out = 16'(-2452);
			3871: out = 16'(-1607);
			3872: out = 16'(8791);
			3873: out = 16'(3086);
			3874: out = 16'(-1184);
			3875: out = 16'(-20625);
			3876: out = 16'(-8629);
			3877: out = 16'(3700);
			3878: out = 16'(9219);
			3879: out = 16'(-3737);
			3880: out = 16'(-24579);
			3881: out = 16'(1832);
			3882: out = 16'(9457);
			3883: out = 16'(19549);
			3884: out = 16'(-12391);
			3885: out = 16'(-21508);
			3886: out = 16'(-21518);
			3887: out = 16'(1447);
			3888: out = 16'(14098);
			3889: out = 16'(13242);
			3890: out = 16'(9039);
			3891: out = 16'(2033);
			3892: out = 16'(-3064);
			3893: out = 16'(-5);
			3894: out = 16'(5648);
			3895: out = 16'(-776);
			3896: out = 16'(3165);
			3897: out = 16'(4202);
			3898: out = 16'(10616);
			3899: out = 16'(4036);
			3900: out = 16'(-4926);
			3901: out = 16'(-420);
			3902: out = 16'(-1544);
			3903: out = 16'(-8189);
			3904: out = 16'(2215);
			3905: out = 16'(5021);
			3906: out = 16'(10457);
			3907: out = 16'(-12343);
			3908: out = 16'(-18710);
			3909: out = 16'(6031);
			3910: out = 16'(12481);
			3911: out = 16'(16028);
			3912: out = 16'(-5812);
			3913: out = 16'(-6789);
			3914: out = 16'(-8791);
			3915: out = 16'(5228);
			3916: out = 16'(3165);
			3917: out = 16'(1389);
			3918: out = 16'(-4150);
			3919: out = 16'(-2791);
			3920: out = 16'(-1823);
			3921: out = 16'(6812);
			3922: out = 16'(5366);
			3923: out = 16'(617);
			3924: out = 16'(-11056);
			3925: out = 16'(-11688);
			3926: out = 16'(4751);
			3927: out = 16'(7851);
			3928: out = 16'(10496);
			3929: out = 16'(8930);
			3930: out = 16'(4900);
			3931: out = 16'(-685);
			3932: out = 16'(-12746);
			3933: out = 16'(-6784);
			3934: out = 16'(5075);
			3935: out = 16'(9252);
			3936: out = 16'(7975);
			3937: out = 16'(-1940);
			3938: out = 16'(4610);
			3939: out = 16'(1268);
			3940: out = 16'(696);
			3941: out = 16'(-15976);
			3942: out = 16'(-16481);
			3943: out = 16'(2060);
			3944: out = 16'(997);
			3945: out = 16'(2096);
			3946: out = 16'(1357);
			3947: out = 16'(-607);
			3948: out = 16'(-2890);
			3949: out = 16'(4675);
			3950: out = 16'(2134);
			3951: out = 16'(415);
			3952: out = 16'(-15781);
			3953: out = 16'(-8742);
			3954: out = 16'(4852);
			3955: out = 16'(8943);
			3956: out = 16'(3581);
			3957: out = 16'(-15797);
			3958: out = 16'(-1285);
			3959: out = 16'(1549);
			3960: out = 16'(9885);
			3961: out = 16'(-13700);
			3962: out = 16'(-16787);
			3963: out = 16'(7256);
			3964: out = 16'(13181);
			3965: out = 16'(12865);
			3966: out = 16'(-15889);
			3967: out = 16'(-12409);
			3968: out = 16'(-6105);
			3969: out = 16'(5548);
			3970: out = 16'(8331);
			3971: out = 16'(7537);
			3972: out = 16'(7903);
			3973: out = 16'(217);
			3974: out = 16'(-10783);
			3975: out = 16'(-3826);
			3976: out = 16'(-3079);
			3977: out = 16'(-5693);
			3978: out = 16'(1348);
			3979: out = 16'(3865);
			3980: out = 16'(4789);
			3981: out = 16'(-1018);
			3982: out = 16'(-4803);
			3983: out = 16'(-6843);
			3984: out = 16'(-1965);
			3985: out = 16'(3119);
			3986: out = 16'(6635);
			3987: out = 16'(7701);
			3988: out = 16'(6713);
			3989: out = 16'(-12622);
			3990: out = 16'(-11264);
			3991: out = 16'(-3847);
			3992: out = 16'(9108);
			3993: out = 16'(7660);
			3994: out = 16'(-3840);
			3995: out = 16'(-4084);
			3996: out = 16'(-3336);
			3997: out = 16'(5694);
			3998: out = 16'(4005);
			3999: out = 16'(2573);
			4000: out = 16'(-10797);
			4001: out = 16'(-2134);
			4002: out = 16'(4133);
			4003: out = 16'(17062);
			4004: out = 16'(8777);
			4005: out = 16'(1401);
			4006: out = 16'(-6705);
			4007: out = 16'(-2020);
			4008: out = 16'(5032);
			4009: out = 16'(5397);
			4010: out = 16'(-733);
			4011: out = 16'(-12808);
			4012: out = 16'(-3095);
			4013: out = 16'(2336);
			4014: out = 16'(10824);
			4015: out = 16'(8385);
			4016: out = 16'(369);
			4017: out = 16'(-29659);
			4018: out = 16'(-10816);
			4019: out = 16'(2146);
			4020: out = 16'(21599);
			4021: out = 16'(-2544);
			4022: out = 16'(-18419);
			4023: out = 16'(-3139);
			4024: out = 16'(9020);
			4025: out = 16'(19886);
			4026: out = 16'(-6497);
			4027: out = 16'(-13522);
			4028: out = 16'(-21228);
			4029: out = 16'(12775);
			4030: out = 16'(18039);
			4031: out = 16'(15781);
			4032: out = 16'(-3579);
			4033: out = 16'(-12374);
			4034: out = 16'(-10481);
			4035: out = 16'(-10617);
			4036: out = 16'(-2543);
			4037: out = 16'(13681);
			4038: out = 16'(11808);
			4039: out = 16'(8374);
			4040: out = 16'(2297);
			4041: out = 16'(-2460);
			4042: out = 16'(-5417);
			4043: out = 16'(4146);
			4044: out = 16'(2061);
			4045: out = 16'(222);
			4046: out = 16'(-4419);
			4047: out = 16'(2688);
			4048: out = 16'(14054);
			4049: out = 16'(3268);
			4050: out = 16'(-2618);
			4051: out = 16'(-12809);
			4052: out = 16'(-328);
			4053: out = 16'(2218);
			4054: out = 16'(-1550);
			4055: out = 16'(-8103);
			4056: out = 16'(-9038);
			4057: out = 16'(9049);
			4058: out = 16'(3180);
			4059: out = 16'(1768);
			4060: out = 16'(-1096);
			4061: out = 16'(8177);
			4062: out = 16'(13225);
			4063: out = 16'(1745);
			4064: out = 16'(-7202);
			4065: out = 16'(-14869);
			4066: out = 16'(-4404);
			4067: out = 16'(4895);
			4068: out = 16'(13327);
			4069: out = 16'(15460);
			4070: out = 16'(7026);
			4071: out = 16'(-14677);
			4072: out = 16'(-12445);
			4073: out = 16'(-8228);
			4074: out = 16'(7098);
			4075: out = 16'(4576);
			4076: out = 16'(3776);
			4077: out = 16'(851);
			4078: out = 16'(1204);
			4079: out = 16'(157);
			4080: out = 16'(-3817);
			4081: out = 16'(-5455);
			4082: out = 16'(-5395);
			4083: out = 16'(-2499);
			4084: out = 16'(2321);
			4085: out = 16'(8130);
			4086: out = 16'(2414);
			4087: out = 16'(-3801);
			4088: out = 16'(-17872);
			4089: out = 16'(2287);
			4090: out = 16'(8131);
			4091: out = 16'(6974);
			4092: out = 16'(-9400);
			4093: out = 16'(-17008);
			4094: out = 16'(1458);
			4095: out = 16'(418);
			4096: out = 16'(2958);
			4097: out = 16'(1006);
			4098: out = 16'(3376);
			4099: out = 16'(2030);
			4100: out = 16'(186);
			4101: out = 16'(-4057);
			4102: out = 16'(-4763);
			4103: out = 16'(-10436);
			4104: out = 16'(-751);
			4105: out = 16'(15606);
			4106: out = 16'(9393);
			4107: out = 16'(5339);
			4108: out = 16'(-47);
			4109: out = 16'(-7098);
			4110: out = 16'(-8389);
			4111: out = 16'(1665);
			4112: out = 16'(5146);
			4113: out = 16'(6810);
			4114: out = 16'(-7479);
			4115: out = 16'(-1996);
			4116: out = 16'(2101);
			4117: out = 16'(1617);
			4118: out = 16'(2768);
			4119: out = 16'(4034);
			4120: out = 16'(-4506);
			4121: out = 16'(-5721);
			4122: out = 16'(-5509);
			4123: out = 16'(1737);
			4124: out = 16'(566);
			4125: out = 16'(-7428);
			4126: out = 16'(-4801);
			4127: out = 16'(189);
			4128: out = 16'(14339);
			4129: out = 16'(7986);
			4130: out = 16'(2617);
			4131: out = 16'(-11546);
			4132: out = 16'(-8134);
			4133: out = 16'(-2707);
			4134: out = 16'(15905);
			4135: out = 16'(11398);
			4136: out = 16'(4705);
			4137: out = 16'(-12719);
			4138: out = 16'(-9661);
			4139: out = 16'(1833);
			4140: out = 16'(11667);
			4141: out = 16'(8922);
			4142: out = 16'(-8060);
			4143: out = 16'(-1423);
			4144: out = 16'(99);
			4145: out = 16'(11725);
			4146: out = 16'(-5251);
			4147: out = 16'(-9120);
			4148: out = 16'(-3605);
			4149: out = 16'(3356);
			4150: out = 16'(7076);
			4151: out = 16'(11690);
			4152: out = 16'(-502);
			4153: out = 16'(-11907);
			4154: out = 16'(-13408);
			4155: out = 16'(-3840);
			4156: out = 16'(10810);
			4157: out = 16'(2727);
			4158: out = 16'(123);
			4159: out = 16'(-8520);
			4160: out = 16'(3899);
			4161: out = 16'(4876);
			4162: out = 16'(5968);
			4163: out = 16'(-5542);
			4164: out = 16'(-6142);
			4165: out = 16'(5737);
			4166: out = 16'(3565);
			4167: out = 16'(1908);
			4168: out = 16'(-1457);
			4169: out = 16'(-921);
			4170: out = 16'(628);
			4171: out = 16'(-634);
			4172: out = 16'(5144);
			4173: out = 16'(10016);
			4174: out = 16'(9661);
			4175: out = 16'(5315);
			4176: out = 16'(-1675);
			4177: out = 16'(-507);
			4178: out = 16'(-941);
			4179: out = 16'(-228);
			4180: out = 16'(4344);
			4181: out = 16'(3410);
			4182: out = 16'(-7549);
			4183: out = 16'(-13);
			4184: out = 16'(2974);
			4185: out = 16'(7636);
			4186: out = 16'(-3839);
			4187: out = 16'(-10945);
			4188: out = 16'(-86);
			4189: out = 16'(-229);
			4190: out = 16'(411);
			4191: out = 16'(-14749);
			4192: out = 16'(-10727);
			4193: out = 16'(-3129);
			4194: out = 16'(7726);
			4195: out = 16'(8145);
			4196: out = 16'(2852);
			4197: out = 16'(-6865);
			4198: out = 16'(-9088);
			4199: out = 16'(1282);
			4200: out = 16'(-5643);
			4201: out = 16'(-3283);
			4202: out = 16'(624);
			4203: out = 16'(10716);
			4204: out = 16'(9854);
			4205: out = 16'(-14348);
			4206: out = 16'(-15578);
			4207: out = 16'(-11406);
			4208: out = 16'(12652);
			4209: out = 16'(11915);
			4210: out = 16'(5546);
			4211: out = 16'(-5806);
			4212: out = 16'(-9778);
			4213: out = 16'(-5664);
			4214: out = 16'(-11239);
			4215: out = 16'(-3027);
			4216: out = 16'(6763);
			4217: out = 16'(18885);
			4218: out = 16'(13007);
			4219: out = 16'(-9167);
			4220: out = 16'(-22420);
			4221: out = 16'(-23324);
			4222: out = 16'(12419);
			4223: out = 16'(10018);
			4224: out = 16'(7730);
			4225: out = 16'(-19705);
			4226: out = 16'(-8265);
			4227: out = 16'(4005);
			4228: out = 16'(9199);
			4229: out = 16'(-1922);
			4230: out = 16'(-20995);
			4231: out = 16'(9032);
			4232: out = 16'(10777);
			4233: out = 16'(10805);
			4234: out = 16'(-13495);
			4235: out = 16'(-18411);
			4236: out = 16'(-12260);
			4237: out = 16'(8231);
			4238: out = 16'(16563);
			4239: out = 16'(10140);
			4240: out = 16'(-4309);
			4241: out = 16'(-13263);
			4242: out = 16'(12270);
			4243: out = 16'(5006);
			4244: out = 16'(2775);
			4245: out = 16'(-15017);
			4246: out = 16'(-808);
			4247: out = 16'(13951);
			4248: out = 16'(7396);
			4249: out = 16'(3356);
			4250: out = 16'(-3346);
			4251: out = 16'(-28);
			4252: out = 16'(606);
			4253: out = 16'(2125);
			4254: out = 16'(4549);
			4255: out = 16'(4337);
			4256: out = 16'(-2104);
			4257: out = 16'(986);
			4258: out = 16'(613);
			4259: out = 16'(555);
			4260: out = 16'(-5539);
			4261: out = 16'(-7621);
			4262: out = 16'(-154);
			4263: out = 16'(7853);
			4264: out = 16'(13896);
			4265: out = 16'(-5840);
			4266: out = 16'(-9367);
			4267: out = 16'(-12846);
			4268: out = 16'(13579);
			4269: out = 16'(11274);
			4270: out = 16'(684);
			4271: out = 16'(-9970);
			4272: out = 16'(-8919);
			4273: out = 16'(7099);
			4274: out = 16'(4602);
			4275: out = 16'(5386);
			4276: out = 16'(381);
			4277: out = 16'(3872);
			4278: out = 16'(1840);
			4279: out = 16'(-8359);
			4280: out = 16'(-3593);
			4281: out = 16'(2989);
			4282: out = 16'(-1187);
			4283: out = 16'(2910);
			4284: out = 16'(4151);
			4285: out = 16'(14155);
			4286: out = 16'(7696);
			4287: out = 16'(-1314);
			4288: out = 16'(-8981);
			4289: out = 16'(-6716);
			4290: out = 16'(3488);
			4291: out = 16'(2184);
			4292: out = 16'(3808);
			4293: out = 16'(7753);
			4294: out = 16'(977);
			4295: out = 16'(-4666);
			4296: out = 16'(-17645);
			4297: out = 16'(-2189);
			4298: out = 16'(8722);
			4299: out = 16'(3764);
			4300: out = 16'(-1417);
			4301: out = 16'(-8598);
			4302: out = 16'(-7017);
			4303: out = 16'(-3923);
			4304: out = 16'(2958);
			4305: out = 16'(2903);
			4306: out = 16'(7154);
			4307: out = 16'(10641);
			4308: out = 16'(334);
			4309: out = 16'(-7542);
			4310: out = 16'(-17128);
			4311: out = 16'(-404);
			4312: out = 16'(8529);
			4313: out = 16'(6881);
			4314: out = 16'(3487);
			4315: out = 16'(-2205);
			4316: out = 16'(-2024);
			4317: out = 16'(-5534);
			4318: out = 16'(-4731);
			4319: out = 16'(-1146);
			4320: out = 16'(1490);
			4321: out = 16'(1048);
			4322: out = 16'(1131);
			4323: out = 16'(-516);
			4324: out = 16'(900);
			4325: out = 16'(-10351);
			4326: out = 16'(-7452);
			4327: out = 16'(772);
			4328: out = 16'(9079);
			4329: out = 16'(8392);
			4330: out = 16'(-1691);
			4331: out = 16'(-4232);
			4332: out = 16'(-5826);
			4333: out = 16'(-7563);
			4334: out = 16'(2970);
			4335: out = 16'(9730);
			4336: out = 16'(8365);
			4337: out = 16'(-3924);
			4338: out = 16'(-17340);
			4339: out = 16'(-562);
			4340: out = 16'(1168);
			4341: out = 16'(3824);
			4342: out = 16'(2932);
			4343: out = 16'(-127);
			4344: out = 16'(-9447);
			4345: out = 16'(7086);
			4346: out = 16'(8533);
			4347: out = 16'(2713);
			4348: out = 16'(-1865);
			4349: out = 16'(-2961);
			4350: out = 16'(6346);
			4351: out = 16'(-1002);
			4352: out = 16'(-4625);
			4353: out = 16'(-5867);
			4354: out = 16'(1112);
			4355: out = 16'(7261);
			4356: out = 16'(-283);
			4357: out = 16'(2847);
			4358: out = 16'(4775);
			4359: out = 16'(-5293);
			4360: out = 16'(-7328);
			4361: out = 16'(-4665);
			4362: out = 16'(-3242);
			4363: out = 16'(5326);
			4364: out = 16'(17750);
			4365: out = 16'(6819);
			4366: out = 16'(-1800);
			4367: out = 16'(-13347);
			4368: out = 16'(-6966);
			4369: out = 16'(-1911);
			4370: out = 16'(-6712);
			4371: out = 16'(4233);
			4372: out = 16'(10650);
			4373: out = 16'(9166);
			4374: out = 16'(1947);
			4375: out = 16'(-7103);
			4376: out = 16'(-2511);
			4377: out = 16'(-1307);
			4378: out = 16'(4123);
			4379: out = 16'(-2209);
			4380: out = 16'(3274);
			4381: out = 16'(9473);
			4382: out = 16'(10867);
			4383: out = 16'(1140);
			4384: out = 16'(-22625);
			4385: out = 16'(-11670);
			4386: out = 16'(-990);
			4387: out = 16'(7908);
			4388: out = 16'(12562);
			4389: out = 16'(11094);
			4390: out = 16'(7945);
			4391: out = 16'(-8083);
			4392: out = 16'(-20747);
			4393: out = 16'(-8556);
			4394: out = 16'(-375);
			4395: out = 16'(8728);
			4396: out = 16'(1668);
			4397: out = 16'(274);
			4398: out = 16'(-1738);
			4399: out = 16'(-57);
			4400: out = 16'(26);
			4401: out = 16'(-1873);
			4402: out = 16'(6392);
			4403: out = 16'(7698);
			4404: out = 16'(2471);
			4405: out = 16'(1367);
			4406: out = 16'(999);
			4407: out = 16'(697);
			4408: out = 16'(3761);
			4409: out = 16'(4139);
			4410: out = 16'(4879);
			4411: out = 16'(-6805);
			4412: out = 16'(-17698);
			4413: out = 16'(-13443);
			4414: out = 16'(-279);
			4415: out = 16'(17923);
			4416: out = 16'(8128);
			4417: out = 16'(3896);
			4418: out = 16'(-6016);
			4419: out = 16'(-5211);
			4420: out = 16'(-3940);
			4421: out = 16'(7755);
			4422: out = 16'(1371);
			4423: out = 16'(-244);
			4424: out = 16'(-12164);
			4425: out = 16'(3002);
			4426: out = 16'(9015);
			4427: out = 16'(4891);
			4428: out = 16'(-5831);
			4429: out = 16'(-14101);
			4430: out = 16'(-11263);
			4431: out = 16'(-3413);
			4432: out = 16'(5070);
			4433: out = 16'(9545);
			4434: out = 16'(6311);
			4435: out = 16'(459);
			4436: out = 16'(-17297);
			4437: out = 16'(-18832);
			4438: out = 16'(-5971);
			4439: out = 16'(4351);
			4440: out = 16'(10563);
			4441: out = 16'(8651);
			4442: out = 16'(4758);
			4443: out = 16'(-1608);
			4444: out = 16'(-16678);
			4445: out = 16'(-4162);
			4446: out = 16'(8355);
			4447: out = 16'(14843);
			4448: out = 16'(7493);
			4449: out = 16'(-4018);
			4450: out = 16'(-13082);
			4451: out = 16'(-11048);
			4452: out = 16'(-800);
			4453: out = 16'(8636);
			4454: out = 16'(6636);
			4455: out = 16'(-9117);
			4456: out = 16'(-496);
			4457: out = 16'(505);
			4458: out = 16'(5330);
			4459: out = 16'(-329);
			4460: out = 16'(-836);
			4461: out = 16'(-526);
			4462: out = 16'(1572);
			4463: out = 16'(612);
			4464: out = 16'(-3661);
			4465: out = 16'(-2239);
			4466: out = 16'(863);
			4467: out = 16'(-5650);
			4468: out = 16'(-7839);
			4469: out = 16'(-13090);
			4470: out = 16'(13942);
			4471: out = 16'(10250);
			4472: out = 16'(3153);
			4473: out = 16'(-19906);
			4474: out = 16'(-14444);
			4475: out = 16'(13487);
			4476: out = 16'(17759);
			4477: out = 16'(14415);
			4478: out = 16'(-7923);
			4479: out = 16'(-14850);
			4480: out = 16'(-16345);
			4481: out = 16'(11192);
			4482: out = 16'(12402);
			4483: out = 16'(13980);
			4484: out = 16'(-15135);
			4485: out = 16'(-1852);
			4486: out = 16'(11263);
			4487: out = 16'(10319);
			4488: out = 16'(284);
			4489: out = 16'(-16285);
			4490: out = 16'(6880);
			4491: out = 16'(12291);
			4492: out = 16'(17536);
			4493: out = 16'(-10312);
			4494: out = 16'(-19973);
			4495: out = 16'(-16016);
			4496: out = 16'(-5090);
			4497: out = 16'(4411);
			4498: out = 16'(4454);
			4499: out = 16'(10785);
			4500: out = 16'(9852);
			4501: out = 16'(-3719);
			4502: out = 16'(-4461);
			4503: out = 16'(-3840);
			4504: out = 16'(1681);
			4505: out = 16'(-2744);
			4506: out = 16'(-8963);
			4507: out = 16'(-1863);
			4508: out = 16'(-1052);
			4509: out = 16'(-947);
			4510: out = 16'(3502);
			4511: out = 16'(3649);
			4512: out = 16'(223);
			4513: out = 16'(-594);
			4514: out = 16'(1157);
			4515: out = 16'(12312);
			4516: out = 16'(1467);
			4517: out = 16'(-2882);
			4518: out = 16'(-251);
			4519: out = 16'(4441);
			4520: out = 16'(6929);
			4521: out = 16'(-5589);
			4522: out = 16'(-2726);
			4523: out = 16'(316);
			4524: out = 16'(-2308);
			4525: out = 16'(-7445);
			4526: out = 16'(-14836);
			4527: out = 16'(5620);
			4528: out = 16'(11132);
			4529: out = 16'(13280);
			4530: out = 16'(-1056);
			4531: out = 16'(-8463);
			4532: out = 16'(-13239);
			4533: out = 16'(-1345);
			4534: out = 16'(5812);
			4535: out = 16'(3654);
			4536: out = 16'(3379);
			4537: out = 16'(-2294);
			4538: out = 16'(-21285);
			4539: out = 16'(-16220);
			4540: out = 16'(-4494);
			4541: out = 16'(5952);
			4542: out = 16'(10009);
			4543: out = 16'(7113);
			4544: out = 16'(9739);
			4545: out = 16'(2285);
			4546: out = 16'(-5474);
			4547: out = 16'(-9342);
			4548: out = 16'(-6081);
			4549: out = 16'(2521);
			4550: out = 16'(1219);
			4551: out = 16'(1768);
			4552: out = 16'(8086);
			4553: out = 16'(-5048);
			4554: out = 16'(-10144);
			4555: out = 16'(153);
			4556: out = 16'(9523);
			4557: out = 16'(17060);
			4558: out = 16'(3682);
			4559: out = 16'(9384);
			4560: out = 16'(11703);
			4561: out = 16'(-4356);
			4562: out = 16'(-12981);
			4563: out = 16'(-19524);
			4564: out = 16'(4907);
			4565: out = 16'(8955);
			4566: out = 16'(-220);
			4567: out = 16'(3950);
			4568: out = 16'(1365);
			4569: out = 16'(3052);
			4570: out = 16'(-15554);
			4571: out = 16'(-16958);
			4572: out = 16'(15327);
			4573: out = 16'(14374);
			4574: out = 16'(12314);
			4575: out = 16'(-16221);
			4576: out = 16'(-11949);
			4577: out = 16'(-6898);
			4578: out = 16'(16328);
			4579: out = 16'(1609);
			4580: out = 16'(-19866);
			4581: out = 16'(-16563);
			4582: out = 16'(-6014);
			4583: out = 16'(15215);
			4584: out = 16'(8961);
			4585: out = 16'(7971);
			4586: out = 16'(-785);
			4587: out = 16'(7874);
			4588: out = 16'(7314);
			4589: out = 16'(3345);
			4590: out = 16'(-1178);
			4591: out = 16'(-2684);
			4592: out = 16'(-449);
			4593: out = 16'(701);
			4594: out = 16'(783);
			4595: out = 16'(-1330);
			4596: out = 16'(235);
			4597: out = 16'(3393);
			4598: out = 16'(-1758);
			4599: out = 16'(219);
			4600: out = 16'(1595);
			4601: out = 16'(13469);
			4602: out = 16'(11624);
			4603: out = 16'(4248);
			4604: out = 16'(-13309);
			4605: out = 16'(-21546);
			4606: out = 16'(-15685);
			4607: out = 16'(-8343);
			4608: out = 16'(-1817);
			4609: out = 16'(-12858);
			4610: out = 16'(-2290);
			4611: out = 16'(3460);
			4612: out = 16'(14409);
			4613: out = 16'(7151);
			4614: out = 16'(563);
			4615: out = 16'(-13483);
			4616: out = 16'(-8223);
			4617: out = 16'(1690);
			4618: out = 16'(5279);
			4619: out = 16'(2777);
			4620: out = 16'(-4355);
			4621: out = 16'(-11969);
			4622: out = 16'(-9345);
			4623: out = 16'(7958);
			4624: out = 16'(1251);
			4625: out = 16'(2564);
			4626: out = 16'(7210);
			4627: out = 16'(5173);
			4628: out = 16'(2561);
			4629: out = 16'(1090);
			4630: out = 16'(1916);
			4631: out = 16'(3836);
			4632: out = 16'(4339);
			4633: out = 16'(1007);
			4634: out = 16'(-5175);
			4635: out = 16'(-1617);
			4636: out = 16'(-5564);
			4637: out = 16'(-7612);
			4638: out = 16'(-6816);
			4639: out = 16'(1320);
			4640: out = 16'(12067);
			4641: out = 16'(14408);
			4642: out = 16'(9658);
			4643: out = 16'(-6293);
			4644: out = 16'(-2460);
			4645: out = 16'(-365);
			4646: out = 16'(3116);
			4647: out = 16'(2165);
			4648: out = 16'(969);
			4649: out = 16'(1869);
			4650: out = 16'(-4525);
			4651: out = 16'(-9933);
			4652: out = 16'(-560);
			4653: out = 16'(2529);
			4654: out = 16'(6264);
			4655: out = 16'(4130);
			4656: out = 16'(3374);
			4657: out = 16'(-308);
			4658: out = 16'(5923);
			4659: out = 16'(5792);
			4660: out = 16'(5541);
			4661: out = 16'(-3763);
			4662: out = 16'(-10573);
			4663: out = 16'(-22500);
			4664: out = 16'(-3603);
			4665: out = 16'(8588);
			4666: out = 16'(2284);
			4667: out = 16'(2251);
			4668: out = 16'(558);
			4669: out = 16'(11106);
			4670: out = 16'(12631);
			4671: out = 16'(14222);
			4672: out = 16'(-7873);
			4673: out = 16'(-11185);
			4674: out = 16'(-11669);
			4675: out = 16'(6678);
			4676: out = 16'(7176);
			4677: out = 16'(-1083);
			4678: out = 16'(-9658);
			4679: out = 16'(-11508);
			4680: out = 16'(1526);
			4681: out = 16'(-7727);
			4682: out = 16'(-6181);
			4683: out = 16'(9325);
			4684: out = 16'(9101);
			4685: out = 16'(8087);
			4686: out = 16'(-1767);
			4687: out = 16'(6479);
			4688: out = 16'(12161);
			4689: out = 16'(-5314);
			4690: out = 16'(-15432);
			4691: out = 16'(-26827);
			4692: out = 16'(1319);
			4693: out = 16'(8731);
			4694: out = 16'(12834);
			4695: out = 16'(-1095);
			4696: out = 16'(-3214);
			4697: out = 16'(32);
			4698: out = 16'(10568);
			4699: out = 16'(12903);
			4700: out = 16'(4746);
			4701: out = 16'(-547);
			4702: out = 16'(-5142);
			4703: out = 16'(210);
			4704: out = 16'(-2433);
			4705: out = 16'(-2239);
			4706: out = 16'(5004);
			4707: out = 16'(-2966);
			4708: out = 16'(-14152);
			4709: out = 16'(6553);
			4710: out = 16'(6172);
			4711: out = 16'(5750);
			4712: out = 16'(701);
			4713: out = 16'(3522);
			4714: out = 16'(5369);
			4715: out = 16'(13527);
			4716: out = 16'(5106);
			4717: out = 16'(-18858);
			4718: out = 16'(-24905);
			4719: out = 16'(-21480);
			4720: out = 16'(3977);
			4721: out = 16'(9947);
			4722: out = 16'(11722);
			4723: out = 16'(-5195);
			4724: out = 16'(-5751);
			4725: out = 16'(-4577);
			4726: out = 16'(5566);
			4727: out = 16'(6189);
			4728: out = 16'(3550);
			4729: out = 16'(10233);
			4730: out = 16'(2354);
			4731: out = 16'(-11303);
			4732: out = 16'(-16693);
			4733: out = 16'(-12182);
			4734: out = 16'(8777);
			4735: out = 16'(-1007);
			4736: out = 16'(-1894);
			4737: out = 16'(-1842);
			4738: out = 16'(5901);
			4739: out = 16'(8463);
			4740: out = 16'(1764);
			4741: out = 16'(-612);
			4742: out = 16'(-2591);
			4743: out = 16'(5407);
			4744: out = 16'(4424);
			4745: out = 16'(3296);
			4746: out = 16'(-14592);
			4747: out = 16'(-10277);
			4748: out = 16'(2949);
			4749: out = 16'(-1600);
			4750: out = 16'(-591);
			4751: out = 16'(-1530);
			4752: out = 16'(4269);
			4753: out = 16'(5341);
			4754: out = 16'(4266);
			4755: out = 16'(1649);
			4756: out = 16'(560);
			4757: out = 16'(4597);
			4758: out = 16'(-2506);
			4759: out = 16'(-7685);
			4760: out = 16'(-3732);
			4761: out = 16'(-3832);
			4762: out = 16'(-1745);
			4763: out = 16'(-745);
			4764: out = 16'(1078);
			4765: out = 16'(381);
			4766: out = 16'(10481);
			4767: out = 16'(6984);
			4768: out = 16'(-50);
			4769: out = 16'(-2218);
			4770: out = 16'(-1903);
			4771: out = 16'(-285);
			4772: out = 16'(6690);
			4773: out = 16'(7690);
			4774: out = 16'(4295);
			4775: out = 16'(-7584);
			4776: out = 16'(-16070);
			4777: out = 16'(-14216);
			4778: out = 16'(-5457);
			4779: out = 16'(6078);
			4780: out = 16'(7578);
			4781: out = 16'(6881);
			4782: out = 16'(260);
			4783: out = 16'(14473);
			4784: out = 16'(7820);
			4785: out = 16'(771);
			4786: out = 16'(-7419);
			4787: out = 16'(-8299);
			4788: out = 16'(-9166);
			4789: out = 16'(6196);
			4790: out = 16'(7740);
			4791: out = 16'(2187);
			4792: out = 16'(-16736);
			4793: out = 16'(-22140);
			4794: out = 16'(6112);
			4795: out = 16'(12763);
			4796: out = 16'(18200);
			4797: out = 16'(635);
			4798: out = 16'(245);
			4799: out = 16'(-3358);
			4800: out = 16'(12134);
			4801: out = 16'(7093);
			4802: out = 16'(3460);
			4803: out = 16'(-17047);
			4804: out = 16'(-14842);
			4805: out = 16'(-3221);
			4806: out = 16'(9220);
			4807: out = 16'(13102);
			4808: out = 16'(11683);
			4809: out = 16'(-4725);
			4810: out = 16'(-9967);
			4811: out = 16'(5904);
			4812: out = 16'(5815);
			4813: out = 16'(5897);
			4814: out = 16'(-6005);
			4815: out = 16'(-7978);
			4816: out = 16'(-9856);
			4817: out = 16'(-871);
			4818: out = 16'(4036);
			4819: out = 16'(9967);
			4820: out = 16'(-4522);
			4821: out = 16'(-6562);
			4822: out = 16'(-8797);
			4823: out = 16'(9409);
			4824: out = 16'(11584);
			4825: out = 16'(6858);
			4826: out = 16'(2888);
			4827: out = 16'(-170);
			4828: out = 16'(-3656);
			4829: out = 16'(-245);
			4830: out = 16'(-773);
			4831: out = 16'(-5134);
			4832: out = 16'(-14142);
			4833: out = 16'(-18104);
			4834: out = 16'(-981);
			4835: out = 16'(5961);
			4836: out = 16'(11616);
			4837: out = 16'(10864);
			4838: out = 16'(4317);
			4839: out = 16'(-7079);
			4840: out = 16'(4000);
			4841: out = 16'(5689);
			4842: out = 16'(8830);
			4843: out = 16'(-1959);
			4844: out = 16'(-5977);
			4845: out = 16'(-9408);
			4846: out = 16'(2494);
			4847: out = 16'(6710);
			4848: out = 16'(-902);
			4849: out = 16'(-5104);
			4850: out = 16'(-8351);
			4851: out = 16'(4283);
			4852: out = 16'(4682);
			4853: out = 16'(6606);
			4854: out = 16'(-19536);
			4855: out = 16'(-7963);
			4856: out = 16'(7674);
			4857: out = 16'(8719);
			4858: out = 16'(262);
			4859: out = 16'(-16278);
			4860: out = 16'(-12119);
			4861: out = 16'(-7336);
			4862: out = 16'(3975);
			4863: out = 16'(1769);
			4864: out = 16'(1938);
			4865: out = 16'(1811);
			4866: out = 16'(-1100);
			4867: out = 16'(-2373);
			4868: out = 16'(395);
			4869: out = 16'(2669);
			4870: out = 16'(4168);
			4871: out = 16'(1750);
			4872: out = 16'(3147);
			4873: out = 16'(4432);
			4874: out = 16'(-19185);
			4875: out = 16'(-13376);
			4876: out = 16'(2402);
			4877: out = 16'(7759);
			4878: out = 16'(9235);
			4879: out = 16'(3150);
			4880: out = 16'(3994);
			4881: out = 16'(1773);
			4882: out = 16'(1590);
			4883: out = 16'(563);
			4884: out = 16'(3037);
			4885: out = 16'(9601);
			4886: out = 16'(4634);
			4887: out = 16'(-3078);
			4888: out = 16'(-21580);
			4889: out = 16'(-16449);
			4890: out = 16'(-5506);
			4891: out = 16'(-1664);
			4892: out = 16'(5868);
			4893: out = 16'(8933);
			4894: out = 16'(13829);
			4895: out = 16'(3928);
			4896: out = 16'(-12819);
			4897: out = 16'(-755);
			4898: out = 16'(1932);
			4899: out = 16'(3048);
			4900: out = 16'(-3213);
			4901: out = 16'(-5781);
			4902: out = 16'(-3691);
			4903: out = 16'(-1730);
			4904: out = 16'(1128);
			4905: out = 16'(1481);
			4906: out = 16'(-938);
			4907: out = 16'(-2775);
			4908: out = 16'(15682);
			4909: out = 16'(10313);
			4910: out = 16'(6444);
			4911: out = 16'(-18378);
			4912: out = 16'(-7141);
			4913: out = 16'(12911);
			4914: out = 16'(13335);
			4915: out = 16'(5829);
			4916: out = 16'(-13623);
			4917: out = 16'(-5486);
			4918: out = 16'(-2999);
			4919: out = 16'(1424);
			4920: out = 16'(6255);
			4921: out = 16'(7868);
			4922: out = 16'(739);
			4923: out = 16'(1631);
			4924: out = 16'(747);
			4925: out = 16'(-481);
			4926: out = 16'(1794);
			4927: out = 16'(3352);
			4928: out = 16'(402);
			4929: out = 16'(-10933);
			4930: out = 16'(-25416);
			4931: out = 16'(-2890);
			4932: out = 16'(7204);
			4933: out = 16'(20896);
			4934: out = 16'(-12129);
			4935: out = 16'(-15285);
			4936: out = 16'(-6631);
			4937: out = 16'(13254);
			4938: out = 16'(16174);
			4939: out = 16'(-935);
			4940: out = 16'(-4755);
			4941: out = 16'(-9032);
			4942: out = 16'(-2039);
			4943: out = 16'(-1709);
			4944: out = 16'(1910);
			4945: out = 16'(4608);
			4946: out = 16'(2159);
			4947: out = 16'(-3406);
			4948: out = 16'(10100);
			4949: out = 16'(4152);
			4950: out = 16'(-1445);
			4951: out = 16'(-1197);
			4952: out = 16'(7094);
			4953: out = 16'(18223);
			4954: out = 16'(6377);
			4955: out = 16'(-5064);
			4956: out = 16'(-22080);
			4957: out = 16'(-12758);
			4958: out = 16'(-2345);
			4959: out = 16'(6470);
			4960: out = 16'(12581);
			4961: out = 16'(11239);
			4962: out = 16'(4121);
			4963: out = 16'(-12171);
			4964: out = 16'(-24792);
			4965: out = 16'(-8510);
			4966: out = 16'(2158);
			4967: out = 16'(14060);
			4968: out = 16'(-8170);
			4969: out = 16'(-4524);
			4970: out = 16'(4861);
			4971: out = 16'(-3663);
			4972: out = 16'(-6480);
			4973: out = 16'(-8256);
			4974: out = 16'(263);
			4975: out = 16'(1808);
			4976: out = 16'(-9156);
			4977: out = 16'(3985);
			4978: out = 16'(9408);
			4979: out = 16'(5587);
			4980: out = 16'(-1857);
			4981: out = 16'(-7083);
			4982: out = 16'(16790);
			4983: out = 16'(7932);
			4984: out = 16'(219);
			4985: out = 16'(-16520);
			4986: out = 16'(-9489);
			4987: out = 16'(4833);
			4988: out = 16'(7693);
			4989: out = 16'(6853);
			4990: out = 16'(486);
			4991: out = 16'(-4762);
			4992: out = 16'(-5519);
			4993: out = 16'(2091);
			4994: out = 16'(4534);
			4995: out = 16'(6170);
			4996: out = 16'(-462);
			4997: out = 16'(1590);
			4998: out = 16'(-870);
			4999: out = 16'(-9018);
			5000: out = 16'(-9651);
			5001: out = 16'(-6524);
			5002: out = 16'(3098);
			5003: out = 16'(3484);
			5004: out = 16'(-243);
			5005: out = 16'(2586);
			5006: out = 16'(523);
			5007: out = 16'(613);
			5008: out = 16'(-9639);
			5009: out = 16'(-6498);
			5010: out = 16'(5229);
			5011: out = 16'(4540);
			5012: out = 16'(1886);
			5013: out = 16'(-8531);
			5014: out = 16'(-2658);
			5015: out = 16'(1091);
			5016: out = 16'(-1817);
			5017: out = 16'(8392);
			5018: out = 16'(13817);
			5019: out = 16'(2081);
			5020: out = 16'(-107);
			5021: out = 16'(-2680);
			5022: out = 16'(8590);
			5023: out = 16'(1483);
			5024: out = 16'(-10759);
			5025: out = 16'(4405);
			5026: out = 16'(8139);
			5027: out = 16'(12276);
			5028: out = 16'(-8541);
			5029: out = 16'(-14792);
			5030: out = 16'(-9320);
			5031: out = 16'(2538);
			5032: out = 16'(9480);
			5033: out = 16'(337);
			5034: out = 16'(2642);
			5035: out = 16'(592);
			5036: out = 16'(7917);
			5037: out = 16'(-3051);
			5038: out = 16'(-10295);
			5039: out = 16'(-10745);
			5040: out = 16'(-731);
			5041: out = 16'(11124);
			5042: out = 16'(5397);
			5043: out = 16'(5326);
			5044: out = 16'(4901);
			5045: out = 16'(-2375);
			5046: out = 16'(-3404);
			5047: out = 16'(1656);
			5048: out = 16'(852);
			5049: out = 16'(3006);
			5050: out = 16'(7435);
			5051: out = 16'(4231);
			5052: out = 16'(1412);
			5053: out = 16'(-1800);
			5054: out = 16'(-282);
			5055: out = 16'(2193);
			5056: out = 16'(8966);
			5057: out = 16'(5259);
			5058: out = 16'(-55);
			5059: out = 16'(-1611);
			5060: out = 16'(-828);
			5061: out = 16'(2714);
			5062: out = 16'(2735);
			5063: out = 16'(2813);
			5064: out = 16'(163);
			5065: out = 16'(-128);
			5066: out = 16'(-1553);
			5067: out = 16'(-540);
			5068: out = 16'(-1076);
			5069: out = 16'(-788);
			5070: out = 16'(-5660);
			5071: out = 16'(-897);
			5072: out = 16'(1093);
			5073: out = 16'(3638);
			5074: out = 16'(4021);
			5075: out = 16'(4454);
			5076: out = 16'(-20643);
			5077: out = 16'(-16451);
			5078: out = 16'(-7234);
			5079: out = 16'(13776);
			5080: out = 16'(12496);
			5081: out = 16'(3800);
			5082: out = 16'(-11916);
			5083: out = 16'(-16663);
			5084: out = 16'(-12986);
			5085: out = 16'(5679);
			5086: out = 16'(13749);
			5087: out = 16'(10493);
			5088: out = 16'(-5055);
			5089: out = 16'(-16654);
			5090: out = 16'(-12926);
			5091: out = 16'(3150);
			5092: out = 16'(18545);
			5093: out = 16'(374);
			5094: out = 16'(-263);
			5095: out = 16'(-7430);
			5096: out = 16'(6061);
			5097: out = 16'(1275);
			5098: out = 16'(565);
			5099: out = 16'(-18066);
			5100: out = 16'(-11553);
			5101: out = 16'(4808);
			5102: out = 16'(10094);
			5103: out = 16'(6713);
			5104: out = 16'(-3786);
			5105: out = 16'(-16785);
			5106: out = 16'(-18728);
			5107: out = 16'(1507);
			5108: out = 16'(10160);
			5109: out = 16'(13612);
			5110: out = 16'(-6288);
			5111: out = 16'(-8077);
			5112: out = 16'(-8933);
			5113: out = 16'(-100);
			5114: out = 16'(1768);
			5115: out = 16'(2381);
			5116: out = 16'(11732);
			5117: out = 16'(6516);
			5118: out = 16'(-4953);
			5119: out = 16'(-9530);
			5120: out = 16'(-6360);
			5121: out = 16'(9656);
			5122: out = 16'(1599);
			5123: out = 16'(130);
			5124: out = 16'(-1532);
			5125: out = 16'(2039);
			5126: out = 16'(1791);
			5127: out = 16'(-6621);
			5128: out = 16'(-5238);
			5129: out = 16'(-1462);
			5130: out = 16'(13595);
			5131: out = 16'(11359);
			5132: out = 16'(5876);
			5133: out = 16'(-10082);
			5134: out = 16'(-12619);
			5135: out = 16'(-8254);
			5136: out = 16'(4450);
			5137: out = 16'(7456);
			5138: out = 16'(147);
			5139: out = 16'(9381);
			5140: out = 16'(5110);
			5141: out = 16'(-8757);
			5142: out = 16'(-5615);
			5143: out = 16'(-1773);
			5144: out = 16'(5547);
			5145: out = 16'(3150);
			5146: out = 16'(1035);
			5147: out = 16'(1994);
			5148: out = 16'(1298);
			5149: out = 16'(1308);
			5150: out = 16'(-137);
			5151: out = 16'(281);
			5152: out = 16'(434);
			5153: out = 16'(3581);
			5154: out = 16'(5599);
			5155: out = 16'(9078);
			5156: out = 16'(863);
			5157: out = 16'(1802);
			5158: out = 16'(7361);
			5159: out = 16'(9871);
			5160: out = 16'(5330);
			5161: out = 16'(-14301);
			5162: out = 16'(-8901);
			5163: out = 16'(-3234);
			5164: out = 16'(9278);
			5165: out = 16'(6091);
			5166: out = 16'(2945);
			5167: out = 16'(2490);
			5168: out = 16'(1955);
			5169: out = 16'(1597);
			5170: out = 16'(-9677);
			5171: out = 16'(-2083);
			5172: out = 16'(14146);
			5173: out = 16'(-5616);
			5174: out = 16'(-7685);
			5175: out = 16'(-10032);
			5176: out = 16'(5176);
			5177: out = 16'(7253);
			5178: out = 16'(7014);
			5179: out = 16'(-15209);
			5180: out = 16'(-21859);
			5181: out = 16'(64);
			5182: out = 16'(11422);
			5183: out = 16'(18105);
			5184: out = 16'(-636);
			5185: out = 16'(-7035);
			5186: out = 16'(-15307);
			5187: out = 16'(10445);
			5188: out = 16'(2032);
			5189: out = 16'(-7648);
			5190: out = 16'(-4444);
			5191: out = 16'(3464);
			5192: out = 16'(14050);
			5193: out = 16'(-474);
			5194: out = 16'(-8883);
			5195: out = 16'(-16490);
			5196: out = 16'(-4816);
			5197: out = 16'(4065);
			5198: out = 16'(3797);
			5199: out = 16'(8877);
			5200: out = 16'(5946);
			5201: out = 16'(3027);
			5202: out = 16'(-16975);
			5203: out = 16'(-27447);
			5204: out = 16'(-2897);
			5205: out = 16'(12263);
			5206: out = 16'(21317);
			5207: out = 16'(3328);
			5208: out = 16'(-11872);
			5209: out = 16'(-30020);
			5210: out = 16'(-7200);
			5211: out = 16'(6417);
			5212: out = 16'(17753);
			5213: out = 16'(6802);
			5214: out = 16'(-1959);
			5215: out = 16'(-14780);
			5216: out = 16'(-5648);
			5217: out = 16'(-988);
			5218: out = 16'(-10562);
			5219: out = 16'(646);
			5220: out = 16'(7293);
			5221: out = 16'(14001);
			5222: out = 16'(4275);
			5223: out = 16'(-4650);
			5224: out = 16'(-2716);
			5225: out = 16'(2619);
			5226: out = 16'(9726);
			5227: out = 16'(4475);
			5228: out = 16'(7331);
			5229: out = 16'(14613);
			5230: out = 16'(-4589);
			5231: out = 16'(-9623);
			5232: out = 16'(-12236);
			5233: out = 16'(7640);
			5234: out = 16'(11802);
			5235: out = 16'(1248);
			5236: out = 16'(-10860);
			5237: out = 16'(-17302);
			5238: out = 16'(-7577);
			5239: out = 16'(6695);
			5240: out = 16'(18126);
			5241: out = 16'(11040);
			5242: out = 16'(-860);
			5243: out = 16'(-18678);
			5244: out = 16'(-5452);
			5245: out = 16'(-4222);
			5246: out = 16'(2060);
			5247: out = 16'(-4477);
			5248: out = 16'(-604);
			5249: out = 16'(2533);
			5250: out = 16'(6022);
			5251: out = 16'(1787);
			5252: out = 16'(-6162);
			5253: out = 16'(-13557);
			5254: out = 16'(-11353);
			5255: out = 16'(9134);
			5256: out = 16'(12482);
			5257: out = 16'(12208);
			5258: out = 16'(-4356);
			5259: out = 16'(-11920);
			5260: out = 16'(-18245);
			5261: out = 16'(12896);
			5262: out = 16'(8206);
			5263: out = 16'(-150);
			5264: out = 16'(-157);
			5265: out = 16'(3736);
			5266: out = 16'(8976);
			5267: out = 16'(6689);
			5268: out = 16'(2994);
			5269: out = 16'(978);
			5270: out = 16'(-9635);
			5271: out = 16'(-11663);
			5272: out = 16'(-7637);
			5273: out = 16'(7752);
			5274: out = 16'(14022);
			5275: out = 16'(925);
			5276: out = 16'(-8168);
			5277: out = 16'(-15746);
			5278: out = 16'(-936);
			5279: out = 16'(6827);
			5280: out = 16'(14713);
			5281: out = 16'(3025);
			5282: out = 16'(-2937);
			5283: out = 16'(-12232);
			5284: out = 16'(-3969);
			5285: out = 16'(1156);
			5286: out = 16'(11153);
			5287: out = 16'(2320);
			5288: out = 16'(-1740);
			5289: out = 16'(-12430);
			5290: out = 16'(4311);
			5291: out = 16'(10738);
			5292: out = 16'(4398);
			5293: out = 16'(-4551);
			5294: out = 16'(-9900);
			5295: out = 16'(11648);
			5296: out = 16'(12946);
			5297: out = 16'(13901);
			5298: out = 16'(-7244);
			5299: out = 16'(-4969);
			5300: out = 16'(1839);
			5301: out = 16'(10877);
			5302: out = 16'(8617);
			5303: out = 16'(-2142);
			5304: out = 16'(-1997);
			5305: out = 16'(-3871);
			5306: out = 16'(421);
			5307: out = 16'(-7706);
			5308: out = 16'(-4450);
			5309: out = 16'(12533);
			5310: out = 16'(9508);
			5311: out = 16'(3119);
			5312: out = 16'(-14012);
			5313: out = 16'(-14571);
			5314: out = 16'(-9658);
			5315: out = 16'(-537);
			5316: out = 16'(1945);
			5317: out = 16'(-1152);
			5318: out = 16'(8026);
			5319: out = 16'(4253);
			5320: out = 16'(3207);
			5321: out = 16'(-19099);
			5322: out = 16'(-15775);
			5323: out = 16'(1952);
			5324: out = 16'(13544);
			5325: out = 16'(12923);
			5326: out = 16'(-1892);
			5327: out = 16'(-9143);
			5328: out = 16'(-14185);
			5329: out = 16'(-18827);
			5330: out = 16'(1315);
			5331: out = 16'(16116);
			5332: out = 16'(12279);
			5333: out = 16'(-1184);
			5334: out = 16'(-17604);
			5335: out = 16'(-743);
			5336: out = 16'(4014);
			5337: out = 16'(11036);
			5338: out = 16'(8700);
			5339: out = 16'(5162);
			5340: out = 16'(-4190);
			5341: out = 16'(-6785);
			5342: out = 16'(-7215);
			5343: out = 16'(1492);
			5344: out = 16'(-698);
			5345: out = 16'(-512);
			5346: out = 16'(-8054);
			5347: out = 16'(1697);
			5348: out = 16'(3849);
			5349: out = 16'(-7747);
			5350: out = 16'(-10138);
			5351: out = 16'(-8657);
			5352: out = 16'(10759);
			5353: out = 16'(14153);
			5354: out = 16'(13701);
			5355: out = 16'(-10645);
			5356: out = 16'(-12498);
			5357: out = 16'(-3822);
			5358: out = 16'(-5344);
			5359: out = 16'(-518);
			5360: out = 16'(3031);
			5361: out = 16'(9878);
			5362: out = 16'(9463);
			5363: out = 16'(4408);
			5364: out = 16'(-5087);
			5365: out = 16'(-7199);
			5366: out = 16'(13197);
			5367: out = 16'(5120);
			5368: out = 16'(-512);
			5369: out = 16'(-17929);
			5370: out = 16'(-4480);
			5371: out = 16'(10481);
			5372: out = 16'(-1193);
			5373: out = 16'(-4039);
			5374: out = 16'(-9981);
			5375: out = 16'(11765);
			5376: out = 16'(12984);
			5377: out = 16'(10755);
			5378: out = 16'(-3485);
			5379: out = 16'(-5722);
			5380: out = 16'(1568);
			5381: out = 16'(4740);
			5382: out = 16'(4541);
			5383: out = 16'(-4723);
			5384: out = 16'(-7631);
			5385: out = 16'(-8685);
			5386: out = 16'(5996);
			5387: out = 16'(-1127);
			5388: out = 16'(-5358);
			5389: out = 16'(-716);
			5390: out = 16'(4290);
			5391: out = 16'(9110);
			5392: out = 16'(1995);
			5393: out = 16'(1012);
			5394: out = 16'(-633);
			5395: out = 16'(5958);
			5396: out = 16'(749);
			5397: out = 16'(-12565);
			5398: out = 16'(-9537);
			5399: out = 16'(-2464);
			5400: out = 16'(18660);
			5401: out = 16'(4662);
			5402: out = 16'(-1881);
			5403: out = 16'(-12455);
			5404: out = 16'(2939);
			5405: out = 16'(12586);
			5406: out = 16'(8860);
			5407: out = 16'(-2797);
			5408: out = 16'(-15737);
			5409: out = 16'(4734);
			5410: out = 16'(1752);
			5411: out = 16'(-1822);
			5412: out = 16'(-9181);
			5413: out = 16'(-4183);
			5414: out = 16'(8945);
			5415: out = 16'(-9165);
			5416: out = 16'(-9931);
			5417: out = 16'(1458);
			5418: out = 16'(809);
			5419: out = 16'(2503);
			5420: out = 16'(716);
			5421: out = 16'(8778);
			5422: out = 16'(8470);
			5423: out = 16'(-17716);
			5424: out = 16'(-9032);
			5425: out = 16'(958);
			5426: out = 16'(5769);
			5427: out = 16'(4507);
			5428: out = 16'(-617);
			5429: out = 16'(1346);
			5430: out = 16'(-2327);
			5431: out = 16'(-5116);
			5432: out = 16'(-220);
			5433: out = 16'(1869);
			5434: out = 16'(-496);
			5435: out = 16'(8784);
			5436: out = 16'(11788);
			5437: out = 16'(15524);
			5438: out = 16'(-3661);
			5439: out = 16'(-14857);
			5440: out = 16'(-9231);
			5441: out = 16'(-4585);
			5442: out = 16'(3209);
			5443: out = 16'(-1766);
			5444: out = 16'(6892);
			5445: out = 16'(10177);
			5446: out = 16'(10257);
			5447: out = 16'(-2916);
			5448: out = 16'(-18799);
			5449: out = 16'(-2979);
			5450: out = 16'(6714);
			5451: out = 16'(17252);
			5452: out = 16'(4937);
			5453: out = 16'(-4410);
			5454: out = 16'(-18665);
			5455: out = 16'(-11891);
			5456: out = 16'(-3735);
			5457: out = 16'(12568);
			5458: out = 16'(5290);
			5459: out = 16'(731);
			5460: out = 16'(-1567);
			5461: out = 16'(3924);
			5462: out = 16'(9050);
			5463: out = 16'(3697);
			5464: out = 16'(2395);
			5465: out = 16'(-975);
			5466: out = 16'(330);
			5467: out = 16'(-2713);
			5468: out = 16'(-4268);
			5469: out = 16'(-8647);
			5470: out = 16'(-4466);
			5471: out = 16'(5861);
			5472: out = 16'(-1109);
			5473: out = 16'(-567);
			5474: out = 16'(10551);
			5475: out = 16'(4316);
			5476: out = 16'(374);
			5477: out = 16'(-14209);
			5478: out = 16'(-2707);
			5479: out = 16'(4295);
			5480: out = 16'(4759);
			5481: out = 16'(-5441);
			5482: out = 16'(-15717);
			5483: out = 16'(-18073);
			5484: out = 16'(-7602);
			5485: out = 16'(8916);
			5486: out = 16'(10356);
			5487: out = 16'(3869);
			5488: out = 16'(-16558);
			5489: out = 16'(-2086);
			5490: out = 16'(1480);
			5491: out = 16'(6628);
			5492: out = 16'(-3453);
			5493: out = 16'(-4188);
			5494: out = 16'(8562);
			5495: out = 16'(4095);
			5496: out = 16'(332);
			5497: out = 16'(-8073);
			5498: out = 16'(-3876);
			5499: out = 16'(1565);
			5500: out = 16'(6369);
			5501: out = 16'(2490);
			5502: out = 16'(-4197);
			5503: out = 16'(9900);
			5504: out = 16'(9395);
			5505: out = 16'(5977);
			5506: out = 16'(2627);
			5507: out = 16'(-2879);
			5508: out = 16'(-12116);
			5509: out = 16'(-3109);
			5510: out = 16'(1196);
			5511: out = 16'(2977);
			5512: out = 16'(185);
			5513: out = 16'(-1404);
			5514: out = 16'(-60);
			5515: out = 16'(3568);
			5516: out = 16'(7114);
			5517: out = 16'(4682);
			5518: out = 16'(5608);
			5519: out = 16'(4031);
			5520: out = 16'(2246);
			5521: out = 16'(-5410);
			5522: out = 16'(-13543);
			5523: out = 16'(-3697);
			5524: out = 16'(1269);
			5525: out = 16'(5253);
			5526: out = 16'(-1634);
			5527: out = 16'(-6749);
			5528: out = 16'(-11200);
			5529: out = 16'(-4157);
			5530: out = 16'(2577);
			5531: out = 16'(3155);
			5532: out = 16'(11951);
			5533: out = 16'(13987);
			5534: out = 16'(9259);
			5535: out = 16'(1993);
			5536: out = 16'(-4319);
			5537: out = 16'(-7099);
			5538: out = 16'(-4301);
			5539: out = 16'(595);
			5540: out = 16'(6233);
			5541: out = 16'(5656);
			5542: out = 16'(1836);
			5543: out = 16'(-1847);
			5544: out = 16'(-3504);
			5545: out = 16'(-3030);
			5546: out = 16'(1775);
			5547: out = 16'(5008);
			5548: out = 16'(8381);
			5549: out = 16'(811);
			5550: out = 16'(-6373);
			5551: out = 16'(-17843);
			5552: out = 16'(-12160);
			5553: out = 16'(-3954);
			5554: out = 16'(9784);
			5555: out = 16'(9666);
			5556: out = 16'(6800);
			5557: out = 16'(-17014);
			5558: out = 16'(-11639);
			5559: out = 16'(3537);
			5560: out = 16'(13015);
			5561: out = 16'(11789);
			5562: out = 16'(-492);
			5563: out = 16'(-5080);
			5564: out = 16'(-9486);
			5565: out = 16'(-4296);
			5566: out = 16'(-7619);
			5567: out = 16'(-4500);
			5568: out = 16'(-167);
			5569: out = 16'(3323);
			5570: out = 16'(4305);
			5571: out = 16'(6949);
			5572: out = 16'(1200);
			5573: out = 16'(-1932);
			5574: out = 16'(10747);
			5575: out = 16'(12003);
			5576: out = 16'(11503);
			5577: out = 16'(-123);
			5578: out = 16'(-3474);
			5579: out = 16'(-4778);
			5580: out = 16'(-202);
			5581: out = 16'(-1557);
			5582: out = 16'(-7893);
			5583: out = 16'(-3208);
			5584: out = 16'(-752);
			5585: out = 16'(1242);
			5586: out = 16'(1265);
			5587: out = 16'(1240);
			5588: out = 16'(1180);
			5589: out = 16'(2571);
			5590: out = 16'(3052);
			5591: out = 16'(-4535);
			5592: out = 16'(-2286);
			5593: out = 16'(-759);
			5594: out = 16'(-2261);
			5595: out = 16'(-7968);
			5596: out = 16'(-14462);
			5597: out = 16'(-1584);
			5598: out = 16'(4296);
			5599: out = 16'(7507);
			5600: out = 16'(10340);
			5601: out = 16'(7490);
			5602: out = 16'(-306);
			5603: out = 16'(-8825);
			5604: out = 16'(-10837);
			5605: out = 16'(6383);
			5606: out = 16'(3153);
			5607: out = 16'(2615);
			5608: out = 16'(-17474);
			5609: out = 16'(-25);
			5610: out = 16'(12526);
			5611: out = 16'(10052);
			5612: out = 16'(940);
			5613: out = 16'(-9463);
			5614: out = 16'(-6572);
			5615: out = 16'(1557);
			5616: out = 16'(13506);
			5617: out = 16'(11641);
			5618: out = 16'(5265);
			5619: out = 16'(-10183);
			5620: out = 16'(-11601);
			5621: out = 16'(-10784);
			5622: out = 16'(2669);
			5623: out = 16'(-4940);
			5624: out = 16'(-5658);
			5625: out = 16'(12);
			5626: out = 16'(3264);
			5627: out = 16'(4355);
			5628: out = 16'(-6821);
			5629: out = 16'(-2802);
			5630: out = 16'(2328);
			5631: out = 16'(8958);
			5632: out = 16'(5877);
			5633: out = 16'(-892);
			5634: out = 16'(-1889);
			5635: out = 16'(-3851);
			5636: out = 16'(-4033);
			5637: out = 16'(-6461);
			5638: out = 16'(-5611);
			5639: out = 16'(-752);
			5640: out = 16'(-408);
			5641: out = 16'(-4);
			5642: out = 16'(-7757);
			5643: out = 16'(3092);
			5644: out = 16'(8993);
			5645: out = 16'(15522);
			5646: out = 16'(4143);
			5647: out = 16'(-6281);
			5648: out = 16'(-17039);
			5649: out = 16'(-7503);
			5650: out = 16'(7564);
			5651: out = 16'(9801);
			5652: out = 16'(4090);
			5653: out = 16'(-11612);
			5654: out = 16'(-1897);
			5655: out = 16'(-526);
			5656: out = 16'(3853);
			5657: out = 16'(245);
			5658: out = 16'(1987);
			5659: out = 16'(4888);
			5660: out = 16'(4141);
			5661: out = 16'(662);
			5662: out = 16'(-4975);
			5663: out = 16'(-6784);
			5664: out = 16'(-6601);
			5665: out = 16'(-8534);
			5666: out = 16'(-3721);
			5667: out = 16'(1231);
			5668: out = 16'(2709);
			5669: out = 16'(4870);
			5670: out = 16'(6905);
			5671: out = 16'(4328);
			5672: out = 16'(5120);
			5673: out = 16'(6192);
			5674: out = 16'(4873);
			5675: out = 16'(2212);
			5676: out = 16'(87);
			5677: out = 16'(-9151);
			5678: out = 16'(-12017);
			5679: out = 16'(-5174);
			5680: out = 16'(960);
			5681: out = 16'(5522);
			5682: out = 16'(-4654);
			5683: out = 16'(2256);
			5684: out = 16'(7514);
			5685: out = 16'(12435);
			5686: out = 16'(8263);
			5687: out = 16'(1332);
			5688: out = 16'(3416);
			5689: out = 16'(-2122);
			5690: out = 16'(-8994);
			5691: out = 16'(-6583);
			5692: out = 16'(-1742);
			5693: out = 16'(8179);
			5694: out = 16'(-1474);
			5695: out = 16'(-4083);
			5696: out = 16'(-1350);
			5697: out = 16'(251);
			5698: out = 16'(1828);
			5699: out = 16'(757);
			5700: out = 16'(2825);
			5701: out = 16'(4319);
			5702: out = 16'(8478);
			5703: out = 16'(406);
			5704: out = 16'(-9441);
			5705: out = 16'(7962);
			5706: out = 16'(3477);
			5707: out = 16'(-2509);
			5708: out = 16'(-21836);
			5709: out = 16'(-19278);
			5710: out = 16'(1184);
			5711: out = 16'(-771);
			5712: out = 16'(7936);
			5713: out = 16'(18546);
			5714: out = 16'(18089);
			5715: out = 16'(8004);
			5716: out = 16'(-25647);
			5717: out = 16'(-18107);
			5718: out = 16'(-6127);
			5719: out = 16'(14435);
			5720: out = 16'(12463);
			5721: out = 16'(5486);
			5722: out = 16'(-11701);
			5723: out = 16'(-14950);
			5724: out = 16'(-10798);
			5725: out = 16'(2968);
			5726: out = 16'(8443);
			5727: out = 16'(6667);
			5728: out = 16'(10140);
			5729: out = 16'(6370);
			5730: out = 16'(945);
			5731: out = 16'(1122);
			5732: out = 16'(-1803);
			5733: out = 16'(-17379);
			5734: out = 16'(-5158);
			5735: out = 16'(-76);
			5736: out = 16'(-482);
			5737: out = 16'(-10513);
			5738: out = 16'(-15729);
			5739: out = 16'(1703);
			5740: out = 16'(9019);
			5741: out = 16'(14394);
			5742: out = 16'(12262);
			5743: out = 16'(6426);
			5744: out = 16'(-2819);
			5745: out = 16'(-6748);
			5746: out = 16'(-7476);
			5747: out = 16'(-1817);
			5748: out = 16'(-5386);
			5749: out = 16'(-3397);
			5750: out = 16'(1945);
			5751: out = 16'(-1107);
			5752: out = 16'(-3628);
			5753: out = 16'(-8394);
			5754: out = 16'(739);
			5755: out = 16'(7986);
			5756: out = 16'(6062);
			5757: out = 16'(3865);
			5758: out = 16'(-540);
			5759: out = 16'(9267);
			5760: out = 16'(1427);
			5761: out = 16'(-7535);
			5762: out = 16'(-1072);
			5763: out = 16'(1512);
			5764: out = 16'(3984);
			5765: out = 16'(-4345);
			5766: out = 16'(-8820);
			5767: out = 16'(-10747);
			5768: out = 16'(-5830);
			5769: out = 16'(2842);
			5770: out = 16'(15934);
			5771: out = 16'(10274);
			5772: out = 16'(3900);
			5773: out = 16'(-385);
			5774: out = 16'(-5240);
			5775: out = 16'(-7717);
			5776: out = 16'(-17686);
			5777: out = 16'(-8140);
			5778: out = 16'(3840);
			5779: out = 16'(6005);
			5780: out = 16'(2357);
			5781: out = 16'(-7491);
			5782: out = 16'(8189);
			5783: out = 16'(8537);
			5784: out = 16'(5252);
			5785: out = 16'(4443);
			5786: out = 16'(3104);
			5787: out = 16'(-552);
			5788: out = 16'(2292);
			5789: out = 16'(1019);
			5790: out = 16'(-5341);
			5791: out = 16'(-7452);
			5792: out = 16'(-7415);
			5793: out = 16'(-1736);
			5794: out = 16'(3499);
			5795: out = 16'(8665);
			5796: out = 16'(8287);
			5797: out = 16'(4300);
			5798: out = 16'(-3838);
			5799: out = 16'(12974);
			5800: out = 16'(8974);
			5801: out = 16'(3502);
			5802: out = 16'(-11828);
			5803: out = 16'(-9241);
			5804: out = 16'(7018);
			5805: out = 16'(5971);
			5806: out = 16'(2704);
			5807: out = 16'(-8925);
			5808: out = 16'(-11737);
			5809: out = 16'(-10054);
			5810: out = 16'(6112);
			5811: out = 16'(9854);
			5812: out = 16'(11849);
			5813: out = 16'(-379);
			5814: out = 16'(2239);
			5815: out = 16'(4722);
			5816: out = 16'(1277);
			5817: out = 16'(511);
			5818: out = 16'(-599);
			5819: out = 16'(878);
			5820: out = 16'(-763);
			5821: out = 16'(-1665);
			5822: out = 16'(-9108);
			5823: out = 16'(-4129);
			5824: out = 16'(14401);
			5825: out = 16'(8461);
			5826: out = 16'(3673);
			5827: out = 16'(-11140);
			5828: out = 16'(2289);
			5829: out = 16'(9709);
			5830: out = 16'(-5680);
			5831: out = 16'(-1559);
			5832: out = 16'(-735);
			5833: out = 16'(6663);
			5834: out = 16'(-3593);
			5835: out = 16'(-14057);
			5836: out = 16'(-12617);
			5837: out = 16'(-6976);
			5838: out = 16'(232);
			5839: out = 16'(12273);
			5840: out = 16'(10582);
			5841: out = 16'(502);
			5842: out = 16'(-9171);
			5843: out = 16'(-11648);
			5844: out = 16'(-1055);
			5845: out = 16'(31);
			5846: out = 16'(2349);
			5847: out = 16'(6640);
			5848: out = 16'(-4578);
			5849: out = 16'(-15411);
			5850: out = 16'(-22921);
			5851: out = 16'(-12325);
			5852: out = 16'(5634);
			5853: out = 16'(8368);
			5854: out = 16'(13466);
			5855: out = 16'(10238);
			5856: out = 16'(13904);
			5857: out = 16'(964);
			5858: out = 16'(-18388);
			5859: out = 16'(-10944);
			5860: out = 16'(-3302);
			5861: out = 16'(8187);
			5862: out = 16'(887);
			5863: out = 16'(-5087);
			5864: out = 16'(-12181);
			5865: out = 16'(-4908);
			5866: out = 16'(2609);
			5867: out = 16'(-539);
			5868: out = 16'(5742);
			5869: out = 16'(7802);
			5870: out = 16'(11630);
			5871: out = 16'(7424);
			5872: out = 16'(4589);
			5873: out = 16'(-16728);
			5874: out = 16'(-12768);
			5875: out = 16'(108);
			5876: out = 16'(13267);
			5877: out = 16'(7951);
			5878: out = 16'(-15861);
			5879: out = 16'(-11506);
			5880: out = 16'(-5101);
			5881: out = 16'(16422);
			5882: out = 16'(10357);
			5883: out = 16'(5947);
			5884: out = 16'(-11529);
			5885: out = 16'(-3373);
			5886: out = 16'(1743);
			5887: out = 16'(-4919);
			5888: out = 16'(-5832);
			5889: out = 16'(-5280);
			5890: out = 16'(9360);
			5891: out = 16'(11696);
			5892: out = 16'(11146);
			5893: out = 16'(-5915);
			5894: out = 16'(-7651);
			5895: out = 16'(1446);
			5896: out = 16'(3047);
			5897: out = 16'(6564);
			5898: out = 16'(4007);
			5899: out = 16'(10708);
			5900: out = 16'(8940);
			5901: out = 16'(3389);
			5902: out = 16'(-10046);
			5903: out = 16'(-17017);
			5904: out = 16'(183);
			5905: out = 16'(-981);
			5906: out = 16'(-1657);
			5907: out = 16'(-8337);
			5908: out = 16'(-1754);
			5909: out = 16'(7515);
			5910: out = 16'(635);
			5911: out = 16'(-2357);
			5912: out = 16'(-10634);
			5913: out = 16'(8943);
			5914: out = 16'(9278);
			5915: out = 16'(4329);
			5916: out = 16'(-13996);
			5917: out = 16'(-18071);
			5918: out = 16'(-132);
			5919: out = 16'(322);
			5920: out = 16'(3640);
			5921: out = 16'(9155);
			5922: out = 16'(-979);
			5923: out = 16'(-10342);
			5924: out = 16'(-3580);
			5925: out = 16'(3781);
			5926: out = 16'(14477);
			5927: out = 16'(178);
			5928: out = 16'(-1835);
			5929: out = 16'(-9282);
			5930: out = 16'(16735);
			5931: out = 16'(12889);
			5932: out = 16'(2640);
			5933: out = 16'(-15523);
			5934: out = 16'(-17071);
			5935: out = 16'(-561);
			5936: out = 16'(5988);
			5937: out = 16'(11462);
			5938: out = 16'(14886);
			5939: out = 16'(5569);
			5940: out = 16'(-2983);
			5941: out = 16'(-14604);
			5942: out = 16'(-1645);
			5943: out = 16'(12169);
			5944: out = 16'(7167);
			5945: out = 16'(-244);
			5946: out = 16'(-13426);
			5947: out = 16'(-9321);
			5948: out = 16'(-6990);
			5949: out = 16'(1947);
			5950: out = 16'(1287);
			5951: out = 16'(3729);
			5952: out = 16'(480);
			5953: out = 16'(5370);
			5954: out = 16'(2371);
			5955: out = 16'(-3394);
			5956: out = 16'(-8599);
			5957: out = 16'(-5389);
			5958: out = 16'(14196);
			5959: out = 16'(14026);
			5960: out = 16'(8564);
			5961: out = 16'(-16531);
			5962: out = 16'(-21951);
			5963: out = 16'(-19274);
			5964: out = 16'(3261);
			5965: out = 16'(13966);
			5966: out = 16'(17244);
			5967: out = 16'(6674);
			5968: out = 16'(-4036);
			5969: out = 16'(-14154);
			5970: out = 16'(-9867);
			5971: out = 16'(-331);
			5972: out = 16'(12757);
			5973: out = 16'(12289);
			5974: out = 16'(5894);
			5975: out = 16'(-8765);
			5976: out = 16'(-15247);
			5977: out = 16'(-14895);
			5978: out = 16'(-1002);
			5979: out = 16'(9577);
			5980: out = 16'(15146);
			5981: out = 16'(2205);
			5982: out = 16'(-7458);
			5983: out = 16'(-18056);
			5984: out = 16'(-6803);
			5985: out = 16'(-2133);
			5986: out = 16'(2554);
			5987: out = 16'(-209);
			5988: out = 16'(-683);
			5989: out = 16'(887);
			5990: out = 16'(-4662);
			5991: out = 16'(-5854);
			5992: out = 16'(-5085);
			5993: out = 16'(3958);
			5994: out = 16'(8134);
			5995: out = 16'(2109);
			5996: out = 16'(2194);
			5997: out = 16'(573);
			5998: out = 16'(-10118);
			5999: out = 16'(-7168);
			6000: out = 16'(-1726);
			6001: out = 16'(10994);
			6002: out = 16'(10879);
			6003: out = 16'(7202);
			6004: out = 16'(-9879);
			6005: out = 16'(-12327);
			6006: out = 16'(-5191);
			6007: out = 16'(8488);
			6008: out = 16'(12677);
			6009: out = 16'(3371);
			6010: out = 16'(2829);
			6011: out = 16'(-50);
			6012: out = 16'(2621);
			6013: out = 16'(595);
			6014: out = 16'(844);
			6015: out = 16'(50);
			6016: out = 16'(-1599);
			6017: out = 16'(-3873);
			6018: out = 16'(1924);
			6019: out = 16'(1573);
			6020: out = 16'(1873);
			6021: out = 16'(-7244);
			6022: out = 16'(-2855);
			6023: out = 16'(7796);
			6024: out = 16'(2592);
			6025: out = 16'(-2384);
			6026: out = 16'(-16974);
			6027: out = 16'(502);
			6028: out = 16'(8095);
			6029: out = 16'(14980);
			6030: out = 16'(361);
			6031: out = 16'(-6566);
			6032: out = 16'(686);
			6033: out = 16'(2606);
			6034: out = 16'(4901);
			6035: out = 16'(8913);
			6036: out = 16'(4772);
			6037: out = 16'(620);
			6038: out = 16'(-5597);
			6039: out = 16'(1692);
			6040: out = 16'(12624);
			6041: out = 16'(15041);
			6042: out = 16'(7299);
			6043: out = 16'(-12044);
			6044: out = 16'(-6333);
			6045: out = 16'(-4477);
			6046: out = 16'(1939);
			6047: out = 16'(1447);
			6048: out = 16'(3890);
			6049: out = 16'(6789);
			6050: out = 16'(3770);
			6051: out = 16'(-13);
			6052: out = 16'(1400);
			6053: out = 16'(-3467);
			6054: out = 16'(-5227);
			6055: out = 16'(3581);
			6056: out = 16'(6489);
			6057: out = 16'(7030);
			6058: out = 16'(-5997);
			6059: out = 16'(-14967);
			6060: out = 16'(-24481);
			6061: out = 16'(-4127);
			6062: out = 16'(5215);
			6063: out = 16'(9475);
			6064: out = 16'(-896);
			6065: out = 16'(-7200);
			6066: out = 16'(-6103);
			6067: out = 16'(-6789);
			6068: out = 16'(-2431);
			6069: out = 16'(5715);
			6070: out = 16'(11328);
			6071: out = 16'(10945);
			6072: out = 16'(-14365);
			6073: out = 16'(-11625);
			6074: out = 16'(-3075);
			6075: out = 16'(7803);
			6076: out = 16'(5561);
			6077: out = 16'(-5616);
			6078: out = 16'(7100);
			6079: out = 16'(8719);
			6080: out = 16'(16093);
			6081: out = 16'(-9793);
			6082: out = 16'(-18050);
			6083: out = 16'(-25255);
			6084: out = 16'(5780);
			6085: out = 16'(17440);
			6086: out = 16'(10154);
			6087: out = 16'(-9877);
			6088: out = 16'(-23520);
			6089: out = 16'(-2525);
			6090: out = 16'(4358);
			6091: out = 16'(12561);
			6092: out = 16'(9332);
			6093: out = 16'(6765);
			6094: out = 16'(-209);
			6095: out = 16'(-7010);
			6096: out = 16'(-13737);
			6097: out = 16'(-18529);
			6098: out = 16'(4005);
			6099: out = 16'(13316);
			6100: out = 16'(15777);
			6101: out = 16'(-2043);
			6102: out = 16'(-10527);
			6103: out = 16'(-4177);
			6104: out = 16'(-1840);
			6105: out = 16'(3689);
			6106: out = 16'(5818);
			6107: out = 16'(9067);
			6108: out = 16'(7153);
			6109: out = 16'(-13165);
			6110: out = 16'(-7942);
			6111: out = 16'(2454);
			6112: out = 16'(10149);
			6113: out = 16'(9115);
			6114: out = 16'(1485);
			6115: out = 16'(6744);
			6116: out = 16'(4633);
			6117: out = 16'(4096);
			6118: out = 16'(-7038);
			6119: out = 16'(-8408);
			6120: out = 16'(-924);
			6121: out = 16'(-126);
			6122: out = 16'(608);
			6123: out = 16'(-6343);
			6124: out = 16'(970);
			6125: out = 16'(3814);
			6126: out = 16'(1997);
			6127: out = 16'(-1664);
			6128: out = 16'(-4168);
			6129: out = 16'(-4417);
			6130: out = 16'(-1297);
			6131: out = 16'(1447);
			6132: out = 16'(5473);
			6133: out = 16'(-667);
			6134: out = 16'(-11866);
			6135: out = 16'(-6359);
			6136: out = 16'(-3656);
			6137: out = 16'(-995);
			6138: out = 16'(1413);
			6139: out = 16'(2110);
			6140: out = 16'(3749);
			6141: out = 16'(-2509);
			6142: out = 16'(-4765);
			6143: out = 16'(-4380);
			6144: out = 16'(6962);
			6145: out = 16'(14356);
			6146: out = 16'(10546);
			6147: out = 16'(-4566);
			6148: out = 16'(-23111);
			6149: out = 16'(2640);
			6150: out = 16'(6813);
			6151: out = 16'(12877);
			6152: out = 16'(-7005);
			6153: out = 16'(-5747);
			6154: out = 16'(2036);
			6155: out = 16'(9905);
			6156: out = 16'(8915);
			6157: out = 16'(-323);
			6158: out = 16'(-7684);
			6159: out = 16'(-8160);
			6160: out = 16'(10317);
			6161: out = 16'(9058);
			6162: out = 16'(6724);
			6163: out = 16'(-17230);
			6164: out = 16'(-12865);
			6165: out = 16'(-5711);
			6166: out = 16'(14219);
			6167: out = 16'(11370);
			6168: out = 16'(3666);
			6169: out = 16'(-6132);
			6170: out = 16'(-5845);
			6171: out = 16'(2874);
			6172: out = 16'(-493);
			6173: out = 16'(2601);
			6174: out = 16'(6008);
			6175: out = 16'(4144);
			6176: out = 16'(68);
			6177: out = 16'(-7014);
			6178: out = 16'(-461);
			6179: out = 16'(3956);
			6180: out = 16'(-6835);
			6181: out = 16'(3673);
			6182: out = 16'(9489);
			6183: out = 16'(7951);
			6184: out = 16'(-1640);
			6185: out = 16'(-11733);
			6186: out = 16'(6522);
			6187: out = 16'(8028);
			6188: out = 16'(6699);
			6189: out = 16'(6285);
			6190: out = 16'(3051);
			6191: out = 16'(-2679);
			6192: out = 16'(-5694);
			6193: out = 16'(-9528);
			6194: out = 16'(-12927);
			6195: out = 16'(-9806);
			6196: out = 16'(-3706);
			6197: out = 16'(5813);
			6198: out = 16'(5909);
			6199: out = 16'(4030);
			6200: out = 16'(1567);
			6201: out = 16'(-2163);
			6202: out = 16'(-4177);
			6203: out = 16'(-653);
			6204: out = 16'(4085);
			6205: out = 16'(9298);
			6206: out = 16'(-4916);
			6207: out = 16'(-9577);
			6208: out = 16'(-13134);
			6209: out = 16'(1277);
			6210: out = 16'(5725);
			6211: out = 16'(3448);
			6212: out = 16'(2318);
			6213: out = 16'(-548);
			6214: out = 16'(-4154);
			6215: out = 16'(-2844);
			6216: out = 16'(360);
			6217: out = 16'(8314);
			6218: out = 16'(6029);
			6219: out = 16'(1553);
			6220: out = 16'(-13293);
			6221: out = 16'(-11108);
			6222: out = 16'(-3873);
			6223: out = 16'(2636);
			6224: out = 16'(-6);
			6225: out = 16'(-10850);
			6226: out = 16'(7582);
			6227: out = 16'(9935);
			6228: out = 16'(12482);
			6229: out = 16'(-10803);
			6230: out = 16'(-14576);
			6231: out = 16'(2421);
			6232: out = 16'(973);
			6233: out = 16'(1686);
			6234: out = 16'(-1680);
			6235: out = 16'(560);
			6236: out = 16'(-126);
			6237: out = 16'(-10674);
			6238: out = 16'(-8944);
			6239: out = 16'(-4382);
			6240: out = 16'(12548);
			6241: out = 16'(12179);
			6242: out = 16'(7779);
			6243: out = 16'(404);
			6244: out = 16'(-2725);
			6245: out = 16'(-4103);
			6246: out = 16'(4415);
			6247: out = 16'(6145);
			6248: out = 16'(5186);
			6249: out = 16'(-1703);
			6250: out = 16'(-5256);
			6251: out = 16'(-9162);
			6252: out = 16'(4237);
			6253: out = 16'(10471);
			6254: out = 16'(4107);
			6255: out = 16'(-3039);
			6256: out = 16'(-8148);
			6257: out = 16'(1746);
			6258: out = 16'(9121);
			6259: out = 16'(15408);
			6260: out = 16'(8453);
			6261: out = 16'(-4780);
			6262: out = 16'(-26156);
			6263: out = 16'(-2679);
			6264: out = 16'(6025);
			6265: out = 16'(16546);
			6266: out = 16'(-7837);
			6267: out = 16'(-13034);
			6268: out = 16'(-540);
			6269: out = 16'(445);
			6270: out = 16'(3136);
			6271: out = 16'(-2805);
			6272: out = 16'(5963);
			6273: out = 16'(8622);
			6274: out = 16'(4214);
			6275: out = 16'(2377);
			6276: out = 16'(1742);
			6277: out = 16'(-11470);
			6278: out = 16'(-6289);
			6279: out = 16'(776);
			6280: out = 16'(9431);
			6281: out = 16'(6651);
			6282: out = 16'(275);
			6283: out = 16'(-7280);
			6284: out = 16'(-6834);
			6285: out = 16'(-1874);
			6286: out = 16'(9663);
			6287: out = 16'(13457);
			6288: out = 16'(15021);
			6289: out = 16'(-9442);
			6290: out = 16'(-23468);
			6291: out = 16'(-10141);
			6292: out = 16'(2072);
			6293: out = 16'(12957);
			6294: out = 16'(-6068);
			6295: out = 16'(-6974);
			6296: out = 16'(-9891);
			6297: out = 16'(7444);
			6298: out = 16'(6390);
			6299: out = 16'(3675);
			6300: out = 16'(1583);
			6301: out = 16'(877);
			6302: out = 16'(-407);
			6303: out = 16'(-3902);
			6304: out = 16'(-6902);
			6305: out = 16'(-6465);
			6306: out = 16'(-7648);
			6307: out = 16'(-5330);
			6308: out = 16'(-3355);
			6309: out = 16'(3589);
			6310: out = 16'(5831);
			6311: out = 16'(712);
			6312: out = 16'(-4570);
			6313: out = 16'(-6912);
			6314: out = 16'(7083);
			6315: out = 16'(12808);
			6316: out = 16'(15894);
			6317: out = 16'(6110);
			6318: out = 16'(-4708);
			6319: out = 16'(-20636);
			6320: out = 16'(-504);
			6321: out = 16'(3615);
			6322: out = 16'(-700);
			6323: out = 16'(-2842);
			6324: out = 16'(-1384);
			6325: out = 16'(12922);
			6326: out = 16'(3184);
			6327: out = 16'(-2078);
			6328: out = 16'(-13456);
			6329: out = 16'(-1586);
			6330: out = 16'(6819);
			6331: out = 16'(4277);
			6332: out = 16'(-1995);
			6333: out = 16'(-9138);
			6334: out = 16'(-10914);
			6335: out = 16'(-5912);
			6336: out = 16'(2825);
			6337: out = 16'(5706);
			6338: out = 16'(2796);
			6339: out = 16'(-7440);
			6340: out = 16'(-1400);
			6341: out = 16'(2612);
			6342: out = 16'(8888);
			6343: out = 16'(4853);
			6344: out = 16'(1565);
			6345: out = 16'(966);
			6346: out = 16'(-2818);
			6347: out = 16'(-5307);
			6348: out = 16'(-21238);
			6349: out = 16'(-2429);
			6350: out = 16'(15963);
			6351: out = 16'(9411);
			6352: out = 16'(1730);
			6353: out = 16'(-12479);
			6354: out = 16'(5267);
			6355: out = 16'(5842);
			6356: out = 16'(6778);
			6357: out = 16'(-2479);
			6358: out = 16'(-1928);
			6359: out = 16'(4313);
			6360: out = 16'(1641);
			6361: out = 16'(3041);
			6362: out = 16'(11884);
			6363: out = 16'(3957);
			6364: out = 16'(-3702);
			6365: out = 16'(-20407);
			6366: out = 16'(-14649);
			6367: out = 16'(-5100);
			6368: out = 16'(5953);
			6369: out = 16'(8289);
			6370: out = 16'(6581);
			6371: out = 16'(1431);
			6372: out = 16'(157);
			6373: out = 16'(1574);
			6374: out = 16'(6166);
			6375: out = 16'(3115);
			6376: out = 16'(-10012);
			6377: out = 16'(-246);
			6378: out = 16'(526);
			6379: out = 16'(2459);
			6380: out = 16'(-8745);
			6381: out = 16'(-10339);
			6382: out = 16'(865);
			6383: out = 16'(6412);
			6384: out = 16'(10228);
			6385: out = 16'(13631);
			6386: out = 16'(5446);
			6387: out = 16'(-3445);
			6388: out = 16'(-8157);
			6389: out = 16'(-1136);
			6390: out = 16'(11631);
			6391: out = 16'(-46);
			6392: out = 16'(-1391);
			6393: out = 16'(-5218);
			6394: out = 16'(6244);
			6395: out = 16'(5032);
			6396: out = 16'(-3779);
			6397: out = 16'(1629);
			6398: out = 16'(3313);
			6399: out = 16'(49);
			6400: out = 16'(2082);
			6401: out = 16'(1121);
			6402: out = 16'(691);
			6403: out = 16'(-12337);
			6404: out = 16'(-21193);
			6405: out = 16'(3673);
			6406: out = 16'(9389);
			6407: out = 16'(14586);
			6408: out = 16'(-18390);
			6409: out = 16'(-19953);
			6410: out = 16'(-14668);
			6411: out = 16'(11299);
			6412: out = 16'(15064);
			6413: out = 16'(8669);
			6414: out = 16'(-7653);
			6415: out = 16'(-15074);
			6416: out = 16'(-10344);
			6417: out = 16'(-559);
			6418: out = 16'(6222);
			6419: out = 16'(-816);
			6420: out = 16'(971);
			6421: out = 16'(-1228);
			6422: out = 16'(-5889);
			6423: out = 16'(-4842);
			6424: out = 16'(-828);
			6425: out = 16'(6776);
			6426: out = 16'(4101);
			6427: out = 16'(-3261);
			6428: out = 16'(4901);
			6429: out = 16'(7136);
			6430: out = 16'(12253);
			6431: out = 16'(-3274);
			6432: out = 16'(-7696);
			6433: out = 16'(-8300);
			6434: out = 16'(-1111);
			6435: out = 16'(2314);
			6436: out = 16'(1591);
			6437: out = 16'(970);
			6438: out = 16'(425);
			6439: out = 16'(-114);
			6440: out = 16'(1870);
			6441: out = 16'(2579);
			6442: out = 16'(2023);
			6443: out = 16'(-5876);
			6444: out = 16'(-13959);
			6445: out = 16'(2332);
			6446: out = 16'(5896);
			6447: out = 16'(7543);
			6448: out = 16'(510);
			6449: out = 16'(-2543);
			6450: out = 16'(-3621);
			6451: out = 16'(-543);
			6452: out = 16'(4560);
			6453: out = 16'(11531);
			6454: out = 16'(11094);
			6455: out = 16'(7532);
			6456: out = 16'(-2804);
			6457: out = 16'(-4847);
			6458: out = 16'(-4493);
			6459: out = 16'(5729);
			6460: out = 16'(4124);
			6461: out = 16'(1724);
			6462: out = 16'(-2655);
			6463: out = 16'(-159);
			6464: out = 16'(5555);
			6465: out = 16'(-783);
			6466: out = 16'(3224);
			6467: out = 16'(8904);
			6468: out = 16'(8647);
			6469: out = 16'(757);
			6470: out = 16'(-19221);
			6471: out = 16'(-4961);
			6472: out = 16'(3486);
			6473: out = 16'(8662);
			6474: out = 16'(3453);
			6475: out = 16'(-1283);
			6476: out = 16'(2973);
			6477: out = 16'(-1010);
			6478: out = 16'(-2321);
			6479: out = 16'(-9446);
			6480: out = 16'(-3708);
			6481: out = 16'(1549);
			6482: out = 16'(10940);
			6483: out = 16'(637);
			6484: out = 16'(-17647);
			6485: out = 16'(-4402);
			6486: out = 16'(1837);
			6487: out = 16'(8335);
			6488: out = 16'(3099);
			6489: out = 16'(-1093);
			6490: out = 16'(-3942);
			6491: out = 16'(-9763);
			6492: out = 16'(-9536);
			6493: out = 16'(-2280);
			6494: out = 16'(6576);
			6495: out = 16'(11432);
			6496: out = 16'(8634);
			6497: out = 16'(-919);
			6498: out = 16'(-11422);
			6499: out = 16'(-6899);
			6500: out = 16'(-5274);
			6501: out = 16'(-524);
			6502: out = 16'(1484);
			6503: out = 16'(3180);
			6504: out = 16'(2046);
			6505: out = 16'(-2162);
			6506: out = 16'(-5719);
			6507: out = 16'(-6443);
			6508: out = 16'(-5506);
			6509: out = 16'(-696);
			6510: out = 16'(8566);
			6511: out = 16'(6609);
			6512: out = 16'(2084);
			6513: out = 16'(-13917);
			6514: out = 16'(-6568);
			6515: out = 16'(1514);
			6516: out = 16'(-4437);
			6517: out = 16'(-672);
			6518: out = 16'(1911);
			6519: out = 16'(1577);
			6520: out = 16'(814);
			6521: out = 16'(450);
			6522: out = 16'(9648);
			6523: out = 16'(9175);
			6524: out = 16'(-362);
			6525: out = 16'(5230);
			6526: out = 16'(1826);
			6527: out = 16'(-3623);
			6528: out = 16'(-9637);
			6529: out = 16'(-9591);
			6530: out = 16'(-4913);
			6531: out = 16'(7073);
			6532: out = 16'(13202);
			6533: out = 16'(4279);
			6534: out = 16'(-2771);
			6535: out = 16'(-10272);
			6536: out = 16'(-131);
			6537: out = 16'(1034);
			6538: out = 16'(3340);
			6539: out = 16'(5501);
			6540: out = 16'(2756);
			6541: out = 16'(-6948);
			6542: out = 16'(1931);
			6543: out = 16'(1594);
			6544: out = 16'(2180);
			6545: out = 16'(-9236);
			6546: out = 16'(-10408);
			6547: out = 16'(0);
			6548: out = 16'(4740);
			6549: out = 16'(7597);
			6550: out = 16'(4976);
			6551: out = 16'(2462);
			6552: out = 16'(-539);
			6553: out = 16'(-1371);
			6554: out = 16'(213);
			6555: out = 16'(2866);
			6556: out = 16'(1082);
			6557: out = 16'(-1041);
			6558: out = 16'(-4511);
			6559: out = 16'(-705);
			6560: out = 16'(2726);
			6561: out = 16'(8734);
			6562: out = 16'(2783);
			6563: out = 16'(-643);
			6564: out = 16'(-6127);
			6565: out = 16'(-1069);
			6566: out = 16'(3314);
			6567: out = 16'(11515);
			6568: out = 16'(1061);
			6569: out = 16'(-6563);
			6570: out = 16'(1554);
			6571: out = 16'(2644);
			6572: out = 16'(5078);
			6573: out = 16'(-20050);
			6574: out = 16'(-11641);
			6575: out = 16'(3352);
			6576: out = 16'(11542);
			6577: out = 16'(6999);
			6578: out = 16'(-9128);
			6579: out = 16'(-2830);
			6580: out = 16'(-523);
			6581: out = 16'(10943);
			6582: out = 16'(-3523);
			6583: out = 16'(-8146);
			6584: out = 16'(-15564);
			6585: out = 16'(3021);
			6586: out = 16'(11853);
			6587: out = 16'(7587);
			6588: out = 16'(-2765);
			6589: out = 16'(-11728);
			6590: out = 16'(-1582);
			6591: out = 16'(-787);
			6592: out = 16'(1280);
			6593: out = 16'(10113);
			6594: out = 16'(10714);
			6595: out = 16'(8209);
			6596: out = 16'(-4992);
			6597: out = 16'(-11193);
			6598: out = 16'(-14311);
			6599: out = 16'(-994);
			6600: out = 16'(6473);
			6601: out = 16'(10431);
			6602: out = 16'(-902);
			6603: out = 16'(-10142);
			6604: out = 16'(-18838);
			6605: out = 16'(-5390);
			6606: out = 16'(8574);
			6607: out = 16'(9000);
			6608: out = 16'(11183);
			6609: out = 16'(7183);
			6610: out = 16'(773);
			6611: out = 16'(-9015);
			6612: out = 16'(-17382);
			6613: out = 16'(-2428);
			6614: out = 16'(1482);
			6615: out = 16'(1513);
			6616: out = 16'(-3593);
			6617: out = 16'(-3720);
			6618: out = 16'(2432);
			6619: out = 16'(3089);
			6620: out = 16'(3861);
			6621: out = 16'(-375);
			6622: out = 16'(-1971);
			6623: out = 16'(-3017);
			6624: out = 16'(8204);
			6625: out = 16'(4201);
			6626: out = 16'(1651);
			6627: out = 16'(-15182);
			6628: out = 16'(-8197);
			6629: out = 16'(1700);
			6630: out = 16'(11575);
			6631: out = 16'(8132);
			6632: out = 16'(-644);
			6633: out = 16'(-6449);
			6634: out = 16'(-5242);
			6635: out = 16'(3691);
			6636: out = 16'(7601);
			6637: out = 16'(7206);
			6638: out = 16'(-3501);
			6639: out = 16'(-5844);
			6640: out = 16'(-7729);
			6641: out = 16'(1143);
			6642: out = 16'(-1177);
			6643: out = 16'(-958);
			6644: out = 16'(-4440);
			6645: out = 16'(668);
			6646: out = 16'(4156);
			6647: out = 16'(1036);
			6648: out = 16'(-1470);
			6649: out = 16'(-3717);
			6650: out = 16'(-903);
			6651: out = 16'(4311);
			6652: out = 16'(12170);
			6653: out = 16'(1590);
			6654: out = 16'(-4654);
			6655: out = 16'(-12911);
			6656: out = 16'(-2854);
			6657: out = 16'(2214);
			6658: out = 16'(127);
			6659: out = 16'(841);
			6660: out = 16'(810);
			6661: out = 16'(4370);
			6662: out = 16'(2529);
			6663: out = 16'(987);
			6664: out = 16'(578);
			6665: out = 16'(-1572);
			6666: out = 16'(-3957);
			6667: out = 16'(3193);
			6668: out = 16'(4815);
			6669: out = 16'(6316);
			6670: out = 16'(-3493);
			6671: out = 16'(-3874);
			6672: out = 16'(2078);
			6673: out = 16'(1880);
			6674: out = 16'(3997);
			6675: out = 16'(7170);
			6676: out = 16'(4167);
			6677: out = 16'(1090);
			6678: out = 16'(-3042);
			6679: out = 16'(561);
			6680: out = 16'(4067);
			6681: out = 16'(2100);
			6682: out = 16'(-1227);
			6683: out = 16'(-6136);
			6684: out = 16'(7842);
			6685: out = 16'(4061);
			6686: out = 16'(-627);
			6687: out = 16'(-6431);
			6688: out = 16'(-7161);
			6689: out = 16'(-7277);
			6690: out = 16'(6627);
			6691: out = 16'(11558);
			6692: out = 16'(14403);
			6693: out = 16'(-3003);
			6694: out = 16'(-11435);
			6695: out = 16'(-8578);
			6696: out = 16'(-1491);
			6697: out = 16'(4716);
			6698: out = 16'(3073);
			6699: out = 16'(1839);
			6700: out = 16'(-1062);
			6701: out = 16'(-4165);
			6702: out = 16'(-2104);
			6703: out = 16'(2114);
			6704: out = 16'(8961);
			6705: out = 16'(7265);
			6706: out = 16'(1035);
			6707: out = 16'(-6464);
			6708: out = 16'(-7452);
			6709: out = 16'(435);
			6710: out = 16'(1599);
			6711: out = 16'(3760);
			6712: out = 16'(-397);
			6713: out = 16'(-126);
			6714: out = 16'(-4476);
			6715: out = 16'(-9102);
			6716: out = 16'(-8022);
			6717: out = 16'(-1870);
			6718: out = 16'(-1199);
			6719: out = 16'(7481);
			6720: out = 16'(9004);
			6721: out = 16'(12474);
			6722: out = 16'(-5221);
			6723: out = 16'(-24891);
			6724: out = 16'(-19860);
			6725: out = 16'(-7049);
			6726: out = 16'(10612);
			6727: out = 16'(14258);
			6728: out = 16'(7642);
			6729: out = 16'(-10057);
			6730: out = 16'(-20729);
			6731: out = 16'(-19676);
			6732: out = 16'(7594);
			6733: out = 16'(10268);
			6734: out = 16'(11806);
			6735: out = 16'(-1467);
			6736: out = 16'(158);
			6737: out = 16'(-779);
			6738: out = 16'(-11596);
			6739: out = 16'(-8591);
			6740: out = 16'(-2020);
			6741: out = 16'(8407);
			6742: out = 16'(6692);
			6743: out = 16'(-661);
			6744: out = 16'(-2867);
			6745: out = 16'(-448);
			6746: out = 16'(8628);
			6747: out = 16'(7199);
			6748: out = 16'(6358);
			6749: out = 16'(557);
			6750: out = 16'(2781);
			6751: out = 16'(96);
			6752: out = 16'(-10944);
			6753: out = 16'(-12066);
			6754: out = 16'(-9173);
			6755: out = 16'(15495);
			6756: out = 16'(11528);
			6757: out = 16'(6115);
			6758: out = 16'(-26263);
			6759: out = 16'(-14564);
			6760: out = 16'(9789);
			6761: out = 16'(19421);
			6762: out = 16'(9015);
			6763: out = 16'(-22249);
			6764: out = 16'(-3375);
			6765: out = 16'(1794);
			6766: out = 16'(13720);
			6767: out = 16'(-6285);
			6768: out = 16'(-10921);
			6769: out = 16'(-2143);
			6770: out = 16'(1059);
			6771: out = 16'(4196);
			6772: out = 16'(4998);
			6773: out = 16'(9814);
			6774: out = 16'(10294);
			6775: out = 16'(-16898);
			6776: out = 16'(-15622);
			6777: out = 16'(-8131);
			6778: out = 16'(13665);
			6779: out = 16'(12054);
			6780: out = 16'(-606);
			6781: out = 16'(3307);
			6782: out = 16'(-1521);
			6783: out = 16'(-4583);
			6784: out = 16'(-8041);
			6785: out = 16'(-5309);
			6786: out = 16'(619);
			6787: out = 16'(908);
			6788: out = 16'(3022);
			6789: out = 16'(16774);
			6790: out = 16'(6721);
			6791: out = 16'(-1031);
			6792: out = 16'(-20284);
			6793: out = 16'(-8006);
			6794: out = 16'(6301);
			6795: out = 16'(7481);
			6796: out = 16'(-1193);
			6797: out = 16'(-16815);
			6798: out = 16'(-2294);
			6799: out = 16'(987);
			6800: out = 16'(5331);
			6801: out = 16'(5861);
			6802: out = 16'(6049);
			6803: out = 16'(1116);
			6804: out = 16'(2273);
			6805: out = 16'(1235);
			6806: out = 16'(5151);
			6807: out = 16'(-2275);
			6808: out = 16'(-5525);
			6809: out = 16'(-8669);
			6810: out = 16'(3745);
			6811: out = 16'(12389);
			6812: out = 16'(-10081);
			6813: out = 16'(-5723);
			6814: out = 16'(1791);
			6815: out = 16'(9129);
			6816: out = 16'(10308);
			6817: out = 16'(6322);
			6818: out = 16'(6690);
			6819: out = 16'(-1033);
			6820: out = 16'(-12956);
			6821: out = 16'(-5741);
			6822: out = 16'(-906);
			6823: out = 16'(-784);
			6824: out = 16'(4332);
			6825: out = 16'(4618);
			6826: out = 16'(6177);
			6827: out = 16'(-3326);
			6828: out = 16'(-7999);
			6829: out = 16'(-6432);
			6830: out = 16'(5765);
			6831: out = 16'(16247);
			6832: out = 16'(11768);
			6833: out = 16'(4786);
			6834: out = 16'(-5737);
			6835: out = 16'(-5227);
			6836: out = 16'(-3896);
			6837: out = 16'(1572);
			6838: out = 16'(1833);
			6839: out = 16'(2664);
			6840: out = 16'(2365);
			6841: out = 16'(-1183);
			6842: out = 16'(-5352);
			6843: out = 16'(-14801);
			6844: out = 16'(-3076);
			6845: out = 16'(6952);
			6846: out = 16'(16074);
			6847: out = 16'(4877);
			6848: out = 16'(-8154);
			6849: out = 16'(-7282);
			6850: out = 16'(-7642);
			6851: out = 16'(-2835);
			6852: out = 16'(-4033);
			6853: out = 16'(648);
			6854: out = 16'(3856);
			6855: out = 16'(3378);
			6856: out = 16'(1155);
			6857: out = 16'(-1329);
			6858: out = 16'(-882);
			6859: out = 16'(2261);
			6860: out = 16'(9675);
			6861: out = 16'(1331);
			6862: out = 16'(-4031);
			6863: out = 16'(-2413);
			6864: out = 16'(-941);
			6865: out = 16'(511);
			6866: out = 16'(-15859);
			6867: out = 16'(-10267);
			6868: out = 16'(-3751);
			6869: out = 16'(7635);
			6870: out = 16'(9392);
			6871: out = 16'(10323);
			6872: out = 16'(-11884);
			6873: out = 16'(-13905);
			6874: out = 16'(-8840);
			6875: out = 16'(12814);
			6876: out = 16'(12651);
			6877: out = 16'(-8073);
			6878: out = 16'(-11925);
			6879: out = 16'(-13474);
			6880: out = 16'(1971);
			6881: out = 16'(610);
			6882: out = 16'(2281);
			6883: out = 16'(-1351);
			6884: out = 16'(-877);
			6885: out = 16'(-2416);
			6886: out = 16'(689);
			6887: out = 16'(5184);
			6888: out = 16'(12922);
			6889: out = 16'(-8052);
			6890: out = 16'(-2975);
			6891: out = 16'(5787);
			6892: out = 16'(11003);
			6893: out = 16'(1600);
			6894: out = 16'(-21535);
			6895: out = 16'(-12358);
			6896: out = 16'(-4559);
			6897: out = 16'(5813);
			6898: out = 16'(10405);
			6899: out = 16'(10769);
			6900: out = 16'(3447);
			6901: out = 16'(-2284);
			6902: out = 16'(-5743);
			6903: out = 16'(6602);
			6904: out = 16'(4695);
			6905: out = 16'(2769);
			6906: out = 16'(1882);
			6907: out = 16'(3381);
			6908: out = 16'(6333);
			6909: out = 16'(-11170);
			6910: out = 16'(-10825);
			6911: out = 16'(-1253);
			6912: out = 16'(4003);
			6913: out = 16'(7528);
			6914: out = 16'(5870);
			6915: out = 16'(5315);
			6916: out = 16'(2626);
			6917: out = 16'(179);
			6918: out = 16'(1251);
			6919: out = 16'(3705);
			6920: out = 16'(5594);
			6921: out = 16'(5295);
			6922: out = 16'(1757);
			6923: out = 16'(-6737);
			6924: out = 16'(-12575);
			6925: out = 16'(-14432);
			6926: out = 16'(3921);
			6927: out = 16'(9930);
			6928: out = 16'(9733);
			6929: out = 16'(9555);
			6930: out = 16'(4769);
			6931: out = 16'(-413);
			6932: out = 16'(-4789);
			6933: out = 16'(-5363);
			6934: out = 16'(-4830);
			6935: out = 16'(4333);
			6936: out = 16'(7261);
			6937: out = 16'(103);
			6938: out = 16'(-8063);
			6939: out = 16'(-13825);
			6940: out = 16'(3792);
			6941: out = 16'(4326);
			6942: out = 16'(6137);
			6943: out = 16'(-8150);
			6944: out = 16'(-2429);
			6945: out = 16'(5624);
			6946: out = 16'(9914);
			6947: out = 16'(4120);
			6948: out = 16'(-9866);
			6949: out = 16'(-1772);
			6950: out = 16'(-157);
			6951: out = 16'(87);
			6952: out = 16'(-211);
			6953: out = 16'(-429);
			6954: out = 16'(-210);
			6955: out = 16'(-1269);
			6956: out = 16'(-1294);
			6957: out = 16'(-676);
			6958: out = 16'(3382);
			6959: out = 16'(5742);
			6960: out = 16'(196);
			6961: out = 16'(-3486);
			6962: out = 16'(-7144);
			6963: out = 16'(488);
			6964: out = 16'(1891);
			6965: out = 16'(2433);
			6966: out = 16'(-6282);
			6967: out = 16'(-6411);
			6968: out = 16'(2329);
			6969: out = 16'(-2756);
			6970: out = 16'(-1194);
			6971: out = 16'(-540);
			6972: out = 16'(8582);
			6973: out = 16'(10037);
			6974: out = 16'(4280);
			6975: out = 16'(-2785);
			6976: out = 16'(-8242);
			6977: out = 16'(-12730);
			6978: out = 16'(-8993);
			6979: out = 16'(-3502);
			6980: out = 16'(13588);
			6981: out = 16'(6885);
			6982: out = 16'(-5642);
			6983: out = 16'(-15147);
			6984: out = 16'(-8631);
			6985: out = 16'(13470);
			6986: out = 16'(4807);
			6987: out = 16'(7123);
			6988: out = 16'(7706);
			6989: out = 16'(5171);
			6990: out = 16'(981);
			6991: out = 16'(2363);
			6992: out = 16'(-3081);
			6993: out = 16'(-4010);
			6994: out = 16'(-6565);
			6995: out = 16'(1488);
			6996: out = 16'(5975);
			6997: out = 16'(3434);
			6998: out = 16'(-4622);
			6999: out = 16'(-13150);
			7000: out = 16'(-5404);
			7001: out = 16'(2193);
			7002: out = 16'(12518);
			7003: out = 16'(2877);
			7004: out = 16'(-1324);
			7005: out = 16'(-9252);
			7006: out = 16'(1463);
			7007: out = 16'(2326);
			7008: out = 16'(-4239);
			7009: out = 16'(-4097);
			7010: out = 16'(-2968);
			7011: out = 16'(1110);
			7012: out = 16'(2982);
			7013: out = 16'(3954);
			7014: out = 16'(1191);
			7015: out = 16'(1386);
			7016: out = 16'(1748);
			7017: out = 16'(4700);
			7018: out = 16'(4087);
			7019: out = 16'(2003);
			7020: out = 16'(1691);
			7021: out = 16'(-2682);
			7022: out = 16'(-8748);
			7023: out = 16'(-2386);
			7024: out = 16'(2694);
			7025: out = 16'(8430);
			7026: out = 16'(7587);
			7027: out = 16'(4178);
			7028: out = 16'(-7635);
			7029: out = 16'(369);
			7030: out = 16'(6312);
			7031: out = 16'(9757);
			7032: out = 16'(3928);
			7033: out = 16'(-3352);
			7034: out = 16'(1420);
			7035: out = 16'(-881);
			7036: out = 16'(-8);
			7037: out = 16'(-12770);
			7038: out = 16'(-6261);
			7039: out = 16'(4350);
			7040: out = 16'(10953);
			7041: out = 16'(7347);
			7042: out = 16'(-4076);
			7043: out = 16'(-10481);
			7044: out = 16'(-9195);
			7045: out = 16'(8197);
			7046: out = 16'(3925);
			7047: out = 16'(2401);
			7048: out = 16'(-6550);
			7049: out = 16'(121);
			7050: out = 16'(2451);
			7051: out = 16'(-8025);
			7052: out = 16'(-9363);
			7053: out = 16'(-8363);
			7054: out = 16'(6707);
			7055: out = 16'(7324);
			7056: out = 16'(4203);
			7057: out = 16'(3365);
			7058: out = 16'(-1724);
			7059: out = 16'(-10407);
			7060: out = 16'(6185);
			7061: out = 16'(10233);
			7062: out = 16'(7713);
			7063: out = 16'(-2344);
			7064: out = 16'(-7703);
			7065: out = 16'(-929);
			7066: out = 16'(-3446);
			7067: out = 16'(-1950);
			7068: out = 16'(74);
			7069: out = 16'(2846);
			7070: out = 16'(3077);
			7071: out = 16'(1349);
			7072: out = 16'(-834);
			7073: out = 16'(-1795);
			7074: out = 16'(-3208);
			7075: out = 16'(-3207);
			7076: out = 16'(-4536);
			7077: out = 16'(6440);
			7078: out = 16'(5301);
			7079: out = 16'(-2269);
			7080: out = 16'(-9603);
			7081: out = 16'(-11571);
			7082: out = 16'(-1917);
			7083: out = 16'(96);
			7084: out = 16'(3061);
			7085: out = 16'(-5369);
			7086: out = 16'(5395);
			7087: out = 16'(9828);
			7088: out = 16'(4626);
			7089: out = 16'(-3038);
			7090: out = 16'(-10133);
			7091: out = 16'(-2040);
			7092: out = 16'(-1448);
			7093: out = 16'(-1189);
			7094: out = 16'(893);
			7095: out = 16'(4481);
			7096: out = 16'(11040);
			7097: out = 16'(-451);
			7098: out = 16'(-2297);
			7099: out = 16'(-105);
			7100: out = 16'(8129);
			7101: out = 16'(9076);
			7102: out = 16'(-2199);
			7103: out = 16'(-2599);
			7104: out = 16'(-2743);
			7105: out = 16'(299);
			7106: out = 16'(6316);
			7107: out = 16'(9901);
			7108: out = 16'(-8779);
			7109: out = 16'(-10863);
			7110: out = 16'(-10778);
			7111: out = 16'(3987);
			7112: out = 16'(2358);
			7113: out = 16'(-6676);
			7114: out = 16'(3321);
			7115: out = 16'(6699);
			7116: out = 16'(12740);
			7117: out = 16'(-7414);
			7118: out = 16'(-15707);
			7119: out = 16'(-13842);
			7120: out = 16'(-5757);
			7121: out = 16'(3229);
			7122: out = 16'(9636);
			7123: out = 16'(7168);
			7124: out = 16'(1759);
			7125: out = 16'(-3074);
			7126: out = 16'(-4315);
			7127: out = 16'(-1977);
			7128: out = 16'(-2522);
			7129: out = 16'(2698);
			7130: out = 16'(7347);
			7131: out = 16'(7160);
			7132: out = 16'(4054);
			7133: out = 16'(-2416);
			7134: out = 16'(2725);
			7135: out = 16'(2663);
			7136: out = 16'(1064);
			7137: out = 16'(-2889);
			7138: out = 16'(-3751);
			7139: out = 16'(1410);
			7140: out = 16'(-185);
			7141: out = 16'(-79);
			7142: out = 16'(2107);
			7143: out = 16'(2294);
			7144: out = 16'(1952);
			7145: out = 16'(826);
			7146: out = 16'(-661);
			7147: out = 16'(-2033);
			7148: out = 16'(418);
			7149: out = 16'(-384);
			7150: out = 16'(-1991);
			7151: out = 16'(27);
			7152: out = 16'(1939);
			7153: out = 16'(4578);
			7154: out = 16'(2787);
			7155: out = 16'(-156);
			7156: out = 16'(-7750);
			7157: out = 16'(-3635);
			7158: out = 16'(-1126);
			7159: out = 16'(983);
			7160: out = 16'(2386);
			7161: out = 16'(1720);
			7162: out = 16'(-15647);
			7163: out = 16'(-8267);
			7164: out = 16'(1954);
			7165: out = 16'(9448);
			7166: out = 16'(12396);
			7167: out = 16'(11724);
			7168: out = 16'(-348);
			7169: out = 16'(-8175);
			7170: out = 16'(-16245);
			7171: out = 16'(5978);
			7172: out = 16'(12490);
			7173: out = 16'(8983);
			7174: out = 16'(939);
			7175: out = 16'(-4222);
			7176: out = 16'(325);
			7177: out = 16'(-590);
			7178: out = 16'(77);
			7179: out = 16'(-6664);
			7180: out = 16'(-2718);
			7181: out = 16'(-673);
			7182: out = 16'(819);
			7183: out = 16'(-2619);
			7184: out = 16'(-5926);
			7185: out = 16'(-2546);
			7186: out = 16'(1638);
			7187: out = 16'(7351);
			7188: out = 16'(2659);
			7189: out = 16'(707);
			7190: out = 16'(-3977);
			7191: out = 16'(96);
			7192: out = 16'(1200);
			7193: out = 16'(6634);
			7194: out = 16'(-7436);
			7195: out = 16'(-12403);
			7196: out = 16'(-5928);
			7197: out = 16'(1113);
			7198: out = 16'(7039);
			7199: out = 16'(7531);
			7200: out = 16'(6360);
			7201: out = 16'(2857);
			7202: out = 16'(-8520);
			7203: out = 16'(-9298);
			7204: out = 16'(-6246);
			7205: out = 16'(1784);
			7206: out = 16'(5035);
			7207: out = 16'(6980);
			7208: out = 16'(-3480);
			7209: out = 16'(-3435);
			7210: out = 16'(3817);
			7211: out = 16'(9582);
			7212: out = 16'(8928);
			7213: out = 16'(-3765);
			7214: out = 16'(-7190);
			7215: out = 16'(-9207);
			7216: out = 16'(1032);
			7217: out = 16'(1113);
			7218: out = 16'(2286);
			7219: out = 16'(-4591);
			7220: out = 16'(-1412);
			7221: out = 16'(1029);
			7222: out = 16'(-2454);
			7223: out = 16'(-2341);
			7224: out = 16'(236);
			7225: out = 16'(1425);
			7226: out = 16'(2593);
			7227: out = 16'(11);
			7228: out = 16'(2771);
			7229: out = 16'(1112);
			7230: out = 16'(2064);
			7231: out = 16'(-7984);
			7232: out = 16'(-9863);
			7233: out = 16'(-4993);
			7234: out = 16'(6192);
			7235: out = 16'(11598);
			7236: out = 16'(4096);
			7237: out = 16'(-2672);
			7238: out = 16'(-8911);
			7239: out = 16'(-4700);
			7240: out = 16'(-1578);
			7241: out = 16'(1951);
			7242: out = 16'(11941);
			7243: out = 16'(6522);
			7244: out = 16'(-6955);
			7245: out = 16'(-7735);
			7246: out = 16'(-3766);
			7247: out = 16'(11389);
			7248: out = 16'(1714);
			7249: out = 16'(759);
			7250: out = 16'(7098);
			7251: out = 16'(2792);
			7252: out = 16'(-2398);
			7253: out = 16'(-19022);
			7254: out = 16'(-10463);
			7255: out = 16'(33);
			7256: out = 16'(12038);
			7257: out = 16'(7827);
			7258: out = 16'(-503);
			7259: out = 16'(-6836);
			7260: out = 16'(-5890);
			7261: out = 16'(1190);
			7262: out = 16'(57);
			7263: out = 16'(2239);
			7264: out = 16'(3542);
			7265: out = 16'(3574);
			7266: out = 16'(3000);
			7267: out = 16'(304);
			7268: out = 16'(4459);
			7269: out = 16'(4552);
			7270: out = 16'(939);
			7271: out = 16'(-2135);
			7272: out = 16'(-3499);
			7273: out = 16'(-9545);
			7274: out = 16'(3386);
			7275: out = 16'(14521);
			7276: out = 16'(11245);
			7277: out = 16'(-2068);
			7278: out = 16'(-22916);
			7279: out = 16'(-1394);
			7280: out = 16'(4378);
			7281: out = 16'(12927);
			7282: out = 16'(-5346);
			7283: out = 16'(-6238);
			7284: out = 16'(1043);
			7285: out = 16'(6004);
			7286: out = 16'(5334);
			7287: out = 16'(-4774);
			7288: out = 16'(-8674);
			7289: out = 16'(-10535);
			7290: out = 16'(184);
			7291: out = 16'(44);
			7292: out = 16'(927);
			7293: out = 16'(-11356);
			7294: out = 16'(-2272);
			7295: out = 16'(7678);
			7296: out = 16'(981);
			7297: out = 16'(-5575);
			7298: out = 16'(-16214);
			7299: out = 16'(3416);
			7300: out = 16'(8239);
			7301: out = 16'(7943);
			7302: out = 16'(3244);
			7303: out = 16'(517);
			7304: out = 16'(1630);
			7305: out = 16'(-4416);
			7306: out = 16'(-6331);
			7307: out = 16'(531);
			7308: out = 16'(-2007);
			7309: out = 16'(-2242);
			7310: out = 16'(-900);
			7311: out = 16'(5355);
			7312: out = 16'(9529);
			7313: out = 16'(-5637);
			7314: out = 16'(-5572);
			7315: out = 16'(-1954);
			7316: out = 16'(4393);
			7317: out = 16'(4260);
			7318: out = 16'(-2769);
			7319: out = 16'(6316);
			7320: out = 16'(4266);
			7321: out = 16'(25);
			7322: out = 16'(-10801);
			7323: out = 16'(-9962);
			7324: out = 16'(8614);
			7325: out = 16'(7305);
			7326: out = 16'(5204);
			7327: out = 16'(-3885);
			7328: out = 16'(-5960);
			7329: out = 16'(-6571);
			7330: out = 16'(-3423);
			7331: out = 16'(-37);
			7332: out = 16'(3113);
			7333: out = 16'(6684);
			7334: out = 16'(4840);
			7335: out = 16'(693);
			7336: out = 16'(-997);
			7337: out = 16'(-2198);
			7338: out = 16'(-3051);
			7339: out = 16'(5315);
			7340: out = 16'(8124);
			7341: out = 16'(6570);
			7342: out = 16'(2184);
			7343: out = 16'(-2011);
			7344: out = 16'(-7324);
			7345: out = 16'(-1864);
			7346: out = 16'(3595);
			7347: out = 16'(7416);
			7348: out = 16'(4273);
			7349: out = 16'(-733);
			7350: out = 16'(-3941);
			7351: out = 16'(-3890);
			7352: out = 16'(-1358);
			7353: out = 16'(3309);
			7354: out = 16'(3424);
			7355: out = 16'(-130);
			7356: out = 16'(-2115);
			7357: out = 16'(-4468);
			7358: out = 16'(-5710);
			7359: out = 16'(-2321);
			7360: out = 16'(3205);
			7361: out = 16'(13920);
			7362: out = 16'(4908);
			7363: out = 16'(-3954);
			7364: out = 16'(-16902);
			7365: out = 16'(-11321);
			7366: out = 16'(-2121);
			7367: out = 16'(-597);
			7368: out = 16'(3135);
			7369: out = 16'(3143);
			7370: out = 16'(4149);
			7371: out = 16'(1993);
			7372: out = 16'(1054);
			7373: out = 16'(2568);
			7374: out = 16'(2884);
			7375: out = 16'(-1606);
			7376: out = 16'(6628);
			7377: out = 16'(5701);
			7378: out = 16'(2680);
			7379: out = 16'(-11359);
			7380: out = 16'(-15896);
			7381: out = 16'(-209);
			7382: out = 16'(-177);
			7383: out = 16'(1719);
			7384: out = 16'(4126);
			7385: out = 16'(7875);
			7386: out = 16'(9304);
			7387: out = 16'(-15233);
			7388: out = 16'(-15962);
			7389: out = 16'(-11258);
			7390: out = 16'(10391);
			7391: out = 16'(12145);
			7392: out = 16'(6033);
			7393: out = 16'(-9264);
			7394: out = 16'(-12191);
			7395: out = 16'(-359);
			7396: out = 16'(4787);
			7397: out = 16'(5963);
			7398: out = 16'(-11011);
			7399: out = 16'(-2823);
			7400: out = 16'(130);
			7401: out = 16'(3125);
			7402: out = 16'(-1245);
			7403: out = 16'(-3941);
			7404: out = 16'(-338);
			7405: out = 16'(-97);
			7406: out = 16'(-181);
			7407: out = 16'(-1325);
			7408: out = 16'(199);
			7409: out = 16'(3152);
			7410: out = 16'(4373);
			7411: out = 16'(3396);
			7412: out = 16'(-2289);
			7413: out = 16'(4676);
			7414: out = 16'(5244);
			7415: out = 16'(3745);
			7416: out = 16'(650);
			7417: out = 16'(-780);
			7418: out = 16'(-2045);
			7419: out = 16'(-96);
			7420: out = 16'(1523);
			7421: out = 16'(9222);
			7422: out = 16'(2956);
			7423: out = 16'(-3442);
			7424: out = 16'(-16489);
			7425: out = 16'(-9384);
			7426: out = 16'(4530);
			7427: out = 16'(7542);
			7428: out = 16'(4935);
			7429: out = 16'(-7321);
			7430: out = 16'(407);
			7431: out = 16'(2619);
			7432: out = 16'(11402);
			7433: out = 16'(-1424);
			7434: out = 16'(-3692);
			7435: out = 16'(-2695);
			7436: out = 16'(8981);
			7437: out = 16'(10563);
			7438: out = 16'(-9398);
			7439: out = 16'(-13359);
			7440: out = 16'(-14696);
			7441: out = 16'(-796);
			7442: out = 16'(170);
			7443: out = 16'(454);
			7444: out = 16'(9174);
			7445: out = 16'(9015);
			7446: out = 16'(6203);
			7447: out = 16'(-2254);
			7448: out = 16'(-3540);
			7449: out = 16'(1354);
			7450: out = 16'(4236);
			7451: out = 16'(2427);
			7452: out = 16'(-12781);
			7453: out = 16'(-4128);
			7454: out = 16'(152);
			7455: out = 16'(11039);
			7456: out = 16'(1332);
			7457: out = 16'(-3621);
			7458: out = 16'(-7922);
			7459: out = 16'(1800);
			7460: out = 16'(9523);
			7461: out = 16'(11364);
			7462: out = 16'(1588);
			7463: out = 16'(-11271);
			7464: out = 16'(-8816);
			7465: out = 16'(-5116);
			7466: out = 16'(1714);
			7467: out = 16'(3130);
			7468: out = 16'(2212);
			7469: out = 16'(-249);
			7470: out = 16'(-8666);
			7471: out = 16'(-8408);
			7472: out = 16'(2435);
			7473: out = 16'(8987);
			7474: out = 16'(10480);
			7475: out = 16'(1259);
			7476: out = 16'(-6771);
			7477: out = 16'(-12965);
			7478: out = 16'(-7240);
			7479: out = 16'(-2990);
			7480: out = 16'(2194);
			7481: out = 16'(7449);
			7482: out = 16'(8457);
			7483: out = 16'(8725);
			7484: out = 16'(-10295);
			7485: out = 16'(-12829);
			7486: out = 16'(-7709);
			7487: out = 16'(8109);
			7488: out = 16'(13924);
			7489: out = 16'(12959);
			7490: out = 16'(-1331);
			7491: out = 16'(-11202);
			7492: out = 16'(-17445);
			7493: out = 16'(-2206);
			7494: out = 16'(10282);
			7495: out = 16'(8697);
			7496: out = 16'(2105);
			7497: out = 16'(-7566);
			7498: out = 16'(-14504);
			7499: out = 16'(-5553);
			7500: out = 16'(11794);
			7501: out = 16'(5253);
			7502: out = 16'(3748);
			7503: out = 16'(-5630);
			7504: out = 16'(5089);
			7505: out = 16'(5529);
			7506: out = 16'(7790);
			7507: out = 16'(-3555);
			7508: out = 16'(-6783);
			7509: out = 16'(-4362);
			7510: out = 16'(-837);
			7511: out = 16'(985);
			7512: out = 16'(-217);
			7513: out = 16'(-415);
			7514: out = 16'(-285);
			7515: out = 16'(-2964);
			7516: out = 16'(-1851);
			7517: out = 16'(-1132);
			7518: out = 16'(8560);
			7519: out = 16'(5689);
			7520: out = 16'(296);
			7521: out = 16'(-11412);
			7522: out = 16'(-10368);
			7523: out = 16'(1410);
			7524: out = 16'(1490);
			7525: out = 16'(3240);
			7526: out = 16'(2403);
			7527: out = 16'(254);
			7528: out = 16'(-2226);
			7529: out = 16'(-4009);
			7530: out = 16'(2438);
			7531: out = 16'(7548);
			7532: out = 16'(709);
			7533: out = 16'(-917);
			7534: out = 16'(-4420);
			7535: out = 16'(7503);
			7536: out = 16'(-1875);
			7537: out = 16'(-14599);
			7538: out = 16'(-626);
			7539: out = 16'(3481);
			7540: out = 16'(6251);
			7541: out = 16'(-1698);
			7542: out = 16'(-3436);
			7543: out = 16'(910);
			7544: out = 16'(-410);
			7545: out = 16'(107);
			7546: out = 16'(-1872);
			7547: out = 16'(2295);
			7548: out = 16'(4359);
			7549: out = 16'(7346);
			7550: out = 16'(4967);
			7551: out = 16'(1924);
			7552: out = 16'(-16084);
			7553: out = 16'(-10933);
			7554: out = 16'(-845);
			7555: out = 16'(6825);
			7556: out = 16'(5352);
			7557: out = 16'(-2433);
			7558: out = 16'(-2074);
			7559: out = 16'(92);
			7560: out = 16'(9412);
			7561: out = 16'(1373);
			7562: out = 16'(767);
			7563: out = 16'(2076);
			7564: out = 16'(5198);
			7565: out = 16'(2273);
			7566: out = 16'(-15687);
			7567: out = 16'(-9545);
			7568: out = 16'(-1025);
			7569: out = 16'(8858);
			7570: out = 16'(12283);
			7571: out = 16'(11751);
			7572: out = 16'(1996);
			7573: out = 16'(633);
			7574: out = 16'(2492);
			7575: out = 16'(319);
			7576: out = 16'(-42);
			7577: out = 16'(-2606);
			7578: out = 16'(5288);
			7579: out = 16'(4461);
			7580: out = 16'(-1045);
			7581: out = 16'(-4681);
			7582: out = 16'(-4976);
			7583: out = 16'(1087);
			7584: out = 16'(-151);
			7585: out = 16'(401);
			7586: out = 16'(5528);
			7587: out = 16'(2857);
			7588: out = 16'(-904);
			7589: out = 16'(-11944);
			7590: out = 16'(-13361);
			7591: out = 16'(-11257);
			7592: out = 16'(8226);
			7593: out = 16'(11164);
			7594: out = 16'(9084);
			7595: out = 16'(-5027);
			7596: out = 16'(-8390);
			7597: out = 16'(-3696);
			7598: out = 16'(1937);
			7599: out = 16'(4346);
			7600: out = 16'(-905);
			7601: out = 16'(-2227);
			7602: out = 16'(-5938);
			7603: out = 16'(-7952);
			7604: out = 16'(-3648);
			7605: out = 16'(2613);
			7606: out = 16'(189);
			7607: out = 16'(2374);
			7608: out = 16'(334);
			7609: out = 16'(10042);
			7610: out = 16'(2181);
			7611: out = 16'(-4617);
			7612: out = 16'(-16373);
			7613: out = 16'(-9995);
			7614: out = 16'(3734);
			7615: out = 16'(12208);
			7616: out = 16'(10305);
			7617: out = 16'(-409);
			7618: out = 16'(-10982);
			7619: out = 16'(-13285);
			7620: out = 16'(778);
			7621: out = 16'(8407);
			7622: out = 16'(10600);
			7623: out = 16'(-14401);
			7624: out = 16'(-10299);
			7625: out = 16'(-6851);
			7626: out = 16'(2541);
			7627: out = 16'(2264);
			7628: out = 16'(1527);
			7629: out = 16'(3958);
			7630: out = 16'(2168);
			7631: out = 16'(-1829);
			7632: out = 16'(-1994);
			7633: out = 16'(-2461);
			7634: out = 16'(-753);
			7635: out = 16'(364);
			7636: out = 16'(1695);
			7637: out = 16'(-7);
			7638: out = 16'(2522);
			7639: out = 16'(2775);
			7640: out = 16'(4485);
			7641: out = 16'(397);
			7642: out = 16'(-1317);
			7643: out = 16'(-1843);
			7644: out = 16'(3469);
			7645: out = 16'(7129);
			7646: out = 16'(1917);
			7647: out = 16'(402);
			7648: out = 16'(-411);
			7649: out = 16'(-7764);
			7650: out = 16'(-2291);
			7651: out = 16'(9514);
			7652: out = 16'(8441);
			7653: out = 16'(6845);
			7654: out = 16'(-1592);
			7655: out = 16'(1137);
			7656: out = 16'(-47);
			7657: out = 16'(1439);
			7658: out = 16'(-3312);
			7659: out = 16'(-3235);
			7660: out = 16'(-7);
			7661: out = 16'(6582);
			7662: out = 16'(8593);
			7663: out = 16'(-2042);
			7664: out = 16'(-8702);
			7665: out = 16'(-13803);
			7666: out = 16'(1835);
			7667: out = 16'(5358);
			7668: out = 16'(6966);
			7669: out = 16'(5185);
			7670: out = 16'(923);
			7671: out = 16'(-8018);
			7672: out = 16'(-1592);
			7673: out = 16'(518);
			7674: out = 16'(5468);
			7675: out = 16'(-4790);
			7676: out = 16'(-8222);
			7677: out = 16'(-5828);
			7678: out = 16'(2156);
			7679: out = 16'(8134);
			7680: out = 16'(7640);
			7681: out = 16'(6435);
			7682: out = 16'(3274);
			7683: out = 16'(-3628);
			7684: out = 16'(-2973);
			7685: out = 16'(622);
			7686: out = 16'(5549);
			7687: out = 16'(4996);
			7688: out = 16'(9);
			7689: out = 16'(-941);
			7690: out = 16'(-2172);
			7691: out = 16'(163);
			7692: out = 16'(-1885);
			7693: out = 16'(-2969);
			7694: out = 16'(-9432);
			7695: out = 16'(2443);
			7696: out = 16'(7687);
			7697: out = 16'(269);
			7698: out = 16'(-1764);
			7699: out = 16'(-4973);
			7700: out = 16'(342);
			7701: out = 16'(-1099);
			7702: out = 16'(25);
			7703: out = 16'(-4963);
			7704: out = 16'(-1695);
			7705: out = 16'(-446);
			7706: out = 16'(10378);
			7707: out = 16'(5586);
			7708: out = 16'(-3157);
			7709: out = 16'(-13535);
			7710: out = 16'(-10370);
			7711: out = 16'(6296);
			7712: out = 16'(9683);
			7713: out = 16'(8591);
			7714: out = 16'(340);
			7715: out = 16'(-7977);
			7716: out = 16'(-13779);
			7717: out = 16'(-19498);
			7718: out = 16'(-4365);
			7719: out = 16'(10854);
			7720: out = 16'(13654);
			7721: out = 16'(5432);
			7722: out = 16'(-8704);
			7723: out = 16'(-6324);
			7724: out = 16'(-1849);
			7725: out = 16'(9743);
			7726: out = 16'(6582);
			7727: out = 16'(5089);
			7728: out = 16'(-2672);
			7729: out = 16'(-4794);
			7730: out = 16'(-6349);
			7731: out = 16'(2114);
			7732: out = 16'(-3234);
			7733: out = 16'(-2753);
			7734: out = 16'(261);
			7735: out = 16'(5087);
			7736: out = 16'(5982);
			7737: out = 16'(-1978);
			7738: out = 16'(-4525);
			7739: out = 16'(-4869);
			7740: out = 16'(310);
			7741: out = 16'(2427);
			7742: out = 16'(2163);
			7743: out = 16'(4204);
			7744: out = 16'(332);
			7745: out = 16'(-5591);
			7746: out = 16'(-9008);
			7747: out = 16'(-5068);
			7748: out = 16'(9054);
			7749: out = 16'(5813);
			7750: out = 16'(1591);
			7751: out = 16'(-14494);
			7752: out = 16'(-5484);
			7753: out = 16'(2532);
			7754: out = 16'(7731);
			7755: out = 16'(5275);
			7756: out = 16'(685);
			7757: out = 16'(6526);
			7758: out = 16'(3654);
			7759: out = 16'(2075);
			7760: out = 16'(-12312);
			7761: out = 16'(-11196);
			7762: out = 16'(-4572);
			7763: out = 16'(8066);
			7764: out = 16'(9210);
			7765: out = 16'(54);
			7766: out = 16'(551);
			7767: out = 16'(-108);
			7768: out = 16'(2888);
			7769: out = 16'(1266);
			7770: out = 16'(782);
			7771: out = 16'(960);
			7772: out = 16'(-682);
			7773: out = 16'(-2046);
			7774: out = 16'(-5802);
			7775: out = 16'(585);
			7776: out = 16'(7766);
			7777: out = 16'(3684);
			7778: out = 16'(737);
			7779: out = 16'(-4987);
			7780: out = 16'(540);
			7781: out = 16'(4026);
			7782: out = 16'(11778);
			7783: out = 16'(-2372);
			7784: out = 16'(-6570);
			7785: out = 16'(-7341);
			7786: out = 16'(-555);
			7787: out = 16'(3025);
			7788: out = 16'(3556);
			7789: out = 16'(-383);
			7790: out = 16'(-3977);
			7791: out = 16'(-7017);
			7792: out = 16'(-463);
			7793: out = 16'(7208);
			7794: out = 16'(5054);
			7795: out = 16'(4925);
			7796: out = 16'(1306);
			7797: out = 16'(6196);
			7798: out = 16'(855);
			7799: out = 16'(-6216);
			7800: out = 16'(-4003);
			7801: out = 16'(-2031);
			7802: out = 16'(-297);
			7803: out = 16'(-1184);
			7804: out = 16'(-895);
			7805: out = 16'(5422);
			7806: out = 16'(-1117);
			7807: out = 16'(-3035);
			7808: out = 16'(-5335);
			7809: out = 16'(6078);
			7810: out = 16'(12877);
			7811: out = 16'(9254);
			7812: out = 16'(-2372);
			7813: out = 16'(-15651);
			7814: out = 16'(1216);
			7815: out = 16'(1358);
			7816: out = 16'(998);
			7817: out = 16'(-1582);
			7818: out = 16'(-2762);
			7819: out = 16'(-4677);
			7820: out = 16'(-1164);
			7821: out = 16'(621);
			7822: out = 16'(2247);
			7823: out = 16'(643);
			7824: out = 16'(-235);
			7825: out = 16'(2908);
			7826: out = 16'(-8669);
			7827: out = 16'(-15252);
			7828: out = 16'(-69);
			7829: out = 16'(2268);
			7830: out = 16'(6013);
			7831: out = 16'(-14211);
			7832: out = 16'(-3347);
			7833: out = 16'(8950);
			7834: out = 16'(4812);
			7835: out = 16'(-1935);
			7836: out = 16'(-11316);
			7837: out = 16'(-5921);
			7838: out = 16'(648);
			7839: out = 16'(8346);
			7840: out = 16'(10431);
			7841: out = 16'(6849);
			7842: out = 16'(-994);
			7843: out = 16'(-12087);
			7844: out = 16'(-15294);
			7845: out = 16'(-1673);
			7846: out = 16'(4465);
			7847: out = 16'(8485);
			7848: out = 16'(4238);
			7849: out = 16'(-88);
			7850: out = 16'(-4338);
			7851: out = 16'(-4515);
			7852: out = 16'(2214);
			7853: out = 16'(10923);
			7854: out = 16'(9562);
			7855: out = 16'(2432);
			7856: out = 16'(-12385);
			7857: out = 16'(-8715);
			7858: out = 16'(-6138);
			7859: out = 16'(779);
			7860: out = 16'(-33);
			7861: out = 16'(-369);
			7862: out = 16'(-928);
			7863: out = 16'(-7223);
			7864: out = 16'(-8456);
			7865: out = 16'(8201);
			7866: out = 16'(11584);
			7867: out = 16'(13541);
			7868: out = 16'(460);
			7869: out = 16'(-1753);
			7870: out = 16'(-4835);
			7871: out = 16'(245);
			7872: out = 16'(-5531);
			7873: out = 16'(-13967);
			7874: out = 16'(-2304);
			7875: out = 16'(6091);
			7876: out = 16'(13317);
			7877: out = 16'(8487);
			7878: out = 16'(2788);
			7879: out = 16'(-3736);
			7880: out = 16'(-8171);
			7881: out = 16'(-6852);
			7882: out = 16'(7216);
			7883: out = 16'(3891);
			7884: out = 16'(711);
			7885: out = 16'(399);
			7886: out = 16'(3004);
			7887: out = 16'(6848);
			7888: out = 16'(-13034);
			7889: out = 16'(-8297);
			7890: out = 16'(895);
			7891: out = 16'(10586);
			7892: out = 16'(8323);
			7893: out = 16'(-860);
			7894: out = 16'(-7106);
			7895: out = 16'(-7981);
			7896: out = 16'(554);
			7897: out = 16'(1262);
			7898: out = 16'(3546);
			7899: out = 16'(4679);
			7900: out = 16'(2184);
			7901: out = 16'(-2029);
			7902: out = 16'(-12190);
			7903: out = 16'(-6136);
			7904: out = 16'(2600);
			7905: out = 16'(8841);
			7906: out = 16'(9282);
			7907: out = 16'(5710);
			7908: out = 16'(1055);
			7909: out = 16'(-1003);
			7910: out = 16'(418);
			7911: out = 16'(181);
			7912: out = 16'(419);
			7913: out = 16'(-2283);
			7914: out = 16'(1744);
			7915: out = 16'(930);
			7916: out = 16'(-2947);
			7917: out = 16'(-3974);
			7918: out = 16'(-3480);
			7919: out = 16'(-15);
			7920: out = 16'(487);
			7921: out = 16'(1101);
			7922: out = 16'(967);
			7923: out = 16'(3980);
			7924: out = 16'(6764);
			7925: out = 16'(218);
			7926: out = 16'(-54);
			7927: out = 16'(-888);
			7928: out = 16'(435);
			7929: out = 16'(-2737);
			7930: out = 16'(-6786);
			7931: out = 16'(-6115);
			7932: out = 16'(-3742);
			7933: out = 16'(-1725);
			7934: out = 16'(7653);
			7935: out = 16'(10524);
			7936: out = 16'(6671);
			7937: out = 16'(338);
			7938: out = 16'(-5815);
			7939: out = 16'(-6037);
			7940: out = 16'(-9374);
			7941: out = 16'(-8785);
			7942: out = 16'(8767);
			7943: out = 16'(6903);
			7944: out = 16'(1283);
			7945: out = 16'(-6387);
			7946: out = 16'(-4899);
			7947: out = 16'(3976);
			7948: out = 16'(-689);
			7949: out = 16'(2299);
			7950: out = 16'(5578);
			7951: out = 16'(7861);
			7952: out = 16'(4665);
			7953: out = 16'(-5808);
			7954: out = 16'(-4557);
			7955: out = 16'(-4002);
			7956: out = 16'(-2678);
			7957: out = 16'(-3641);
			7958: out = 16'(-3352);
			7959: out = 16'(-753);
			7960: out = 16'(4451);
			7961: out = 16'(9082);
			7962: out = 16'(206);
			7963: out = 16'(841);
			7964: out = 16'(2471);
			7965: out = 16'(4290);
			7966: out = 16'(2911);
			7967: out = 16'(-935);
			7968: out = 16'(-2238);
			7969: out = 16'(-2676);
			7970: out = 16'(351);
			7971: out = 16'(-725);
			7972: out = 16'(-427);
			7973: out = 16'(-3634);
			7974: out = 16'(4057);
			7975: out = 16'(7089);
			7976: out = 16'(-230);
			7977: out = 16'(-2593);
			7978: out = 16'(-3465);
			7979: out = 16'(6752);
			7980: out = 16'(6963);
			7981: out = 16'(4570);
			7982: out = 16'(1860);
			7983: out = 16'(-3388);
			7984: out = 16'(-8648);
			7985: out = 16'(-8855);
			7986: out = 16'(-4843);
			7987: out = 16'(3954);
			7988: out = 16'(1629);
			7989: out = 16'(762);
			7990: out = 16'(-483);
			7991: out = 16'(1127);
			7992: out = 16'(2480);
			7993: out = 16'(153);
			7994: out = 16'(3818);
			7995: out = 16'(4741);
			7996: out = 16'(1589);
			7997: out = 16'(-7129);
			7998: out = 16'(-15518);
			7999: out = 16'(306);
			8000: out = 16'(4407);
			8001: out = 16'(6781);
			8002: out = 16'(2984);
			8003: out = 16'(1865);
			8004: out = 16'(2234);
			8005: out = 16'(-2847);
			8006: out = 16'(-4049);
			8007: out = 16'(-1777);
			8008: out = 16'(5127);
			8009: out = 16'(6556);
			8010: out = 16'(-9359);
			8011: out = 16'(-6277);
			8012: out = 16'(-4820);
			8013: out = 16'(7197);
			8014: out = 16'(2181);
			8015: out = 16'(-1243);
			8016: out = 16'(-16903);
			8017: out = 16'(-4954);
			8018: out = 16'(12753);
			8019: out = 16'(12958);
			8020: out = 16'(6434);
			8021: out = 16'(-10414);
			8022: out = 16'(-2496);
			8023: out = 16'(-681);
			8024: out = 16'(5322);
			8025: out = 16'(-4279);
			8026: out = 16'(-5926);
			8027: out = 16'(1023);
			8028: out = 16'(-1039);
			8029: out = 16'(-2872);
			8030: out = 16'(-11393);
			8031: out = 16'(-1055);
			8032: out = 16'(8091);
			8033: out = 16'(3038);
			8034: out = 16'(2844);
			8035: out = 16'(412);
			8036: out = 16'(7682);
			8037: out = 16'(5152);
			8038: out = 16'(1683);
			8039: out = 16'(-4456);
			8040: out = 16'(-4524);
			8041: out = 16'(298);
			8042: out = 16'(-4669);
			8043: out = 16'(-4251);
			8044: out = 16'(1641);
			8045: out = 16'(-1350);
			8046: out = 16'(1134);
			8047: out = 16'(12591);
			8048: out = 16'(10784);
			8049: out = 16'(6073);
			8050: out = 16'(-15028);
			8051: out = 16'(-8809);
			8052: out = 16'(855);
			8053: out = 16'(-4156);
			8054: out = 16'(-302);
			8055: out = 16'(608);
			8056: out = 16'(7185);
			8057: out = 16'(-1959);
			8058: out = 16'(-18112);
			8059: out = 16'(-10409);
			8060: out = 16'(-2439);
			8061: out = 16'(10949);
			8062: out = 16'(7397);
			8063: out = 16'(6011);
			8064: out = 16'(1956);
			8065: out = 16'(935);
			8066: out = 16'(-1456);
			8067: out = 16'(-1184);
			8068: out = 16'(-3655);
			8069: out = 16'(-4696);
			8070: out = 16'(-12588);
			8071: out = 16'(-5636);
			8072: out = 16'(2771);
			8073: out = 16'(5320);
			8074: out = 16'(3062);
			8075: out = 16'(-3358);
			8076: out = 16'(6839);
			8077: out = 16'(7258);
			8078: out = 16'(5503);
			8079: out = 16'(1273);
			8080: out = 16'(-2700);
			8081: out = 16'(-6891);
			8082: out = 16'(-9031);
			8083: out = 16'(-5303);
			8084: out = 16'(13556);
			8085: out = 16'(9232);
			8086: out = 16'(4969);
			8087: out = 16'(-18936);
			8088: out = 16'(-4055);
			8089: out = 16'(10983);
			8090: out = 16'(10040);
			8091: out = 16'(6382);
			8092: out = 16'(-1741);
			8093: out = 16'(240);
			8094: out = 16'(-2647);
			8095: out = 16'(-4321);
			8096: out = 16'(-355);
			8097: out = 16'(-2215);
			8098: out = 16'(-12039);
			8099: out = 16'(-3827);
			8100: out = 16'(81);
			8101: out = 16'(5090);
			8102: out = 16'(2948);
			8103: out = 16'(1928);
			8104: out = 16'(-1953);
			8105: out = 16'(18);
			8106: out = 16'(1279);
			8107: out = 16'(7002);
			8108: out = 16'(3009);
			8109: out = 16'(-1223);
			8110: out = 16'(-12848);
			8111: out = 16'(-8089);
			8112: out = 16'(2744);
			8113: out = 16'(2875);
			8114: out = 16'(625);
			8115: out = 16'(-9264);
			8116: out = 16'(59);
			8117: out = 16'(1823);
			8118: out = 16'(4407);
			8119: out = 16'(343);
			8120: out = 16'(1729);
			8121: out = 16'(7699);
			8122: out = 16'(5709);
			8123: out = 16'(2051);
			8124: out = 16'(2230);
			8125: out = 16'(-3957);
			8126: out = 16'(-7234);
			8127: out = 16'(-14194);
			8128: out = 16'(-6747);
			8129: out = 16'(2471);
			8130: out = 16'(12676);
			8131: out = 16'(8274);
			8132: out = 16'(-2693);
			8133: out = 16'(-7694);
			8134: out = 16'(-5758);
			8135: out = 16'(5790);
			8136: out = 16'(4457);
			8137: out = 16'(2700);
			8138: out = 16'(-5660);
			8139: out = 16'(-10399);
			8140: out = 16'(-12419);
			8141: out = 16'(576);
			8142: out = 16'(354);
			8143: out = 16'(2543);
			8144: out = 16'(-538);
			8145: out = 16'(6401);
			8146: out = 16'(10746);
			8147: out = 16'(2282);
			8148: out = 16'(-925);
			8149: out = 16'(-2533);
			8150: out = 16'(2487);
			8151: out = 16'(3066);
			8152: out = 16'(-642);
			8153: out = 16'(5178);
			8154: out = 16'(3544);
			8155: out = 16'(-1501);
			8156: out = 16'(-5546);
			8157: out = 16'(-5348);
			8158: out = 16'(691);
			8159: out = 16'(5911);
			8160: out = 16'(8658);
			8161: out = 16'(4638);
			8162: out = 16'(72);
			8163: out = 16'(-4640);
			8164: out = 16'(3423);
			8165: out = 16'(845);
			8166: out = 16'(-2391);
			8167: out = 16'(-7333);
			8168: out = 16'(-7289);
			8169: out = 16'(-3318);
			8170: out = 16'(-3813);
			8171: out = 16'(-50);
			8172: out = 16'(3436);
			8173: out = 16'(5807);
			8174: out = 16'(4728);
			8175: out = 16'(4319);
			8176: out = 16'(-7143);
			8177: out = 16'(-10589);
			8178: out = 16'(3683);
			8179: out = 16'(3574);
			8180: out = 16'(3244);
			8181: out = 16'(1301);
			8182: out = 16'(-1202);
			8183: out = 16'(-3318);
			8184: out = 16'(-10322);
			8185: out = 16'(-6358);
			8186: out = 16'(1255);
			8187: out = 16'(4940);
			8188: out = 16'(4439);
			8189: out = 16'(-242);
			8190: out = 16'(-3912);
			8191: out = 16'(-2271);
			8192: out = 16'(8964);
			8193: out = 16'(6858);
			8194: out = 16'(4527);
			8195: out = 16'(-8982);
			8196: out = 16'(-2077);
			8197: out = 16'(1802);
			8198: out = 16'(3702);
			8199: out = 16'(-461);
			8200: out = 16'(-4595);
			8201: out = 16'(-1546);
			8202: out = 16'(-504);
			8203: out = 16'(1851);
			8204: out = 16'(464);
			8205: out = 16'(2362);
			8206: out = 16'(3294);
			8207: out = 16'(6844);
			8208: out = 16'(1258);
			8209: out = 16'(-13390);
			8210: out = 16'(-5335);
			8211: out = 16'(-1606);
			8212: out = 16'(1048);
			8213: out = 16'(-1470);
			8214: out = 16'(-1408);
			8215: out = 16'(7224);
			8216: out = 16'(5977);
			8217: out = 16'(4983);
			8218: out = 16'(-4175);
			8219: out = 16'(-1335);
			8220: out = 16'(1642);
			8221: out = 16'(8461);
			8222: out = 16'(4245);
			8223: out = 16'(-2641);
			8224: out = 16'(-8444);
			8225: out = 16'(-6114);
			8226: out = 16'(3285);
			8227: out = 16'(3626);
			8228: out = 16'(3717);
			8229: out = 16'(-1043);
			8230: out = 16'(-1957);
			8231: out = 16'(-2122);
			8232: out = 16'(5156);
			8233: out = 16'(1207);
			8234: out = 16'(-514);
			8235: out = 16'(-3222);
			8236: out = 16'(-1296);
			8237: out = 16'(-68);
			8238: out = 16'(1012);
			8239: out = 16'(-2712);
			8240: out = 16'(-7062);
			8241: out = 16'(-827);
			8242: out = 16'(1766);
			8243: out = 16'(4896);
			8244: out = 16'(-2513);
			8245: out = 16'(-4113);
			8246: out = 16'(-2554);
			8247: out = 16'(-220);
			8248: out = 16'(4290);
			8249: out = 16'(12967);
			8250: out = 16'(4479);
			8251: out = 16'(-2907);
			8252: out = 16'(-8795);
			8253: out = 16'(-11029);
			8254: out = 16'(-8994);
			8255: out = 16'(1394);
			8256: out = 16'(5680);
			8257: out = 16'(7517);
			8258: out = 16'(-2834);
			8259: out = 16'(-3841);
			8260: out = 16'(-2204);
			8261: out = 16'(4277);
			8262: out = 16'(6002);
			8263: out = 16'(4069);
			8264: out = 16'(2548);
			8265: out = 16'(-1518);
			8266: out = 16'(-6789);
			8267: out = 16'(-7220);
			8268: out = 16'(-4095);
			8269: out = 16'(6078);
			8270: out = 16'(3670);
			8271: out = 16'(2043);
			8272: out = 16'(-510);
			8273: out = 16'(4554);
			8274: out = 16'(8110);
			8275: out = 16'(-5981);
			8276: out = 16'(-8587);
			8277: out = 16'(-10554);
			8278: out = 16'(6126);
			8279: out = 16'(5611);
			8280: out = 16'(340);
			8281: out = 16'(-3074);
			8282: out = 16'(-3159);
			8283: out = 16'(453);
			8284: out = 16'(-236);
			8285: out = 16'(2493);
			8286: out = 16'(11508);
			8287: out = 16'(3329);
			8288: out = 16'(-2498);
			8289: out = 16'(-14520);
			8290: out = 16'(-1225);
			8291: out = 16'(9022);
			8292: out = 16'(5838);
			8293: out = 16'(-4597);
			8294: out = 16'(-17842);
			8295: out = 16'(3738);
			8296: out = 16'(5853);
			8297: out = 16'(9252);
			8298: out = 16'(-12126);
			8299: out = 16'(-12009);
			8300: out = 16'(-3112);
			8301: out = 16'(1890);
			8302: out = 16'(4389);
			8303: out = 16'(3700);
			8304: out = 16'(-462);
			8305: out = 16'(-2712);
			8306: out = 16'(232);
			8307: out = 16'(309);
			8308: out = 16'(2005);
			8309: out = 16'(4561);
			8310: out = 16'(5002);
			8311: out = 16'(3561);
			8312: out = 16'(-5846);
			8313: out = 16'(-5328);
			8314: out = 16'(-1947);
			8315: out = 16'(614);
			8316: out = 16'(1259);
			8317: out = 16'(-446);
			8318: out = 16'(3240);
			8319: out = 16'(3677);
			8320: out = 16'(3652);
			8321: out = 16'(2705);
			8322: out = 16'(1656);
			8323: out = 16'(-485);
			8324: out = 16'(-2881);
			8325: out = 16'(-2589);
			8326: out = 16'(9608);
			8327: out = 16'(18);
			8328: out = 16'(-5923);
			8329: out = 16'(-3366);
			8330: out = 16'(4762);
			8331: out = 16'(12832);
			8332: out = 16'(-4890);
			8333: out = 16'(-3137);
			8334: out = 16'(-348);
			8335: out = 16'(577);
			8336: out = 16'(-6746);
			8337: out = 16'(-20978);
			8338: out = 16'(-3600);
			8339: out = 16'(5269);
			8340: out = 16'(11044);
			8341: out = 16'(3542);
			8342: out = 16'(-2153);
			8343: out = 16'(-3317);
			8344: out = 16'(-4741);
			8345: out = 16'(-2280);
			8346: out = 16'(1775);
			8347: out = 16'(5128);
			8348: out = 16'(5067);
			8349: out = 16'(3664);
			8350: out = 16'(-4142);
			8351: out = 16'(-10641);
			8352: out = 16'(-1675);
			8353: out = 16'(5048);
			8354: out = 16'(10952);
			8355: out = 16'(3464);
			8356: out = 16'(-1728);
			8357: out = 16'(-5019);
			8358: out = 16'(-9382);
			8359: out = 16'(-3519);
			8360: out = 16'(13181);
			8361: out = 16'(12422);
			8362: out = 16'(7770);
			8363: out = 16'(-7885);
			8364: out = 16'(-11216);
			8365: out = 16'(-10820);
			8366: out = 16'(-227);
			8367: out = 16'(6952);
			8368: out = 16'(11559);
			8369: out = 16'(1876);
			8370: out = 16'(-3687);
			8371: out = 16'(-10036);
			8372: out = 16'(-375);
			8373: out = 16'(-44);
			8374: out = 16'(-3023);
			8375: out = 16'(1715);
			8376: out = 16'(2816);
			8377: out = 16'(3933);
			8378: out = 16'(-1004);
			8379: out = 16'(-3378);
			8380: out = 16'(-5558);
			8381: out = 16'(-1904);
			8382: out = 16'(1647);
			8383: out = 16'(12555);
			8384: out = 16'(2165);
			8385: out = 16'(-6934);
			8386: out = 16'(-13397);
			8387: out = 16'(-3781);
			8388: out = 16'(9911);
			8389: out = 16'(3395);
			8390: out = 16'(3375);
			8391: out = 16'(643);
			8392: out = 16'(-2536);
			8393: out = 16'(-3436);
			8394: out = 16'(542);
			8395: out = 16'(5434);
			8396: out = 16'(7196);
			8397: out = 16'(-1172);
			8398: out = 16'(827);
			8399: out = 16'(-506);
			8400: out = 16'(8513);
			8401: out = 16'(-6928);
			8402: out = 16'(-14664);
			8403: out = 16'(-5276);
			8404: out = 16'(5523);
			8405: out = 16'(13729);
			8406: out = 16'(2639);
			8407: out = 16'(-6051);
			8408: out = 16'(-17784);
			8409: out = 16'(-8006);
			8410: out = 16'(-1271);
			8411: out = 16'(10540);
			8412: out = 16'(-2520);
			8413: out = 16'(-5649);
			8414: out = 16'(-8217);
			8415: out = 16'(989);
			8416: out = 16'(4037);
			8417: out = 16'(1870);
			8418: out = 16'(-123);
			8419: out = 16'(-758);
			8420: out = 16'(-405);
			8421: out = 16'(5408);
			8422: out = 16'(9124);
			8423: out = 16'(6776);
			8424: out = 16'(-2585);
			8425: out = 16'(-14381);
			8426: out = 16'(-331);
			8427: out = 16'(4423);
			8428: out = 16'(10836);
			8429: out = 16'(-1694);
			8430: out = 16'(-3625);
			8431: out = 16'(-2695);
			8432: out = 16'(3775);
			8433: out = 16'(6253);
			8434: out = 16'(5823);
			8435: out = 16'(2666);
			8436: out = 16'(-66);
			8437: out = 16'(-3004);
			8438: out = 16'(1990);
			8439: out = 16'(5764);
			8440: out = 16'(919);
			8441: out = 16'(-3822);
			8442: out = 16'(-9495);
			8443: out = 16'(7732);
			8444: out = 16'(6340);
			8445: out = 16'(2964);
			8446: out = 16'(-6356);
			8447: out = 16'(-7742);
			8448: out = 16'(-5123);
			8449: out = 16'(2106);
			8450: out = 16'(5528);
			8451: out = 16'(5545);
			8452: out = 16'(-671);
			8453: out = 16'(-5109);
			8454: out = 16'(-3650);
			8455: out = 16'(-2094);
			8456: out = 16'(1012);
			8457: out = 16'(619);
			8458: out = 16'(1108);
			8459: out = 16'(-271);
			8460: out = 16'(4767);
			8461: out = 16'(3941);
			8462: out = 16'(4643);
			8463: out = 16'(-5013);
			8464: out = 16'(-3152);
			8465: out = 16'(752);
			8466: out = 16'(9121);
			8467: out = 16'(7687);
			8468: out = 16'(545);
			8469: out = 16'(-5108);
			8470: out = 16'(-6191);
			8471: out = 16'(-795);
			8472: out = 16'(4784);
			8473: out = 16'(6425);
			8474: out = 16'(-1911);
			8475: out = 16'(-4972);
			8476: out = 16'(-6955);
			8477: out = 16'(-927);
			8478: out = 16'(-2200);
			8479: out = 16'(-3891);
			8480: out = 16'(11703);
			8481: out = 16'(7504);
			8482: out = 16'(-223);
			8483: out = 16'(-15415);
			8484: out = 16'(-15646);
			8485: out = 16'(-4223);
			8486: out = 16'(-29);
			8487: out = 16'(3860);
			8488: out = 16'(4670);
			8489: out = 16'(-2906);
			8490: out = 16'(-6164);
			8491: out = 16'(1399);
			8492: out = 16'(4293);
			8493: out = 16'(6914);
			8494: out = 16'(569);
			8495: out = 16'(576);
			8496: out = 16'(-1619);
			8497: out = 16'(-8462);
			8498: out = 16'(-7114);
			8499: out = 16'(-1460);
			8500: out = 16'(-1383);
			8501: out = 16'(2205);
			8502: out = 16'(3615);
			8503: out = 16'(11117);
			8504: out = 16'(6645);
			8505: out = 16'(-7956);
			8506: out = 16'(241);
			8507: out = 16'(4339);
			8508: out = 16'(11243);
			8509: out = 16'(2484);
			8510: out = 16'(-5205);
			8511: out = 16'(-18503);
			8512: out = 16'(-12460);
			8513: out = 16'(-3528);
			8514: out = 16'(8936);
			8515: out = 16'(9018);
			8516: out = 16'(5739);
			8517: out = 16'(-2849);
			8518: out = 16'(-2787);
			8519: out = 16'(576);
			8520: out = 16'(4162);
			8521: out = 16'(-1226);
			8522: out = 16'(-16797);
			8523: out = 16'(943);
			8524: out = 16'(5363);
			8525: out = 16'(4812);
			8526: out = 16'(-2012);
			8527: out = 16'(-5517);
			8528: out = 16'(-649);
			8529: out = 16'(-4379);
			8530: out = 16'(-3732);
			8531: out = 16'(2085);
			8532: out = 16'(5500);
			8533: out = 16'(6385);
			8534: out = 16'(-670);
			8535: out = 16'(-783);
			8536: out = 16'(1521);
			8537: out = 16'(-532);
			8538: out = 16'(-1837);
			8539: out = 16'(-7503);
			8540: out = 16'(10722);
			8541: out = 16'(8604);
			8542: out = 16'(42);
			8543: out = 16'(-13951);
			8544: out = 16'(-13617);
			8545: out = 16'(7065);
			8546: out = 16'(7552);
			8547: out = 16'(9272);
			8548: out = 16'(7908);
			8549: out = 16'(2589);
			8550: out = 16'(-4334);
			8551: out = 16'(-17901);
			8552: out = 16'(-7162);
			8553: out = 16'(8379);
			8554: out = 16'(-64);
			8555: out = 16'(1995);
			8556: out = 16'(-629);
			8557: out = 16'(10816);
			8558: out = 16'(4063);
			8559: out = 16'(-8805);
			8560: out = 16'(167);
			8561: out = 16'(2863);
			8562: out = 16'(673);
			8563: out = 16'(1768);
			8564: out = 16'(2113);
			8565: out = 16'(11208);
			8566: out = 16'(-5602);
			8567: out = 16'(-13480);
			8568: out = 16'(-3226);
			8569: out = 16'(4185);
			8570: out = 16'(9369);
			8571: out = 16'(-5896);
			8572: out = 16'(-8525);
			8573: out = 16'(-9952);
			8574: out = 16'(5815);
			8575: out = 16'(9763);
			8576: out = 16'(10446);
			8577: out = 16'(3483);
			8578: out = 16'(-3025);
			8579: out = 16'(-11211);
			8580: out = 16'(-3027);
			8581: out = 16'(1516);
			8582: out = 16'(1995);
			8583: out = 16'(1989);
			8584: out = 16'(609);
			8585: out = 16'(4494);
			8586: out = 16'(-2961);
			8587: out = 16'(-7471);
			8588: out = 16'(-12590);
			8589: out = 16'(-3549);
			8590: out = 16'(7001);
			8591: out = 16'(12658);
			8592: out = 16'(11331);
			8593: out = 16'(5050);
			8594: out = 16'(-5886);
			8595: out = 16'(-13138);
			8596: out = 16'(-16230);
			8597: out = 16'(-4903);
			8598: out = 16'(5040);
			8599: out = 16'(12861);
			8600: out = 16'(7061);
			8601: out = 16'(7);
			8602: out = 16'(-10465);
			8603: out = 16'(-6968);
			8604: out = 16'(-1807);
			8605: out = 16'(4466);
			8606: out = 16'(3356);
			8607: out = 16'(-140);
			8608: out = 16'(-5469);
			8609: out = 16'(-6889);
			8610: out = 16'(-5712);
			8611: out = 16'(-2123);
			8612: out = 16'(883);
			8613: out = 16'(3100);
			8614: out = 16'(-321);
			8615: out = 16'(57);
			8616: out = 16'(3281);
			8617: out = 16'(5924);
			8618: out = 16'(6709);
			8619: out = 16'(2063);
			8620: out = 16'(3189);
			8621: out = 16'(1504);
			8622: out = 16'(927);
			8623: out = 16'(-5568);
			8624: out = 16'(-8610);
			8625: out = 16'(-594);
			8626: out = 16'(1962);
			8627: out = 16'(3972);
			8628: out = 16'(-1191);
			8629: out = 16'(3233);
			8630: out = 16'(10613);
			8631: out = 16'(-1141);
			8632: out = 16'(-4643);
			8633: out = 16'(-9958);
			8634: out = 16'(7942);
			8635: out = 16'(9555);
			8636: out = 16'(506);
			8637: out = 16'(-6816);
			8638: out = 16'(-10660);
			8639: out = 16'(-4824);
			8640: out = 16'(-1656);
			8641: out = 16'(1965);
			8642: out = 16'(125);
			8643: out = 16'(-1350);
			8644: out = 16'(-3888);
			8645: out = 16'(1619);
			8646: out = 16'(2352);
			8647: out = 16'(4232);
			8648: out = 16'(-1053);
			8649: out = 16'(381);
			8650: out = 16'(2648);
			8651: out = 16'(1118);
			8652: out = 16'(-2595);
			8653: out = 16'(-9391);
			8654: out = 16'(-3496);
			8655: out = 16'(464);
			8656: out = 16'(2643);
			8657: out = 16'(5895);
			8658: out = 16'(6902);
			8659: out = 16'(3693);
			8660: out = 16'(2009);
			8661: out = 16'(-263);
			8662: out = 16'(4519);
			8663: out = 16'(-4960);
			8664: out = 16'(-13470);
			8665: out = 16'(4201);
			8666: out = 16'(9009);
			8667: out = 16'(12636);
			8668: out = 16'(-7028);
			8669: out = 16'(-10833);
			8670: out = 16'(-7286);
			8671: out = 16'(-1657);
			8672: out = 16'(3758);
			8673: out = 16'(6836);
			8674: out = 16'(7418);
			8675: out = 16'(5309);
			8676: out = 16'(112);
			8677: out = 16'(-1664);
			8678: out = 16'(-2632);
			8679: out = 16'(2955);
			8680: out = 16'(-4606);
			8681: out = 16'(-11197);
			8682: out = 16'(-4094);
			8683: out = 16'(-1263);
			8684: out = 16'(3541);
			8685: out = 16'(-5149);
			8686: out = 16'(964);
			8687: out = 16'(10861);
			8688: out = 16'(5708);
			8689: out = 16'(3249);
			8690: out = 16'(-589);
			8691: out = 16'(5156);
			8692: out = 16'(4602);
			8693: out = 16'(-6460);
			8694: out = 16'(-1548);
			8695: out = 16'(-61);
			8696: out = 16'(5610);
			8697: out = 16'(-6304);
			8698: out = 16'(-13111);
			8699: out = 16'(-3553);
			8700: out = 16'(4713);
			8701: out = 16'(12675);
			8702: out = 16'(9504);
			8703: out = 16'(5814);
			8704: out = 16'(-1943);
			8705: out = 16'(-647);
			8706: out = 16'(-4238);
			8707: out = 16'(-6522);
			8708: out = 16'(-6258);
			8709: out = 16'(-3137);
			8710: out = 16'(1290);
			8711: out = 16'(621);
			8712: out = 16'(-147);
			8713: out = 16'(-29);
			8714: out = 16'(-444);
			8715: out = 16'(12);
			8716: out = 16'(-48);
			8717: out = 16'(188);
			8718: out = 16'(-512);
			8719: out = 16'(2);
			8720: out = 16'(-35);
			8721: out = 16'(1114);
			8722: out = 16'(-4852);
			8723: out = 16'(-4777);
			8724: out = 16'(-5200);
			8725: out = 16'(8536);
			8726: out = 16'(8095);
			8727: out = 16'(1023);
			8728: out = 16'(-8536);
			8729: out = 16'(-8083);
			8730: out = 16'(10001);
			8731: out = 16'(8720);
			8732: out = 16'(7802);
			8733: out = 16'(-7652);
			8734: out = 16'(-129);
			8735: out = 16'(3143);
			8736: out = 16'(1851);
			8737: out = 16'(-5471);
			8738: out = 16'(-12106);
			8739: out = 16'(305);
			8740: out = 16'(1471);
			8741: out = 16'(1368);
			8742: out = 16'(328);
			8743: out = 16'(98);
			8744: out = 16'(-269);
			8745: out = 16'(758);
			8746: out = 16'(1114);
			8747: out = 16'(1350);
			8748: out = 16'(1378);
			8749: out = 16'(-196);
			8750: out = 16'(-6674);
			8751: out = 16'(-7249);
			8752: out = 16'(-5194);
			8753: out = 16'(13158);
			8754: out = 16'(6678);
			8755: out = 16'(502);
			8756: out = 16'(-18467);
			8757: out = 16'(-10508);
			8758: out = 16'(3701);
			8759: out = 16'(11972);
			8760: out = 16'(8501);
			8761: out = 16'(-4373);
			8762: out = 16'(-782);
			8763: out = 16'(1969);
			8764: out = 16'(14216);
			8765: out = 16'(-1495);
			8766: out = 16'(-8597);
			8767: out = 16'(-21749);
			8768: out = 16'(-2719);
			8769: out = 16'(9227);
			8770: out = 16'(15279);
			8771: out = 16'(8652);
			8772: out = 16'(655);
			8773: out = 16'(-12578);
			8774: out = 16'(-8702);
			8775: out = 16'(-443);
			8776: out = 16'(9370);
			8777: out = 16'(6861);
			8778: out = 16'(-1729);
			8779: out = 16'(-466);
			8780: out = 16'(-2572);
			8781: out = 16'(-2205);
			8782: out = 16'(1823);
			8783: out = 16'(4205);
			8784: out = 16'(3094);
			8785: out = 16'(-2243);
			8786: out = 16'(-3892);
			8787: out = 16'(9216);
			8788: out = 16'(873);
			8789: out = 16'(-2914);
			8790: out = 16'(-16056);
			8791: out = 16'(-273);
			8792: out = 16'(11385);
			8793: out = 16'(2823);
			8794: out = 16'(-2206);
			8795: out = 16'(-8512);
			8796: out = 16'(-3125);
			8797: out = 16'(-1373);
			8798: out = 16'(705);
			8799: out = 16'(9857);
			8800: out = 16'(8610);
			8801: out = 16'(-1041);
			8802: out = 16'(259);
			8803: out = 16'(-283);
			8804: out = 16'(2735);
			8805: out = 16'(986);
			8806: out = 16'(-205);
			8807: out = 16'(-5718);
			8808: out = 16'(-3784);
			8809: out = 16'(-2167);
			8810: out = 16'(2402);
			8811: out = 16'(364);
			8812: out = 16'(-1514);
			8813: out = 16'(449);
			8814: out = 16'(4162);
			8815: out = 16'(8694);
			8816: out = 16'(-3575);
			8817: out = 16'(-6942);
			8818: out = 16'(-9410);
			8819: out = 16'(4412);
			8820: out = 16'(6361);
			8821: out = 16'(-1131);
			8822: out = 16'(-655);
			8823: out = 16'(-1465);
			8824: out = 16'(1938);
			8825: out = 16'(-2464);
			8826: out = 16'(-2147);
			8827: out = 16'(7495);
			8828: out = 16'(8306);
			8829: out = 16'(6676);
			8830: out = 16'(-9362);
			8831: out = 16'(-10387);
			8832: out = 16'(-8204);
			8833: out = 16'(2044);
			8834: out = 16'(2788);
			8835: out = 16'(-233);
			8836: out = 16'(119);
			8837: out = 16'(179);
			8838: out = 16'(1564);
			8839: out = 16'(4480);
			8840: out = 16'(4949);
			8841: out = 16'(382);
			8842: out = 16'(-434);
			8843: out = 16'(-1033);
			8844: out = 16'(6295);
			8845: out = 16'(154);
			8846: out = 16'(-3705);
			8847: out = 16'(-9538);
			8848: out = 16'(-1205);
			8849: out = 16'(7411);
			8850: out = 16'(50);
			8851: out = 16'(-4125);
			8852: out = 16'(-10964);
			8853: out = 16'(5536);
			8854: out = 16'(8781);
			8855: out = 16'(10747);
			8856: out = 16'(-4022);
			8857: out = 16'(-7853);
			8858: out = 16'(-3620);
			8859: out = 16'(-945);
			8860: out = 16'(1405);
			8861: out = 16'(-406);
			8862: out = 16'(5591);
			8863: out = 16'(6747);
			8864: out = 16'(-10787);
			8865: out = 16'(-6165);
			8866: out = 16'(-1068);
			8867: out = 16'(12852);
			8868: out = 16'(8481);
			8869: out = 16'(2126);
			8870: out = 16'(-12945);
			8871: out = 16'(-9165);
			8872: out = 16'(3845);
			8873: out = 16'(8743);
			8874: out = 16'(5926);
			8875: out = 16'(-9678);
			8876: out = 16'(-6150);
			8877: out = 16'(-6618);
			8878: out = 16'(-3291);
			8879: out = 16'(432);
			8880: out = 16'(4374);
			8881: out = 16'(-675);
			8882: out = 16'(-1044);
			8883: out = 16'(-3353);
			8884: out = 16'(14468);
			8885: out = 16'(4360);
			8886: out = 16'(-3758);
			8887: out = 16'(-18810);
			8888: out = 16'(-8737);
			8889: out = 16'(8601);
			8890: out = 16'(8685);
			8891: out = 16'(2094);
			8892: out = 16'(-14469);
			8893: out = 16'(-9040);
			8894: out = 16'(-1608);
			8895: out = 16'(15642);
			8896: out = 16'(10328);
			8897: out = 16'(5456);
			8898: out = 16'(-9317);
			8899: out = 16'(-5892);
			8900: out = 16'(-2842);
			8901: out = 16'(-99);
			8902: out = 16'(2824);
			8903: out = 16'(4607);
			8904: out = 16'(-876);
			8905: out = 16'(-791);
			8906: out = 16'(466);
			8907: out = 16'(-150);
			8908: out = 16'(23);
			8909: out = 16'(-1705);
			8910: out = 16'(8673);
			8911: out = 16'(10308);
			8912: out = 16'(9540);
			8913: out = 16'(-2274);
			8914: out = 16'(-8994);
			8915: out = 16'(-12363);
			8916: out = 16'(-4921);
			8917: out = 16'(1387);
			8918: out = 16'(4400);
			8919: out = 16'(2653);
			8920: out = 16'(-809);
			8921: out = 16'(-14596);
			8922: out = 16'(-5741);
			8923: out = 16'(6827);
			8924: out = 16'(7820);
			8925: out = 16'(6315);
			8926: out = 16'(-478);
			8927: out = 16'(-3633);
			8928: out = 16'(-4267);
			8929: out = 16'(2045);
			8930: out = 16'(102);
			8931: out = 16'(598);
			8932: out = 16'(-5096);
			8933: out = 16'(3707);
			8934: out = 16'(4593);
			8935: out = 16'(1549);
			8936: out = 16'(-5740);
			8937: out = 16'(-7582);
			8938: out = 16'(4049);
			8939: out = 16'(8620);
			8940: out = 16'(11042);
			8941: out = 16'(3053);
			8942: out = 16'(-2874);
			8943: out = 16'(-10210);
			8944: out = 16'(-590);
			8945: out = 16'(-1288);
			8946: out = 16'(-2684);
			8947: out = 16'(-5212);
			8948: out = 16'(-3274);
			8949: out = 16'(1237);
			8950: out = 16'(3579);
			8951: out = 16'(5847);
			8952: out = 16'(8718);
			8953: out = 16'(3900);
			8954: out = 16'(-1732);
			8955: out = 16'(-11922);
			8956: out = 16'(-8777);
			8957: out = 16'(-3154);
			8958: out = 16'(4968);
			8959: out = 16'(4119);
			8960: out = 16'(305);
			8961: out = 16'(-509);
			8962: out = 16'(-3093);
			8963: out = 16'(-3545);
			8964: out = 16'(-3368);
			8965: out = 16'(-691);
			8966: out = 16'(1408);
			8967: out = 16'(6828);
			8968: out = 16'(6012);
			8969: out = 16'(-392);
			8970: out = 16'(1149);
			8971: out = 16'(119);
			8972: out = 16'(-4089);
			8973: out = 16'(-4752);
			8974: out = 16'(-4133);
			8975: out = 16'(5073);
			8976: out = 16'(1764);
			8977: out = 16'(305);
			8978: out = 16'(-2155);
			8979: out = 16'(4698);
			8980: out = 16'(10856);
			8981: out = 16'(8284);
			8982: out = 16'(3599);
			8983: out = 16'(-2279);
			8984: out = 16'(-3190);
			8985: out = 16'(-1730);
			8986: out = 16'(233);
			8987: out = 16'(5652);
			8988: out = 16'(3396);
			8989: out = 16'(-3976);
			8990: out = 16'(-14093);
			8991: out = 16'(-16026);
			8992: out = 16'(-1883);
			8993: out = 16'(6414);
			8994: out = 16'(12191);
			8995: out = 16'(8580);
			8996: out = 16'(2923);
			8997: out = 16'(-4121);
			8998: out = 16'(-1652);
			8999: out = 16'(1356);
			9000: out = 16'(6743);
			9001: out = 16'(-6405);
			9002: out = 16'(-7859);
			9003: out = 16'(-4921);
			9004: out = 16'(-5033);
			9005: out = 16'(-2232);
			9006: out = 16'(-787);
			9007: out = 16'(9651);
			9008: out = 16'(10426);
			9009: out = 16'(2346);
			9010: out = 16'(-5033);
			9011: out = 16'(-9048);
			9012: out = 16'(-1539);
			9013: out = 16'(-54);
			9014: out = 16'(1369);
			9015: out = 16'(1525);
			9016: out = 16'(-2485);
			9017: out = 16'(-6715);
			9018: out = 16'(-3341);
			9019: out = 16'(181);
			9020: out = 16'(4082);
			9021: out = 16'(9727);
			9022: out = 16'(8001);
			9023: out = 16'(1729);
			9024: out = 16'(-7246);
			9025: out = 16'(-9052);
			9026: out = 16'(1862);
			9027: out = 16'(472);
			9028: out = 16'(1197);
			9029: out = 16'(-3331);
			9030: out = 16'(-781);
			9031: out = 16'(-716);
			9032: out = 16'(-943);
			9033: out = 16'(-3655);
			9034: out = 16'(-4575);
			9035: out = 16'(113);
			9036: out = 16'(4715);
			9037: out = 16'(8908);
			9038: out = 16'(1226);
			9039: out = 16'(-601);
			9040: out = 16'(-1626);
			9041: out = 16'(-138);
			9042: out = 16'(-35);
			9043: out = 16'(184);
			9044: out = 16'(-2738);
			9045: out = 16'(-4821);
			9046: out = 16'(-8030);
			9047: out = 16'(-1283);
			9048: out = 16'(3460);
			9049: out = 16'(903);
			9050: out = 16'(4240);
			9051: out = 16'(5896);
			9052: out = 16'(5893);
			9053: out = 16'(2451);
			9054: out = 16'(-2317);
			9055: out = 16'(366);
			9056: out = 16'(201);
			9057: out = 16'(2806);
			9058: out = 16'(-11419);
			9059: out = 16'(-8492);
			9060: out = 16'(4658);
			9061: out = 16'(8612);
			9062: out = 16'(8320);
			9063: out = 16'(-4021);
			9064: out = 16'(2125);
			9065: out = 16'(2542);
			9066: out = 16'(175);
			9067: out = 16'(-485);
			9068: out = 16'(479);
			9069: out = 16'(1707);
			9070: out = 16'(1896);
			9071: out = 16'(-100);
			9072: out = 16'(1972);
			9073: out = 16'(-4495);
			9074: out = 16'(-10860);
			9075: out = 16'(-8046);
			9076: out = 16'(779);
			9077: out = 16'(14370);
			9078: out = 16'(3341);
			9079: out = 16'(-2260);
			9080: out = 16'(-9678);
			9081: out = 16'(-2240);
			9082: out = 16'(1805);
			9083: out = 16'(691);
			9084: out = 16'(3894);
			9085: out = 16'(2425);
			9086: out = 16'(-8472);
			9087: out = 16'(-10360);
			9088: out = 16'(-8629);
			9089: out = 16'(3372);
			9090: out = 16'(7366);
			9091: out = 16'(8447);
			9092: out = 16'(4533);
			9093: out = 16'(2082);
			9094: out = 16'(1231);
			9095: out = 16'(-4576);
			9096: out = 16'(-3434);
			9097: out = 16'(1423);
			9098: out = 16'(2084);
			9099: out = 16'(1656);
			9100: out = 16'(-308);
			9101: out = 16'(-1312);
			9102: out = 16'(-2574);
			9103: out = 16'(-9772);
			9104: out = 16'(-2057);
			9105: out = 16'(4025);
			9106: out = 16'(10694);
			9107: out = 16'(5588);
			9108: out = 16'(-526);
			9109: out = 16'(-8407);
			9110: out = 16'(-7163);
			9111: out = 16'(-3284);
			9112: out = 16'(6493);
			9113: out = 16'(5442);
			9114: out = 16'(550);
			9115: out = 16'(-15653);
			9116: out = 16'(-17909);
			9117: out = 16'(-5118);
			9118: out = 16'(6074);
			9119: out = 16'(13501);
			9120: out = 16'(8909);
			9121: out = 16'(5571);
			9122: out = 16'(-2302);
			9123: out = 16'(-9072);
			9124: out = 16'(-9450);
			9125: out = 16'(-3968);
			9126: out = 16'(1023);
			9127: out = 16'(5050);
			9128: out = 16'(4244);
			9129: out = 16'(8907);
			9130: out = 16'(3476);
			9131: out = 16'(-1337);
			9132: out = 16'(-10986);
			9133: out = 16'(-3619);
			9134: out = 16'(15935);
			9135: out = 16'(10508);
			9136: out = 16'(5084);
			9137: out = 16'(-11786);
			9138: out = 16'(-5876);
			9139: out = 16'(-1820);
			9140: out = 16'(9277);
			9141: out = 16'(4506);
			9142: out = 16'(127);
			9143: out = 16'(-17831);
			9144: out = 16'(-9822);
			9145: out = 16'(1203);
			9146: out = 16'(12111);
			9147: out = 16'(10330);
			9148: out = 16'(3110);
			9149: out = 16'(-831);
			9150: out = 16'(-5739);
			9151: out = 16'(-9054);
			9152: out = 16'(-1597);
			9153: out = 16'(3980);
			9154: out = 16'(10144);
			9155: out = 16'(-3597);
			9156: out = 16'(-9385);
			9157: out = 16'(-3246);
			9158: out = 16'(365);
			9159: out = 16'(3667);
			9160: out = 16'(-5879);
			9161: out = 16'(-1677);
			9162: out = 16'(814);
			9163: out = 16'(10928);
			9164: out = 16'(5976);
			9165: out = 16'(549);
			9166: out = 16'(-4793);
			9167: out = 16'(-1131);
			9168: out = 16'(6353);
			9169: out = 16'(1555);
			9170: out = 16'(-1491);
			9171: out = 16'(-7094);
			9172: out = 16'(-1538);
			9173: out = 16'(1776);
			9174: out = 16'(5835);
			9175: out = 16'(4163);
			9176: out = 16'(2809);
			9177: out = 16'(694);
			9178: out = 16'(1558);
			9179: out = 16'(1961);
			9180: out = 16'(-625);
			9181: out = 16'(-1008);
			9182: out = 16'(-2166);
			9183: out = 16'(482);
			9184: out = 16'(-6049);
			9185: out = 16'(-13959);
			9186: out = 16'(-4332);
			9187: out = 16'(673);
			9188: out = 16'(6413);
			9189: out = 16'(-191);
			9190: out = 16'(-146);
			9191: out = 16'(3991);
			9192: out = 16'(773);
			9193: out = 16'(-938);
			9194: out = 16'(-2754);
			9195: out = 16'(-2639);
			9196: out = 16'(-2270);
			9197: out = 16'(368);
			9198: out = 16'(496);
			9199: out = 16'(1093);
			9200: out = 16'(-2886);
			9201: out = 16'(187);
			9202: out = 16'(3426);
			9203: out = 16'(12486);
			9204: out = 16'(12151);
			9205: out = 16'(9647);
			9206: out = 16'(-3926);
			9207: out = 16'(-7356);
			9208: out = 16'(-5315);
			9209: out = 16'(132);
			9210: out = 16'(2663);
			9211: out = 16'(3521);
			9212: out = 16'(-8259);
			9213: out = 16'(-12295);
			9214: out = 16'(1390);
			9215: out = 16'(6640);
			9216: out = 16'(11474);
			9217: out = 16'(-2785);
			9218: out = 16'(2033);
			9219: out = 16'(2626);
			9220: out = 16'(8609);
			9221: out = 16'(-1508);
			9222: out = 16'(-11567);
			9223: out = 16'(-12923);
			9224: out = 16'(-5062);
			9225: out = 16'(7546);
			9226: out = 16'(4277);
			9227: out = 16'(-1048);
			9228: out = 16'(-12608);
			9229: out = 16'(-7508);
			9230: out = 16'(-1444);
			9231: out = 16'(7679);
			9232: out = 16'(11587);
			9233: out = 16'(8117);
			9234: out = 16'(-14216);
			9235: out = 16'(-17201);
			9236: out = 16'(-14827);
			9237: out = 16'(7247);
			9238: out = 16'(12832);
			9239: out = 16'(14294);
			9240: out = 16'(-360);
			9241: out = 16'(-7411);
			9242: out = 16'(-13466);
			9243: out = 16'(-94);
			9244: out = 16'(4057);
			9245: out = 16'(4675);
			9246: out = 16'(2453);
			9247: out = 16'(1042);
			9248: out = 16'(1559);
			9249: out = 16'(2882);
			9250: out = 16'(559);
			9251: out = 16'(-17193);
			9252: out = 16'(-9978);
			9253: out = 16'(-3148);
			9254: out = 16'(16113);
			9255: out = 16'(5502);
			9256: out = 16'(-4193);
			9257: out = 16'(-15640);
			9258: out = 16'(-6295);
			9259: out = 16'(7921);
			9260: out = 16'(6808);
			9261: out = 16'(4370);
			9262: out = 16'(-1858);
			9263: out = 16'(-8367);
			9264: out = 16'(-7488);
			9265: out = 16'(1313);
			9266: out = 16'(6159);
			9267: out = 16'(6917);
			9268: out = 16'(-26);
			9269: out = 16'(-9034);
			9270: out = 16'(-13071);
			9271: out = 16'(2419);
			9272: out = 16'(7185);
			9273: out = 16'(11871);
			9274: out = 16'(-7771);
			9275: out = 16'(-1494);
			9276: out = 16'(3693);
			9277: out = 16'(13504);
			9278: out = 16'(8462);
			9279: out = 16'(454);
			9280: out = 16'(-9361);
			9281: out = 16'(-9063);
			9282: out = 16'(32);
			9283: out = 16'(3845);
			9284: out = 16'(4552);
			9285: out = 16'(-6303);
			9286: out = 16'(4356);
			9287: out = 16'(6687);
			9288: out = 16'(6537);
			9289: out = 16'(-1849);
			9290: out = 16'(-5462);
			9291: out = 16'(5778);
			9292: out = 16'(2978);
			9293: out = 16'(-925);
			9294: out = 16'(-4125);
			9295: out = 16'(-4791);
			9296: out = 16'(-1676);
			9297: out = 16'(-9181);
			9298: out = 16'(-2695);
			9299: out = 16'(6451);
			9300: out = 16'(9031);
			9301: out = 16'(4058);
			9302: out = 16'(-8065);
			9303: out = 16'(-6906);
			9304: out = 16'(-4203);
			9305: out = 16'(23);
			9306: out = 16'(7221);
			9307: out = 16'(9036);
			9308: out = 16'(4529);
			9309: out = 16'(-4977);
			9310: out = 16'(-12245);
			9311: out = 16'(-9238);
			9312: out = 16'(-1076);
			9313: out = 16'(8781);
			9314: out = 16'(10345);
			9315: out = 16'(7180);
			9316: out = 16'(-1017);
			9317: out = 16'(-4587);
			9318: out = 16'(-5077);
			9319: out = 16'(1365);
			9320: out = 16'(636);
			9321: out = 16'(1019);
			9322: out = 16'(-4454);
			9323: out = 16'(197);
			9324: out = 16'(1063);
			9325: out = 16'(1604);
			9326: out = 16'(-1233);
			9327: out = 16'(-1712);
			9328: out = 16'(2320);
			9329: out = 16'(5016);
			9330: out = 16'(6588);
			9331: out = 16'(-692);
			9332: out = 16'(-1477);
			9333: out = 16'(-1158);
			9334: out = 16'(1915);
			9335: out = 16'(3319);
			9336: out = 16'(4647);
			9337: out = 16'(-2966);
			9338: out = 16'(-5770);
			9339: out = 16'(-4780);
			9340: out = 16'(-2022);
			9341: out = 16'(1510);
			9342: out = 16'(3244);
			9343: out = 16'(6773);
			9344: out = 16'(6026);
			9345: out = 16'(-5047);
			9346: out = 16'(-2650);
			9347: out = 16'(744);
			9348: out = 16'(5419);
			9349: out = 16'(1);
			9350: out = 16'(-8737);
			9351: out = 16'(5158);
			9352: out = 16'(5278);
			9353: out = 16'(7222);
			9354: out = 16'(-11944);
			9355: out = 16'(-10374);
			9356: out = 16'(1942);
			9357: out = 16'(8400);
			9358: out = 16'(8353);
			9359: out = 16'(-811);
			9360: out = 16'(-4516);
			9361: out = 16'(-7125);
			9362: out = 16'(-6898);
			9363: out = 16'(653);
			9364: out = 16'(6858);
			9365: out = 16'(7682);
			9366: out = 16'(1991);
			9367: out = 16'(-5339);
			9368: out = 16'(-5007);
			9369: out = 16'(-2464);
			9370: out = 16'(3368);
			9371: out = 16'(3832);
			9372: out = 16'(3297);
			9373: out = 16'(-1162);
			9374: out = 16'(-964);
			9375: out = 16'(-1507);
			9376: out = 16'(1307);
			9377: out = 16'(-324);
			9378: out = 16'(1474);
			9379: out = 16'(5291);
			9380: out = 16'(6464);
			9381: out = 16'(3586);
			9382: out = 16'(-11997);
			9383: out = 16'(-10962);
			9384: out = 16'(-7400);
			9385: out = 16'(6942);
			9386: out = 16'(5343);
			9387: out = 16'(1688);
			9388: out = 16'(-2315);
			9389: out = 16'(-932);
			9390: out = 16'(2501);
			9391: out = 16'(568);
			9392: out = 16'(-2738);
			9393: out = 16'(-8302);
			9394: out = 16'(-10088);
			9395: out = 16'(-7648);
			9396: out = 16'(2128);
			9397: out = 16'(2771);
			9398: out = 16'(3932);
			9399: out = 16'(1123);
			9400: out = 16'(1764);
			9401: out = 16'(1779);
			9402: out = 16'(7155);
			9403: out = 16'(3584);
			9404: out = 16'(-163);
			9405: out = 16'(-7276);
			9406: out = 16'(-5001);
			9407: out = 16'(892);
			9408: out = 16'(1528);
			9409: out = 16'(3205);
			9410: out = 16'(1833);
			9411: out = 16'(3142);
			9412: out = 16'(965);
			9413: out = 16'(679);
			9414: out = 16'(-7292);
			9415: out = 16'(-6615);
			9416: out = 16'(2474);
			9417: out = 16'(5595);
			9418: out = 16'(5494);
			9419: out = 16'(-1061);
			9420: out = 16'(-5373);
			9421: out = 16'(-7349);
			9422: out = 16'(-862);
			9423: out = 16'(3495);
			9424: out = 16'(7532);
			9425: out = 16'(9336);
			9426: out = 16'(7618);
			9427: out = 16'(3288);
			9428: out = 16'(-4219);
			9429: out = 16'(-11632);
			9430: out = 16'(-20106);
			9431: out = 16'(-6202);
			9432: out = 16'(3209);
			9433: out = 16'(12292);
			9434: out = 16'(3488);
			9435: out = 16'(-2231);
			9436: out = 16'(-9562);
			9437: out = 16'(2708);
			9438: out = 16'(10965);
			9439: out = 16'(9707);
			9440: out = 16'(147);
			9441: out = 16'(-10244);
			9442: out = 16'(2416);
			9443: out = 16'(3560);
			9444: out = 16'(6992);
			9445: out = 16'(-8175);
			9446: out = 16'(-5018);
			9447: out = 16'(3009);
			9448: out = 16'(2209);
			9449: out = 16'(766);
			9450: out = 16'(-4630);
			9451: out = 16'(5084);
			9452: out = 16'(5582);
			9453: out = 16'(-4768);
			9454: out = 16'(-6254);
			9455: out = 16'(-6032);
			9456: out = 16'(10950);
			9457: out = 16'(929);
			9458: out = 16'(-5054);
			9459: out = 16'(-15430);
			9460: out = 16'(-1763);
			9461: out = 16'(12174);
			9462: out = 16'(7240);
			9463: out = 16'(-1451);
			9464: out = 16'(-16358);
			9465: out = 16'(-2766);
			9466: out = 16'(1020);
			9467: out = 16'(6841);
			9468: out = 16'(-1176);
			9469: out = 16'(-1375);
			9470: out = 16'(1468);
			9471: out = 16'(1734);
			9472: out = 16'(-128);
			9473: out = 16'(-6399);
			9474: out = 16'(-2627);
			9475: out = 16'(1258);
			9476: out = 16'(3489);
			9477: out = 16'(1624);
			9478: out = 16'(-1241);
			9479: out = 16'(9302);
			9480: out = 16'(2647);
			9481: out = 16'(-4296);
			9482: out = 16'(-4320);
			9483: out = 16'(2483);
			9484: out = 16'(13166);
			9485: out = 16'(3180);
			9486: out = 16'(-3096);
			9487: out = 16'(-14093);
			9488: out = 16'(-5135);
			9489: out = 16'(-1230);
			9490: out = 16'(1751);
			9491: out = 16'(-472);
			9492: out = 16'(-556);
			9493: out = 16'(1155);
			9494: out = 16'(6403);
			9495: out = 16'(9187);
			9496: out = 16'(1473);
			9497: out = 16'(-1003);
			9498: out = 16'(-4305);
			9499: out = 16'(2505);
			9500: out = 16'(-537);
			9501: out = 16'(-3995);
			9502: out = 16'(-6302);
			9503: out = 16'(-3759);
			9504: out = 16'(1450);
			9505: out = 16'(515);
			9506: out = 16'(77);
			9507: out = 16'(215);
			9508: out = 16'(-2828);
			9509: out = 16'(-2704);
			9510: out = 16'(116);
			9511: out = 16'(5676);
			9512: out = 16'(8909);
			9513: out = 16'(6707);
			9514: out = 16'(1936);
			9515: out = 16'(-3873);
			9516: out = 16'(-1999);
			9517: out = 16'(-3808);
			9518: out = 16'(-3275);
			9519: out = 16'(-3476);
			9520: out = 16'(2035);
			9521: out = 16'(9019);
			9522: out = 16'(1326);
			9523: out = 16'(-630);
			9524: out = 16'(-206);
			9525: out = 16'(861);
			9526: out = 16'(-502);
			9527: out = 16'(-8318);
			9528: out = 16'(-2592);
			9529: out = 16'(442);
			9530: out = 16'(1447);
			9531: out = 16'(-796);
			9532: out = 16'(-2572);
			9533: out = 16'(-47);
			9534: out = 16'(-769);
			9535: out = 16'(-255);
			9536: out = 16'(11078);
			9537: out = 16'(11340);
			9538: out = 16'(8267);
			9539: out = 16'(-3750);
			9540: out = 16'(-5100);
			9541: out = 16'(3455);
			9542: out = 16'(-8684);
			9543: out = 16'(-8771);
			9544: out = 16'(-4196);
			9545: out = 16'(3910);
			9546: out = 16'(3722);
			9547: out = 16'(-12205);
			9548: out = 16'(-6922);
			9549: out = 16'(-554);
			9550: out = 16'(12815);
			9551: out = 16'(10109);
			9552: out = 16'(4914);
			9553: out = 16'(1375);
			9554: out = 16'(-4767);
			9555: out = 16'(-9003);
			9556: out = 16'(-5135);
			9557: out = 16'(918);
			9558: out = 16'(8156);
			9559: out = 16'(4361);
			9560: out = 16'(-263);
			9561: out = 16'(-9711);
			9562: out = 16'(-4344);
			9563: out = 16'(771);
			9564: out = 16'(12232);
			9565: out = 16'(3507);
			9566: out = 16'(-1463);
			9567: out = 16'(-6729);
			9568: out = 16'(-1373);
			9569: out = 16'(3004);
			9570: out = 16'(3374);
			9571: out = 16'(-100);
			9572: out = 16'(-4444);
			9573: out = 16'(-1714);
			9574: out = 16'(2085);
			9575: out = 16'(8243);
			9576: out = 16'(584);
			9577: out = 16'(-1118);
			9578: out = 16'(-4633);
			9579: out = 16'(2072);
			9580: out = 16'(4629);
			9581: out = 16'(10089);
			9582: out = 16'(-4962);
			9583: out = 16'(-11829);
			9584: out = 16'(-12049);
			9585: out = 16'(-579);
			9586: out = 16'(7449);
			9587: out = 16'(-1117);
			9588: out = 16'(1111);
			9589: out = 16'(275);
			9590: out = 16'(1500);
			9591: out = 16'(-1257);
			9592: out = 16'(-2327);
			9593: out = 16'(557);
			9594: out = 16'(336);
			9595: out = 16'(-3274);
			9596: out = 16'(3884);
			9597: out = 16'(4357);
			9598: out = 16'(6081);
			9599: out = 16'(-9705);
			9600: out = 16'(-14009);
			9601: out = 16'(-7288);
			9602: out = 16'(-386);
			9603: out = 16'(4906);
			9604: out = 16'(3280);
			9605: out = 16'(1993);
			9606: out = 16'(-456);
			9607: out = 16'(1595);
			9608: out = 16'(4265);
			9609: out = 16'(7853);
			9610: out = 16'(-954);
			9611: out = 16'(-5165);
			9612: out = 16'(-12414);
			9613: out = 16'(7734);
			9614: out = 16'(6323);
			9615: out = 16'(825);
			9616: out = 16'(-13800);
			9617: out = 16'(-12442);
			9618: out = 16'(6362);
			9619: out = 16'(910);
			9620: out = 16'(1939);
			9621: out = 16'(7040);
			9622: out = 16'(3447);
			9623: out = 16'(-66);
			9624: out = 16'(-7773);
			9625: out = 16'(338);
			9626: out = 16'(6979);
			9627: out = 16'(-2124);
			9628: out = 16'(-6393);
			9629: out = 16'(-11675);
			9630: out = 16'(2562);
			9631: out = 16'(3075);
			9632: out = 16'(1663);
			9633: out = 16'(1065);
			9634: out = 16'(4183);
			9635: out = 16'(11256);
			9636: out = 16'(3190);
			9637: out = 16'(-768);
			9638: out = 16'(-5507);
			9639: out = 16'(900);
			9640: out = 16'(3330);
			9641: out = 16'(4);
			9642: out = 16'(571);
			9643: out = 16'(353);
			9644: out = 16'(-6827);
			9645: out = 16'(928);
			9646: out = 16'(9132);
			9647: out = 16'(12434);
			9648: out = 16'(7787);
			9649: out = 16'(-1914);
			9650: out = 16'(2923);
			9651: out = 16'(-3094);
			9652: out = 16'(-10969);
			9653: out = 16'(-6013);
			9654: out = 16'(-228);
			9655: out = 16'(8918);
			9656: out = 16'(-1530);
			9657: out = 16'(-5273);
			9658: out = 16'(110);
			9659: out = 16'(-230);
			9660: out = 16'(883);
			9661: out = 16'(-3576);
			9662: out = 16'(3408);
			9663: out = 16'(7228);
			9664: out = 16'(1468);
			9665: out = 16'(-2013);
			9666: out = 16'(-5721);
			9667: out = 16'(-854);
			9668: out = 16'(49);
			9669: out = 16'(1225);
			9670: out = 16'(-3300);
			9671: out = 16'(-3692);
			9672: out = 16'(-2651);
			9673: out = 16'(2698);
			9674: out = 16'(4186);
			9675: out = 16'(635);
			9676: out = 16'(1475);
			9677: out = 16'(853);
			9678: out = 16'(2657);
			9679: out = 16'(-1192);
			9680: out = 16'(-2750);
			9681: out = 16'(-2115);
			9682: out = 16'(3273);
			9683: out = 16'(7269);
			9684: out = 16'(-1055);
			9685: out = 16'(-3916);
			9686: out = 16'(-6789);
			9687: out = 16'(1212);
			9688: out = 16'(1830);
			9689: out = 16'(638);
			9690: out = 16'(1003);
			9691: out = 16'(996);
			9692: out = 16'(589);
			9693: out = 16'(197);
			9694: out = 16'(36);
			9695: out = 16'(2531);
			9696: out = 16'(-4412);
			9697: out = 16'(-7978);
			9698: out = 16'(-2490);
			9699: out = 16'(-1770);
			9700: out = 16'(-253);
			9701: out = 16'(-6692);
			9702: out = 16'(-3095);
			9703: out = 16'(325);
			9704: out = 16'(2243);
			9705: out = 16'(4428);
			9706: out = 16'(8153);
			9707: out = 16'(-1433);
			9708: out = 16'(-3527);
			9709: out = 16'(-7198);
			9710: out = 16'(8206);
			9711: out = 16'(8721);
			9712: out = 16'(922);
			9713: out = 16'(-10001);
			9714: out = 16'(-13445);
			9715: out = 16'(-3963);
			9716: out = 16'(7153);
			9717: out = 16'(15162);
			9718: out = 16'(10945);
			9719: out = 16'(4428);
			9720: out = 16'(-4250);
			9721: out = 16'(2705);
			9722: out = 16'(1766);
			9723: out = 16'(3256);
			9724: out = 16'(-7936);
			9725: out = 16'(-9255);
			9726: out = 16'(-8933);
			9727: out = 16'(-1932);
			9728: out = 16'(2776);
			9729: out = 16'(7928);
			9730: out = 16'(5269);
			9731: out = 16'(2145);
			9732: out = 16'(-7214);
			9733: out = 16'(-1122);
			9734: out = 16'(1377);
			9735: out = 16'(4178);
			9736: out = 16'(-8308);
			9737: out = 16'(-16924);
			9738: out = 16'(2937);
			9739: out = 16'(7515);
			9740: out = 16'(11839);
			9741: out = 16'(-14791);
			9742: out = 16'(-14892);
			9743: out = 16'(-8836);
			9744: out = 16'(8130);
			9745: out = 16'(9899);
			9746: out = 16'(1562);
			9747: out = 16'(4232);
			9748: out = 16'(2026);
			9749: out = 16'(-1156);
			9750: out = 16'(-1554);
			9751: out = 16'(574);
			9752: out = 16'(8939);
			9753: out = 16'(2574);
			9754: out = 16'(-3231);
			9755: out = 16'(-9840);
			9756: out = 16'(-5295);
			9757: out = 16'(1849);
			9758: out = 16'(2588);
			9759: out = 16'(4797);
			9760: out = 16'(3918);
			9761: out = 16'(1268);
			9762: out = 16'(-182);
			9763: out = 16'(1791);
			9764: out = 16'(-3146);
			9765: out = 16'(-5461);
			9766: out = 16'(-12581);
			9767: out = 16'(904);
			9768: out = 16'(4365);
			9769: out = 16'(1965);
			9770: out = 16'(-6806);
			9771: out = 16'(-10690);
			9772: out = 16'(-3839);
			9773: out = 16'(5679);
			9774: out = 16'(12937);
			9775: out = 16'(1240);
			9776: out = 16'(1270);
			9777: out = 16'(-207);
			9778: out = 16'(972);
			9779: out = 16'(-3733);
			9780: out = 16'(-10358);
			9781: out = 16'(-212);
			9782: out = 16'(3153);
			9783: out = 16'(6453);
			9784: out = 16'(-2477);
			9785: out = 16'(-3329);
			9786: out = 16'(1590);
			9787: out = 16'(9194);
			9788: out = 16'(10905);
			9789: out = 16'(948);
			9790: out = 16'(-5286);
			9791: out = 16'(-9427);
			9792: out = 16'(6994);
			9793: out = 16'(3502);
			9794: out = 16'(1087);
			9795: out = 16'(-2462);
			9796: out = 16'(-1467);
			9797: out = 16'(-147);
			9798: out = 16'(260);
			9799: out = 16'(716);
			9800: out = 16'(2813);
			9801: out = 16'(-3779);
			9802: out = 16'(-3644);
			9803: out = 16'(310);
			9804: out = 16'(6807);
			9805: out = 16'(8242);
			9806: out = 16'(-1180);
			9807: out = 16'(467);
			9808: out = 16'(-814);
			9809: out = 16'(353);
			9810: out = 16'(-5011);
			9811: out = 16'(-7645);
			9812: out = 16'(-4477);
			9813: out = 16'(-1635);
			9814: out = 16'(689);
			9815: out = 16'(7312);
			9816: out = 16'(3396);
			9817: out = 16'(-4644);
			9818: out = 16'(-1882);
			9819: out = 16'(2704);
			9820: out = 16'(13234);
			9821: out = 16'(2419);
			9822: out = 16'(-4280);
			9823: out = 16'(-17225);
			9824: out = 16'(-5326);
			9825: out = 16'(1137);
			9826: out = 16'(2492);
			9827: out = 16'(1091);
			9828: out = 16'(289);
			9829: out = 16'(-490);
			9830: out = 16'(2133);
			9831: out = 16'(3808);
			9832: out = 16'(9901);
			9833: out = 16'(1351);
			9834: out = 16'(-10296);
			9835: out = 16'(-9057);
			9836: out = 16'(-3707);
			9837: out = 16'(7993);
			9838: out = 16'(-1015);
			9839: out = 16'(-4589);
			9840: out = 16'(-10692);
			9841: out = 16'(-2994);
			9842: out = 16'(3310);
			9843: out = 16'(11826);
			9844: out = 16'(10449);
			9845: out = 16'(6555);
			9846: out = 16'(-10402);
			9847: out = 16'(-5444);
			9848: out = 16'(-449);
			9849: out = 16'(2377);
			9850: out = 16'(-2011);
			9851: out = 16'(-8094);
			9852: out = 16'(1066);
			9853: out = 16'(820);
			9854: out = 16'(580);
			9855: out = 16'(-1323);
			9856: out = 16'(921);
			9857: out = 16'(4954);
			9858: out = 16'(2267);
			9859: out = 16'(1047);
			9860: out = 16'(1620);
			9861: out = 16'(294);
			9862: out = 16'(-300);
			9863: out = 16'(-4251);
			9864: out = 16'(-969);
			9865: out = 16'(180);
			9866: out = 16'(1912);
			9867: out = 16'(-2346);
			9868: out = 16'(-4802);
			9869: out = 16'(-4493);
			9870: out = 16'(2039);
			9871: out = 16'(8364);
			9872: out = 16'(9988);
			9873: out = 16'(2808);
			9874: out = 16'(-10137);
			9875: out = 16'(-8966);
			9876: out = 16'(-3710);
			9877: out = 16'(11071);
			9878: out = 16'(6192);
			9879: out = 16'(2532);
			9880: out = 16'(-13073);
			9881: out = 16'(-380);
			9882: out = 16'(4890);
			9883: out = 16'(2572);
			9884: out = 16'(827);
			9885: out = 16'(4);
			9886: out = 16'(925);
			9887: out = 16'(3170);
			9888: out = 16'(4427);
			9889: out = 16'(7051);
			9890: out = 16'(-1011);
			9891: out = 16'(-13096);
			9892: out = 16'(-6001);
			9893: out = 16'(-2103);
			9894: out = 16'(5606);
			9895: out = 16'(-1496);
			9896: out = 16'(-2713);
			9897: out = 16'(-4127);
			9898: out = 16'(-1818);
			9899: out = 16'(866);
			9900: out = 16'(11496);
			9901: out = 16'(5574);
			9902: out = 16'(917);
			9903: out = 16'(-19794);
			9904: out = 16'(-6531);
			9905: out = 16'(5785);
			9906: out = 16'(13434);
			9907: out = 16'(1089);
			9908: out = 16'(-16353);
			9909: out = 16'(-8874);
			9910: out = 16'(-4616);
			9911: out = 16'(4184);
			9912: out = 16'(4024);
			9913: out = 16'(4850);
			9914: out = 16'(2357);
			9915: out = 16'(-885);
			9916: out = 16'(606);
			9917: out = 16'(13468);
			9918: out = 16'(6271);
			9919: out = 16'(-190);
			9920: out = 16'(-17331);
			9921: out = 16'(-15904);
			9922: out = 16'(-11247);
			9923: out = 16'(8225);
			9924: out = 16'(8203);
			9925: out = 16'(6243);
			9926: out = 16'(-6184);
			9927: out = 16'(-3851);
			9928: out = 16'(2228);
			9929: out = 16'(7263);
			9930: out = 16'(3039);
			9931: out = 16'(-9866);
			9932: out = 16'(-3120);
			9933: out = 16'(479);
			9934: out = 16'(10130);
			9935: out = 16'(-233);
			9936: out = 16'(-5047);
			9937: out = 16'(-11796);
			9938: out = 16'(-2313);
			9939: out = 16'(5055);
			9940: out = 16'(10723);
			9941: out = 16'(8367);
			9942: out = 16'(4129);
			9943: out = 16'(-8824);
			9944: out = 16'(-8538);
			9945: out = 16'(-4848);
			9946: out = 16'(7257);
			9947: out = 16'(7367);
			9948: out = 16'(3142);
			9949: out = 16'(-7089);
			9950: out = 16'(-9128);
			9951: out = 16'(-3901);
			9952: out = 16'(7085);
			9953: out = 16'(12962);
			9954: out = 16'(9862);
			9955: out = 16'(6002);
			9956: out = 16'(1356);
			9957: out = 16'(5471);
			9958: out = 16'(1578);
			9959: out = 16'(-116);
			9960: out = 16'(-10577);
			9961: out = 16'(-6411);
			9962: out = 16'(-1440);
			9963: out = 16'(7635);
			9964: out = 16'(6971);
			9965: out = 16'(3780);
			9966: out = 16'(-3526);
			9967: out = 16'(-5673);
			9968: out = 16'(-4989);
			9969: out = 16'(-602);
			9970: out = 16'(2138);
			9971: out = 16'(4859);
			9972: out = 16'(-3212);
			9973: out = 16'(-5474);
			9974: out = 16'(1569);
			9975: out = 16'(3230);
			9976: out = 16'(3108);
			9977: out = 16'(-8718);
			9978: out = 16'(-8214);
			9979: out = 16'(-6517);
			9980: out = 16'(1956);
			9981: out = 16'(2891);
			9982: out = 16'(2562);
			9983: out = 16'(1424);
			9984: out = 16'(1946);
			9985: out = 16'(3864);
			9986: out = 16'(-2425);
			9987: out = 16'(-3832);
			9988: out = 16'(-3612);
			9989: out = 16'(1715);
			9990: out = 16'(4598);
			9991: out = 16'(5687);
			9992: out = 16'(2795);
			9993: out = 16'(-875);
			9994: out = 16'(-7732);
			9995: out = 16'(-2952);
			9996: out = 16'(2922);
			9997: out = 16'(8986);
			9998: out = 16'(6415);
			9999: out = 16'(1003);
			10000: out = 16'(-500);
			10001: out = 16'(-1842);
			10002: out = 16'(67);
			10003: out = 16'(-7334);
			10004: out = 16'(-5506);
			10005: out = 16'(-1110);
			10006: out = 16'(2569);
			10007: out = 16'(3211);
			10008: out = 16'(1126);
			10009: out = 16'(650);
			10010: out = 16'(-1422);
			10011: out = 16'(-7931);
			10012: out = 16'(-3737);
			10013: out = 16'(404);
			10014: out = 16'(7834);
			10015: out = 16'(3687);
			10016: out = 16'(-1014);
			10017: out = 16'(-7143);
			10018: out = 16'(-3768);
			10019: out = 16'(2253);
			10020: out = 16'(-128);
			10021: out = 16'(-1610);
			10022: out = 16'(-5130);
			10023: out = 16'(3030);
			10024: out = 16'(7206);
			10025: out = 16'(11709);
			10026: out = 16'(6325);
			10027: out = 16'(1779);
			10028: out = 16'(-5527);
			10029: out = 16'(-4438);
			10030: out = 16'(-2891);
			10031: out = 16'(2429);
			10032: out = 16'(3374);
			10033: out = 16'(3585);
			10034: out = 16'(-7888);
			10035: out = 16'(-4986);
			10036: out = 16'(-1736);
			10037: out = 16'(8882);
			10038: out = 16'(7489);
			10039: out = 16'(4990);
			10040: out = 16'(-9746);
			10041: out = 16'(-7878);
			10042: out = 16'(1589);
			10043: out = 16'(6304);
			10044: out = 16'(4334);
			10045: out = 16'(-5755);
			10046: out = 16'(-10736);
			10047: out = 16'(-11197);
			10048: out = 16'(347);
			10049: out = 16'(3968);
			10050: out = 16'(6917);
			10051: out = 16'(1014);
			10052: out = 16'(379);
			10053: out = 16'(-1790);
			10054: out = 16'(1312);
			10055: out = 16'(284);
			10056: out = 16'(601);
			10057: out = 16'(2899);
			10058: out = 16'(2939);
			10059: out = 16'(129);
			10060: out = 16'(-1397);
			10061: out = 16'(-4195);
			10062: out = 16'(-4533);
			10063: out = 16'(-5957);
			10064: out = 16'(-754);
			10065: out = 16'(9696);
			10066: out = 16'(9877);
			10067: out = 16'(7359);
			10068: out = 16'(-54);
			10069: out = 16'(-4206);
			10070: out = 16'(-6560);
			10071: out = 16'(-2893);
			10072: out = 16'(-764);
			10073: out = 16'(1652);
			10074: out = 16'(810);
			10075: out = 16'(-417);
			10076: out = 16'(-2874);
			10077: out = 16'(2929);
			10078: out = 16'(2662);
			10079: out = 16'(1138);
			10080: out = 16'(-88);
			10081: out = 16'(881);
			10082: out = 16'(4690);
			10083: out = 16'(1184);
			10084: out = 16'(-2036);
			10085: out = 16'(-9482);
			10086: out = 16'(-2592);
			10087: out = 16'(1477);
			10088: out = 16'(-3043);
			10089: out = 16'(-1089);
			10090: out = 16'(298);
			10091: out = 16'(4461);
			10092: out = 16'(2879);
			10093: out = 16'(769);
			10094: out = 16'(4293);
			10095: out = 16'(2703);
			10096: out = 16'(-520);
			10097: out = 16'(-144);
			10098: out = 16'(-14);
			10099: out = 16'(2663);
			10100: out = 16'(-3877);
			10101: out = 16'(-4158);
			10102: out = 16'(49);
			10103: out = 16'(2967);
			10104: out = 16'(3685);
			10105: out = 16'(-1877);
			10106: out = 16'(-108);
			10107: out = 16'(375);
			10108: out = 16'(-2860);
			10109: out = 16'(-860);
			10110: out = 16'(2035);
			10111: out = 16'(6632);
			10112: out = 16'(7656);
			10113: out = 16'(6513);
			10114: out = 16'(1206);
			10115: out = 16'(-4420);
			10116: out = 16'(-11308);
			10117: out = 16'(-4522);
			10118: out = 16'(-2164);
			10119: out = 16'(-151);
			10120: out = 16'(-4320);
			10121: out = 16'(-3140);
			10122: out = 16'(4522);
			10123: out = 16'(7581);
			10124: out = 16'(8358);
			10125: out = 16'(724);
			10126: out = 16'(396);
			10127: out = 16'(-1996);
			10128: out = 16'(-7146);
			10129: out = 16'(-10352);
			10130: out = 16'(-10974);
			10131: out = 16'(584);
			10132: out = 16'(3061);
			10133: out = 16'(2113);
			10134: out = 16'(2603);
			10135: out = 16'(3080);
			10136: out = 16'(5963);
			10137: out = 16'(1795);
			10138: out = 16'(528);
			10139: out = 16'(-2144);
			10140: out = 16'(2158);
			10141: out = 16'(2452);
			10142: out = 16'(163);
			10143: out = 16'(-3486);
			10144: out = 16'(-5943);
			10145: out = 16'(-9325);
			10146: out = 16'(-4216);
			10147: out = 16'(1678);
			10148: out = 16'(9763);
			10149: out = 16'(6575);
			10150: out = 16'(111);
			10151: out = 16'(-876);
			10152: out = 16'(-1537);
			10153: out = 16'(-180);
			10154: out = 16'(2595);
			10155: out = 16'(2017);
			10156: out = 16'(-1969);
			10157: out = 16'(-6139);
			10158: out = 16'(-6297);
			10159: out = 16'(3092);
			10160: out = 16'(-590);
			10161: out = 16'(-1504);
			10162: out = 16'(-3060);
			10163: out = 16'(2216);
			10164: out = 16'(4906);
			10165: out = 16'(-7592);
			10166: out = 16'(-3544);
			10167: out = 16'(2024);
			10168: out = 16'(6951);
			10169: out = 16'(4394);
			10170: out = 16'(-2802);
			10171: out = 16'(-3835);
			10172: out = 16'(-5730);
			10173: out = 16'(-2953);
			10174: out = 16'(-7658);
			10175: out = 16'(-5265);
			10176: out = 16'(-1465);
			10177: out = 16'(7653);
			10178: out = 16'(10328);
			10179: out = 16'(6878);
			10180: out = 16'(1840);
			10181: out = 16'(-1772);
			10182: out = 16'(243);
			10183: out = 16'(629);
			10184: out = 16'(1557);
			10185: out = 16'(4400);
			10186: out = 16'(2856);
			10187: out = 16'(646);
			10188: out = 16'(-5488);
			10189: out = 16'(-6517);
			10190: out = 16'(-6164);
			10191: out = 16'(6464);
			10192: out = 16'(10116);
			10193: out = 16'(10297);
			10194: out = 16'(-2882);
			10195: out = 16'(-7697);
			10196: out = 16'(-1185);
			10197: out = 16'(2626);
			10198: out = 16'(5105);
			10199: out = 16'(-577);
			10200: out = 16'(-4404);
			10201: out = 16'(-7595);
			10202: out = 16'(1919);
			10203: out = 16'(5798);
			10204: out = 16'(10206);
			10205: out = 16'(-5502);
			10206: out = 16'(-5134);
			10207: out = 16'(-2430);
			10208: out = 16'(8242);
			10209: out = 16'(7246);
			10210: out = 16'(-1682);
			10211: out = 16'(2056);
			10212: out = 16'(622);
			10213: out = 16'(-1646);
			10214: out = 16'(-3676);
			10215: out = 16'(-4373);
			10216: out = 16'(-5622);
			10217: out = 16'(-3074);
			10218: out = 16'(-467);
			10219: out = 16'(5276);
			10220: out = 16'(5190);
			10221: out = 16'(5072);
			10222: out = 16'(-1751);
			10223: out = 16'(1944);
			10224: out = 16'(6351);
			10225: out = 16'(6488);
			10226: out = 16'(1353);
			10227: out = 16'(-7779);
			10228: out = 16'(-6727);
			10229: out = 16'(-6575);
			10230: out = 16'(-5352);
			10231: out = 16'(-1241);
			10232: out = 16'(2071);
			10233: out = 16'(5514);
			10234: out = 16'(826);
			10235: out = 16'(-1731);
			10236: out = 16'(407);
			10237: out = 16'(4868);
			10238: out = 16'(7106);
			10239: out = 16'(-5744);
			10240: out = 16'(-9951);
			10241: out = 16'(-13094);
			10242: out = 16'(-900);
			10243: out = 16'(2605);
			10244: out = 16'(4570);
			10245: out = 16'(499);
			10246: out = 16'(-381);
			10247: out = 16'(77);
			10248: out = 16'(-20);
			10249: out = 16'(-778);
			10250: out = 16'(-4184);
			10251: out = 16'(240);
			10252: out = 16'(4067);
			10253: out = 16'(10359);
			10254: out = 16'(4171);
			10255: out = 16'(-2801);
			10256: out = 16'(-9434);
			10257: out = 16'(-10531);
			10258: out = 16'(-7080);
			10259: out = 16'(3539);
			10260: out = 16'(7425);
			10261: out = 16'(6910);
			10262: out = 16'(7303);
			10263: out = 16'(3406);
			10264: out = 16'(-305);
			10265: out = 16'(-5679);
			10266: out = 16'(-5183);
			10267: out = 16'(-11);
			10268: out = 16'(2242);
			10269: out = 16'(1519);
			10270: out = 16'(-7111);
			10271: out = 16'(-2854);
			10272: out = 16'(469);
			10273: out = 16'(1806);
			10274: out = 16'(2428);
			10275: out = 16'(1983);
			10276: out = 16'(4426);
			10277: out = 16'(2747);
			10278: out = 16'(1756);
			10279: out = 16'(-4972);
			10280: out = 16'(-3845);
			10281: out = 16'(-1660);
			10282: out = 16'(5262);
			10283: out = 16'(3980);
			10284: out = 16'(-329);
			10285: out = 16'(-8143);
			10286: out = 16'(-8662);
			10287: out = 16'(-1504);
			10288: out = 16'(5778);
			10289: out = 16'(8247);
			10290: out = 16'(468);
			10291: out = 16'(-2786);
			10292: out = 16'(-5057);
			10293: out = 16'(800);
			10294: out = 16'(3607);
			10295: out = 16'(6528);
			10296: out = 16'(5160);
			10297: out = 16'(2593);
			10298: out = 16'(-1726);
			10299: out = 16'(-10269);
			10300: out = 16'(-7884);
			10301: out = 16'(3687);
			10302: out = 16'(1860);
			10303: out = 16'(2668);
			10304: out = 16'(-4405);
			10305: out = 16'(6310);
			10306: out = 16'(5344);
			10307: out = 16'(-1102);
			10308: out = 16'(-10631);
			10309: out = 16'(-12491);
			10310: out = 16'(1621);
			10311: out = 16'(6885);
			10312: out = 16'(9146);
			10313: out = 16'(-723);
			10314: out = 16'(-7792);
			10315: out = 16'(-14612);
			10316: out = 16'(662);
			10317: out = 16'(4767);
			10318: out = 16'(8677);
			10319: out = 16'(-412);
			10320: out = 16'(170);
			10321: out = 16'(4482);
			10322: out = 16'(628);
			10323: out = 16'(-1197);
			10324: out = 16'(-1563);
			10325: out = 16'(-2598);
			10326: out = 16'(-3587);
			10327: out = 16'(-8153);
			10328: out = 16'(-1564);
			10329: out = 16'(2771);
			10330: out = 16'(-106);
			10331: out = 16'(-1052);
			10332: out = 16'(-2249);
			10333: out = 16'(6139);
			10334: out = 16'(6230);
			10335: out = 16'(6034);
			10336: out = 16'(-3957);
			10337: out = 16'(-3806);
			10338: out = 16'(-85);
			10339: out = 16'(363);
			10340: out = 16'(561);
			10341: out = 16'(-107);
			10342: out = 16'(-1168);
			10343: out = 16'(-2073);
			10344: out = 16'(-4226);
			10345: out = 16'(1634);
			10346: out = 16'(4470);
			10347: out = 16'(2101);
			10348: out = 16'(102);
			10349: out = 16'(-1371);
			10350: out = 16'(3000);
			10351: out = 16'(5547);
			10352: out = 16'(7569);
			10353: out = 16'(-2920);
			10354: out = 16'(-7882);
			10355: out = 16'(-13411);
			10356: out = 16'(2656);
			10357: out = 16'(7181);
			10358: out = 16'(10332);
			10359: out = 16'(-3211);
			10360: out = 16'(-4965);
			10361: out = 16'(2555);
			10362: out = 16'(6146);
			10363: out = 16'(5371);
			10364: out = 16'(-9937);
			10365: out = 16'(-4864);
			10366: out = 16'(-2130);
			10367: out = 16'(2295);
			10368: out = 16'(661);
			10369: out = 16'(92);
			10370: out = 16'(718);
			10371: out = 16'(702);
			10372: out = 16'(-958);
			10373: out = 16'(931);
			10374: out = 16'(1676);
			10375: out = 16'(6011);
			10376: out = 16'(-8369);
			10377: out = 16'(-7304);
			10378: out = 16'(-435);
			10379: out = 16'(7242);
			10380: out = 16'(6058);
			10381: out = 16'(-3963);
			10382: out = 16'(-9293);
			10383: out = 16'(-10408);
			10384: out = 16'(-4498);
			10385: out = 16'(5865);
			10386: out = 16'(12029);
			10387: out = 16'(7115);
			10388: out = 16'(-4925);
			10389: out = 16'(-18205);
			10390: out = 16'(-1192);
			10391: out = 16'(4889);
			10392: out = 16'(12878);
			10393: out = 16'(885);
			10394: out = 16'(-1006);
			10395: out = 16'(-3343);
			10396: out = 16'(-392);
			10397: out = 16'(-1386);
			10398: out = 16'(-2279);
			10399: out = 16'(-5653);
			10400: out = 16'(-4592);
			10401: out = 16'(1085);
			10402: out = 16'(5907);
			10403: out = 16'(6519);
			10404: out = 16'(-10075);
			10405: out = 16'(-4866);
			10406: out = 16'(925);
			10407: out = 16'(1898);
			10408: out = 16'(2344);
			10409: out = 16'(920);
			10410: out = 16'(3906);
			10411: out = 16'(-2010);
			10412: out = 16'(-12132);
			10413: out = 16'(-2130);
			10414: out = 16'(2455);
			10415: out = 16'(8248);
			10416: out = 16'(-1791);
			10417: out = 16'(-4394);
			10418: out = 16'(253);
			10419: out = 16'(1383);
			10420: out = 16'(2704);
			10421: out = 16'(642);
			10422: out = 16'(3825);
			10423: out = 16'(5042);
			10424: out = 16'(-1344);
			10425: out = 16'(419);
			10426: out = 16'(2823);
			10427: out = 16'(6895);
			10428: out = 16'(4735);
			10429: out = 16'(-116);
			10430: out = 16'(-219);
			10431: out = 16'(1808);
			10432: out = 16'(8893);
			10433: out = 16'(1418);
			10434: out = 16'(-218);
			10435: out = 16'(-3937);
			10436: out = 16'(3210);
			10437: out = 16'(4543);
			10438: out = 16'(5697);
			10439: out = 16'(-5143);
			10440: out = 16'(-11258);
			10441: out = 16'(-11241);
			10442: out = 16'(1514);
			10443: out = 16'(12613);
			10444: out = 16'(4097);
			10445: out = 16'(-2431);
			10446: out = 16'(-12977);
			10447: out = 16'(5879);
			10448: out = 16'(4719);
			10449: out = 16'(1696);
			10450: out = 16'(-8491);
			10451: out = 16'(-7910);
			10452: out = 16'(1473);
			10453: out = 16'(-1712);
			10454: out = 16'(-689);
			10455: out = 16'(724);
			10456: out = 16'(2739);
			10457: out = 16'(2174);
			10458: out = 16'(-1381);
			10459: out = 16'(-4052);
			10460: out = 16'(-4133);
			10461: out = 16'(4775);
			10462: out = 16'(4912);
			10463: out = 16'(3385);
			10464: out = 16'(-828);
			10465: out = 16'(-3205);
			10466: out = 16'(-3927);
			10467: out = 16'(-3408);
			10468: out = 16'(-1693);
			10469: out = 16'(-550);
			10470: out = 16'(2715);
			10471: out = 16'(3013);
			10472: out = 16'(3513);
			10473: out = 16'(-4664);
			10474: out = 16'(-8041);
			10475: out = 16'(-6507);
			10476: out = 16'(321);
			10477: out = 16'(4240);
			10478: out = 16'(-4032);
			10479: out = 16'(-3497);
			10480: out = 16'(-3269);
			10481: out = 16'(3290);
			10482: out = 16'(2505);
			10483: out = 16'(1045);
			10484: out = 16'(156);
			10485: out = 16'(-1260);
			10486: out = 16'(-2701);
			10487: out = 16'(-4515);
			10488: out = 16'(-3948);
			10489: out = 16'(-824);
			10490: out = 16'(1353);
			10491: out = 16'(2604);
			10492: out = 16'(-272);
			10493: out = 16'(2968);
			10494: out = 16'(2726);
			10495: out = 16'(228);
			10496: out = 16'(-1932);
			10497: out = 16'(-1423);
			10498: out = 16'(3826);
			10499: out = 16'(7326);
			10500: out = 16'(8563);
			10501: out = 16'(1879);
			10502: out = 16'(-2756);
			10503: out = 16'(-6606);
			10504: out = 16'(-3704);
			10505: out = 16'(1328);
			10506: out = 16'(8813);
			10507: out = 16'(3308);
			10508: out = 16'(323);
			10509: out = 16'(-4358);
			10510: out = 16'(-1553);
			10511: out = 16'(910);
			10512: out = 16'(5345);
			10513: out = 16'(3977);
			10514: out = 16'(864);
			10515: out = 16'(-11596);
			10516: out = 16'(-7854);
			10517: out = 16'(-1533);
			10518: out = 16'(9735);
			10519: out = 16'(10600);
			10520: out = 16'(7597);
			10521: out = 16'(-968);
			10522: out = 16'(-5736);
			10523: out = 16'(-7843);
			10524: out = 16'(-4083);
			10525: out = 16'(-3063);
			10526: out = 16'(-5627);
			10527: out = 16'(-1021);
			10528: out = 16'(1542);
			10529: out = 16'(7020);
			10530: out = 16'(2183);
			10531: out = 16'(359);
			10532: out = 16'(-2122);
			10533: out = 16'(1656);
			10534: out = 16'(3557);
			10535: out = 16'(8645);
			10536: out = 16'(1297);
			10537: out = 16'(-4978);
			10538: out = 16'(-8105);
			10539: out = 16'(-2536);
			10540: out = 16'(5155);
			10541: out = 16'(10088);
			10542: out = 16'(6412);
			10543: out = 16'(-2919);
			10544: out = 16'(-7538);
			10545: out = 16'(-6442);
			10546: out = 16'(4023);
			10547: out = 16'(4836);
			10548: out = 16'(3654);
			10549: out = 16'(-10240);
			10550: out = 16'(-4685);
			10551: out = 16'(-1774);
			10552: out = 16'(5648);
			10553: out = 16'(1594);
			10554: out = 16'(-328);
			10555: out = 16'(1574);
			10556: out = 16'(3278);
			10557: out = 16'(3351);
			10558: out = 16'(-1807);
			10559: out = 16'(-4227);
			10560: out = 16'(-3803);
			10561: out = 16'(-10107);
			10562: out = 16'(-6454);
			10563: out = 16'(1608);
			10564: out = 16'(6640);
			10565: out = 16'(6418);
			10566: out = 16'(-934);
			10567: out = 16'(-3480);
			10568: out = 16'(-4831);
			10569: out = 16'(287);
			10570: out = 16'(1565);
			10571: out = 16'(3428);
			10572: out = 16'(-811);
			10573: out = 16'(182);
			10574: out = 16'(-269);
			10575: out = 16'(3463);
			10576: out = 16'(756);
			10577: out = 16'(-1726);
			10578: out = 16'(-1931);
			10579: out = 16'(-401);
			10580: out = 16'(1012);
			10581: out = 16'(5483);
			10582: out = 16'(4557);
			10583: out = 16'(327);
			10584: out = 16'(-5659);
			10585: out = 16'(-5559);
			10586: out = 16'(7201);
			10587: out = 16'(1396);
			10588: out = 16'(-567);
			10589: out = 16'(-3283);
			10590: out = 16'(122);
			10591: out = 16'(2003);
			10592: out = 16'(717);
			10593: out = 16'(303);
			10594: out = 16'(846);
			10595: out = 16'(1571);
			10596: out = 16'(955);
			10597: out = 16'(-2498);
			10598: out = 16'(5826);
			10599: out = 16'(1807);
			10600: out = 16'(-5697);
			10601: out = 16'(-11820);
			10602: out = 16'(-10035);
			10603: out = 16'(392);
			10604: out = 16'(5565);
			10605: out = 16'(7747);
			10606: out = 16'(1646);
			10607: out = 16'(2332);
			10608: out = 16'(1189);
			10609: out = 16'(-2854);
			10610: out = 16'(-1504);
			10611: out = 16'(445);
			10612: out = 16'(7017);
			10613: out = 16'(2522);
			10614: out = 16'(-4128);
			10615: out = 16'(-10696);
			10616: out = 16'(-7700);
			10617: out = 16'(2356);
			10618: out = 16'(434);
			10619: out = 16'(318);
			10620: out = 16'(-4675);
			10621: out = 16'(2621);
			10622: out = 16'(4647);
			10623: out = 16'(5480);
			10624: out = 16'(741);
			10625: out = 16'(-2011);
			10626: out = 16'(-177);
			10627: out = 16'(147);
			10628: out = 16'(951);
			10629: out = 16'(-4151);
			10630: out = 16'(-2407);
			10631: out = 16'(-1208);
			10632: out = 16'(6200);
			10633: out = 16'(2836);
			10634: out = 16'(-2217);
			10635: out = 16'(-12430);
			10636: out = 16'(-9917);
			10637: out = 16'(2378);
			10638: out = 16'(2248);
			10639: out = 16'(3705);
			10640: out = 16'(222);
			10641: out = 16'(1991);
			10642: out = 16'(-687);
			10643: out = 16'(-5734);
			10644: out = 16'(-5905);
			10645: out = 16'(-3184);
			10646: out = 16'(1894);
			10647: out = 16'(3581);
			10648: out = 16'(3583);
			10649: out = 16'(6748);
			10650: out = 16'(5661);
			10651: out = 16'(5297);
			10652: out = 16'(-2016);
			10653: out = 16'(-2101);
			10654: out = 16'(-1603);
			10655: out = 16'(9040);
			10656: out = 16'(8561);
			10657: out = 16'(2857);
			10658: out = 16'(-8646);
			10659: out = 16'(-10776);
			10660: out = 16'(4167);
			10661: out = 16'(3807);
			10662: out = 16'(4761);
			10663: out = 16'(-3504);
			10664: out = 16'(-279);
			10665: out = 16'(2003);
			10666: out = 16'(12264);
			10667: out = 16'(9009);
			10668: out = 16'(4597);
			10669: out = 16'(-4134);
			10670: out = 16'(-8010);
			10671: out = 16'(-10760);
			10672: out = 16'(-2051);
			10673: out = 16'(511);
			10674: out = 16'(2146);
			10675: out = 16'(-8410);
			10676: out = 16'(-11375);
			10677: out = 16'(-7389);
			10678: out = 16'(1602);
			10679: out = 16'(7319);
			10680: out = 16'(2515);
			10681: out = 16'(2178);
			10682: out = 16'(-774);
			10683: out = 16'(4316);
			10684: out = 16'(-2395);
			10685: out = 16'(-6907);
			10686: out = 16'(-12968);
			10687: out = 16'(-5336);
			10688: out = 16'(5944);
			10689: out = 16'(2174);
			10690: out = 16'(2444);
			10691: out = 16'(635);
			10692: out = 16'(4082);
			10693: out = 16'(4074);
			10694: out = 16'(3382);
			10695: out = 16'(3244);
			10696: out = 16'(2348);
			10697: out = 16'(-1876);
			10698: out = 16'(-709);
			10699: out = 16'(-243);
			10700: out = 16'(2357);
			10701: out = 16'(1092);
			10702: out = 16'(64);
			10703: out = 16'(-7685);
			10704: out = 16'(-4052);
			10705: out = 16'(942);
			10706: out = 16'(7214);
			10707: out = 16'(6822);
			10708: out = 16'(3349);
			10709: out = 16'(-5216);
			10710: out = 16'(-10225);
			10711: out = 16'(-13131);
			10712: out = 16'(-3808);
			10713: out = 16'(363);
			10714: out = 16'(-1630);
			10715: out = 16'(-5189);
			10716: out = 16'(-5177);
			10717: out = 16'(10412);
			10718: out = 16'(3567);
			10719: out = 16'(-1169);
			10720: out = 16'(-9848);
			10721: out = 16'(-4415);
			10722: out = 16'(3181);
			10723: out = 16'(6467);
			10724: out = 16'(8727);
			10725: out = 16'(7374);
			10726: out = 16'(794);
			10727: out = 16'(-4266);
			10728: out = 16'(-5899);
			10729: out = 16'(-9045);
			10730: out = 16'(-5381);
			10731: out = 16'(1441);
			10732: out = 16'(7599);
			10733: out = 16'(7127);
			10734: out = 16'(-4116);
			10735: out = 16'(-1237);
			10736: out = 16'(1625);
			10737: out = 16'(7216);
			10738: out = 16'(6632);
			10739: out = 16'(4370);
			10740: out = 16'(3063);
			10741: out = 16'(-3006);
			10742: out = 16'(-8132);
			10743: out = 16'(-5829);
			10744: out = 16'(-1607);
			10745: out = 16'(3700);
			10746: out = 16'(587);
			10747: out = 16'(-3551);
			10748: out = 16'(-10458);
			10749: out = 16'(-4709);
			10750: out = 16'(818);
			10751: out = 16'(7671);
			10752: out = 16'(8009);
			10753: out = 16'(4528);
			10754: out = 16'(-7440);
			10755: out = 16'(-8467);
			10756: out = 16'(-7535);
			10757: out = 16'(-36);
			10758: out = 16'(894);
			10759: out = 16'(1493);
			10760: out = 16'(3418);
			10761: out = 16'(5323);
			10762: out = 16'(7627);
			10763: out = 16'(-2620);
			10764: out = 16'(-1997);
			10765: out = 16'(1626);
			10766: out = 16'(7756);
			10767: out = 16'(7486);
			10768: out = 16'(1571);
			10769: out = 16'(-1175);
			10770: out = 16'(-2755);
			10771: out = 16'(1072);
			10772: out = 16'(247);
			10773: out = 16'(825);
			10774: out = 16'(-439);
			10775: out = 16'(1202);
			10776: out = 16'(2070);
			10777: out = 16'(715);
			10778: out = 16'(4291);
			10779: out = 16'(7922);
			10780: out = 16'(-1210);
			10781: out = 16'(-2801);
			10782: out = 16'(-4680);
			10783: out = 16'(594);
			10784: out = 16'(-2247);
			10785: out = 16'(-8220);
			10786: out = 16'(-10078);
			10787: out = 16'(-6896);
			10788: out = 16'(4149);
			10789: out = 16'(3014);
			10790: out = 16'(2779);
			10791: out = 16'(-3362);
			10792: out = 16'(3392);
			10793: out = 16'(5927);
			10794: out = 16'(1388);
			10795: out = 16'(-3513);
			10796: out = 16'(-7629);
			10797: out = 16'(4127);
			10798: out = 16'(2016);
			10799: out = 16'(-815);
			10800: out = 16'(-8040);
			10801: out = 16'(-5012);
			10802: out = 16'(3385);
			10803: out = 16'(-11);
			10804: out = 16'(573);
			10805: out = 16'(-237);
			10806: out = 16'(6628);
			10807: out = 16'(5956);
			10808: out = 16'(-4590);
			10809: out = 16'(408);
			10810: out = 16'(2954);
			10811: out = 16'(6631);
			10812: out = 16'(-323);
			10813: out = 16'(-5799);
			10814: out = 16'(-200);
			10815: out = 16'(-635);
			10816: out = 16'(77);
			10817: out = 16'(-3918);
			10818: out = 16'(-3568);
			10819: out = 16'(-3845);
			10820: out = 16'(2712);
			10821: out = 16'(3184);
			10822: out = 16'(3658);
			10823: out = 16'(-9434);
			10824: out = 16'(-10239);
			10825: out = 16'(716);
			10826: out = 16'(4363);
			10827: out = 16'(4764);
			10828: out = 16'(-9644);
			10829: out = 16'(-2369);
			10830: out = 16'(947);
			10831: out = 16'(5217);
			10832: out = 16'(-1271);
			10833: out = 16'(-5552);
			10834: out = 16'(3989);
			10835: out = 16'(6187);
			10836: out = 16'(7290);
			10837: out = 16'(-127);
			10838: out = 16'(-1763);
			10839: out = 16'(-1142);
			10840: out = 16'(-2639);
			10841: out = 16'(-1279);
			10842: out = 16'(1011);
			10843: out = 16'(3736);
			10844: out = 16'(3576);
			10845: out = 16'(-416);
			10846: out = 16'(-988);
			10847: out = 16'(-745);
			10848: out = 16'(3507);
			10849: out = 16'(3172);
			10850: out = 16'(3754);
			10851: out = 16'(6070);
			10852: out = 16'(4387);
			10853: out = 16'(1047);
			10854: out = 16'(386);
			10855: out = 16'(-4584);
			10856: out = 16'(-9153);
			10857: out = 16'(-6308);
			10858: out = 16'(-123);
			10859: out = 16'(10005);
			10860: out = 16'(1675);
			10861: out = 16'(-1813);
			10862: out = 16'(-6911);
			10863: out = 16'(-333);
			10864: out = 16'(3893);
			10865: out = 16'(9304);
			10866: out = 16'(4629);
			10867: out = 16'(-177);
			10868: out = 16'(-11675);
			10869: out = 16'(-5962);
			10870: out = 16'(1242);
			10871: out = 16'(7432);
			10872: out = 16'(4608);
			10873: out = 16'(-1621);
			10874: out = 16'(-2149);
			10875: out = 16'(-2338);
			10876: out = 16'(488);
			10877: out = 16'(2039);
			10878: out = 16'(3615);
			10879: out = 16'(2626);
			10880: out = 16'(833);
			10881: out = 16'(-1594);
			10882: out = 16'(-1319);
			10883: out = 16'(-1331);
			10884: out = 16'(500);
			10885: out = 16'(-1163);
			10886: out = 16'(5173);
			10887: out = 16'(6611);
			10888: out = 16'(-1925);
			10889: out = 16'(-8418);
			10890: out = 16'(-12679);
			10891: out = 16'(264);
			10892: out = 16'(5464);
			10893: out = 16'(8944);
			10894: out = 16'(1023);
			10895: out = 16'(-1141);
			10896: out = 16'(-33);
			10897: out = 16'(-7317);
			10898: out = 16'(-9077);
			10899: out = 16'(-7802);
			10900: out = 16'(-1724);
			10901: out = 16'(2505);
			10902: out = 16'(4263);
			10903: out = 16'(3164);
			10904: out = 16'(1808);
			10905: out = 16'(-247);
			10906: out = 16'(3454);
			10907: out = 16'(6009);
			10908: out = 16'(1583);
			10909: out = 16'(-4663);
			10910: out = 16'(-12294);
			10911: out = 16'(-454);
			10912: out = 16'(1338);
			10913: out = 16'(2478);
			10914: out = 16'(-1021);
			10915: out = 16'(-843);
			10916: out = 16'(888);
			10917: out = 16'(903);
			10918: out = 16'(2711);
			10919: out = 16'(8461);
			10920: out = 16'(6041);
			10921: out = 16'(2656);
			10922: out = 16'(-10916);
			10923: out = 16'(-4615);
			10924: out = 16'(693);
			10925: out = 16'(7325);
			10926: out = 16'(-167);
			10927: out = 16'(-8680);
			10928: out = 16'(-1982);
			10929: out = 16'(-167);
			10930: out = 16'(2445);
			10931: out = 16'(1183);
			10932: out = 16'(-984);
			10933: out = 16'(-5635);
			10934: out = 16'(-4240);
			10935: out = 16'(-1250);
			10936: out = 16'(7120);
			10937: out = 16'(3112);
			10938: out = 16'(693);
			10939: out = 16'(-7093);
			10940: out = 16'(545);
			10941: out = 16'(4249);
			10942: out = 16'(-139);
			10943: out = 16'(-173);
			10944: out = 16'(-590);
			10945: out = 16'(-1567);
			10946: out = 16'(-829);
			10947: out = 16'(319);
			10948: out = 16'(4793);
			10949: out = 16'(2943);
			10950: out = 16'(-2322);
			10951: out = 16'(647);
			10952: out = 16'(113);
			10953: out = 16'(81);
			10954: out = 16'(-5946);
			10955: out = 16'(-6204);
			10956: out = 16'(1857);
			10957: out = 16'(-1839);
			10958: out = 16'(-1978);
			10959: out = 16'(-737);
			10960: out = 16'(5507);
			10961: out = 16'(9213);
			10962: out = 16'(2948);
			10963: out = 16'(5401);
			10964: out = 16'(5882);
			10965: out = 16'(-8581);
			10966: out = 16'(-12177);
			10967: out = 16'(-12350);
			10968: out = 16'(1388);
			10969: out = 16'(6015);
			10970: out = 16'(5995);
			10971: out = 16'(682);
			10972: out = 16'(-2670);
			10973: out = 16'(-2247);
			10974: out = 16'(-1399);
			10975: out = 16'(2011);
			10976: out = 16'(5928);
			10977: out = 16'(6197);
			10978: out = 16'(3051);
			10979: out = 16'(-4456);
			10980: out = 16'(-8602);
			10981: out = 16'(-9096);
			10982: out = 16'(2321);
			10983: out = 16'(2319);
			10984: out = 16'(-620);
			10985: out = 16'(1648);
			10986: out = 16'(469);
			10987: out = 16'(1572);
			10988: out = 16'(-9950);
			10989: out = 16'(-8006);
			10990: out = 16'(264);
			10991: out = 16'(7276);
			10992: out = 16'(7204);
			10993: out = 16'(-1749);
			10994: out = 16'(-6098);
			10995: out = 16'(-7748);
			10996: out = 16'(1412);
			10997: out = 16'(996);
			10998: out = 16'(1530);
			10999: out = 16'(-173);
			11000: out = 16'(169);
			11001: out = 16'(283);
			11002: out = 16'(-196);
			11003: out = 16'(490);
			11004: out = 16'(1141);
			11005: out = 16'(6090);
			11006: out = 16'(4507);
			11007: out = 16'(533);
			11008: out = 16'(-2995);
			11009: out = 16'(-2024);
			11010: out = 16'(3761);
			11011: out = 16'(4657);
			11012: out = 16'(4622);
			11013: out = 16'(812);
			11014: out = 16'(829);
			11015: out = 16'(569);
			11016: out = 16'(344);
			11017: out = 16'(4272);
			11018: out = 16'(7119);
			11019: out = 16'(3001);
			11020: out = 16'(1407);
			11021: out = 16'(-1110);
			11022: out = 16'(-2578);
			11023: out = 16'(-3076);
			11024: out = 16'(-1565);
			11025: out = 16'(-3294);
			11026: out = 16'(-1267);
			11027: out = 16'(2082);
			11028: out = 16'(1999);
			11029: out = 16'(205);
			11030: out = 16'(-5836);
			11031: out = 16'(-2940);
			11032: out = 16'(444);
			11033: out = 16'(10267);
			11034: out = 16'(6026);
			11035: out = 16'(1821);
			11036: out = 16'(-13386);
			11037: out = 16'(-6048);
			11038: out = 16'(1765);
			11039: out = 16'(2083);
			11040: out = 16'(-3732);
			11041: out = 16'(-12621);
			11042: out = 16'(-8316);
			11043: out = 16'(-2045);
			11044: out = 16'(9755);
			11045: out = 16'(2898);
			11046: out = 16'(428);
			11047: out = 16'(-7437);
			11048: out = 16'(1474);
			11049: out = 16'(3153);
			11050: out = 16'(4038);
			11051: out = 16'(-5548);
			11052: out = 16'(-10028);
			11053: out = 16'(-5069);
			11054: out = 16'(-214);
			11055: out = 16'(4452);
			11056: out = 16'(3267);
			11057: out = 16'(2191);
			11058: out = 16'(-830);
			11059: out = 16'(-847);
			11060: out = 16'(-639);
			11061: out = 16'(1796);
			11062: out = 16'(-1058);
			11063: out = 16'(-3149);
			11064: out = 16'(-9169);
			11065: out = 16'(-476);
			11066: out = 16'(3605);
			11067: out = 16'(11247);
			11068: out = 16'(-597);
			11069: out = 16'(-6162);
			11070: out = 16'(-11826);
			11071: out = 16'(2261);
			11072: out = 16'(11305);
			11073: out = 16'(8289);
			11074: out = 16'(1769);
			11075: out = 16'(-5861);
			11076: out = 16'(-2166);
			11077: out = 16'(-580);
			11078: out = 16'(3181);
			11079: out = 16'(3896);
			11080: out = 16'(3503);
			11081: out = 16'(713);
			11082: out = 16'(-4509);
			11083: out = 16'(-3149);
			11084: out = 16'(7578);
			11085: out = 16'(4103);
			11086: out = 16'(3076);
			11087: out = 16'(-6208);
			11088: out = 16'(5414);
			11089: out = 16'(9350);
			11090: out = 16'(5391);
			11091: out = 16'(-821);
			11092: out = 16'(-5439);
			11093: out = 16'(368);
			11094: out = 16'(2531);
			11095: out = 16'(4943);
			11096: out = 16'(-3395);
			11097: out = 16'(-3234);
			11098: out = 16'(-1432);
			11099: out = 16'(1238);
			11100: out = 16'(1766);
			11101: out = 16'(233);
			11102: out = 16'(985);
			11103: out = 16'(1030);
			11104: out = 16'(3345);
			11105: out = 16'(-3560);
			11106: out = 16'(-7635);
			11107: out = 16'(-10135);
			11108: out = 16'(-4586);
			11109: out = 16'(1795);
			11110: out = 16'(7428);
			11111: out = 16'(4831);
			11112: out = 16'(-702);
			11113: out = 16'(-468);
			11114: out = 16'(-3881);
			11115: out = 16'(-4737);
			11116: out = 16'(-8885);
			11117: out = 16'(-3316);
			11118: out = 16'(6146);
			11119: out = 16'(3613);
			11120: out = 16'(2119);
			11121: out = 16'(-1714);
			11122: out = 16'(319);
			11123: out = 16'(846);
			11124: out = 16'(796);
			11125: out = 16'(375);
			11126: out = 16'(-120);
			11127: out = 16'(143);
			11128: out = 16'(-318);
			11129: out = 16'(56);
			11130: out = 16'(664);
			11131: out = 16'(4172);
			11132: out = 16'(6891);
			11133: out = 16'(902);
			11134: out = 16'(-3592);
			11135: out = 16'(-9112);
			11136: out = 16'(-1550);
			11137: out = 16'(1826);
			11138: out = 16'(5548);
			11139: out = 16'(1646);
			11140: out = 16'(604);
			11141: out = 16'(482);
			11142: out = 16'(2460);
			11143: out = 16'(2362);
			11144: out = 16'(-311);
			11145: out = 16'(-4058);
			11146: out = 16'(-5732);
			11147: out = 16'(3069);
			11148: out = 16'(1367);
			11149: out = 16'(-474);
			11150: out = 16'(-2488);
			11151: out = 16'(-1717);
			11152: out = 16'(190);
			11153: out = 16'(-1447);
			11154: out = 16'(-1789);
			11155: out = 16'(-2754);
			11156: out = 16'(1271);
			11157: out = 16'(2496);
			11158: out = 16'(3279);
			11159: out = 16'(465);
			11160: out = 16'(-426);
			11161: out = 16'(532);
			11162: out = 16'(2182);
			11163: out = 16'(3076);
			11164: out = 16'(3031);
			11165: out = 16'(1120);
			11166: out = 16'(-844);
			11167: out = 16'(-2822);
			11168: out = 16'(-1834);
			11169: out = 16'(271);
			11170: out = 16'(4224);
			11171: out = 16'(4690);
			11172: out = 16'(3422);
			11173: out = 16'(-2745);
			11174: out = 16'(-2971);
			11175: out = 16'(2421);
			11176: out = 16'(1387);
			11177: out = 16'(-291);
			11178: out = 16'(-10138);
			11179: out = 16'(-2281);
			11180: out = 16'(2163);
			11181: out = 16'(10237);
			11182: out = 16'(1734);
			11183: out = 16'(-4682);
			11184: out = 16'(-11755);
			11185: out = 16'(-5413);
			11186: out = 16'(2428);
			11187: out = 16'(7202);
			11188: out = 16'(3625);
			11189: out = 16'(-4184);
			11190: out = 16'(-3360);
			11191: out = 16'(-4148);
			11192: out = 16'(-2339);
			11193: out = 16'(-446);
			11194: out = 16'(790);
			11195: out = 16'(-799);
			11196: out = 16'(417);
			11197: out = 16'(2127);
			11198: out = 16'(8279);
			11199: out = 16'(4639);
			11200: out = 16'(859);
			11201: out = 16'(-8930);
			11202: out = 16'(-6437);
			11203: out = 16'(-2711);
			11204: out = 16'(3593);
			11205: out = 16'(2353);
			11206: out = 16'(-518);
			11207: out = 16'(3006);
			11208: out = 16'(3195);
			11209: out = 16'(4024);
			11210: out = 16'(-1898);
			11211: out = 16'(-4508);
			11212: out = 16'(-8188);
			11213: out = 16'(3117);
			11214: out = 16'(5760);
			11215: out = 16'(2815);
			11216: out = 16'(-3303);
			11217: out = 16'(-6335);
			11218: out = 16'(43);
			11219: out = 16'(-1051);
			11220: out = 16'(-16);
			11221: out = 16'(-993);
			11222: out = 16'(1291);
			11223: out = 16'(1529);
			11224: out = 16'(-931);
			11225: out = 16'(-3585);
			11226: out = 16'(-4843);
			11227: out = 16'(-1376);
			11228: out = 16'(1082);
			11229: out = 16'(2068);
			11230: out = 16'(5816);
			11231: out = 16'(4180);
			11232: out = 16'(-390);
			11233: out = 16'(-2976);
			11234: out = 16'(-3190);
			11235: out = 16'(802);
			11236: out = 16'(2194);
			11237: out = 16'(2757);
			11238: out = 16'(-206);
			11239: out = 16'(-2899);
			11240: out = 16'(-4641);
			11241: out = 16'(5210);
			11242: out = 16'(3256);
			11243: out = 16'(1978);
			11244: out = 16'(-831);
			11245: out = 16'(3088);
			11246: out = 16'(7880);
			11247: out = 16'(1709);
			11248: out = 16'(-3106);
			11249: out = 16'(-9509);
			11250: out = 16'(-4505);
			11251: out = 16'(18);
			11252: out = 16'(7506);
			11253: out = 16'(3163);
			11254: out = 16'(1094);
			11255: out = 16'(-2160);
			11256: out = 16'(2554);
			11257: out = 16'(4398);
			11258: out = 16'(-706);
			11259: out = 16'(-3129);
			11260: out = 16'(-5572);
			11261: out = 16'(-565);
			11262: out = 16'(-1426);
			11263: out = 16'(-1585);
			11264: out = 16'(-4095);
			11265: out = 16'(-2054);
			11266: out = 16'(844);
			11267: out = 16'(943);
			11268: out = 16'(1498);
			11269: out = 16'(3383);
			11270: out = 16'(411);
			11271: out = 16'(-1294);
			11272: out = 16'(-7262);
			11273: out = 16'(3834);
			11274: out = 16'(6278);
			11275: out = 16'(-3601);
			11276: out = 16'(-11488);
			11277: out = 16'(-14860);
			11278: out = 16'(9419);
			11279: out = 16'(10534);
			11280: out = 16'(11246);
			11281: out = 16'(23);
			11282: out = 16'(140);
			11283: out = 16'(23);
			11284: out = 16'(1441);
			11285: out = 16'(-769);
			11286: out = 16'(-1238);
			11287: out = 16'(-7256);
			11288: out = 16'(-5249);
			11289: out = 16'(-890);
			11290: out = 16'(8770);
			11291: out = 16'(9200);
			11292: out = 16'(881);
			11293: out = 16'(-8888);
			11294: out = 16'(-13374);
			11295: out = 16'(-1989);
			11296: out = 16'(5200);
			11297: out = 16'(10859);
			11298: out = 16'(2276);
			11299: out = 16'(-1101);
			11300: out = 16'(-5921);
			11301: out = 16'(-2889);
			11302: out = 16'(-789);
			11303: out = 16'(3778);
			11304: out = 16'(717);
			11305: out = 16'(154);
			11306: out = 16'(-2025);
			11307: out = 16'(2159);
			11308: out = 16'(2363);
			11309: out = 16'(-738);
			11310: out = 16'(467);
			11311: out = 16'(1681);
			11312: out = 16'(6258);
			11313: out = 16'(1883);
			11314: out = 16'(-1071);
			11315: out = 16'(-844);
			11316: out = 16'(1621);
			11317: out = 16'(3806);
			11318: out = 16'(819);
			11319: out = 16'(-3172);
			11320: out = 16'(-8194);
			11321: out = 16'(468);
			11322: out = 16'(3723);
			11323: out = 16'(7081);
			11324: out = 16'(694);
			11325: out = 16'(-1002);
			11326: out = 16'(-450);
			11327: out = 16'(1110);
			11328: out = 16'(-26);
			11329: out = 16'(-8416);
			11330: out = 16'(-4692);
			11331: out = 16'(-2297);
			11332: out = 16'(1061);
			11333: out = 16'(-3141);
			11334: out = 16'(-6252);
			11335: out = 16'(288);
			11336: out = 16'(1788);
			11337: out = 16'(3237);
			11338: out = 16'(-249);
			11339: out = 16'(-70);
			11340: out = 16'(573);
			11341: out = 16'(-303);
			11342: out = 16'(-516);
			11343: out = 16'(-27);
			11344: out = 16'(205);
			11345: out = 16'(769);
			11346: out = 16'(243);
			11347: out = 16'(2487);
			11348: out = 16'(1853);
			11349: out = 16'(-2725);
			11350: out = 16'(-5828);
			11351: out = 16'(-7066);
			11352: out = 16'(972);
			11353: out = 16'(299);
			11354: out = 16'(331);
			11355: out = 16'(1559);
			11356: out = 16'(4499);
			11357: out = 16'(6917);
			11358: out = 16'(583);
			11359: out = 16'(-576);
			11360: out = 16'(1092);
			11361: out = 16'(-6130);
			11362: out = 16'(-7622);
			11363: out = 16'(-6262);
			11364: out = 16'(993);
			11365: out = 16'(5162);
			11366: out = 16'(3638);
			11367: out = 16'(5219);
			11368: out = 16'(4094);
			11369: out = 16'(809);
			11370: out = 16'(-125);
			11371: out = 16'(-304);
			11372: out = 16'(-678);
			11373: out = 16'(-1616);
			11374: out = 16'(-3112);
			11375: out = 16'(439);
			11376: out = 16'(-535);
			11377: out = 16'(-1557);
			11378: out = 16'(-1187);
			11379: out = 16'(2388);
			11380: out = 16'(8087);
			11381: out = 16'(2531);
			11382: out = 16'(-148);
			11383: out = 16'(-35);
			11384: out = 16'(-2494);
			11385: out = 16'(-3006);
			11386: out = 16'(-4693);
			11387: out = 16'(2883);
			11388: out = 16'(6611);
			11389: out = 16'(1151);
			11390: out = 16'(-6068);
			11391: out = 16'(-12911);
			11392: out = 16'(4144);
			11393: out = 16'(7115);
			11394: out = 16'(10550);
			11395: out = 16'(-10338);
			11396: out = 16'(-10659);
			11397: out = 16'(-4524);
			11398: out = 16'(5968);
			11399: out = 16'(7955);
			11400: out = 16'(2291);
			11401: out = 16'(1022);
			11402: out = 16'(-3387);
			11403: out = 16'(-11760);
			11404: out = 16'(-4028);
			11405: out = 16'(2744);
			11406: out = 16'(6852);
			11407: out = 16'(2000);
			11408: out = 16'(-3382);
			11409: out = 16'(3552);
			11410: out = 16'(1487);
			11411: out = 16'(798);
			11412: out = 16'(-4958);
			11413: out = 16'(-3157);
			11414: out = 16'(166);
			11415: out = 16'(-282);
			11416: out = 16'(888);
			11417: out = 16'(3326);
			11418: out = 16'(-1390);
			11419: out = 16'(-3853);
			11420: out = 16'(-6566);
			11421: out = 16'(-421);
			11422: out = 16'(1754);
			11423: out = 16'(-4180);
			11424: out = 16'(-1460);
			11425: out = 16'(340);
			11426: out = 16'(3327);
			11427: out = 16'(1647);
			11428: out = 16'(-232);
			11429: out = 16'(1014);
			11430: out = 16'(-898);
			11431: out = 16'(-2586);
			11432: out = 16'(503);
			11433: out = 16'(3078);
			11434: out = 16'(6421);
			11435: out = 16'(-1059);
			11436: out = 16'(-2207);
			11437: out = 16'(1107);
			11438: out = 16'(1427);
			11439: out = 16'(1324);
			11440: out = 16'(-4711);
			11441: out = 16'(3763);
			11442: out = 16'(6639);
			11443: out = 16'(1999);
			11444: out = 16'(-692);
			11445: out = 16'(-3474);
			11446: out = 16'(-2557);
			11447: out = 16'(-4695);
			11448: out = 16'(-5762);
			11449: out = 16'(5111);
			11450: out = 16'(5457);
			11451: out = 16'(3689);
			11452: out = 16'(-3754);
			11453: out = 16'(-3279);
			11454: out = 16'(2708);
			11455: out = 16'(587);
			11456: out = 16'(707);
			11457: out = 16'(461);
			11458: out = 16'(138);
			11459: out = 16'(-334);
			11460: out = 16'(-570);
			11461: out = 16'(189);
			11462: out = 16'(-34);
			11463: out = 16'(-3836);
			11464: out = 16'(-2935);
			11465: out = 16'(-937);
			11466: out = 16'(-745);
			11467: out = 16'(3168);
			11468: out = 16'(6209);
			11469: out = 16'(6477);
			11470: out = 16'(1305);
			11471: out = 16'(-7373);
			11472: out = 16'(-4315);
			11473: out = 16'(-2694);
			11474: out = 16'(1512);
			11475: out = 16'(2013);
			11476: out = 16'(4518);
			11477: out = 16'(6636);
			11478: out = 16'(4796);
			11479: out = 16'(456);
			11480: out = 16'(-5945);
			11481: out = 16'(-8054);
			11482: out = 16'(-6073);
			11483: out = 16'(1925);
			11484: out = 16'(5631);
			11485: out = 16'(6467);
			11486: out = 16'(3784);
			11487: out = 16'(381);
			11488: out = 16'(-2057);
			11489: out = 16'(-8309);
			11490: out = 16'(-6608);
			11491: out = 16'(-1297);
			11492: out = 16'(4432);
			11493: out = 16'(4425);
			11494: out = 16'(-2189);
			11495: out = 16'(-3909);
			11496: out = 16'(-5145);
			11497: out = 16'(-2564);
			11498: out = 16'(-569);
			11499: out = 16'(1390);
			11500: out = 16'(-616);
			11501: out = 16'(46);
			11502: out = 16'(-97);
			11503: out = 16'(1251);
			11504: out = 16'(-1591);
			11505: out = 16'(-5012);
			11506: out = 16'(6297);
			11507: out = 16'(4488);
			11508: out = 16'(-627);
			11509: out = 16'(-4085);
			11510: out = 16'(-3293);
			11511: out = 16'(2821);
			11512: out = 16'(-898);
			11513: out = 16'(-504);
			11514: out = 16'(3532);
			11515: out = 16'(583);
			11516: out = 16'(-578);
			11517: out = 16'(-2053);
			11518: out = 16'(5356);
			11519: out = 16'(8681);
			11520: out = 16'(-4711);
			11521: out = 16'(-8276);
			11522: out = 16'(-10847);
			11523: out = 16'(4145);
			11524: out = 16'(5684);
			11525: out = 16'(6277);
			11526: out = 16'(-658);
			11527: out = 16'(-938);
			11528: out = 16'(-207);
			11529: out = 16'(4380);
			11530: out = 16'(2950);
			11531: out = 16'(-2934);
			11532: out = 16'(-7024);
			11533: out = 16'(-6743);
			11534: out = 16'(3756);
			11535: out = 16'(1675);
			11536: out = 16'(397);
			11537: out = 16'(-4977);
			11538: out = 16'(-3076);
			11539: out = 16'(-522);
			11540: out = 16'(2769);
			11541: out = 16'(4914);
			11542: out = 16'(5965);
			11543: out = 16'(1690);
			11544: out = 16'(-2540);
			11545: out = 16'(-7903);
			11546: out = 16'(-1341);
			11547: out = 16'(1985);
			11548: out = 16'(6731);
			11549: out = 16'(242);
			11550: out = 16'(-1452);
			11551: out = 16'(-536);
			11552: out = 16'(2754);
			11553: out = 16'(3544);
			11554: out = 16'(0);
			11555: out = 16'(-2982);
			11556: out = 16'(-5095);
			11557: out = 16'(-1667);
			11558: out = 16'(716);
			11559: out = 16'(3605);
			11560: out = 16'(613);
			11561: out = 16'(930);
			11562: out = 16'(402);
			11563: out = 16'(2272);
			11564: out = 16'(-426);
			11565: out = 16'(-5383);
			11566: out = 16'(-2456);
			11567: out = 16'(135);
			11568: out = 16'(4443);
			11569: out = 16'(1224);
			11570: out = 16'(-1185);
			11571: out = 16'(-5155);
			11572: out = 16'(-1573);
			11573: out = 16'(1450);
			11574: out = 16'(1999);
			11575: out = 16'(516);
			11576: out = 16'(-1892);
			11577: out = 16'(306);
			11578: out = 16'(-488);
			11579: out = 16'(-320);
			11580: out = 16'(-6915);
			11581: out = 16'(-4644);
			11582: out = 16'(774);
			11583: out = 16'(4241);
			11584: out = 16'(3984);
			11585: out = 16'(-2126);
			11586: out = 16'(1821);
			11587: out = 16'(1501);
			11588: out = 16'(307);
			11589: out = 16'(-2595);
			11590: out = 16'(-3058);
			11591: out = 16'(1155);
			11592: out = 16'(1159);
			11593: out = 16'(1406);
			11594: out = 16'(3161);
			11595: out = 16'(3183);
			11596: out = 16'(2903);
			11597: out = 16'(-1080);
			11598: out = 16'(-1642);
			11599: out = 16'(-1458);
			11600: out = 16'(2477);
			11601: out = 16'(2208);
			11602: out = 16'(-361);
			11603: out = 16'(-139);
			11604: out = 16'(623);
			11605: out = 16'(3153);
			11606: out = 16'(2402);
			11607: out = 16'(677);
			11608: out = 16'(-3932);
			11609: out = 16'(-6424);
			11610: out = 16'(-6451);
			11611: out = 16'(3817);
			11612: out = 16'(5977);
			11613: out = 16'(7123);
			11614: out = 16'(-8004);
			11615: out = 16'(-6851);
			11616: out = 16'(-3127);
			11617: out = 16'(7204);
			11618: out = 16'(8104);
			11619: out = 16'(5406);
			11620: out = 16'(-6563);
			11621: out = 16'(-11033);
			11622: out = 16'(-8215);
			11623: out = 16'(-2307);
			11624: out = 16'(2376);
			11625: out = 16'(287);
			11626: out = 16'(3263);
			11627: out = 16'(2180);
			11628: out = 16'(668);
			11629: out = 16'(-4592);
			11630: out = 16'(-7056);
			11631: out = 16'(-347);
			11632: out = 16'(1251);
			11633: out = 16'(2315);
			11634: out = 16'(-14);
			11635: out = 16'(-729);
			11636: out = 16'(-1467);
			11637: out = 16'(-395);
			11638: out = 16'(219);
			11639: out = 16'(1384);
			11640: out = 16'(276);
			11641: out = 16'(-693);
			11642: out = 16'(-4062);
			11643: out = 16'(-337);
			11644: out = 16'(1959);
			11645: out = 16'(6922);
			11646: out = 16'(-702);
			11647: out = 16'(-5211);
			11648: out = 16'(-1338);
			11649: out = 16'(-67);
			11650: out = 16'(1431);
			11651: out = 16'(-230);
			11652: out = 16'(846);
			11653: out = 16'(2256);
			11654: out = 16'(-6599);
			11655: out = 16'(-3504);
			11656: out = 16'(4288);
			11657: out = 16'(5735);
			11658: out = 16'(2928);
			11659: out = 16'(-8671);
			11660: out = 16'(-676);
			11661: out = 16'(1355);
			11662: out = 16'(3931);
			11663: out = 16'(-211);
			11664: out = 16'(-740);
			11665: out = 16'(652);
			11666: out = 16'(6185);
			11667: out = 16'(7931);
			11668: out = 16'(-705);
			11669: out = 16'(-7270);
			11670: out = 16'(-12271);
			11671: out = 16'(4676);
			11672: out = 16'(8058);
			11673: out = 16'(9729);
			11674: out = 16'(55);
			11675: out = 16'(-2402);
			11676: out = 16'(-2770);
			11677: out = 16'(2549);
			11678: out = 16'(3639);
			11679: out = 16'(447);
			11680: out = 16'(1159);
			11681: out = 16'(462);
			11682: out = 16'(784);
			11683: out = 16'(-569);
			11684: out = 16'(96);
			11685: out = 16'(2594);
			11686: out = 16'(3223);
			11687: out = 16'(2088);
			11688: out = 16'(402);
			11689: out = 16'(-4234);
			11690: out = 16'(-7971);
			11691: out = 16'(-4819);
			11692: out = 16'(-1432);
			11693: out = 16'(2236);
			11694: out = 16'(319);
			11695: out = 16'(-818);
			11696: out = 16'(-1443);
			11697: out = 16'(-4532);
			11698: out = 16'(-3913);
			11699: out = 16'(-413);
			11700: out = 16'(3616);
			11701: out = 16'(4568);
			11702: out = 16'(-88);
			11703: out = 16'(-1541);
			11704: out = 16'(-2943);
			11705: out = 16'(-2696);
			11706: out = 16'(-1502);
			11707: out = 16'(153);
			11708: out = 16'(3134);
			11709: out = 16'(1902);
			11710: out = 16'(-387);
			11711: out = 16'(-5263);
			11712: out = 16'(-4742);
			11713: out = 16'(-775);
			11714: out = 16'(2252);
			11715: out = 16'(2960);
			11716: out = 16'(-280);
			11717: out = 16'(241);
			11718: out = 16'(-708);
			11719: out = 16'(-1160);
			11720: out = 16'(-796);
			11721: out = 16'(582);
			11722: out = 16'(3276);
			11723: out = 16'(2151);
			11724: out = 16'(148);
			11725: out = 16'(-3399);
			11726: out = 16'(-1132);
			11727: out = 16'(2903);
			11728: out = 16'(-88);
			11729: out = 16'(-437);
			11730: out = 16'(-3134);
			11731: out = 16'(357);
			11732: out = 16'(-889);
			11733: out = 16'(-692);
			11734: out = 16'(-9368);
			11735: out = 16'(-7231);
			11736: out = 16'(4873);
			11737: out = 16'(9190);
			11738: out = 16'(8219);
			11739: out = 16'(-7444);
			11740: out = 16'(-8614);
			11741: out = 16'(-7608);
			11742: out = 16'(9979);
			11743: out = 16'(8592);
			11744: out = 16'(6504);
			11745: out = 16'(-5203);
			11746: out = 16'(-3554);
			11747: out = 16'(666);
			11748: out = 16'(2970);
			11749: out = 16'(1142);
			11750: out = 16'(-4107);
			11751: out = 16'(-638);
			11752: out = 16'(2670);
			11753: out = 16'(9622);
			11754: out = 16'(3221);
			11755: out = 16'(-258);
			11756: out = 16'(-3921);
			11757: out = 16'(-1732);
			11758: out = 16'(273);
			11759: out = 16'(2051);
			11760: out = 16'(1642);
			11761: out = 16'(741);
			11762: out = 16'(-132);
			11763: out = 16'(-2026);
			11764: out = 16'(-3881);
			11765: out = 16'(369);
			11766: out = 16'(1241);
			11767: out = 16'(2343);
			11768: out = 16'(-2987);
			11769: out = 16'(-2604);
			11770: out = 16'(153);
			11771: out = 16'(3326);
			11772: out = 16'(2810);
			11773: out = 16'(-2930);
			11774: out = 16'(-3286);
			11775: out = 16'(-3360);
			11776: out = 16'(-126);
			11777: out = 16'(-110);
			11778: out = 16'(345);
			11779: out = 16'(788);
			11780: out = 16'(874);
			11781: out = 16'(1123);
			11782: out = 16'(3992);
			11783: out = 16'(3504);
			11784: out = 16'(1663);
			11785: out = 16'(484);
			11786: out = 16'(149);
			11787: out = 16'(2515);
			11788: out = 16'(-2987);
			11789: out = 16'(-4593);
			11790: out = 16'(-8266);
			11791: out = 16'(2826);
			11792: out = 16'(5701);
			11793: out = 16'(2415);
			11794: out = 16'(-4163);
			11795: out = 16'(-6764);
			11796: out = 16'(287);
			11797: out = 16'(6557);
			11798: out = 16'(10121);
			11799: out = 16'(479);
			11800: out = 16'(-6748);
			11801: out = 16'(-14612);
			11802: out = 16'(-1230);
			11803: out = 16'(272);
			11804: out = 16'(113);
			11805: out = 16'(-1897);
			11806: out = 16'(-2047);
			11807: out = 16'(349);
			11808: out = 16'(-4089);
			11809: out = 16'(-2796);
			11810: out = 16'(2451);
			11811: out = 16'(6566);
			11812: out = 16'(7634);
			11813: out = 16'(3347);
			11814: out = 16'(1252);
			11815: out = 16'(-1472);
			11816: out = 16'(-7314);
			11817: out = 16'(-5098);
			11818: out = 16'(-1256);
			11819: out = 16'(7355);
			11820: out = 16'(7051);
			11821: out = 16'(4629);
			11822: out = 16'(-5801);
			11823: out = 16'(-4954);
			11824: out = 16'(2024);
			11825: out = 16'(6970);
			11826: out = 16'(8251);
			11827: out = 16'(3328);
			11828: out = 16'(3064);
			11829: out = 16'(-304);
			11830: out = 16'(-6671);
			11831: out = 16'(-1932);
			11832: out = 16'(1328);
			11833: out = 16'(564);
			11834: out = 16'(-3912);
			11835: out = 16'(-6672);
			11836: out = 16'(9263);
			11837: out = 16'(8624);
			11838: out = 16'(7022);
			11839: out = 16'(-2966);
			11840: out = 16'(-3269);
			11841: out = 16'(-458);
			11842: out = 16'(-2834);
			11843: out = 16'(-3278);
			11844: out = 16'(-4257);
			11845: out = 16'(670);
			11846: out = 16'(826);
			11847: out = 16'(-4387);
			11848: out = 16'(-4602);
			11849: out = 16'(-3980);
			11850: out = 16'(3784);
			11851: out = 16'(704);
			11852: out = 16'(426);
			11853: out = 16'(357);
			11854: out = 16'(3688);
			11855: out = 16'(4637);
			11856: out = 16'(6804);
			11857: out = 16'(-1514);
			11858: out = 16'(-10949);
			11859: out = 16'(-12513);
			11860: out = 16'(-6998);
			11861: out = 16'(4591);
			11862: out = 16'(3522);
			11863: out = 16'(3608);
			11864: out = 16'(-634);
			11865: out = 16'(607);
			11866: out = 16'(-1363);
			11867: out = 16'(-4736);
			11868: out = 16'(-1498);
			11869: out = 16'(1849);
			11870: out = 16'(1787);
			11871: out = 16'(1939);
			11872: out = 16'(173);
			11873: out = 16'(700);
			11874: out = 16'(-1633);
			11875: out = 16'(-2699);
			11876: out = 16'(-9301);
			11877: out = 16'(-6696);
			11878: out = 16'(-1384);
			11879: out = 16'(6352);
			11880: out = 16'(8141);
			11881: out = 16'(5780);
			11882: out = 16'(1644);
			11883: out = 16'(-1017);
			11884: out = 16'(89);
			11885: out = 16'(329);
			11886: out = 16'(1273);
			11887: out = 16'(-740);
			11888: out = 16'(16);
			11889: out = 16'(-650);
			11890: out = 16'(397);
			11891: out = 16'(-53);
			11892: out = 16'(1196);
			11893: out = 16'(-2104);
			11894: out = 16'(1695);
			11895: out = 16'(4212);
			11896: out = 16'(10442);
			11897: out = 16'(4743);
			11898: out = 16'(-4739);
			11899: out = 16'(-7960);
			11900: out = 16'(-5179);
			11901: out = 16'(4770);
			11902: out = 16'(6025);
			11903: out = 16'(4089);
			11904: out = 16'(-8330);
			11905: out = 16'(-5689);
			11906: out = 16'(-3239);
			11907: out = 16'(7459);
			11908: out = 16'(2389);
			11909: out = 16'(-499);
			11910: out = 16'(1774);
			11911: out = 16'(3867);
			11912: out = 16'(5710);
			11913: out = 16'(129);
			11914: out = 16'(-1349);
			11915: out = 16'(-3368);
			11916: out = 16'(-2593);
			11917: out = 16'(-2644);
			11918: out = 16'(43);
			11919: out = 16'(-7424);
			11920: out = 16'(-6891);
			11921: out = 16'(-2764);
			11922: out = 16'(6879);
			11923: out = 16'(10012);
			11924: out = 16'(4896);
			11925: out = 16'(-2399);
			11926: out = 16'(-7762);
			11927: out = 16'(1486);
			11928: out = 16'(145);
			11929: out = 16'(944);
			11930: out = 16'(-2026);
			11931: out = 16'(-597);
			11932: out = 16'(-1027);
			11933: out = 16'(-727);
			11934: out = 16'(-3863);
			11935: out = 16'(-5722);
			11936: out = 16'(-5012);
			11937: out = 16'(970);
			11938: out = 16'(8976);
			11939: out = 16'(9345);
			11940: out = 16'(4621);
			11941: out = 16'(-7609);
			11942: out = 16'(-8503);
			11943: out = 16'(-6409);
			11944: out = 16'(3001);
			11945: out = 16'(4604);
			11946: out = 16'(4288);
			11947: out = 16'(-694);
			11948: out = 16'(-6386);
			11949: out = 16'(-10761);
			11950: out = 16'(15);
			11951: out = 16'(4691);
			11952: out = 16'(9224);
			11953: out = 16'(858);
			11954: out = 16'(-170);
			11955: out = 16'(829);
			11956: out = 16'(-220);
			11957: out = 16'(-131);
			11958: out = 16'(728);
			11959: out = 16'(20);
			11960: out = 16'(-1383);
			11961: out = 16'(-5028);
			11962: out = 16'(-1287);
			11963: out = 16'(1691);
			11964: out = 16'(-537);
			11965: out = 16'(2695);
			11966: out = 16'(4479);
			11967: out = 16'(8974);
			11968: out = 16'(3218);
			11969: out = 16'(-3730);
			11970: out = 16'(-2545);
			11971: out = 16'(-1880);
			11972: out = 16'(96);
			11973: out = 16'(-1104);
			11974: out = 16'(-3942);
			11975: out = 16'(-10089);
			11976: out = 16'(-3514);
			11977: out = 16'(917);
			11978: out = 16'(5353);
			11979: out = 16'(5975);
			11980: out = 16'(5383);
			11981: out = 16'(863);
			11982: out = 16'(2941);
			11983: out = 16'(3321);
			11984: out = 16'(-2376);
			11985: out = 16'(-4404);
			11986: out = 16'(-5695);
			11987: out = 16'(5403);
			11988: out = 16'(3342);
			11989: out = 16'(-905);
			11990: out = 16'(-3311);
			11991: out = 16'(-1602);
			11992: out = 16'(3662);
			11993: out = 16'(1993);
			11994: out = 16'(1607);
			11995: out = 16'(-434);
			11996: out = 16'(2172);
			11997: out = 16'(2884);
			11998: out = 16'(1749);
			11999: out = 16'(760);
			12000: out = 16'(-1137);
			12001: out = 16'(-2201);
			12002: out = 16'(-6285);
			12003: out = 16'(-8037);
			12004: out = 16'(-2318);
			12005: out = 16'(2294);
			12006: out = 16'(6261);
			12007: out = 16'(1401);
			12008: out = 16'(-1475);
			12009: out = 16'(-5261);
			12010: out = 16'(-747);
			12011: out = 16'(316);
			12012: out = 16'(890);
			12013: out = 16'(-1888);
			12014: out = 16'(-355);
			12015: out = 16'(8470);
			12016: out = 16'(2439);
			12017: out = 16'(-2098);
			12018: out = 16'(-11212);
			12019: out = 16'(-5045);
			12020: out = 16'(1470);
			12021: out = 16'(5500);
			12022: out = 16'(6421);
			12023: out = 16'(5415);
			12024: out = 16'(627);
			12025: out = 16'(-1281);
			12026: out = 16'(-2883);
			12027: out = 16'(1648);
			12028: out = 16'(268);
			12029: out = 16'(-2729);
			12030: out = 16'(-7432);
			12031: out = 16'(-6110);
			12032: out = 16'(1558);
			12033: out = 16'(5081);
			12034: out = 16'(7030);
			12035: out = 16'(3704);
			12036: out = 16'(3022);
			12037: out = 16'(1478);
			12038: out = 16'(2140);
			12039: out = 16'(928);
			12040: out = 16'(702);
			12041: out = 16'(3583);
			12042: out = 16'(2882);
			12043: out = 16'(917);
			12044: out = 16'(-7087);
			12045: out = 16'(-9812);
			12046: out = 16'(-9416);
			12047: out = 16'(-1694);
			12048: out = 16'(3856);
			12049: out = 16'(7687);
			12050: out = 16'(2350);
			12051: out = 16'(-1467);
			12052: out = 16'(-2313);
			12053: out = 16'(-2449);
			12054: out = 16'(-535);
			12055: out = 16'(1545);
			12056: out = 16'(2297);
			12057: out = 16'(1274);
			12058: out = 16'(-22);
			12059: out = 16'(-1633);
			12060: out = 16'(-1400);
			12061: out = 16'(-4482);
			12062: out = 16'(1149);
			12063: out = 16'(8097);
			12064: out = 16'(4596);
			12065: out = 16'(753);
			12066: out = 16'(-5752);
			12067: out = 16'(-606);
			12068: out = 16'(875);
			12069: out = 16'(-782);
			12070: out = 16'(2935);
			12071: out = 16'(2955);
			12072: out = 16'(783);
			12073: out = 16'(-6242);
			12074: out = 16'(-9413);
			12075: out = 16'(298);
			12076: out = 16'(3276);
			12077: out = 16'(6053);
			12078: out = 16'(483);
			12079: out = 16'(348);
			12080: out = 16'(-626);
			12081: out = 16'(1924);
			12082: out = 16'(-158);
			12083: out = 16'(-3199);
			12084: out = 16'(-5842);
			12085: out = 16'(-4488);
			12086: out = 16'(1538);
			12087: out = 16'(461);
			12088: out = 16'(-1727);
			12089: out = 16'(-13710);
			12090: out = 16'(-1623);
			12091: out = 16'(4833);
			12092: out = 16'(10202);
			12093: out = 16'(452);
			12094: out = 16'(-7477);
			12095: out = 16'(-8396);
			12096: out = 16'(-2866);
			12097: out = 16'(4233);
			12098: out = 16'(-7);
			12099: out = 16'(-606);
			12100: out = 16'(-2857);
			12101: out = 16'(-3281);
			12102: out = 16'(-1712);
			12103: out = 16'(3027);
			12104: out = 16'(2811);
			12105: out = 16'(2933);
			12106: out = 16'(-404);
			12107: out = 16'(2743);
			12108: out = 16'(2679);
			12109: out = 16'(1297);
			12110: out = 16'(-1269);
			12111: out = 16'(-2361);
			12112: out = 16'(869);
			12113: out = 16'(85);
			12114: out = 16'(-280);
			12115: out = 16'(48);
			12116: out = 16'(-538);
			12117: out = 16'(-1417);
			12118: out = 16'(848);
			12119: out = 16'(3581);
			12120: out = 16'(8265);
			12121: out = 16'(-4954);
			12122: out = 16'(-8683);
			12123: out = 16'(-11354);
			12124: out = 16'(4281);
			12125: out = 16'(8980);
			12126: out = 16'(4893);
			12127: out = 16'(-2736);
			12128: out = 16'(-7764);
			12129: out = 16'(-1768);
			12130: out = 16'(-1210);
			12131: out = 16'(2127);
			12132: out = 16'(1419);
			12133: out = 16'(4996);
			12134: out = 16'(5414);
			12135: out = 16'(943);
			12136: out = 16'(-762);
			12137: out = 16'(112);
			12138: out = 16'(-2077);
			12139: out = 16'(767);
			12140: out = 16'(2826);
			12141: out = 16'(6990);
			12142: out = 16'(2241);
			12143: out = 16'(-9036);
			12144: out = 16'(-9066);
			12145: out = 16'(-4463);
			12146: out = 16'(9091);
			12147: out = 16'(10434);
			12148: out = 16'(9550);
			12149: out = 16'(-621);
			12150: out = 16'(-2416);
			12151: out = 16'(-3877);
			12152: out = 16'(2920);
			12153: out = 16'(1607);
			12154: out = 16'(153);
			12155: out = 16'(-8964);
			12156: out = 16'(-8354);
			12157: out = 16'(-4149);
			12158: out = 16'(-307);
			12159: out = 16'(2152);
			12160: out = 16'(1802);
			12161: out = 16'(3444);
			12162: out = 16'(1653);
			12163: out = 16'(-1247);
			12164: out = 16'(-5746);
			12165: out = 16'(-5414);
			12166: out = 16'(4532);
			12167: out = 16'(2944);
			12168: out = 16'(570);
			12169: out = 16'(-10667);
			12170: out = 16'(-7332);
			12171: out = 16'(-1942);
			12172: out = 16'(3476);
			12173: out = 16'(4535);
			12174: out = 16'(2920);
			12175: out = 16'(2838);
			12176: out = 16'(2500);
			12177: out = 16'(4676);
			12178: out = 16'(-3470);
			12179: out = 16'(-3541);
			12180: out = 16'(-244);
			12181: out = 16'(5367);
			12182: out = 16'(5112);
			12183: out = 16'(-4115);
			12184: out = 16'(-3551);
			12185: out = 16'(-2752);
			12186: out = 16'(3448);
			12187: out = 16'(1118);
			12188: out = 16'(276);
			12189: out = 16'(5757);
			12190: out = 16'(6878);
			12191: out = 16'(7017);
			12192: out = 16'(-3776);
			12193: out = 16'(-6259);
			12194: out = 16'(-7462);
			12195: out = 16'(2421);
			12196: out = 16'(3152);
			12197: out = 16'(504);
			12198: out = 16'(-5551);
			12199: out = 16'(-6238);
			12200: out = 16'(-1162);
			12201: out = 16'(4349);
			12202: out = 16'(6478);
			12203: out = 16'(-529);
			12204: out = 16'(-430);
			12205: out = 16'(-2092);
			12206: out = 16'(-929);
			12207: out = 16'(-4762);
			12208: out = 16'(-6675);
			12209: out = 16'(2553);
			12210: out = 16'(3382);
			12211: out = 16'(2902);
			12212: out = 16'(-4720);
			12213: out = 16'(-5422);
			12214: out = 16'(-3069);
			12215: out = 16'(1711);
			12216: out = 16'(4665);
			12217: out = 16'(6178);
			12218: out = 16'(2786);
			12219: out = 16'(-1136);
			12220: out = 16'(-8733);
			12221: out = 16'(-938);
			12222: out = 16'(4573);
			12223: out = 16'(5915);
			12224: out = 16'(2871);
			12225: out = 16'(-1646);
			12226: out = 16'(-4181);
			12227: out = 16'(-4782);
			12228: out = 16'(-2946);
			12229: out = 16'(-966);
			12230: out = 16'(825);
			12231: out = 16'(1085);
			12232: out = 16'(524);
			12233: out = 16'(203);
			12234: out = 16'(1172);
			12235: out = 16'(108);
			12236: out = 16'(523);
			12237: out = 16'(698);
			12238: out = 16'(1134);
			12239: out = 16'(-377);
			12240: out = 16'(-4676);
			12241: out = 16'(-2988);
			12242: out = 16'(-370);
			12243: out = 16'(791);
			12244: out = 16'(1014);
			12245: out = 16'(-167);
			12246: out = 16'(7346);
			12247: out = 16'(4805);
			12248: out = 16'(2891);
			12249: out = 16'(-11004);
			12250: out = 16'(-6885);
			12251: out = 16'(4324);
			12252: out = 16'(9245);
			12253: out = 16'(6305);
			12254: out = 16'(-7271);
			12255: out = 16'(-4131);
			12256: out = 16'(-1346);
			12257: out = 16'(8558);
			12258: out = 16'(4384);
			12259: out = 16'(3058);
			12260: out = 16'(3940);
			12261: out = 16'(3342);
			12262: out = 16'(2029);
			12263: out = 16'(-3758);
			12264: out = 16'(-3544);
			12265: out = 16'(-2403);
			12266: out = 16'(4369);
			12267: out = 16'(2737);
			12268: out = 16'(-911);
			12269: out = 16'(-9417);
			12270: out = 16'(-9521);
			12271: out = 16'(-2891);
			12272: out = 16'(220);
			12273: out = 16'(3461);
			12274: out = 16'(3762);
			12275: out = 16'(4525);
			12276: out = 16'(2148);
			12277: out = 16'(-5055);
			12278: out = 16'(-4233);
			12279: out = 16'(-3332);
			12280: out = 16'(189);
			12281: out = 16'(-1520);
			12282: out = 16'(-2609);
			12283: out = 16'(-6185);
			12284: out = 16'(-2877);
			12285: out = 16'(878);
			12286: out = 16'(8967);
			12287: out = 16'(7692);
			12288: out = 16'(3777);
			12289: out = 16'(-5192);
			12290: out = 16'(-6039);
			12291: out = 16'(-1116);
			12292: out = 16'(5505);
			12293: out = 16'(6769);
			12294: out = 16'(816);
			12295: out = 16'(-3485);
			12296: out = 16'(-6323);
			12297: out = 16'(-3759);
			12298: out = 16'(759);
			12299: out = 16'(5046);
			12300: out = 16'(5996);
			12301: out = 16'(2532);
			12302: out = 16'(-2486);
			12303: out = 16'(-5716);
			12304: out = 16'(-2290);
			12305: out = 16'(5067);
			12306: out = 16'(2128);
			12307: out = 16'(-592);
			12308: out = 16'(-8311);
			12309: out = 16'(-2348);
			12310: out = 16'(-574);
			12311: out = 16'(2768);
			12312: out = 16'(-1389);
			12313: out = 16'(-1720);
			12314: out = 16'(1062);
			12315: out = 16'(3232);
			12316: out = 16'(2745);
			12317: out = 16'(-8220);
			12318: out = 16'(-4822);
			12319: out = 16'(-272);
			12320: out = 16'(695);
			12321: out = 16'(1661);
			12322: out = 16'(541);
			12323: out = 16'(2860);
			12324: out = 16'(-1461);
			12325: out = 16'(-7333);
			12326: out = 16'(-2783);
			12327: out = 16'(2627);
			12328: out = 16'(10297);
			12329: out = 16'(7173);
			12330: out = 16'(4442);
			12331: out = 16'(-592);
			12332: out = 16'(320);
			12333: out = 16'(810);
			12334: out = 16'(2170);
			12335: out = 16'(-1964);
			12336: out = 16'(-4795);
			12337: out = 16'(4305);
			12338: out = 16'(1411);
			12339: out = 16'(-950);
			12340: out = 16'(-9481);
			12341: out = 16'(-4918);
			12342: out = 16'(3106);
			12343: out = 16'(3664);
			12344: out = 16'(3335);
			12345: out = 16'(722);
			12346: out = 16'(-1634);
			12347: out = 16'(-2831);
			12348: out = 16'(-2588);
			12349: out = 16'(2169);
			12350: out = 16'(3771);
			12351: out = 16'(-237);
			12352: out = 16'(-1389);
			12353: out = 16'(-3203);
			12354: out = 16'(-4847);
			12355: out = 16'(-677);
			12356: out = 16'(3960);
			12357: out = 16'(844);
			12358: out = 16'(461);
			12359: out = 16'(-1909);
			12360: out = 16'(1389);
			12361: out = 16'(540);
			12362: out = 16'(1231);
			12363: out = 16'(-3547);
			12364: out = 16'(-915);
			12365: out = 16'(4215);
			12366: out = 16'(6816);
			12367: out = 16'(2844);
			12368: out = 16'(-11641);
			12369: out = 16'(-7259);
			12370: out = 16'(-2008);
			12371: out = 16'(7723);
			12372: out = 16'(7200);
			12373: out = 16'(4955);
			12374: out = 16'(1843);
			12375: out = 16'(-4056);
			12376: out = 16'(-8868);
			12377: out = 16'(-5409);
			12378: out = 16'(-645);
			12379: out = 16'(5839);
			12380: out = 16'(-2443);
			12381: out = 16'(-5882);
			12382: out = 16'(-11328);
			12383: out = 16'(2770);
			12384: out = 16'(8048);
			12385: out = 16'(9879);
			12386: out = 16'(2965);
			12387: out = 16'(-2182);
			12388: out = 16'(-5967);
			12389: out = 16'(-1753);
			12390: out = 16'(1593);
			12391: out = 16'(-1588);
			12392: out = 16'(-2781);
			12393: out = 16'(-4343);
			12394: out = 16'(6325);
			12395: out = 16'(3141);
			12396: out = 16'(-7);
			12397: out = 16'(-1438);
			12398: out = 16'(659);
			12399: out = 16'(3393);
			12400: out = 16'(4161);
			12401: out = 16'(3585);
			12402: out = 16'(3262);
			12403: out = 16'(-3929);
			12404: out = 16'(-6273);
			12405: out = 16'(-4932);
			12406: out = 16'(492);
			12407: out = 16'(4101);
			12408: out = 16'(5177);
			12409: out = 16'(1342);
			12410: out = 16'(-1806);
			12411: out = 16'(-72);
			12412: out = 16'(2427);
			12413: out = 16'(5054);
			12414: out = 16'(251);
			12415: out = 16'(-1764);
			12416: out = 16'(-3963);
			12417: out = 16'(-194);
			12418: out = 16'(2411);
			12419: out = 16'(5042);
			12420: out = 16'(3640);
			12421: out = 16'(-40);
			12422: out = 16'(-7939);
			12423: out = 16'(-3306);
			12424: out = 16'(-690);
			12425: out = 16'(-345);
			12426: out = 16'(2244);
			12427: out = 16'(2882);
			12428: out = 16'(2402);
			12429: out = 16'(-1860);
			12430: out = 16'(-5201);
			12431: out = 16'(-2659);
			12432: out = 16'(-2014);
			12433: out = 16'(-1378);
			12434: out = 16'(-2277);
			12435: out = 16'(-1828);
			12436: out = 16'(250);
			12437: out = 16'(-4339);
			12438: out = 16'(-2957);
			12439: out = 16'(-116);
			12440: out = 16'(5777);
			12441: out = 16'(6517);
			12442: out = 16'(4520);
			12443: out = 16'(-3458);
			12444: out = 16'(-7009);
			12445: out = 16'(-2519);
			12446: out = 16'(2239);
			12447: out = 16'(4378);
			12448: out = 16'(-6453);
			12449: out = 16'(-9671);
			12450: out = 16'(-11161);
			12451: out = 16'(16);
			12452: out = 16'(5315);
			12453: out = 16'(9451);
			12454: out = 16'(5238);
			12455: out = 16'(3797);
			12456: out = 16'(3434);
			12457: out = 16'(-3035);
			12458: out = 16'(-3785);
			12459: out = 16'(111);
			12460: out = 16'(3644);
			12461: out = 16'(4870);
			12462: out = 16'(600);
			12463: out = 16'(373);
			12464: out = 16'(-894);
			12465: out = 16'(-3601);
			12466: out = 16'(-11);
			12467: out = 16'(4283);
			12468: out = 16'(6575);
			12469: out = 16'(4130);
			12470: out = 16'(-1386);
			12471: out = 16'(3548);
			12472: out = 16'(-71);
			12473: out = 16'(-3869);
			12474: out = 16'(-6181);
			12475: out = 16'(-2724);
			12476: out = 16'(5696);
			12477: out = 16'(1766);
			12478: out = 16'(-643);
			12479: out = 16'(-5186);
			12480: out = 16'(938);
			12481: out = 16'(5074);
			12482: out = 16'(4490);
			12483: out = 16'(5365);
			12484: out = 16'(4459);
			12485: out = 16'(6247);
			12486: out = 16'(2263);
			12487: out = 16'(-1139);
			12488: out = 16'(-7178);
			12489: out = 16'(-6315);
			12490: out = 16'(-3506);
			12491: out = 16'(3577);
			12492: out = 16'(3439);
			12493: out = 16'(-679);
			12494: out = 16'(-462);
			12495: out = 16'(-300);
			12496: out = 16'(298);
			12497: out = 16'(4298);
			12498: out = 16'(5357);
			12499: out = 16'(3919);
			12500: out = 16'(-2555);
			12501: out = 16'(-6843);
			12502: out = 16'(-3003);
			12503: out = 16'(418);
			12504: out = 16'(3639);
			12505: out = 16'(-4907);
			12506: out = 16'(-5803);
			12507: out = 16'(-6264);
			12508: out = 16'(-84);
			12509: out = 16'(1119);
			12510: out = 16'(767);
			12511: out = 16'(1834);
			12512: out = 16'(1729);
			12513: out = 16'(1960);
			12514: out = 16'(-3288);
			12515: out = 16'(-5577);
			12516: out = 16'(-5048);
			12517: out = 16'(-2171);
			12518: out = 16'(-652);
			12519: out = 16'(-5266);
			12520: out = 16'(-2130);
			12521: out = 16'(167);
			12522: out = 16'(686);
			12523: out = 16'(-35);
			12524: out = 16'(-1327);
			12525: out = 16'(4172);
			12526: out = 16'(2323);
			12527: out = 16'(-223);
			12528: out = 16'(-4249);
			12529: out = 16'(-3255);
			12530: out = 16'(416);
			12531: out = 16'(2673);
			12532: out = 16'(1105);
			12533: out = 16'(-6574);
			12534: out = 16'(-3366);
			12535: out = 16'(-1128);
			12536: out = 16'(3651);
			12537: out = 16'(1282);
			12538: out = 16'(172);
			12539: out = 16'(1285);
			12540: out = 16'(1708);
			12541: out = 16'(2162);
			12542: out = 16'(-1403);
			12543: out = 16'(437);
			12544: out = 16'(2154);
			12545: out = 16'(592);
			12546: out = 16'(-3204);
			12547: out = 16'(-8691);
			12548: out = 16'(-788);
			12549: out = 16'(2163);
			12550: out = 16'(3385);
			12551: out = 16'(5553);
			12552: out = 16'(6093);
			12553: out = 16'(4959);
			12554: out = 16'(3211);
			12555: out = 16'(1057);
			12556: out = 16'(-223);
			12557: out = 16'(-2794);
			12558: out = 16'(-3325);
			12559: out = 16'(1754);
			12560: out = 16'(2939);
			12561: out = 16'(3658);
			12562: out = 16'(-3581);
			12563: out = 16'(-1897);
			12564: out = 16'(1244);
			12565: out = 16'(1672);
			12566: out = 16'(1528);
			12567: out = 16'(464);
			12568: out = 16'(3976);
			12569: out = 16'(3996);
			12570: out = 16'(-276);
			12571: out = 16'(3990);
			12572: out = 16'(4466);
			12573: out = 16'(6235);
			12574: out = 16'(-4834);
			12575: out = 16'(-10832);
			12576: out = 16'(-6497);
			12577: out = 16'(-2737);
			12578: out = 16'(1635);
			12579: out = 16'(293);
			12580: out = 16'(2096);
			12581: out = 16'(2366);
			12582: out = 16'(-4296);
			12583: out = 16'(-4586);
			12584: out = 16'(-2401);
			12585: out = 16'(-857);
			12586: out = 16'(1007);
			12587: out = 16'(3143);
			12588: out = 16'(-1340);
			12589: out = 16'(-4288);
			12590: out = 16'(-9045);
			12591: out = 16'(289);
			12592: out = 16'(5003);
			12593: out = 16'(5118);
			12594: out = 16'(-157);
			12595: out = 16'(-4090);
			12596: out = 16'(79);
			12597: out = 16'(1389);
			12598: out = 16'(3016);
			12599: out = 16'(-2418);
			12600: out = 16'(-2682);
			12601: out = 16'(-2653);
			12602: out = 16'(-2671);
			12603: out = 16'(-2054);
			12604: out = 16'(-1275);
			12605: out = 16'(2628);
			12606: out = 16'(1492);
			12607: out = 16'(-3998);
			12608: out = 16'(-2649);
			12609: out = 16'(-1103);
			12610: out = 16'(3624);
			12611: out = 16'(2550);
			12612: out = 16'(1713);
			12613: out = 16'(-1278);
			12614: out = 16'(-2581);
			12615: out = 16'(-2648);
			12616: out = 16'(6974);
			12617: out = 16'(6033);
			12618: out = 16'(4213);
			12619: out = 16'(-8442);
			12620: out = 16'(-6809);
			12621: out = 16'(-188);
			12622: out = 16'(4507);
			12623: out = 16'(5963);
			12624: out = 16'(2344);
			12625: out = 16'(4540);
			12626: out = 16'(2319);
			12627: out = 16'(-240);
			12628: out = 16'(-2460);
			12629: out = 16'(-2290);
			12630: out = 16'(-2000);
			12631: out = 16'(2159);
			12632: out = 16'(4085);
			12633: out = 16'(4213);
			12634: out = 16'(264);
			12635: out = 16'(-3100);
			12636: out = 16'(-680);
			12637: out = 16'(-96);
			12638: out = 16'(832);
			12639: out = 16'(4292);
			12640: out = 16'(5800);
			12641: out = 16'(7382);
			12642: out = 16'(-4841);
			12643: out = 16'(-8298);
			12644: out = 16'(-7474);
			12645: out = 16'(1361);
			12646: out = 16'(5475);
			12647: out = 16'(3423);
			12648: out = 16'(584);
			12649: out = 16'(-2697);
			12650: out = 16'(-2545);
			12651: out = 16'(-1384);
			12652: out = 16'(1202);
			12653: out = 16'(1390);
			12654: out = 16'(1540);
			12655: out = 16'(-72);
			12656: out = 16'(789);
			12657: out = 16'(-261);
			12658: out = 16'(-171);
			12659: out = 16'(-3758);
			12660: out = 16'(-2453);
			12661: out = 16'(699);
			12662: out = 16'(3838);
			12663: out = 16'(4251);
			12664: out = 16'(1405);
			12665: out = 16'(528);
			12666: out = 16'(-1336);
			12667: out = 16'(-2670);
			12668: out = 16'(-3885);
			12669: out = 16'(-3417);
			12670: out = 16'(-843);
			12671: out = 16'(-421);
			12672: out = 16'(-464);
			12673: out = 16'(1976);
			12674: out = 16'(697);
			12675: out = 16'(-898);
			12676: out = 16'(-5643);
			12677: out = 16'(-3974);
			12678: out = 16'(1357);
			12679: out = 16'(205);
			12680: out = 16'(930);
			12681: out = 16'(-580);
			12682: out = 16'(3518);
			12683: out = 16'(888);
			12684: out = 16'(-10090);
			12685: out = 16'(-7455);
			12686: out = 16'(-4166);
			12687: out = 16'(3302);
			12688: out = 16'(1310);
			12689: out = 16'(296);
			12690: out = 16'(6008);
			12691: out = 16'(5563);
			12692: out = 16'(4106);
			12693: out = 16'(-6168);
			12694: out = 16'(-6420);
			12695: out = 16'(-2969);
			12696: out = 16'(-480);
			12697: out = 16'(2558);
			12698: out = 16'(4015);
			12699: out = 16'(5911);
			12700: out = 16'(4212);
			12701: out = 16'(-766);
			12702: out = 16'(-202);
			12703: out = 16'(288);
			12704: out = 16'(3138);
			12705: out = 16'(783);
			12706: out = 16'(-277);
			12707: out = 16'(449);
			12708: out = 16'(696);
			12709: out = 16'(691);
			12710: out = 16'(628);
			12711: out = 16'(-719);
			12712: out = 16'(-1760);
			12713: out = 16'(-2020);
			12714: out = 16'(1525);
			12715: out = 16'(7202);
			12716: out = 16'(407);
			12717: out = 16'(-1483);
			12718: out = 16'(-3183);
			12719: out = 16'(797);
			12720: out = 16'(830);
			12721: out = 16'(-3091);
			12722: out = 16'(-2881);
			12723: out = 16'(-1902);
			12724: out = 16'(3021);
			12725: out = 16'(1587);
			12726: out = 16'(255);
			12727: out = 16'(-2635);
			12728: out = 16'(-3473);
			12729: out = 16'(-3092);
			12730: out = 16'(6644);
			12731: out = 16'(7684);
			12732: out = 16'(7073);
			12733: out = 16'(1422);
			12734: out = 16'(-1507);
			12735: out = 16'(-4547);
			12736: out = 16'(-245);
			12737: out = 16'(1468);
			12738: out = 16'(5224);
			12739: out = 16'(-4551);
			12740: out = 16'(-7695);
			12741: out = 16'(-5497);
			12742: out = 16'(662);
			12743: out = 16'(3731);
			12744: out = 16'(762);
			12745: out = 16'(-5302);
			12746: out = 16'(-9765);
			12747: out = 16'(-1200);
			12748: out = 16'(4684);
			12749: out = 16'(10610);
			12750: out = 16'(368);
			12751: out = 16'(-2771);
			12752: out = 16'(-7012);
			12753: out = 16'(-4906);
			12754: out = 16'(-4639);
			12755: out = 16'(-1971);
			12756: out = 16'(-1195);
			12757: out = 16'(896);
			12758: out = 16'(-786);
			12759: out = 16'(5571);
			12760: out = 16'(5408);
			12761: out = 16'(147);
			12762: out = 16'(-4981);
			12763: out = 16'(-6701);
			12764: out = 16'(-2152);
			12765: out = 16'(3367);
			12766: out = 16'(7194);
			12767: out = 16'(6514);
			12768: out = 16'(93);
			12769: out = 16'(-8175);
			12770: out = 16'(-3434);
			12771: out = 16'(1428);
			12772: out = 16'(9454);
			12773: out = 16'(5312);
			12774: out = 16'(3468);
			12775: out = 16'(-1239);
			12776: out = 16'(1428);
			12777: out = 16'(1101);
			12778: out = 16'(-382);
			12779: out = 16'(-490);
			12780: out = 16'(-606);
			12781: out = 16'(-1782);
			12782: out = 16'(-3007);
			12783: out = 16'(-4056);
			12784: out = 16'(-1606);
			12785: out = 16'(-2313);
			12786: out = 16'(-2427);
			12787: out = 16'(29);
			12788: out = 16'(2219);
			12789: out = 16'(3946);
			12790: out = 16'(1598);
			12791: out = 16'(-1510);
			12792: out = 16'(-6669);
			12793: out = 16'(-3498);
			12794: out = 16'(-958);
			12795: out = 16'(4591);
			12796: out = 16'(-699);
			12797: out = 16'(-3796);
			12798: out = 16'(-8791);
			12799: out = 16'(-1965);
			12800: out = 16'(3744);
			12801: out = 16'(7685);
			12802: out = 16'(4313);
			12803: out = 16'(-127);
			12804: out = 16'(-125);
			12805: out = 16'(1213);
			12806: out = 16'(4354);
			12807: out = 16'(-221);
			12808: out = 16'(-1212);
			12809: out = 16'(-3084);
			12810: out = 16'(142);
			12811: out = 16'(616);
			12812: out = 16'(1109);
			12813: out = 16'(-111);
			12814: out = 16'(-39);
			12815: out = 16'(-827);
			12816: out = 16'(2653);
			12817: out = 16'(3335);
			12818: out = 16'(-140);
			12819: out = 16'(-1729);
			12820: out = 16'(-3061);
			12821: out = 16'(-3931);
			12822: out = 16'(-1698);
			12823: out = 16'(803);
			12824: out = 16'(-1272);
			12825: out = 16'(-3780);
			12826: out = 16'(-7476);
			12827: out = 16'(734);
			12828: out = 16'(4280);
			12829: out = 16'(8141);
			12830: out = 16'(-260);
			12831: out = 16'(-3679);
			12832: out = 16'(-4899);
			12833: out = 16'(-1066);
			12834: out = 16'(1062);
			12835: out = 16'(-586);
			12836: out = 16'(548);
			12837: out = 16'(969);
			12838: out = 16'(2148);
			12839: out = 16'(3057);
			12840: out = 16'(4103);
			12841: out = 16'(860);
			12842: out = 16'(1569);
			12843: out = 16'(1860);
			12844: out = 16'(3862);
			12845: out = 16'(3251);
			12846: out = 16'(2881);
			12847: out = 16'(587);
			12848: out = 16'(162);
			12849: out = 16'(-1175);
			12850: out = 16'(1449);
			12851: out = 16'(1840);
			12852: out = 16'(5495);
			12853: out = 16'(-5580);
			12854: out = 16'(-10634);
			12855: out = 16'(-10534);
			12856: out = 16'(-624);
			12857: out = 16'(6966);
			12858: out = 16'(5838);
			12859: out = 16'(68);
			12860: out = 16'(-7237);
			12861: out = 16'(-2871);
			12862: out = 16'(-181);
			12863: out = 16'(4491);
			12864: out = 16'(288);
			12865: out = 16'(-2515);
			12866: out = 16'(-8011);
			12867: out = 16'(-2715);
			12868: out = 16'(75);
			12869: out = 16'(3395);
			12870: out = 16'(3124);
			12871: out = 16'(2552);
			12872: out = 16'(-190);
			12873: out = 16'(531);
			12874: out = 16'(480);
			12875: out = 16'(-355);
			12876: out = 16'(-1596);
			12877: out = 16'(-2239);
			12878: out = 16'(3847);
			12879: out = 16'(3817);
			12880: out = 16'(3595);
			12881: out = 16'(-7212);
			12882: out = 16'(-6910);
			12883: out = 16'(-3022);
			12884: out = 16'(6209);
			12885: out = 16'(9460);
			12886: out = 16'(9070);
			12887: out = 16'(3372);
			12888: out = 16'(-2731);
			12889: out = 16'(-13098);
			12890: out = 16'(-2995);
			12891: out = 16'(2771);
			12892: out = 16'(1905);
			12893: out = 16'(-3139);
			12894: out = 16'(-7808);
			12895: out = 16'(-3611);
			12896: out = 16'(-1020);
			12897: out = 16'(3004);
			12898: out = 16'(2743);
			12899: out = 16'(2170);
			12900: out = 16'(-896);
			12901: out = 16'(1315);
			12902: out = 16'(260);
			12903: out = 16'(-226);
			12904: out = 16'(-3049);
			12905: out = 16'(-3215);
			12906: out = 16'(-1188);
			12907: out = 16'(-3778);
			12908: out = 16'(-3919);
			12909: out = 16'(366);
			12910: out = 16'(2980);
			12911: out = 16'(5582);
			12912: out = 16'(392);
			12913: out = 16'(5322);
			12914: out = 16'(6947);
			12915: out = 16'(1896);
			12916: out = 16'(-4974);
			12917: out = 16'(-11196);
			12918: out = 16'(-3930);
			12919: out = 16'(-220);
			12920: out = 16'(2233);
			12921: out = 16'(4229);
			12922: out = 16'(1741);
			12923: out = 16'(-3695);
			12924: out = 16'(-7282);
			12925: out = 16'(-4763);
			12926: out = 16'(8503);
			12927: out = 16'(8363);
			12928: out = 16'(6375);
			12929: out = 16'(-8471);
			12930: out = 16'(-7504);
			12931: out = 16'(-6049);
			12932: out = 16'(6154);
			12933: out = 16'(1921);
			12934: out = 16'(-2932);
			12935: out = 16'(-5744);
			12936: out = 16'(-1074);
			12937: out = 16'(7206);
			12938: out = 16'(2515);
			12939: out = 16'(1454);
			12940: out = 16'(-1794);
			12941: out = 16'(3313);
			12942: out = 16'(3111);
			12943: out = 16'(-389);
			12944: out = 16'(343);
			12945: out = 16'(1164);
			12946: out = 16'(1972);
			12947: out = 16'(1459);
			12948: out = 16'(130);
			12949: out = 16'(27);
			12950: out = 16'(-2443);
			12951: out = 16'(-3234);
			12952: out = 16'(183);
			12953: out = 16'(4198);
			12954: out = 16'(7891);
			12955: out = 16'(6082);
			12956: out = 16'(3759);
			12957: out = 16'(-134);
			12958: out = 16'(354);
			12959: out = 16'(973);
			12960: out = 16'(3888);
			12961: out = 16'(-1959);
			12962: out = 16'(-6035);
			12963: out = 16'(-10111);
			12964: out = 16'(-6635);
			12965: out = 16'(-2127);
			12966: out = 16'(1254);
			12967: out = 16'(5153);
			12968: out = 16'(6225);
			12969: out = 16'(1272);
			12970: out = 16'(-606);
			12971: out = 16'(-1981);
			12972: out = 16'(-2777);
			12973: out = 16'(-3235);
			12974: out = 16'(-3944);
			12975: out = 16'(1184);
			12976: out = 16'(1300);
			12977: out = 16'(-234);
			12978: out = 16'(-4792);
			12979: out = 16'(-5369);
			12980: out = 16'(-1120);
			12981: out = 16'(761);
			12982: out = 16'(2753);
			12983: out = 16'(2910);
			12984: out = 16'(1884);
			12985: out = 16'(267);
			12986: out = 16'(1255);
			12987: out = 16'(153);
			12988: out = 16'(-488);
			12989: out = 16'(-4738);
			12990: out = 16'(-4025);
			12991: out = 16'(-2261);
			12992: out = 16'(-795);
			12993: out = 16'(268);
			12994: out = 16'(887);
			12995: out = 16'(2677);
			12996: out = 16'(3586);
			12997: out = 16'(4007);
			12998: out = 16'(4807);
			12999: out = 16'(3747);
			13000: out = 16'(-918);
			13001: out = 16'(308);
			13002: out = 16'(91);
			13003: out = 16'(72);
			13004: out = 16'(-3855);
			13005: out = 16'(-6802);
			13006: out = 16'(-7454);
			13007: out = 16'(-3992);
			13008: out = 16'(1315);
			13009: out = 16'(3041);
			13010: out = 16'(6312);
			13011: out = 16'(7411);
			13012: out = 16'(6688);
			13013: out = 16'(2510);
			13014: out = 16'(-3281);
			13015: out = 16'(-2938);
			13016: out = 16'(-2225);
			13017: out = 16'(-159);
			13018: out = 16'(-445);
			13019: out = 16'(-1679);
			13020: out = 16'(-6480);
			13021: out = 16'(-2543);
			13022: out = 16'(1081);
			13023: out = 16'(3592);
			13024: out = 16'(4277);
			13025: out = 16'(3716);
			13026: out = 16'(5148);
			13027: out = 16'(2209);
			13028: out = 16'(-1002);
			13029: out = 16'(-5694);
			13030: out = 16'(-4600);
			13031: out = 16'(-130);
			13032: out = 16'(-4444);
			13033: out = 16'(-6018);
			13034: out = 16'(-8713);
			13035: out = 16'(-635);
			13036: out = 16'(4226);
			13037: out = 16'(7900);
			13038: out = 16'(2626);
			13039: out = 16'(-1275);
			13040: out = 16'(94);
			13041: out = 16'(-101);
			13042: out = 16'(1242);
			13043: out = 16'(-3274);
			13044: out = 16'(330);
			13045: out = 16'(1878);
			13046: out = 16'(4598);
			13047: out = 16'(117);
			13048: out = 16'(-4081);
			13049: out = 16'(-10682);
			13050: out = 16'(-5964);
			13051: out = 16'(4078);
			13052: out = 16'(8359);
			13053: out = 16'(7439);
			13054: out = 16'(183);
			13055: out = 16'(-3980);
			13056: out = 16'(-5448);
			13057: out = 16'(327);
			13058: out = 16'(1803);
			13059: out = 16'(2924);
			13060: out = 16'(-274);
			13061: out = 16'(-4027);
			13062: out = 16'(-7353);
			13063: out = 16'(-1485);
			13064: out = 16'(649);
			13065: out = 16'(4037);
			13066: out = 16'(2608);
			13067: out = 16'(5393);
			13068: out = 16'(7547);
			13069: out = 16'(2393);
			13070: out = 16'(-1336);
			13071: out = 16'(-5232);
			13072: out = 16'(-440);
			13073: out = 16'(-305);
			13074: out = 16'(-6691);
			13075: out = 16'(-4162);
			13076: out = 16'(-3176);
			13077: out = 16'(658);
			13078: out = 16'(-4417);
			13079: out = 16'(-6353);
			13080: out = 16'(-217);
			13081: out = 16'(5244);
			13082: out = 16'(10052);
			13083: out = 16'(1086);
			13084: out = 16'(1121);
			13085: out = 16'(486);
			13086: out = 16'(5138);
			13087: out = 16'(1724);
			13088: out = 16'(-4169);
			13089: out = 16'(-7364);
			13090: out = 16'(-7632);
			13091: out = 16'(-4370);
			13092: out = 16'(746);
			13093: out = 16'(4817);
			13094: out = 16'(5911);
			13095: out = 16'(4028);
			13096: out = 16'(1872);
			13097: out = 16'(5681);
			13098: out = 16'(1766);
			13099: out = 16'(-641);
			13100: out = 16'(-4964);
			13101: out = 16'(-2243);
			13102: out = 16'(730);
			13103: out = 16'(-3111);
			13104: out = 16'(-4772);
			13105: out = 16'(-5660);
			13106: out = 16'(-743);
			13107: out = 16'(3548);
			13108: out = 16'(7124);
			13109: out = 16'(7282);
			13110: out = 16'(5678);
			13111: out = 16'(3087);
			13112: out = 16'(-1657);
			13113: out = 16'(-4732);
			13114: out = 16'(-6221);
			13115: out = 16'(-2280);
			13116: out = 16'(1665);
			13117: out = 16'(2792);
			13118: out = 16'(1614);
			13119: out = 16'(-995);
			13120: out = 16'(-1212);
			13121: out = 16'(90);
			13122: out = 16'(3738);
			13123: out = 16'(-714);
			13124: out = 16'(2779);
			13125: out = 16'(7752);
			13126: out = 16'(6445);
			13127: out = 16'(1329);
			13128: out = 16'(-10973);
			13129: out = 16'(-3079);
			13130: out = 16'(-113);
			13131: out = 16'(643);
			13132: out = 16'(-3804);
			13133: out = 16'(-5669);
			13134: out = 16'(1197);
			13135: out = 16'(548);
			13136: out = 16'(1068);
			13137: out = 16'(1679);
			13138: out = 16'(2261);
			13139: out = 16'(1385);
			13140: out = 16'(511);
			13141: out = 16'(-2540);
			13142: out = 16'(-5080);
			13143: out = 16'(-6501);
			13144: out = 16'(-2428);
			13145: out = 16'(5673);
			13146: out = 16'(1841);
			13147: out = 16'(-1928);
			13148: out = 16'(-10094);
			13149: out = 16'(-4897);
			13150: out = 16'(80);
			13151: out = 16'(7989);
			13152: out = 16'(6320);
			13153: out = 16'(4389);
			13154: out = 16'(1145);
			13155: out = 16'(1486);
			13156: out = 16'(1558);
			13157: out = 16'(-2180);
			13158: out = 16'(-3897);
			13159: out = 16'(-4859);
			13160: out = 16'(-2081);
			13161: out = 16'(-326);
			13162: out = 16'(1254);
			13163: out = 16'(1019);
			13164: out = 16'(1418);
			13165: out = 16'(2126);
			13166: out = 16'(2019);
			13167: out = 16'(1867);
			13168: out = 16'(772);
			13169: out = 16'(2985);
			13170: out = 16'(3389);
			13171: out = 16'(-259);
			13172: out = 16'(-1538);
			13173: out = 16'(-3016);
			13174: out = 16'(-272);
			13175: out = 16'(-2411);
			13176: out = 16'(-3440);
			13177: out = 16'(75);
			13178: out = 16'(4336);
			13179: out = 16'(8679);
			13180: out = 16'(1854);
			13181: out = 16'(-1279);
			13182: out = 16'(-4173);
			13183: out = 16'(-236);
			13184: out = 16'(-1);
			13185: out = 16'(-4430);
			13186: out = 16'(-891);
			13187: out = 16'(-1169);
			13188: out = 16'(-4676);
			13189: out = 16'(-8073);
			13190: out = 16'(-7511);
			13191: out = 16'(7759);
			13192: out = 16'(5459);
			13193: out = 16'(2601);
			13194: out = 16'(227);
			13195: out = 16'(2388);
			13196: out = 16'(6350);
			13197: out = 16'(-1137);
			13198: out = 16'(-623);
			13199: out = 16'(417);
			13200: out = 16'(4577);
			13201: out = 16'(1819);
			13202: out = 16'(-5449);
			13203: out = 16'(-7002);
			13204: out = 16'(-5411);
			13205: out = 16'(2340);
			13206: out = 16'(4463);
			13207: out = 16'(5263);
			13208: out = 16'(-1926);
			13209: out = 16'(-1268);
			13210: out = 16'(-1427);
			13211: out = 16'(4289);
			13212: out = 16'(902);
			13213: out = 16'(-2173);
			13214: out = 16'(-8205);
			13215: out = 16'(-4372);
			13216: out = 16'(2933);
			13217: out = 16'(-11);
			13218: out = 16'(-911);
			13219: out = 16'(-4053);
			13220: out = 16'(249);
			13221: out = 16'(2181);
			13222: out = 16'(5467);
			13223: out = 16'(1404);
			13224: out = 16'(-1563);
			13225: out = 16'(-7662);
			13226: out = 16'(-3565);
			13227: out = 16'(-770);
			13228: out = 16'(1336);
			13229: out = 16'(-1422);
			13230: out = 16'(-3362);
			13231: out = 16'(-664);
			13232: out = 16'(3393);
			13233: out = 16'(7543);
			13234: out = 16'(5273);
			13235: out = 16'(3948);
			13236: out = 16'(1680);
			13237: out = 16'(60);
			13238: out = 16'(-285);
			13239: out = 16'(1008);
			13240: out = 16'(1695);
			13241: out = 16'(-65);
			13242: out = 16'(-7952);
			13243: out = 16'(-3599);
			13244: out = 16'(175);
			13245: out = 16'(5879);
			13246: out = 16'(4925);
			13247: out = 16'(2867);
			13248: out = 16'(-2268);
			13249: out = 16'(-4133);
			13250: out = 16'(-4721);
			13251: out = 16'(339);
			13252: out = 16'(1911);
			13253: out = 16'(3033);
			13254: out = 16'(-954);
			13255: out = 16'(-1673);
			13256: out = 16'(-1625);
			13257: out = 16'(642);
			13258: out = 16'(-817);
			13259: out = 16'(-6478);
			13260: out = 16'(-4393);
			13261: out = 16'(-2173);
			13262: out = 16'(3531);
			13263: out = 16'(1077);
			13264: out = 16'(330);
			13265: out = 16'(1994);
			13266: out = 16'(3846);
			13267: out = 16'(4512);
			13268: out = 16'(-2152);
			13269: out = 16'(-3768);
			13270: out = 16'(-4612);
			13271: out = 16'(3134);
			13272: out = 16'(4559);
			13273: out = 16'(4963);
			13274: out = 16'(-1402);
			13275: out = 16'(-2003);
			13276: out = 16'(883);
			13277: out = 16'(3010);
			13278: out = 16'(3197);
			13279: out = 16'(-978);
			13280: out = 16'(316);
			13281: out = 16'(921);
			13282: out = 16'(4057);
			13283: out = 16'(1778);
			13284: out = 16'(-1043);
			13285: out = 16'(-9649);
			13286: out = 16'(-7814);
			13287: out = 16'(-3644);
			13288: out = 16'(2849);
			13289: out = 16'(5390);
			13290: out = 16'(5554);
			13291: out = 16'(2867);
			13292: out = 16'(-436);
			13293: out = 16'(-4112);
			13294: out = 16'(-1397);
			13295: out = 16'(1081);
			13296: out = 16'(5156);
			13297: out = 16'(-1259);
			13298: out = 16'(-5927);
			13299: out = 16'(-11204);
			13300: out = 16'(-4668);
			13301: out = 16'(1113);
			13302: out = 16'(450);
			13303: out = 16'(2289);
			13304: out = 16'(2407);
			13305: out = 16'(9009);
			13306: out = 16'(4660);
			13307: out = 16'(218);
			13308: out = 16'(-5698);
			13309: out = 16'(-2514);
			13310: out = 16'(4729);
			13311: out = 16'(1123);
			13312: out = 16'(-422);
			13313: out = 16'(-4359);
			13314: out = 16'(-1);
			13315: out = 16'(670);
			13316: out = 16'(-511);
			13317: out = 16'(-439);
			13318: out = 16'(8);
			13319: out = 16'(2158);
			13320: out = 16'(687);
			13321: out = 16'(-107);
			13322: out = 16'(694);
			13323: out = 16'(-425);
			13324: out = 16'(-1724);
			13325: out = 16'(108);
			13326: out = 16'(-917);
			13327: out = 16'(-1434);
			13328: out = 16'(-4741);
			13329: out = 16'(-2713);
			13330: out = 16'(1161);
			13331: out = 16'(5728);
			13332: out = 16'(6641);
			13333: out = 16'(4775);
			13334: out = 16'(-1097);
			13335: out = 16'(-4175);
			13336: out = 16'(-1131);
			13337: out = 16'(-611);
			13338: out = 16'(585);
			13339: out = 16'(-4336);
			13340: out = 16'(407);
			13341: out = 16'(2956);
			13342: out = 16'(-92);
			13343: out = 16'(-2044);
			13344: out = 16'(-3687);
			13345: out = 16'(605);
			13346: out = 16'(706);
			13347: out = 16'(-42);
			13348: out = 16'(1628);
			13349: out = 16'(3009);
			13350: out = 16'(5072);
			13351: out = 16'(-695);
			13352: out = 16'(-3522);
			13353: out = 16'(-3576);
			13354: out = 16'(-1859);
			13355: out = 16'(144);
			13356: out = 16'(-775);
			13357: out = 16'(-623);
			13358: out = 16'(-1221);
			13359: out = 16'(5522);
			13360: out = 16'(2382);
			13361: out = 16'(867);
			13362: out = 16'(-6386);
			13363: out = 16'(-169);
			13364: out = 16'(7342);
			13365: out = 16'(7168);
			13366: out = 16'(2747);
			13367: out = 16'(-4389);
			13368: out = 16'(-9809);
			13369: out = 16'(-8091);
			13370: out = 16'(1578);
			13371: out = 16'(6301);
			13372: out = 16'(7552);
			13373: out = 16'(224);
			13374: out = 16'(-3385);
			13375: out = 16'(-5443);
			13376: out = 16'(5362);
			13377: out = 16'(2848);
			13378: out = 16'(1800);
			13379: out = 16'(-376);
			13380: out = 16'(818);
			13381: out = 16'(1641);
			13382: out = 16'(-1102);
			13383: out = 16'(-3106);
			13384: out = 16'(-5117);
			13385: out = 16'(651);
			13386: out = 16'(2423);
			13387: out = 16'(2966);
			13388: out = 16'(-1347);
			13389: out = 16'(-1798);
			13390: out = 16'(3267);
			13391: out = 16'(2041);
			13392: out = 16'(753);
			13393: out = 16'(-5235);
			13394: out = 16'(-3712);
			13395: out = 16'(-2191);
			13396: out = 16'(774);
			13397: out = 16'(917);
			13398: out = 16'(672);
			13399: out = 16'(-3371);
			13400: out = 16'(-3435);
			13401: out = 16'(-2251);
			13402: out = 16'(4566);
			13403: out = 16'(5342);
			13404: out = 16'(2450);
			13405: out = 16'(3079);
			13406: out = 16'(3463);
			13407: out = 16'(7046);
			13408: out = 16'(-1798);
			13409: out = 16'(-7282);
			13410: out = 16'(-11365);
			13411: out = 16'(-5889);
			13412: out = 16'(12);
			13413: out = 16'(-23);
			13414: out = 16'(5729);
			13415: out = 16'(7952);
			13416: out = 16'(1440);
			13417: out = 16'(-623);
			13418: out = 16'(-1762);
			13419: out = 16'(89);
			13420: out = 16'(-230);
			13421: out = 16'(-2036);
			13422: out = 16'(3157);
			13423: out = 16'(2475);
			13424: out = 16'(-552);
			13425: out = 16'(-3067);
			13426: out = 16'(-4050);
			13427: out = 16'(-2775);
			13428: out = 16'(-823);
			13429: out = 16'(1946);
			13430: out = 16'(6669);
			13431: out = 16'(3206);
			13432: out = 16'(-550);
			13433: out = 16'(-4698);
			13434: out = 16'(-4241);
			13435: out = 16'(-2229);
			13436: out = 16'(69);
			13437: out = 16'(-215);
			13438: out = 16'(-1739);
			13439: out = 16'(181);
			13440: out = 16'(2712);
			13441: out = 16'(7011);
			13442: out = 16'(1653);
			13443: out = 16'(-1867);
			13444: out = 16'(-7977);
			13445: out = 16'(-2159);
			13446: out = 16'(1580);
			13447: out = 16'(7927);
			13448: out = 16'(651);
			13449: out = 16'(-3039);
			13450: out = 16'(-642);
			13451: out = 16'(1310);
			13452: out = 16'(2201);
			13453: out = 16'(-4637);
			13454: out = 16'(-5228);
			13455: out = 16'(-4473);
			13456: out = 16'(-235);
			13457: out = 16'(829);
			13458: out = 16'(-352);
			13459: out = 16'(6175);
			13460: out = 16'(4475);
			13461: out = 16'(333);
			13462: out = 16'(-7508);
			13463: out = 16'(-6866);
			13464: out = 16'(4760);
			13465: out = 16'(3505);
			13466: out = 16'(2484);
			13467: out = 16'(-6717);
			13468: out = 16'(-2369);
			13469: out = 16'(11);
			13470: out = 16'(2054);
			13471: out = 16'(1260);
			13472: out = 16'(979);
			13473: out = 16'(-405);
			13474: out = 16'(2239);
			13475: out = 16'(4837);
			13476: out = 16'(2353);
			13477: out = 16'(-781);
			13478: out = 16'(-5413);
			13479: out = 16'(-539);
			13480: out = 16'(1606);
			13481: out = 16'(4011);
			13482: out = 16'(1209);
			13483: out = 16'(422);
			13484: out = 16'(653);
			13485: out = 16'(2127);
			13486: out = 16'(1521);
			13487: out = 16'(-5142);
			13488: out = 16'(-5180);
			13489: out = 16'(-3572);
			13490: out = 16'(7900);
			13491: out = 16'(6921);
			13492: out = 16'(4339);
			13493: out = 16'(-8370);
			13494: out = 16'(-8888);
			13495: out = 16'(-5561);
			13496: out = 16'(-1339);
			13497: out = 16'(182);
			13498: out = 16'(-571);
			13499: out = 16'(-1203);
			13500: out = 16'(-967);
			13501: out = 16'(817);
			13502: out = 16'(218);
			13503: out = 16'(577);
			13504: out = 16'(4481);
			13505: out = 16'(-2318);
			13506: out = 16'(-6381);
			13507: out = 16'(-4643);
			13508: out = 16'(-1924);
			13509: out = 16'(1811);
			13510: out = 16'(2664);
			13511: out = 16'(4307);
			13512: out = 16'(4700);
			13513: out = 16'(-664);
			13514: out = 16'(-667);
			13515: out = 16'(1403);
			13516: out = 16'(6319);
			13517: out = 16'(5245);
			13518: out = 16'(-2620);
			13519: out = 16'(-208);
			13520: out = 16'(-840);
			13521: out = 16'(1538);
			13522: out = 16'(-4234);
			13523: out = 16'(-6214);
			13524: out = 16'(-7728);
			13525: out = 16'(142);
			13526: out = 16'(5920);
			13527: out = 16'(5732);
			13528: out = 16'(2456);
			13529: out = 16'(-2319);
			13530: out = 16'(-107);
			13531: out = 16'(-676);
			13532: out = 16'(159);
			13533: out = 16'(-1561);
			13534: out = 16'(-1329);
			13535: out = 16'(-1622);
			13536: out = 16'(594);
			13537: out = 16'(1228);
			13538: out = 16'(2109);
			13539: out = 16'(1842);
			13540: out = 16'(1424);
			13541: out = 16'(-1847);
			13542: out = 16'(-689);
			13543: out = 16'(146);
			13544: out = 16'(6149);
			13545: out = 16'(2109);
			13546: out = 16'(-1087);
			13547: out = 16'(-9606);
			13548: out = 16'(-3017);
			13549: out = 16'(6004);
			13550: out = 16'(5391);
			13551: out = 16'(2877);
			13552: out = 16'(-3599);
			13553: out = 16'(-722);
			13554: out = 16'(1326);
			13555: out = 16'(7217);
			13556: out = 16'(2645);
			13557: out = 16'(-496);
			13558: out = 16'(-9349);
			13559: out = 16'(-3000);
			13560: out = 16'(422);
			13561: out = 16'(5174);
			13562: out = 16'(-1080);
			13563: out = 16'(-5767);
			13564: out = 16'(-7370);
			13565: out = 16'(-2742);
			13566: out = 16'(2773);
			13567: out = 16'(797);
			13568: out = 16'(-157);
			13569: out = 16'(-2924);
			13570: out = 16'(433);
			13571: out = 16'(1050);
			13572: out = 16'(2247);
			13573: out = 16'(31);
			13574: out = 16'(-688);
			13575: out = 16'(-1605);
			13576: out = 16'(-642);
			13577: out = 16'(-127);
			13578: out = 16'(1184);
			13579: out = 16'(-593);
			13580: out = 16'(-1363);
			13581: out = 16'(-496);
			13582: out = 16'(1988);
			13583: out = 16'(4019);
			13584: out = 16'(-117);
			13585: out = 16'(408);
			13586: out = 16'(618);
			13587: out = 16'(3708);
			13588: out = 16'(2216);
			13589: out = 16'(-526);
			13590: out = 16'(-445);
			13591: out = 16'(-1255);
			13592: out = 16'(-2973);
			13593: out = 16'(790);
			13594: out = 16'(1993);
			13595: out = 16'(1859);
			13596: out = 16'(223);
			13597: out = 16'(-1047);
			13598: out = 16'(-2902);
			13599: out = 16'(-31);
			13600: out = 16'(2656);
			13601: out = 16'(6505);
			13602: out = 16'(3005);
			13603: out = 16'(-1892);
			13604: out = 16'(-6655);
			13605: out = 16'(-5029);
			13606: out = 16'(767);
			13607: out = 16'(-2111);
			13608: out = 16'(-655);
			13609: out = 16'(-897);
			13610: out = 16'(4208);
			13611: out = 16'(3531);
			13612: out = 16'(892);
			13613: out = 16'(-1128);
			13614: out = 16'(-1789);
			13615: out = 16'(-3162);
			13616: out = 16'(1677);
			13617: out = 16'(3765);
			13618: out = 16'(3117);
			13619: out = 16'(-1622);
			13620: out = 16'(-5316);
			13621: out = 16'(-3000);
			13622: out = 16'(-71);
			13623: out = 16'(3284);
			13624: out = 16'(2761);
			13625: out = 16'(2369);
			13626: out = 16'(1648);
			13627: out = 16'(-3028);
			13628: out = 16'(-2994);
			13629: out = 16'(-517);
			13630: out = 16'(5049);
			13631: out = 16'(3862);
			13632: out = 16'(-6864);
			13633: out = 16'(-6758);
			13634: out = 16'(-6113);
			13635: out = 16'(2447);
			13636: out = 16'(-1015);
			13637: out = 16'(-2065);
			13638: out = 16'(1837);
			13639: out = 16'(2077);
			13640: out = 16'(1619);
			13641: out = 16'(-2206);
			13642: out = 16'(-1860);
			13643: out = 16'(64);
			13644: out = 16'(2257);
			13645: out = 16'(3881);
			13646: out = 16'(4653);
			13647: out = 16'(823);
			13648: out = 16'(-1904);
			13649: out = 16'(-3775);
			13650: out = 16'(-1736);
			13651: out = 16'(644);
			13652: out = 16'(2681);
			13653: out = 16'(3701);
			13654: out = 16'(2527);
			13655: out = 16'(-3615);
			13656: out = 16'(-5241);
			13657: out = 16'(-5153);
			13658: out = 16'(5363);
			13659: out = 16'(3898);
			13660: out = 16'(1344);
			13661: out = 16'(-3287);
			13662: out = 16'(-1396);
			13663: out = 16'(3404);
			13664: out = 16'(1878);
			13665: out = 16'(-394);
			13666: out = 16'(-6859);
			13667: out = 16'(-531);
			13668: out = 16'(1635);
			13669: out = 16'(4149);
			13670: out = 16'(1520);
			13671: out = 16'(668);
			13672: out = 16'(-998);
			13673: out = 16'(2256);
			13674: out = 16'(4062);
			13675: out = 16'(7660);
			13676: out = 16'(138);
			13677: out = 16'(-7550);
			13678: out = 16'(-6070);
			13679: out = 16'(-4155);
			13680: out = 16'(659);
			13681: out = 16'(-1274);
			13682: out = 16'(2116);
			13683: out = 16'(5685);
			13684: out = 16'(1822);
			13685: out = 16'(215);
			13686: out = 16'(546);
			13687: out = 16'(-311);
			13688: out = 16'(-1244);
			13689: out = 16'(-5506);
			13690: out = 16'(-1842);
			13691: out = 16'(320);
			13692: out = 16'(2946);
			13693: out = 16'(-355);
			13694: out = 16'(-3074);
			13695: out = 16'(-1674);
			13696: out = 16'(-536);
			13697: out = 16'(991);
			13698: out = 16'(-1487);
			13699: out = 16'(-1203);
			13700: out = 16'(-483);
			13701: out = 16'(-2410);
			13702: out = 16'(-1656);
			13703: out = 16'(887);
			13704: out = 16'(1556);
			13705: out = 16'(1323);
			13706: out = 16'(-1895);
			13707: out = 16'(-614);
			13708: out = 16'(212);
			13709: out = 16'(4225);
			13710: out = 16'(2403);
			13711: out = 16'(899);
			13712: out = 16'(-7550);
			13713: out = 16'(-3530);
			13714: out = 16'(536);
			13715: out = 16'(8192);
			13716: out = 16'(3857);
			13717: out = 16'(-2525);
			13718: out = 16'(-6721);
			13719: out = 16'(-3160);
			13720: out = 16'(5813);
			13721: out = 16'(1120);
			13722: out = 16'(-1818);
			13723: out = 16'(-9090);
			13724: out = 16'(-1993);
			13725: out = 16'(332);
			13726: out = 16'(-111);
			13727: out = 16'(805);
			13728: out = 16'(996);
			13729: out = 16'(1246);
			13730: out = 16'(-2252);
			13731: out = 16'(-4571);
			13732: out = 16'(1077);
			13733: out = 16'(1453);
			13734: out = 16'(2248);
			13735: out = 16'(-257);
			13736: out = 16'(-169);
			13737: out = 16'(-451);
			13738: out = 16'(129);
			13739: out = 16'(746);
			13740: out = 16'(3504);
			13741: out = 16'(-4173);
			13742: out = 16'(-5726);
			13743: out = 16'(-4765);
			13744: out = 16'(3553);
			13745: out = 16'(6997);
			13746: out = 16'(2724);
			13747: out = 16'(1314);
			13748: out = 16'(-211);
			13749: out = 16'(5297);
			13750: out = 16'(2950);
			13751: out = 16'(1483);
			13752: out = 16'(-2544);
			13753: out = 16'(-2200);
			13754: out = 16'(-1284);
			13755: out = 16'(3238);
			13756: out = 16'(4176);
			13757: out = 16'(4704);
			13758: out = 16'(-1635);
			13759: out = 16'(-1419);
			13760: out = 16'(3113);
			13761: out = 16'(3314);
			13762: out = 16'(1830);
			13763: out = 16'(-5785);
			13764: out = 16'(-2665);
			13765: out = 16'(-1142);
			13766: out = 16'(2055);
			13767: out = 16'(225);
			13768: out = 16'(-1232);
			13769: out = 16'(-7386);
			13770: out = 16'(-3277);
			13771: out = 16'(1576);
			13772: out = 16'(5249);
			13773: out = 16'(4335);
			13774: out = 16'(1241);
			13775: out = 16'(-1747);
			13776: out = 16'(-2761);
			13777: out = 16'(-1248);
			13778: out = 16'(-707);
			13779: out = 16'(295);
			13780: out = 16'(446);
			13781: out = 16'(210);
			13782: out = 16'(-364);
			13783: out = 16'(-380);
			13784: out = 16'(-351);
			13785: out = 16'(275);
			13786: out = 16'(2992);
			13787: out = 16'(-1156);
			13788: out = 16'(-4989);
			13789: out = 16'(2887);
			13790: out = 16'(2513);
			13791: out = 16'(2843);
			13792: out = 16'(-5428);
			13793: out = 16'(-3930);
			13794: out = 16'(-250);
			13795: out = 16'(2606);
			13796: out = 16'(917);
			13797: out = 16'(-3859);
			13798: out = 16'(-7139);
			13799: out = 16'(-6075);
			13800: out = 16'(2547);
			13801: out = 16'(3256);
			13802: out = 16'(3393);
			13803: out = 16'(-2685);
			13804: out = 16'(-1608);
			13805: out = 16'(-1269);
			13806: out = 16'(219);
			13807: out = 16'(-652);
			13808: out = 16'(-1176);
			13809: out = 16'(-50);
			13810: out = 16'(584);
			13811: out = 16'(1010);
			13812: out = 16'(-4530);
			13813: out = 16'(-5038);
			13814: out = 16'(-1653);
			13815: out = 16'(33);
			13816: out = 16'(2308);
			13817: out = 16'(1753);
			13818: out = 16'(6627);
			13819: out = 16'(6385);
			13820: out = 16'(1261);
			13821: out = 16'(-1235);
			13822: out = 16'(-2126);
			13823: out = 16'(756);
			13824: out = 16'(3666);
			13825: out = 16'(5705);
			13826: out = 16'(2348);
			13827: out = 16'(-2031);
			13828: out = 16'(-7687);
			13829: out = 16'(1083);
			13830: out = 16'(2873);
			13831: out = 16'(5250);
			13832: out = 16'(95);
			13833: out = 16'(584);
			13834: out = 16'(2651);
			13835: out = 16'(2491);
			13836: out = 16'(-241);
			13837: out = 16'(-4559);
			13838: out = 16'(-10706);
			13839: out = 16'(-12277);
			13840: out = 16'(-3727);
			13841: out = 16'(742);
			13842: out = 16'(5152);
			13843: out = 16'(4631);
			13844: out = 16'(4557);
			13845: out = 16'(2311);
			13846: out = 16'(723);
			13847: out = 16'(-265);
			13848: out = 16'(1054);
			13849: out = 16'(-1523);
			13850: out = 16'(-2500);
			13851: out = 16'(-6804);
			13852: out = 16'(2298);
			13853: out = 16'(2790);
			13854: out = 16'(419);
			13855: out = 16'(-10333);
			13856: out = 16'(-11717);
			13857: out = 16'(6573);
			13858: out = 16'(8304);
			13859: out = 16'(8963);
			13860: out = 16'(-7396);
			13861: out = 16'(-3067);
			13862: out = 16'(752);
			13863: out = 16'(7418);
			13864: out = 16'(4152);
			13865: out = 16'(-842);
			13866: out = 16'(-3030);
			13867: out = 16'(-3964);
			13868: out = 16'(-3470);
			13869: out = 16'(750);
			13870: out = 16'(3399);
			13871: out = 16'(6035);
			13872: out = 16'(-2639);
			13873: out = 16'(-7085);
			13874: out = 16'(-6950);
			13875: out = 16'(-871);
			13876: out = 16'(4097);
			13877: out = 16'(356);
			13878: out = 16'(1148);
			13879: out = 16'(-943);
			13880: out = 16'(3080);
			13881: out = 16'(-1436);
			13882: out = 16'(-3716);
			13883: out = 16'(-13193);
			13884: out = 16'(-6179);
			13885: out = 16'(4660);
			13886: out = 16'(9456);
			13887: out = 16'(7406);
			13888: out = 16'(-690);
			13889: out = 16'(-1530);
			13890: out = 16'(-1293);
			13891: out = 16'(3629);
			13892: out = 16'(2988);
			13893: out = 16'(2296);
			13894: out = 16'(-1433);
			13895: out = 16'(-3450);
			13896: out = 16'(-4290);
			13897: out = 16'(-52);
			13898: out = 16'(2724);
			13899: out = 16'(5086);
			13900: out = 16'(-148);
			13901: out = 16'(-759);
			13902: out = 16'(-1262);
			13903: out = 16'(3385);
			13904: out = 16'(4471);
			13905: out = 16'(4616);
			13906: out = 16'(-926);
			13907: out = 16'(-4903);
			13908: out = 16'(-8347);
			13909: out = 16'(-4289);
			13910: out = 16'(-1785);
			13911: out = 16'(-2855);
			13912: out = 16'(190);
			13913: out = 16'(1628);
			13914: out = 16'(6709);
			13915: out = 16'(741);
			13916: out = 16'(-3244);
			13917: out = 16'(-8365);
			13918: out = 16'(-1727);
			13919: out = 16'(5460);
			13920: out = 16'(8271);
			13921: out = 16'(5533);
			13922: out = 16'(-434);
			13923: out = 16'(-6402);
			13924: out = 16'(-8823);
			13925: out = 16'(-7570);
			13926: out = 16'(-185);
			13927: out = 16'(2920);
			13928: out = 16'(966);
			13929: out = 16'(586);
			13930: out = 16'(1354);
			13931: out = 16'(8389);
			13932: out = 16'(5227);
			13933: out = 16'(3204);
			13934: out = 16'(-1431);
			13935: out = 16'(-750);
			13936: out = 16'(-949);
			13937: out = 16'(-5570);
			13938: out = 16'(-5004);
			13939: out = 16'(-2826);
			13940: out = 16'(-541);
			13941: out = 16'(1749);
			13942: out = 16'(3370);
			13943: out = 16'(3285);
			13944: out = 16'(2574);
			13945: out = 16'(879);
			13946: out = 16'(1197);
			13947: out = 16'(-1060);
			13948: out = 16'(-6041);
			13949: out = 16'(-4294);
			13950: out = 16'(-2755);
			13951: out = 16'(-1206);
			13952: out = 16'(-436);
			13953: out = 16'(719);
			13954: out = 16'(4178);
			13955: out = 16'(5247);
			13956: out = 16'(5666);
			13957: out = 16'(-1915);
			13958: out = 16'(-1445);
			13959: out = 16'(159);
			13960: out = 16'(6160);
			13961: out = 16'(4905);
			13962: out = 16'(425);
			13963: out = 16'(-1537);
			13964: out = 16'(-2909);
			13965: out = 16'(-2328);
			13966: out = 16'(648);
			13967: out = 16'(2212);
			13968: out = 16'(471);
			13969: out = 16'(-1156);
			13970: out = 16'(-1600);
			13971: out = 16'(7364);
			13972: out = 16'(2434);
			13973: out = 16'(-268);
			13974: out = 16'(-767);
			13975: out = 16'(2662);
			13976: out = 16'(5562);
			13977: out = 16'(-860);
			13978: out = 16'(-2003);
			13979: out = 16'(-1357);
			13980: out = 16'(-224);
			13981: out = 16'(668);
			13982: out = 16'(-1139);
			13983: out = 16'(4854);
			13984: out = 16'(3785);
			13985: out = 16'(-7);
			13986: out = 16'(-7938);
			13987: out = 16'(-9415);
			13988: out = 16'(-227);
			13989: out = 16'(5533);
			13990: out = 16'(8566);
			13991: out = 16'(-1558);
			13992: out = 16'(-3710);
			13993: out = 16'(-6283);
			13994: out = 16'(473);
			13995: out = 16'(-118);
			13996: out = 16'(-214);
			13997: out = 16'(-764);
			13998: out = 16'(1028);
			13999: out = 16'(2909);
			14000: out = 16'(650);
			14001: out = 16'(-1384);
			14002: out = 16'(-3740);
			14003: out = 16'(-837);
			14004: out = 16'(2003);
			14005: out = 16'(4702);
			14006: out = 16'(3262);
			14007: out = 16'(76);
			14008: out = 16'(-5548);
			14009: out = 16'(-8417);
			14010: out = 16'(-8421);
			14011: out = 16'(-148);
			14012: out = 16'(5196);
			14013: out = 16'(9406);
			14014: out = 16'(-525);
			14015: out = 16'(-3544);
			14016: out = 16'(-7510);
			14017: out = 16'(5813);
			14018: out = 16'(6112);
			14019: out = 16'(2873);
			14020: out = 16'(-5685);
			14021: out = 16'(-7611);
			14022: out = 16'(-3445);
			14023: out = 16'(2346);
			14024: out = 16'(4607);
			14025: out = 16'(3);
			14026: out = 16'(-5434);
			14027: out = 16'(-8194);
			14028: out = 16'(7113);
			14029: out = 16'(5547);
			14030: out = 16'(4792);
			14031: out = 16'(-1359);
			14032: out = 16'(727);
			14033: out = 16'(2912);
			14034: out = 16'(1367);
			14035: out = 16'(-3583);
			14036: out = 16'(-11424);
			14037: out = 16'(-2393);
			14038: out = 16'(1396);
			14039: out = 16'(4302);
			14040: out = 16'(3909);
			14041: out = 16'(3364);
			14042: out = 16'(-566);
			14043: out = 16'(2237);
			14044: out = 16'(3628);
			14045: out = 16'(9782);
			14046: out = 16'(2546);
			14047: out = 16'(-3121);
			14048: out = 16'(-11031);
			14049: out = 16'(-4845);
			14050: out = 16'(3107);
			14051: out = 16'(6162);
			14052: out = 16'(2676);
			14053: out = 16'(-4745);
			14054: out = 16'(-2754);
			14055: out = 16'(-406);
			14056: out = 16'(5381);
			14057: out = 16'(4519);
			14058: out = 16'(2987);
			14059: out = 16'(-3442);
			14060: out = 16'(-3279);
			14061: out = 16'(-3745);
			14062: out = 16'(-176);
			14063: out = 16'(-1608);
			14064: out = 16'(-1101);
			14065: out = 16'(-508);
			14066: out = 16'(654);
			14067: out = 16'(863);
			14068: out = 16'(3008);
			14069: out = 16'(1723);
			14070: out = 16'(795);
			14071: out = 16'(-367);
			14072: out = 16'(300);
			14073: out = 16'(532);
			14074: out = 16'(1946);
			14075: out = 16'(383);
			14076: out = 16'(-1547);
			14077: out = 16'(-6945);
			14078: out = 16'(-7545);
			14079: out = 16'(-3759);
			14080: out = 16'(2025);
			14081: out = 16'(5064);
			14082: out = 16'(1803);
			14083: out = 16'(180);
			14084: out = 16'(-1746);
			14085: out = 16'(673);
			14086: out = 16'(668);
			14087: out = 16'(942);
			14088: out = 16'(647);
			14089: out = 16'(193);
			14090: out = 16'(-336);
			14091: out = 16'(-5255);
			14092: out = 16'(-4713);
			14093: out = 16'(-1053);
			14094: out = 16'(1239);
			14095: out = 16'(1186);
			14096: out = 16'(-2862);
			14097: out = 16'(-1620);
			14098: out = 16'(-321);
			14099: out = 16'(4345);
			14100: out = 16'(1417);
			14101: out = 16'(0);
			14102: out = 16'(2095);
			14103: out = 16'(1928);
			14104: out = 16'(938);
			14105: out = 16'(-10007);
			14106: out = 16'(-9327);
			14107: out = 16'(-5860);
			14108: out = 16'(4402);
			14109: out = 16'(6297);
			14110: out = 16'(4697);
			14111: out = 16'(1254);
			14112: out = 16'(-679);
			14113: out = 16'(-1207);
			14114: out = 16'(3165);
			14115: out = 16'(6225);
			14116: out = 16'(8367);
			14117: out = 16'(2720);
			14118: out = 16'(-2634);
			14119: out = 16'(-7064);
			14120: out = 16'(-4521);
			14121: out = 16'(-160);
			14122: out = 16'(2323);
			14123: out = 16'(1282);
			14124: out = 16'(-2153);
			14125: out = 16'(3305);
			14126: out = 16'(2181);
			14127: out = 16'(3371);
			14128: out = 16'(-4771);
			14129: out = 16'(-2008);
			14130: out = 16'(1698);
			14131: out = 16'(9776);
			14132: out = 16'(6642);
			14133: out = 16'(-3055);
			14134: out = 16'(-11661);
			14135: out = 16'(-13842);
			14136: out = 16'(-5958);
			14137: out = 16'(1422);
			14138: out = 16'(7753);
			14139: out = 16'(10770);
			14140: out = 16'(6083);
			14141: out = 16'(701);
			14142: out = 16'(-1457);
			14143: out = 16'(1593);
			14144: out = 16'(5849);
			14145: out = 16'(3125);
			14146: out = 16'(-1441);
			14147: out = 16'(-8353);
			14148: out = 16'(-10491);
			14149: out = 16'(-8051);
			14150: out = 16'(440);
			14151: out = 16'(1796);
			14152: out = 16'(3060);
			14153: out = 16'(573);
			14154: out = 16'(1005);
			14155: out = 16'(475);
			14156: out = 16'(1043);
			14157: out = 16'(219);
			14158: out = 16'(131);
			14159: out = 16'(4005);
			14160: out = 16'(1402);
			14161: out = 16'(-1494);
			14162: out = 16'(-10297);
			14163: out = 16'(-7977);
			14164: out = 16'(-2540);
			14165: out = 16'(5371);
			14166: out = 16'(5934);
			14167: out = 16'(2520);
			14168: out = 16'(-1231);
			14169: out = 16'(-2599);
			14170: out = 16'(-1383);
			14171: out = 16'(3937);
			14172: out = 16'(4240);
			14173: out = 16'(-4147);
			14174: out = 16'(-4284);
			14175: out = 16'(-3959);
			14176: out = 16'(2137);
			14177: out = 16'(2518);
			14178: out = 16'(2872);
			14179: out = 16'(79);
			14180: out = 16'(-1245);
			14181: out = 16'(-2259);
			14182: out = 16'(4067);
			14183: out = 16'(6783);
			14184: out = 16'(9075);
			14185: out = 16'(1042);
			14186: out = 16'(-2844);
			14187: out = 16'(-6546);
			14188: out = 16'(-809);
			14189: out = 16'(540);
			14190: out = 16'(-1920);
			14191: out = 16'(-2240);
			14192: out = 16'(-2118);
			14193: out = 16'(2302);
			14194: out = 16'(-429);
			14195: out = 16'(-2098);
			14196: out = 16'(-6276);
			14197: out = 16'(-1767);
			14198: out = 16'(3261);
			14199: out = 16'(7785);
			14200: out = 16'(6708);
			14201: out = 16'(2680);
			14202: out = 16'(-1246);
			14203: out = 16'(-5514);
			14204: out = 16'(-8448);
			14205: out = 16'(-5921);
			14206: out = 16'(-3505);
			14207: out = 16'(-1356);
			14208: out = 16'(207);
			14209: out = 16'(994);
			14210: out = 16'(685);
			14211: out = 16'(2368);
			14212: out = 16'(3795);
			14213: out = 16'(6910);
			14214: out = 16'(2756);
			14215: out = 16'(-1187);
			14216: out = 16'(-32);
			14217: out = 16'(-661);
			14218: out = 16'(49);
			14219: out = 16'(-3676);
			14220: out = 16'(-1883);
			14221: out = 16'(58);
			14222: out = 16'(1823);
			14223: out = 16'(1437);
			14224: out = 16'(826);
			14225: out = 16'(-238);
			14226: out = 16'(1217);
			14227: out = 16'(3619);
			14228: out = 16'(5323);
			14229: out = 16'(4639);
			14230: out = 16'(3051);
			14231: out = 16'(-2209);
			14232: out = 16'(-6133);
			14233: out = 16'(-12153);
			14234: out = 16'(-5336);
			14235: out = 16'(2053);
			14236: out = 16'(5382);
			14237: out = 16'(945);
			14238: out = 16'(-6606);
			14239: out = 16'(-842);
			14240: out = 16'(3289);
			14241: out = 16'(10668);
			14242: out = 16'(1163);
			14243: out = 16'(-2681);
			14244: out = 16'(-8835);
			14245: out = 16'(-1350);
			14246: out = 16'(372);
			14247: out = 16'(-1302);
			14248: out = 16'(-2251);
			14249: out = 16'(-1320);
			14250: out = 16'(2756);
			14251: out = 16'(5239);
			14252: out = 16'(6327);
			14253: out = 16'(3030);
			14254: out = 16'(1644);
			14255: out = 16'(252);
			14256: out = 16'(-265);
			14257: out = 16'(1572);
			14258: out = 16'(4744);
			14259: out = 16'(163);
			14260: out = 16'(-3117);
			14261: out = 16'(-8886);
			14262: out = 16'(-1412);
			14263: out = 16'(1745);
			14264: out = 16'(4989);
			14265: out = 16'(130);
			14266: out = 16'(-1759);
			14267: out = 16'(-1900);
			14268: out = 16'(3824);
			14269: out = 16'(7096);
			14270: out = 16'(2542);
			14271: out = 16'(508);
			14272: out = 16'(-2439);
			14273: out = 16'(-1539);
			14274: out = 16'(-1036);
			14275: out = 16'(834);
			14276: out = 16'(-3389);
			14277: out = 16'(-6039);
			14278: out = 16'(-11219);
			14279: out = 16'(470);
			14280: out = 16'(3887);
			14281: out = 16'(5994);
			14282: out = 16'(-1366);
			14283: out = 16'(-3218);
			14284: out = 16'(-628);
			14285: out = 16'(4688);
			14286: out = 16'(6681);
			14287: out = 16'(1870);
			14288: out = 16'(-2563);
			14289: out = 16'(-6109);
			14290: out = 16'(-524);
			14291: out = 16'(3509);
			14292: out = 16'(8439);
			14293: out = 16'(916);
			14294: out = 16'(-385);
			14295: out = 16'(-3475);
			14296: out = 16'(2304);
			14297: out = 16'(1470);
			14298: out = 16'(861);
			14299: out = 16'(-5131);
			14300: out = 16'(-4622);
			14301: out = 16'(174);
			14302: out = 16'(2850);
			14303: out = 16'(1995);
			14304: out = 16'(-3561);
			14305: out = 16'(-8335);
			14306: out = 16'(-10231);
			14307: out = 16'(-4175);
			14308: out = 16'(395);
			14309: out = 16'(4691);
			14310: out = 16'(6351);
			14311: out = 16'(3661);
			14312: out = 16'(-1548);
			14313: out = 16'(-4957);
			14314: out = 16'(-4500);
			14315: out = 16'(760);
			14316: out = 16'(-729);
			14317: out = 16'(111);
			14318: out = 16'(-2104);
			14319: out = 16'(780);
			14320: out = 16'(-1425);
			14321: out = 16'(-6741);
			14322: out = 16'(-6686);
			14323: out = 16'(-3755);
			14324: out = 16'(1589);
			14325: out = 16'(5805);
			14326: out = 16'(7416);
			14327: out = 16'(6408);
			14328: out = 16'(5);
			14329: out = 16'(-6427);
			14330: out = 16'(-1780);
			14331: out = 16'(2080);
			14332: out = 16'(7952);
			14333: out = 16'(-3126);
			14334: out = 16'(-5880);
			14335: out = 16'(-8279);
			14336: out = 16'(2112);
			14337: out = 16'(5551);
			14338: out = 16'(4708);
			14339: out = 16'(2345);
			14340: out = 16'(322);
			14341: out = 16'(30);
			14342: out = 16'(241);
			14343: out = 16'(275);
			14344: out = 16'(-2696);
			14345: out = 16'(-859);
			14346: out = 16'(706);
			14347: out = 16'(-1526);
			14348: out = 16'(-846);
			14349: out = 16'(-155);
			14350: out = 16'(4445);
			14351: out = 16'(2524);
			14352: out = 16'(-1962);
			14353: out = 16'(-256);
			14354: out = 16'(1171);
			14355: out = 16'(5138);
			14356: out = 16'(-161);
			14357: out = 16'(-1835);
			14358: out = 16'(-1578);
			14359: out = 16'(1249);
			14360: out = 16'(2904);
			14361: out = 16'(415);
			14362: out = 16'(2167);
			14363: out = 16'(2652);
			14364: out = 16'(3818);
			14365: out = 16'(1718);
			14366: out = 16'(269);
			14367: out = 16'(1351);
			14368: out = 16'(1209);
			14369: out = 16'(-132);
			14370: out = 16'(2604);
			14371: out = 16'(1313);
			14372: out = 16'(606);
			14373: out = 16'(-7878);
			14374: out = 16'(-9033);
			14375: out = 16'(-6178);
			14376: out = 16'(2231);
			14377: out = 16'(5594);
			14378: out = 16'(2573);
			14379: out = 16'(-1957);
			14380: out = 16'(-5057);
			14381: out = 16'(-456);
			14382: out = 16'(1063);
			14383: out = 16'(2949);
			14384: out = 16'(688);
			14385: out = 16'(-270);
			14386: out = 16'(-2031);
			14387: out = 16'(-2618);
			14388: out = 16'(-1075);
			14389: out = 16'(2110);
			14390: out = 16'(96);
			14391: out = 16'(-2571);
			14392: out = 16'(-8806);
			14393: out = 16'(-3066);
			14394: out = 16'(734);
			14395: out = 16'(7177);
			14396: out = 16'(1632);
			14397: out = 16'(-720);
			14398: out = 16'(-512);
			14399: out = 16'(1020);
			14400: out = 16'(1813);
			14401: out = 16'(751);
			14402: out = 16'(-1137);
			14403: out = 16'(-2538);
			14404: out = 16'(-386);
			14405: out = 16'(1619);
			14406: out = 16'(3933);
			14407: out = 16'(1308);
			14408: out = 16'(-1471);
			14409: out = 16'(-6421);
			14410: out = 16'(-320);
			14411: out = 16'(2270);
			14412: out = 16'(6055);
			14413: out = 16'(-1946);
			14414: out = 16'(-5781);
			14415: out = 16'(-7074);
			14416: out = 16'(-2037);
			14417: out = 16'(1803);
			14418: out = 16'(383);
			14419: out = 16'(1013);
			14420: out = 16'(834);
			14421: out = 16'(4001);
			14422: out = 16'(2828);
			14423: out = 16'(1902);
			14424: out = 16'(2757);
			14425: out = 16'(1730);
			14426: out = 16'(-665);
			14427: out = 16'(962);
			14428: out = 16'(51);
			14429: out = 16'(-398);
			14430: out = 16'(-5736);
			14431: out = 16'(-6510);
			14432: out = 16'(-3400);
			14433: out = 16'(-625);
			14434: out = 16'(2347);
			14435: out = 16'(5727);
			14436: out = 16'(2412);
			14437: out = 16'(-751);
			14438: out = 16'(228);
			14439: out = 16'(-418);
			14440: out = 16'(-65);
			14441: out = 16'(-2565);
			14442: out = 16'(-1926);
			14443: out = 16'(-1349);
			14444: out = 16'(1721);
			14445: out = 16'(840);
			14446: out = 16'(-1612);
			14447: out = 16'(-539);
			14448: out = 16'(-323);
			14449: out = 16'(-377);
			14450: out = 16'(-42);
			14451: out = 16'(293);
			14452: out = 16'(2212);
			14453: out = 16'(-945);
			14454: out = 16'(-2430);
			14455: out = 16'(-275);
			14456: out = 16'(-198);
			14457: out = 16'(187);
			14458: out = 16'(591);
			14459: out = 16'(1783);
			14460: out = 16'(2874);
			14461: out = 16'(-2083);
			14462: out = 16'(-2069);
			14463: out = 16'(-1210);
			14464: out = 16'(4716);
			14465: out = 16'(4055);
			14466: out = 16'(-612);
			14467: out = 16'(-939);
			14468: out = 16'(-1158);
			14469: out = 16'(1182);
			14470: out = 16'(1351);
			14471: out = 16'(1527);
			14472: out = 16'(-1805);
			14473: out = 16'(-1286);
			14474: out = 16'(-1358);
			14475: out = 16'(2158);
			14476: out = 16'(849);
			14477: out = 16'(660);
			14478: out = 16'(-3029);
			14479: out = 16'(1776);
			14480: out = 16'(6745);
			14481: out = 16'(5933);
			14482: out = 16'(889);
			14483: out = 16'(-8133);
			14484: out = 16'(-3495);
			14485: out = 16'(-1857);
			14486: out = 16'(738);
			14487: out = 16'(474);
			14488: out = 16'(1728);
			14489: out = 16'(4690);
			14490: out = 16'(1431);
			14491: out = 16'(-643);
			14492: out = 16'(525);
			14493: out = 16'(1422);
			14494: out = 16'(2847);
			14495: out = 16'(1362);
			14496: out = 16'(871);
			14497: out = 16'(-934);
			14498: out = 16'(1869);
			14499: out = 16'(-603);
			14500: out = 16'(-3104);
			14501: out = 16'(-6824);
			14502: out = 16'(-6576);
			14503: out = 16'(-4775);
			14504: out = 16'(310);
			14505: out = 16'(2160);
			14506: out = 16'(1899);
			14507: out = 16'(-1210);
			14508: out = 16'(-2345);
			14509: out = 16'(-127);
			14510: out = 16'(2231);
			14511: out = 16'(3641);
			14512: out = 16'(544);
			14513: out = 16'(-549);
			14514: out = 16'(-1899);
			14515: out = 16'(-2551);
			14516: out = 16'(-1748);
			14517: out = 16'(-85);
			14518: out = 16'(2422);
			14519: out = 16'(1839);
			14520: out = 16'(-859);
			14521: out = 16'(28);
			14522: out = 16'(-971);
			14523: out = 16'(-2676);
			14524: out = 16'(-382);
			14525: out = 16'(1850);
			14526: out = 16'(5896);
			14527: out = 16'(868);
			14528: out = 16'(-2406);
			14529: out = 16'(-3719);
			14530: out = 16'(-669);
			14531: out = 16'(2279);
			14532: out = 16'(596);
			14533: out = 16'(869);
			14534: out = 16'(432);
			14535: out = 16'(1696);
			14536: out = 16'(2462);
			14537: out = 16'(3646);
			14538: out = 16'(256);
			14539: out = 16'(-1563);
			14540: out = 16'(-4145);
			14541: out = 16'(-1188);
			14542: out = 16'(-1127);
			14543: out = 16'(-2723);
			14544: out = 16'(-4230);
			14545: out = 16'(-3471);
			14546: out = 16'(3262);
			14547: out = 16'(846);
			14548: out = 16'(-806);
			14549: out = 16'(-5989);
			14550: out = 16'(-2322);
			14551: out = 16'(1368);
			14552: out = 16'(2865);
			14553: out = 16'(729);
			14554: out = 16'(-3083);
			14555: out = 16'(-3107);
			14556: out = 16'(-2640);
			14557: out = 16'(336);
			14558: out = 16'(-1574);
			14559: out = 16'(-96);
			14560: out = 16'(927);
			14561: out = 16'(4977);
			14562: out = 16'(4491);
			14563: out = 16'(-72);
			14564: out = 16'(-2349);
			14565: out = 16'(-2585);
			14566: out = 16'(4173);
			14567: out = 16'(2551);
			14568: out = 16'(1764);
			14569: out = 16'(-295);
			14570: out = 16'(2336);
			14571: out = 16'(4430);
			14572: out = 16'(-3077);
			14573: out = 16'(-3442);
			14574: out = 16'(-2460);
			14575: out = 16'(-510);
			14576: out = 16'(-719);
			14577: out = 16'(-2705);
			14578: out = 16'(1121);
			14579: out = 16'(1861);
			14580: out = 16'(852);
			14581: out = 16'(-644);
			14582: out = 16'(-869);
			14583: out = 16'(3328);
			14584: out = 16'(1883);
			14585: out = 16'(1731);
			14586: out = 16'(-1945);
			14587: out = 16'(230);
			14588: out = 16'(822);
			14589: out = 16'(5170);
			14590: out = 16'(279);
			14591: out = 16'(-4167);
			14592: out = 16'(-9319);
			14593: out = 16'(-4865);
			14594: out = 16'(2725);
			14595: out = 16'(7288);
			14596: out = 16'(5955);
			14597: out = 16'(105);
			14598: out = 16'(-5989);
			14599: out = 16'(-7122);
			14600: out = 16'(-1126);
			14601: out = 16'(4317);
			14602: out = 16'(7641);
			14603: out = 16'(4419);
			14604: out = 16'(687);
			14605: out = 16'(-3525);
			14606: out = 16'(-1234);
			14607: out = 16'(-764);
			14608: out = 16'(1217);
			14609: out = 16'(-811);
			14610: out = 16'(-120);
			14611: out = 16'(-423);
			14612: out = 16'(-268);
			14613: out = 16'(-1385);
			14614: out = 16'(-2701);
			14615: out = 16'(52);
			14616: out = 16'(-1026);
			14617: out = 16'(-6304);
			14618: out = 16'(-3342);
			14619: out = 16'(-1187);
			14620: out = 16'(3349);
			14621: out = 16'(935);
			14622: out = 16'(437);
			14623: out = 16'(2910);
			14624: out = 16'(3050);
			14625: out = 16'(2133);
			14626: out = 16'(-3098);
			14627: out = 16'(-3409);
			14628: out = 16'(-1987);
			14629: out = 16'(-1061);
			14630: out = 16'(2106);
			14631: out = 16'(4733);
			14632: out = 16'(19);
			14633: out = 16'(-4319);
			14634: out = 16'(-9367);
			14635: out = 16'(-1013);
			14636: out = 16'(4110);
			14637: out = 16'(5283);
			14638: out = 16'(5824);
			14639: out = 16'(3554);
			14640: out = 16'(3855);
			14641: out = 16'(-5149);
			14642: out = 16'(-8867);
			14643: out = 16'(-3270);
			14644: out = 16'(3532);
			14645: out = 16'(8374);
			14646: out = 16'(4463);
			14647: out = 16'(-2018);
			14648: out = 16'(-10242);
			14649: out = 16'(-5235);
			14650: out = 16'(-1945);
			14651: out = 16'(3731);
			14652: out = 16'(323);
			14653: out = 16'(75);
			14654: out = 16'(-392);
			14655: out = 16'(-246);
			14656: out = 16'(-476);
			14657: out = 16'(-1488);
			14658: out = 16'(404);
			14659: out = 16'(1037);
			14660: out = 16'(1348);
			14661: out = 16'(-2227);
			14662: out = 16'(-4661);
			14663: out = 16'(-3495);
			14664: out = 16'(-504);
			14665: out = 16'(2626);
			14666: out = 16'(1077);
			14667: out = 16'(107);
			14668: out = 16'(-1154);
			14669: out = 16'(-354);
			14670: out = 16'(313);
			14671: out = 16'(21);
			14672: out = 16'(3584);
			14673: out = 16'(2889);
			14674: out = 16'(7);
			14675: out = 16'(-4128);
			14676: out = 16'(-4791);
			14677: out = 16'(-1335);
			14678: out = 16'(2833);
			14679: out = 16'(5674);
			14680: out = 16'(7781);
			14681: out = 16'(2843);
			14682: out = 16'(-2376);
			14683: out = 16'(-6493);
			14684: out = 16'(-3906);
			14685: out = 16'(797);
			14686: out = 16'(2783);
			14687: out = 16'(560);
			14688: out = 16'(-4969);
			14689: out = 16'(-5310);
			14690: out = 16'(-3317);
			14691: out = 16'(2794);
			14692: out = 16'(4879);
			14693: out = 16'(5138);
			14694: out = 16'(-208);
			14695: out = 16'(794);
			14696: out = 16'(1181);
			14697: out = 16'(2999);
			14698: out = 16'(4630);
			14699: out = 16'(5076);
			14700: out = 16'(-934);
			14701: out = 16'(-3640);
			14702: out = 16'(-5543);
			14703: out = 16'(2032);
			14704: out = 16'(3882);
			14705: out = 16'(4647);
			14706: out = 16'(825);
			14707: out = 16'(-889);
			14708: out = 16'(-1412);
			14709: out = 16'(-3279);
			14710: out = 16'(-3039);
			14711: out = 16'(-1400);
			14712: out = 16'(2726);
			14713: out = 16'(5516);
			14714: out = 16'(5231);
			14715: out = 16'(5377);
			14716: out = 16'(2990);
			14717: out = 16'(-3032);
			14718: out = 16'(-7062);
			14719: out = 16'(-8506);
			14720: out = 16'(4370);
			14721: out = 16'(6176);
			14722: out = 16'(5832);
			14723: out = 16'(-5192);
			14724: out = 16'(-6576);
			14725: out = 16'(-3100);
			14726: out = 16'(-1429);
			14727: out = 16'(-1009);
			14728: out = 16'(-5269);
			14729: out = 16'(501);
			14730: out = 16'(2718);
			14731: out = 16'(5107);
			14732: out = 16'(1991);
			14733: out = 16'(48);
			14734: out = 16'(-2760);
			14735: out = 16'(650);
			14736: out = 16'(2957);
			14737: out = 16'(2112);
			14738: out = 16'(-1297);
			14739: out = 16'(-4910);
			14740: out = 16'(-39);
			14741: out = 16'(2667);
			14742: out = 16'(5722);
			14743: out = 16'(-279);
			14744: out = 16'(-2876);
			14745: out = 16'(-4828);
			14746: out = 16'(-1727);
			14747: out = 16'(62);
			14748: out = 16'(-517);
			14749: out = 16'(2228);
			14750: out = 16'(1761);
			14751: out = 16'(-2398);
			14752: out = 16'(-4798);
			14753: out = 16'(-5126);
			14754: out = 16'(590);
			14755: out = 16'(3066);
			14756: out = 16'(4843);
			14757: out = 16'(2072);
			14758: out = 16'(891);
			14759: out = 16'(-949);
			14760: out = 16'(-2062);
			14761: out = 16'(-4010);
			14762: out = 16'(-5883);
			14763: out = 16'(-1394);
			14764: out = 16'(1706);
			14765: out = 16'(5039);
			14766: out = 16'(1262);
			14767: out = 16'(-377);
			14768: out = 16'(-369);
			14769: out = 16'(1058);
			14770: out = 16'(2071);
			14771: out = 16'(1846);
			14772: out = 16'(584);
			14773: out = 16'(-592);
			14774: out = 16'(849);
			14775: out = 16'(1224);
			14776: out = 16'(1673);
			14777: out = 16'(-1219);
			14778: out = 16'(-2533);
			14779: out = 16'(-3775);
			14780: out = 16'(-97);
			14781: out = 16'(489);
			14782: out = 16'(-225);
			14783: out = 16'(-1147);
			14784: out = 16'(-562);
			14785: out = 16'(3281);
			14786: out = 16'(558);
			14787: out = 16'(-1097);
			14788: out = 16'(-6395);
			14789: out = 16'(-258);
			14790: out = 16'(3479);
			14791: out = 16'(3894);
			14792: out = 16'(517);
			14793: out = 16'(-3487);
			14794: out = 16'(-5452);
			14795: out = 16'(-5134);
			14796: out = 16'(-2749);
			14797: out = 16'(2043);
			14798: out = 16'(3149);
			14799: out = 16'(1659);
			14800: out = 16'(748);
			14801: out = 16'(-1012);
			14802: out = 16'(-2346);
			14803: out = 16'(-1102);
			14804: out = 16'(1218);
			14805: out = 16'(4990);
			14806: out = 16'(4222);
			14807: out = 16'(2981);
			14808: out = 16'(-1734);
			14809: out = 16'(1200);
			14810: out = 16'(2817);
			14811: out = 16'(1990);
			14812: out = 16'(-473);
			14813: out = 16'(-3131);
			14814: out = 16'(-3554);
			14815: out = 16'(-3747);
			14816: out = 16'(-3384);
			14817: out = 16'(2054);
			14818: out = 16'(2141);
			14819: out = 16'(-430);
			14820: out = 16'(-1668);
			14821: out = 16'(-3909);
			14822: out = 16'(-7099);
			14823: out = 16'(-2117);
			14824: out = 16'(2816);
			14825: out = 16'(11256);
			14826: out = 16'(2547);
			14827: out = 16'(-4640);
			14828: out = 16'(-10165);
			14829: out = 16'(-4723);
			14830: out = 16'(3343);
			14831: out = 16'(6367);
			14832: out = 16'(6867);
			14833: out = 16'(2360);
			14834: out = 16'(1724);
			14835: out = 16'(-4328);
			14836: out = 16'(-7698);
			14837: out = 16'(-12235);
			14838: out = 16'(-5235);
			14839: out = 16'(7670);
			14840: out = 16'(8964);
			14841: out = 16'(6525);
			14842: out = 16'(-2763);
			14843: out = 16'(-4599);
			14844: out = 16'(-4256);
			14845: out = 16'(4340);
			14846: out = 16'(4880);
			14847: out = 16'(5515);
			14848: out = 16'(-166);
			14849: out = 16'(659);
			14850: out = 16'(293);
			14851: out = 16'(24);
			14852: out = 16'(-1148);
			14853: out = 16'(-1320);
			14854: out = 16'(-4539);
			14855: out = 16'(-2629);
			14856: out = 16'(1079);
			14857: out = 16'(1022);
			14858: out = 16'(1020);
			14859: out = 16'(834);
			14860: out = 16'(-2335);
			14861: out = 16'(-2689);
			14862: out = 16'(1385);
			14863: out = 16'(1621);
			14864: out = 16'(1264);
			14865: out = 16'(-5964);
			14866: out = 16'(-1682);
			14867: out = 16'(1720);
			14868: out = 16'(2022);
			14869: out = 16'(1221);
			14870: out = 16'(-584);
			14871: out = 16'(-835);
			14872: out = 16'(-2248);
			14873: out = 16'(-3118);
			14874: out = 16'(1062);
			14875: out = 16'(3769);
			14876: out = 16'(5909);
			14877: out = 16'(3140);
			14878: out = 16'(893);
			14879: out = 16'(-1336);
			14880: out = 16'(-166);
			14881: out = 16'(1423);
			14882: out = 16'(2738);
			14883: out = 16'(3133);
			14884: out = 16'(1907);
			14885: out = 16'(-2100);
			14886: out = 16'(-4502);
			14887: out = 16'(-5609);
			14888: out = 16'(-1864);
			14889: out = 16'(257);
			14890: out = 16'(2307);
			14891: out = 16'(1053);
			14892: out = 16'(707);
			14893: out = 16'(-545);
			14894: out = 16'(971);
			14895: out = 16'(747);
			14896: out = 16'(887);
			14897: out = 16'(-3379);
			14898: out = 16'(-3695);
			14899: out = 16'(897);
			14900: out = 16'(2732);
			14901: out = 16'(3689);
			14902: out = 16'(-255);
			14903: out = 16'(-491);
			14904: out = 16'(-1606);
			14905: out = 16'(1300);
			14906: out = 16'(429);
			14907: out = 16'(834);
			14908: out = 16'(-4836);
			14909: out = 16'(-800);
			14910: out = 16'(4056);
			14911: out = 16'(4461);
			14912: out = 16'(-1294);
			14913: out = 16'(-12413);
			14914: out = 16'(-7440);
			14915: out = 16'(-1573);
			14916: out = 16'(8938);
			14917: out = 16'(7773);
			14918: out = 16'(6415);
			14919: out = 16'(1896);
			14920: out = 16'(575);
			14921: out = 16'(-696);
			14922: out = 16'(-102);
			14923: out = 16'(795);
			14924: out = 16'(1483);
			14925: out = 16'(-4288);
			14926: out = 16'(-5368);
			14927: out = 16'(-5573);
			14928: out = 16'(73);
			14929: out = 16'(1022);
			14930: out = 16'(-212);
			14931: out = 16'(17);
			14932: out = 16'(367);
			14933: out = 16'(3547);
			14934: out = 16'(130);
			14935: out = 16'(-505);
			14936: out = 16'(-3169);
			14937: out = 16'(2804);
			14938: out = 16'(4812);
			14939: out = 16'(6306);
			14940: out = 16'(-1299);
			14941: out = 16'(-6688);
			14942: out = 16'(-9829);
			14943: out = 16'(-549);
			14944: out = 16'(9164);
			14945: out = 16'(3492);
			14946: out = 16'(-2725);
			14947: out = 16'(-12687);
			14948: out = 16'(-1705);
			14949: out = 16'(3317);
			14950: out = 16'(9782);
			14951: out = 16'(2750);
			14952: out = 16'(-522);
			14953: out = 16'(-3661);
			14954: out = 16'(-5180);
			14955: out = 16'(-4738);
			14956: out = 16'(1059);
			14957: out = 16'(773);
			14958: out = 16'(1455);
			14959: out = 16'(704);
			14960: out = 16'(4305);
			14961: out = 16'(6377);
			14962: out = 16'(269);
			14963: out = 16'(-696);
			14964: out = 16'(-1563);
			14965: out = 16'(1697);
			14966: out = 16'(1291);
			14967: out = 16'(412);
			14968: out = 16'(-5615);
			14969: out = 16'(-7346);
			14970: out = 16'(-6801);
			14971: out = 16'(-1157);
			14972: out = 16'(2473);
			14973: out = 16'(3958);
			14974: out = 16'(1486);
			14975: out = 16'(-725);
			14976: out = 16'(55);
			14977: out = 16'(-495);
			14978: out = 16'(142);
			14979: out = 16'(865);
			14980: out = 16'(1743);
			14981: out = 16'(1725);
			14982: out = 16'(-1891);
			14983: out = 16'(-2583);
			14984: out = 16'(-2123);
			14985: out = 16'(580);
			14986: out = 16'(283);
			14987: out = 16'(-2651);
			14988: out = 16'(1350);
			14989: out = 16'(3323);
			14990: out = 16'(7232);
			14991: out = 16'(-3);
			14992: out = 16'(-2224);
			14993: out = 16'(716);
			14994: out = 16'(3819);
			14995: out = 16'(4710);
			14996: out = 16'(-4949);
			14997: out = 16'(-2808);
			14998: out = 16'(-975);
			14999: out = 16'(2814);
			15000: out = 16'(1488);
			15001: out = 16'(-254);
			15002: out = 16'(570);
			15003: out = 16'(389);
			15004: out = 16'(-151);
			15005: out = 16'(3141);
			15006: out = 16'(3248);
			15007: out = 16'(1576);
			15008: out = 16'(392);
			15009: out = 16'(-1014);
			15010: out = 16'(-2666);
			15011: out = 16'(-2610);
			15012: out = 16'(-2482);
			15013: out = 16'(-1335);
			15014: out = 16'(-2245);
			15015: out = 16'(-1985);
			15016: out = 16'(-367);
			15017: out = 16'(1643);
			15018: out = 16'(2974);
			15019: out = 16'(3864);
			15020: out = 16'(1823);
			15021: out = 16'(-1054);
			15022: out = 16'(-6937);
			15023: out = 16'(-5783);
			15024: out = 16'(546);
			15025: out = 16'(-565);
			15026: out = 16'(721);
			15027: out = 16'(392);
			15028: out = 16'(1321);
			15029: out = 16'(652);
			15030: out = 16'(1398);
			15031: out = 16'(-897);
			15032: out = 16'(-588);
			15033: out = 16'(1477);
			15034: out = 16'(5214);
			15035: out = 16'(6157);
			15036: out = 16'(-2820);
			15037: out = 16'(-4974);
			15038: out = 16'(-5532);
			15039: out = 16'(-3113);
			15040: out = 16'(-693);
			15041: out = 16'(1192);
			15042: out = 16'(5115);
			15043: out = 16'(3476);
			15044: out = 16'(-1878);
			15045: out = 16'(-1317);
			15046: out = 16'(-481);
			15047: out = 16'(3151);
			15048: out = 16'(1326);
			15049: out = 16'(1145);
			15050: out = 16'(2852);
			15051: out = 16'(953);
			15052: out = 16'(-1124);
			15053: out = 16'(-5731);
			15054: out = 16'(-3133);
			15055: out = 16'(167);
			15056: out = 16'(-329);
			15057: out = 16'(39);
			15058: out = 16'(-480);
			15059: out = 16'(1075);
			15060: out = 16'(-1014);
			15061: out = 16'(-4826);
			15062: out = 16'(-381);
			15063: out = 16'(3432);
			15064: out = 16'(10336);
			15065: out = 16'(2086);
			15066: out = 16'(-3303);
			15067: out = 16'(-13599);
			15068: out = 16'(-4497);
			15069: out = 16'(1838);
			15070: out = 16'(10274);
			15071: out = 16'(2482);
			15072: out = 16'(-3961);
			15073: out = 16'(-14241);
			15074: out = 16'(-1882);
			15075: out = 16'(12508);
			15076: out = 16'(10119);
			15077: out = 16'(4035);
			15078: out = 16'(-8768);
			15079: out = 16'(-2252);
			15080: out = 16'(-2044);
			15081: out = 16'(1813);
			15082: out = 16'(-3029);
			15083: out = 16'(-3591);
			15084: out = 16'(-6180);
			15085: out = 16'(-466);
			15086: out = 16'(1387);
			15087: out = 16'(2478);
			15088: out = 16'(-1437);
			15089: out = 16'(-2411);
			15090: out = 16'(3817);
			15091: out = 16'(4556);
			15092: out = 16'(4143);
			15093: out = 16'(-1767);
			15094: out = 16'(-2640);
			15095: out = 16'(-2261);
			15096: out = 16'(-4465);
			15097: out = 16'(-2575);
			15098: out = 16'(584);
			15099: out = 16'(4011);
			15100: out = 16'(3467);
			15101: out = 16'(-1825);
			15102: out = 16'(93);
			15103: out = 16'(838);
			15104: out = 16'(5406);
			15105: out = 16'(1044);
			15106: out = 16'(-1146);
			15107: out = 16'(-6131);
			15108: out = 16'(-297);
			15109: out = 16'(3161);
			15110: out = 16'(2278);
			15111: out = 16'(-1791);
			15112: out = 16'(-5831);
			15113: out = 16'(-3532);
			15114: out = 16'(-494);
			15115: out = 16'(3856);
			15116: out = 16'(6634);
			15117: out = 16'(5606);
			15118: out = 16'(196);
			15119: out = 16'(759);
			15120: out = 16'(-648);
			15121: out = 16'(486);
			15122: out = 16'(-5108);
			15123: out = 16'(-5644);
			15124: out = 16'(-53);
			15125: out = 16'(-228);
			15126: out = 16'(-454);
			15127: out = 16'(-3309);
			15128: out = 16'(-993);
			15129: out = 16'(1268);
			15130: out = 16'(106);
			15131: out = 16'(727);
			15132: out = 16'(862);
			15133: out = 16'(995);
			15134: out = 16'(430);
			15135: out = 16'(-93);
			15136: out = 16'(84);
			15137: out = 16'(538);
			15138: out = 16'(1144);
			15139: out = 16'(455);
			15140: out = 16'(165);
			15141: out = 16'(1028);
			15142: out = 16'(164);
			15143: out = 16'(610);
			15144: out = 16'(1797);
			15145: out = 16'(3273);
			15146: out = 16'(3600);
			15147: out = 16'(3175);
			15148: out = 16'(545);
			15149: out = 16'(-1461);
			15150: out = 16'(168);
			15151: out = 16'(2389);
			15152: out = 16'(4491);
			15153: out = 16'(454);
			15154: out = 16'(-1954);
			15155: out = 16'(-3479);
			15156: out = 16'(-1307);
			15157: out = 16'(711);
			15158: out = 16'(282);
			15159: out = 16'(6227);
			15160: out = 16'(7339);
			15161: out = 16'(6590);
			15162: out = 16'(-2186);
			15163: out = 16'(-8059);
			15164: out = 16'(-7108);
			15165: out = 16'(-3081);
			15166: out = 16'(1761);
			15167: out = 16'(3169);
			15168: out = 16'(2402);
			15169: out = 16'(-200);
			15170: out = 16'(-4979);
			15171: out = 16'(-4204);
			15172: out = 16'(242);
			15173: out = 16'(3921);
			15174: out = 16'(6330);
			15175: out = 16'(6744);
			15176: out = 16'(1570);
			15177: out = 16'(-1619);
			15178: out = 16'(-1571);
			15179: out = 16'(275);
			15180: out = 16'(843);
			15181: out = 16'(-5024);
			15182: out = 16'(-5367);
			15183: out = 16'(-5493);
			15184: out = 16'(-351);
			15185: out = 16'(613);
			15186: out = 16'(2149);
			15187: out = 16'(466);
			15188: out = 16'(2560);
			15189: out = 16'(4267);
			15190: out = 16'(608);
			15191: out = 16'(-3126);
			15192: out = 16'(-7134);
			15193: out = 16'(-6304);
			15194: out = 16'(-3862);
			15195: out = 16'(1167);
			15196: out = 16'(848);
			15197: out = 16'(617);
			15198: out = 16'(-1533);
			15199: out = 16'(-747);
			15200: out = 16'(-166);
			15201: out = 16'(947);
			15202: out = 16'(886);
			15203: out = 16'(860);
			15204: out = 16'(-74);
			15205: out = 16'(-557);
			15206: out = 16'(-1642);
			15207: out = 16'(650);
			15208: out = 16'(-1026);
			15209: out = 16'(-3634);
			15210: out = 16'(-4523);
			15211: out = 16'(-2306);
			15212: out = 16'(3485);
			15213: out = 16'(3457);
			15214: out = 16'(2654);
			15215: out = 16'(-4081);
			15216: out = 16'(496);
			15217: out = 16'(2227);
			15218: out = 16'(4102);
			15219: out = 16'(656);
			15220: out = 16'(-2351);
			15221: out = 16'(-7706);
			15222: out = 16'(-6243);
			15223: out = 16'(-3631);
			15224: out = 16'(4235);
			15225: out = 16'(3014);
			15226: out = 16'(-74);
			15227: out = 16'(-1259);
			15228: out = 16'(1569);
			15229: out = 16'(6923);
			15230: out = 16'(7909);
			15231: out = 16'(5444);
			15232: out = 16'(-1900);
			15233: out = 16'(-5347);
			15234: out = 16'(-5212);
			15235: out = 16'(5199);
			15236: out = 16'(3121);
			15237: out = 16'(1530);
			15238: out = 16'(-8184);
			15239: out = 16'(-3420);
			15240: out = 16'(1816);
			15241: out = 16'(4880);
			15242: out = 16'(5465);
			15243: out = 16'(4121);
			15244: out = 16'(5718);
			15245: out = 16'(2695);
			15246: out = 16'(-1055);
			15247: out = 16'(-2629);
			15248: out = 16'(-1022);
			15249: out = 16'(3793);
			15250: out = 16'(960);
			15251: out = 16'(-860);
			15252: out = 16'(-4104);
			15253: out = 16'(-1149);
			15254: out = 16'(618);
			15255: out = 16'(58);
			15256: out = 16'(83);
			15257: out = 16'(-145);
			15258: out = 16'(4534);
			15259: out = 16'(2114);
			15260: out = 16'(55);
			15261: out = 16'(-4800);
			15262: out = 16'(-3134);
			15263: out = 16'(-663);
			15264: out = 16'(518);
			15265: out = 16'(-2788);
			15266: out = 16'(-8442);
			15267: out = 16'(-6712);
			15268: out = 16'(-2284);
			15269: out = 16'(6003);
			15270: out = 16'(7795);
			15271: out = 16'(7697);
			15272: out = 16'(2224);
			15273: out = 16'(948);
			15274: out = 16'(-1000);
			15275: out = 16'(-124);
			15276: out = 16'(-892);
			15277: out = 16'(-458);
			15278: out = 16'(-47);
			15279: out = 16'(472);
			15280: out = 16'(-359);
			15281: out = 16'(-5122);
			15282: out = 16'(-5677);
			15283: out = 16'(-2880);
			15284: out = 16'(-750);
			15285: out = 16'(3641);
			15286: out = 16'(6731);
			15287: out = 16'(5651);
			15288: out = 16'(1809);
			15289: out = 16'(-2462);
			15290: out = 16'(-7708);
			15291: out = 16'(-9374);
			15292: out = 16'(-9819);
			15293: out = 16'(47);
			15294: out = 16'(5830);
			15295: out = 16'(13);
			15296: out = 16'(-3861);
			15297: out = 16'(-7222);
			15298: out = 16'(6555);
			15299: out = 16'(7673);
			15300: out = 16'(7738);
			15301: out = 16'(934);
			15302: out = 16'(-955);
			15303: out = 16'(-1572);
			15304: out = 16'(-2484);
			15305: out = 16'(-1880);
			15306: out = 16'(4);
			15307: out = 16'(-1116);
			15308: out = 16'(-1320);
			15309: out = 16'(-249);
			15310: out = 16'(224);
			15311: out = 16'(1764);
			15312: out = 16'(3267);
			15313: out = 16'(5500);
			15314: out = 16'(5850);
			15315: out = 16'(4808);
			15316: out = 16'(1625);
			15317: out = 16'(-1427);
			15318: out = 16'(-6680);
			15319: out = 16'(-5547);
			15320: out = 16'(-2248);
			15321: out = 16'(1066);
			15322: out = 16'(162);
			15323: out = 16'(-3997);
			15324: out = 16'(-5272);
			15325: out = 16'(-3986);
			15326: out = 16'(2384);
			15327: out = 16'(2346);
			15328: out = 16'(2482);
			15329: out = 16'(-534);
			15330: out = 16'(-4016);
			15331: out = 16'(-6786);
			15332: out = 16'(1197);
			15333: out = 16'(-200);
			15334: out = 16'(-145);
			15335: out = 16'(-11381);
			15336: out = 16'(-5571);
			15337: out = 16'(2020);
			15338: out = 16'(9065);
			15339: out = 16'(6712);
			15340: out = 16'(132);
			15341: out = 16'(-5255);
			15342: out = 16'(-3077);
			15343: out = 16'(8482);
			15344: out = 16'(7337);
			15345: out = 16'(6765);
			15346: out = 16'(-1356);
			15347: out = 16'(1077);
			15348: out = 16'(104);
			15349: out = 16'(1493);
			15350: out = 16'(-2872);
			15351: out = 16'(-4711);
			15352: out = 16'(-6294);
			15353: out = 16'(-1243);
			15354: out = 16'(3575);
			15355: out = 16'(6140);
			15356: out = 16'(4534);
			15357: out = 16'(1275);
			15358: out = 16'(-2751);
			15359: out = 16'(-2191);
			15360: out = 16'(2240);
			15361: out = 16'(1512);
			15362: out = 16'(1289);
			15363: out = 16'(-787);
			15364: out = 16'(-2485);
			15365: out = 16'(-4411);
			15366: out = 16'(-5699);
			15367: out = 16'(-1992);
			15368: out = 16'(2178);
			15369: out = 16'(3116);
			15370: out = 16'(4221);
			15371: out = 16'(3068);
			15372: out = 16'(3352);
			15373: out = 16'(-83);
			15374: out = 16'(-2834);
			15375: out = 16'(-4757);
			15376: out = 16'(-2629);
			15377: out = 16'(1083);
			15378: out = 16'(194);
			15379: out = 16'(-2327);
			15380: out = 16'(-8239);
			15381: out = 16'(-3333);
			15382: out = 16'(1322);
			15383: out = 16'(8236);
			15384: out = 16'(7516);
			15385: out = 16'(5840);
			15386: out = 16'(-325);
			15387: out = 16'(-231);
			15388: out = 16'(-330);
			15389: out = 16'(1749);
			15390: out = 16'(512);
			15391: out = 16'(-950);
			15392: out = 16'(-8418);
			15393: out = 16'(-8592);
			15394: out = 16'(-6208);
			15395: out = 16'(2749);
			15396: out = 16'(4194);
			15397: out = 16'(301);
			15398: out = 16'(476);
			15399: out = 16'(-773);
			15400: out = 16'(447);
			15401: out = 16'(-704);
			15402: out = 16'(99);
			15403: out = 16'(-938);
			15404: out = 16'(2232);
			15405: out = 16'(1766);
			15406: out = 16'(-1621);
			15407: out = 16'(-7049);
			15408: out = 16'(-9396);
			15409: out = 16'(-367);
			15410: out = 16'(3646);
			15411: out = 16'(5951);
			15412: out = 16'(8995);
			15413: out = 16'(5691);
			15414: out = 16'(289);
			15415: out = 16'(-4510);
			15416: out = 16'(-4505);
			15417: out = 16'(353);
			15418: out = 16'(276);
			15419: out = 16'(603);
			15420: out = 16'(796);
			15421: out = 16'(-3686);
			15422: out = 16'(-5212);
			15423: out = 16'(-1525);
			15424: out = 16'(4719);
			15425: out = 16'(8723);
			15426: out = 16'(-74);
			15427: out = 16'(-1989);
			15428: out = 16'(-4827);
			15429: out = 16'(3600);
			15430: out = 16'(2146);
			15431: out = 16'(350);
			15432: out = 16'(-6893);
			15433: out = 16'(-5294);
			15434: out = 16'(1429);
			15435: out = 16'(421);
			15436: out = 16'(-241);
			15437: out = 16'(-5110);
			15438: out = 16'(577);
			15439: out = 16'(2116);
			15440: out = 16'(2279);
			15441: out = 16'(-160);
			15442: out = 16'(-1712);
			15443: out = 16'(-4667);
			15444: out = 16'(-1459);
			15445: out = 16'(1824);
			15446: out = 16'(7967);
			15447: out = 16'(5710);
			15448: out = 16'(1896);
			15449: out = 16'(-7581);
			15450: out = 16'(-7785);
			15451: out = 16'(-3644);
			15452: out = 16'(4441);
			15453: out = 16'(6182);
			15454: out = 16'(2382);
			15455: out = 16'(967);
			15456: out = 16'(1047);
			15457: out = 16'(7021);
			15458: out = 16'(3003);
			15459: out = 16'(694);
			15460: out = 16'(-3729);
			15461: out = 16'(-3031);
			15462: out = 16'(-2153);
			15463: out = 16'(431);
			15464: out = 16'(575);
			15465: out = 16'(545);
			15466: out = 16'(592);
			15467: out = 16'(-336);
			15468: out = 16'(-1568);
			15469: out = 16'(597);
			15470: out = 16'(854);
			15471: out = 16'(850);
			15472: out = 16'(754);
			15473: out = 16'(1332);
			15474: out = 16'(2779);
			15475: out = 16'(-175);
			15476: out = 16'(-3263);
			15477: out = 16'(-8033);
			15478: out = 16'(-5492);
			15479: out = 16'(-1201);
			15480: out = 16'(6844);
			15481: out = 16'(7932);
			15482: out = 16'(6669);
			15483: out = 16'(-2887);
			15484: out = 16'(-4909);
			15485: out = 16'(-5393);
			15486: out = 16'(4501);
			15487: out = 16'(3771);
			15488: out = 16'(187);
			15489: out = 16'(-5499);
			15490: out = 16'(-5520);
			15491: out = 16'(403);
			15492: out = 16'(-985);
			15493: out = 16'(399);
			15494: out = 16'(240);
			15495: out = 16'(3119);
			15496: out = 16'(3767);
			15497: out = 16'(4871);
			15498: out = 16'(2065);
			15499: out = 16'(108);
			15500: out = 16'(-3813);
			15501: out = 16'(-1240);
			15502: out = 16'(853);
			15503: out = 16'(778);
			15504: out = 16'(-2864);
			15505: out = 16'(-7275);
			15506: out = 16'(-3101);
			15507: out = 16'(-1384);
			15508: out = 16'(154);
			15509: out = 16'(3144);
			15510: out = 16'(2801);
			15511: out = 16'(-642);
			15512: out = 16'(-2560);
			15513: out = 16'(-2458);
			15514: out = 16'(3416);
			15515: out = 16'(664);
			15516: out = 16'(-163);
			15517: out = 16'(-1601);
			15518: out = 16'(1137);
			15519: out = 16'(2912);
			15520: out = 16'(882);
			15521: out = 16'(803);
			15522: out = 16'(745);
			15523: out = 16'(4239);
			15524: out = 16'(4152);
			15525: out = 16'(3222);
			15526: out = 16'(-587);
			15527: out = 16'(-3690);
			15528: out = 16'(-7374);
			15529: out = 16'(-1984);
			15530: out = 16'(-236);
			15531: out = 16'(-470);
			15532: out = 16'(-2568);
			15533: out = 16'(-3312);
			15534: out = 16'(-1245);
			15535: out = 16'(-615);
			15536: out = 16'(472);
			15537: out = 16'(1848);
			15538: out = 16'(2002);
			15539: out = 16'(1828);
			15540: out = 16'(713);
			15541: out = 16'(195);
			15542: out = 16'(-479);
			15543: out = 16'(2713);
			15544: out = 16'(1468);
			15545: out = 16'(-568);
			15546: out = 16'(-3211);
			15547: out = 16'(-1463);
			15548: out = 16'(4141);
			15549: out = 16'(2159);
			15550: out = 16'(1479);
			15551: out = 16'(774);
			15552: out = 16'(-99);
			15553: out = 16'(-1258);
			15554: out = 16'(-5055);
			15555: out = 16'(196);
			15556: out = 16'(4149);
			15557: out = 16'(2596);
			15558: out = 16'(294);
			15559: out = 16'(-3231);
			15560: out = 16'(-1209);
			15561: out = 16'(-1270);
			15562: out = 16'(378);
			15563: out = 16'(-810);
			15564: out = 16'(182);
			15565: out = 16'(-442);
			15566: out = 16'(6061);
			15567: out = 16'(5000);
			15568: out = 16'(-696);
			15569: out = 16'(-5125);
			15570: out = 16'(-5003);
			15571: out = 16'(6099);
			15572: out = 16'(2059);
			15573: out = 16'(-690);
			15574: out = 16'(-8096);
			15575: out = 16'(-3195);
			15576: out = 16'(1419);
			15577: out = 16'(-2610);
			15578: out = 16'(-1054);
			15579: out = 16'(302);
			15580: out = 16'(5117);
			15581: out = 16'(2819);
			15582: out = 16'(-3055);
			15583: out = 16'(3663);
			15584: out = 16'(4763);
			15585: out = 16'(5522);
			15586: out = 16'(-1298);
			15587: out = 16'(-4484);
			15588: out = 16'(-4640);
			15589: out = 16'(-1976);
			15590: out = 16'(939);
			15591: out = 16'(3473);
			15592: out = 16'(1618);
			15593: out = 16'(-516);
			15594: out = 16'(1987);
			15595: out = 16'(963);
			15596: out = 16'(511);
			15597: out = 16'(-4421);
			15598: out = 16'(-3840);
			15599: out = 16'(-2430);
			15600: out = 16'(-248);
			15601: out = 16'(-2235);
			15602: out = 16'(-7210);
			15603: out = 16'(-6647);
			15604: out = 16'(-4737);
			15605: out = 16'(1918);
			15606: out = 16'(559);
			15607: out = 16'(1416);
			15608: out = 16'(-411);
			15609: out = 16'(4771);
			15610: out = 16'(5925);
			15611: out = 16'(2613);
			15612: out = 16'(-2201);
			15613: out = 16'(-6023);
			15614: out = 16'(-6732);
			15615: out = 16'(-3241);
			15616: out = 16'(1823);
			15617: out = 16'(4247);
			15618: out = 16'(4558);
			15619: out = 16'(2756);
			15620: out = 16'(2374);
			15621: out = 16'(1607);
			15622: out = 16'(537);
			15623: out = 16'(3137);
			15624: out = 16'(3218);
			15625: out = 16'(2088);
			15626: out = 16'(-4534);
			15627: out = 16'(-7333);
			15628: out = 16'(139);
			15629: out = 16'(1910);
			15630: out = 16'(3744);
			15631: out = 16'(-2514);
			15632: out = 16'(-1216);
			15633: out = 16'(-71);
			15634: out = 16'(3476);
			15635: out = 16'(3379);
			15636: out = 16'(2618);
			15637: out = 16'(180);
			15638: out = 16'(-1313);
			15639: out = 16'(-2608);
			15640: out = 16'(-647);
			15641: out = 16'(148);
			15642: out = 16'(669);
			15643: out = 16'(-926);
			15644: out = 16'(-632);
			15645: out = 16'(3791);
			15646: out = 16'(2466);
			15647: out = 16'(614);
			15648: out = 16'(-5667);
			15649: out = 16'(-4901);
			15650: out = 16'(-2464);
			15651: out = 16'(4632);
			15652: out = 16'(6147);
			15653: out = 16'(5801);
			15654: out = 16'(-510);
			15655: out = 16'(-1390);
			15656: out = 16'(746);
			15657: out = 16'(275);
			15658: out = 16'(600);
			15659: out = 16'(-1143);
			15660: out = 16'(2164);
			15661: out = 16'(963);
			15662: out = 16'(-3797);
			15663: out = 16'(-5417);
			15664: out = 16'(-5105);
			15665: out = 16'(-222);
			15666: out = 16'(-318);
			15667: out = 16'(-366);
			15668: out = 16'(920);
			15669: out = 16'(256);
			15670: out = 16'(-572);
			15671: out = 16'(-6345);
			15672: out = 16'(-5665);
			15673: out = 16'(-2949);
			15674: out = 16'(-662);
			15675: out = 16'(1270);
			15676: out = 16'(3200);
			15677: out = 16'(-418);
			15678: out = 16'(-1024);
			15679: out = 16'(-346);
			15680: out = 16'(4720);
			15681: out = 16'(5756);
			15682: out = 16'(748);
			15683: out = 16'(-1598);
			15684: out = 16'(-3958);
			15685: out = 16'(-2181);
			15686: out = 16'(-1599);
			15687: out = 16'(0);
			15688: out = 16'(-2617);
			15689: out = 16'(-1102);
			15690: out = 16'(-80);
			15691: out = 16'(2816);
			15692: out = 16'(2547);
			15693: out = 16'(2097);
			15694: out = 16'(1706);
			15695: out = 16'(2973);
			15696: out = 16'(4578);
			15697: out = 16'(4739);
			15698: out = 16'(3554);
			15699: out = 16'(1766);
			15700: out = 16'(-1393);
			15701: out = 16'(-2968);
			15702: out = 16'(-2840);
			15703: out = 16'(-637);
			15704: out = 16'(969);
			15705: out = 16'(1868);
			15706: out = 16'(-2137);
			15707: out = 16'(-6068);
			15708: out = 16'(83);
			15709: out = 16'(1801);
			15710: out = 16'(3836);
			15711: out = 16'(-1084);
			15712: out = 16'(-789);
			15713: out = 16'(896);
			15714: out = 16'(531);
			15715: out = 16'(-359);
			15716: out = 16'(-2887);
			15717: out = 16'(624);
			15718: out = 16'(2120);
			15719: out = 16'(2694);
			15720: out = 16'(823);
			15721: out = 16'(-1060);
			15722: out = 16'(-3566);
			15723: out = 16'(-3776);
			15724: out = 16'(-3081);
			15725: out = 16'(1656);
			15726: out = 16'(1203);
			15727: out = 16'(205);
			15728: out = 16'(-5323);
			15729: out = 16'(-3341);
			15730: out = 16'(1194);
			15731: out = 16'(719);
			15732: out = 16'(1079);
			15733: out = 16'(894);
			15734: out = 16'(773);
			15735: out = 16'(-286);
			15736: out = 16'(-3960);
			15737: out = 16'(1223);
			15738: out = 16'(2552);
			15739: out = 16'(928);
			15740: out = 16'(-4104);
			15741: out = 16'(-5910);
			15742: out = 16'(2619);
			15743: out = 16'(5764);
			15744: out = 16'(7433);
			15745: out = 16'(-2550);
			15746: out = 16'(-6086);
			15747: out = 16'(-8904);
			15748: out = 16'(548);
			15749: out = 16'(4255);
			15750: out = 16'(7545);
			15751: out = 16'(2094);
			15752: out = 16'(122);
			15753: out = 16'(-1564);
			15754: out = 16'(345);
			15755: out = 16'(1675);
			15756: out = 16'(4951);
			15757: out = 16'(-184);
			15758: out = 16'(-3095);
			15759: out = 16'(-3645);
			15760: out = 16'(507);
			15761: out = 16'(3844);
			15762: out = 16'(-1563);
			15763: out = 16'(-1726);
			15764: out = 16'(-2385);
			15765: out = 16'(4315);
			15766: out = 16'(2903);
			15767: out = 16'(270);
			15768: out = 16'(-334);
			15769: out = 16'(-409);
			15770: out = 16'(-222);
			15771: out = 16'(418);
			15772: out = 16'(484);
			15773: out = 16'(951);
			15774: out = 16'(-969);
			15775: out = 16'(-1494);
			15776: out = 16'(-1771);
			15777: out = 16'(1293);
			15778: out = 16'(2672);
			15779: out = 16'(2006);
			15780: out = 16'(-2247);
			15781: out = 16'(-6162);
			15782: out = 16'(-2660);
			15783: out = 16'(-277);
			15784: out = 16'(3411);
			15785: out = 16'(721);
			15786: out = 16'(845);
			15787: out = 16'(-525);
			15788: out = 16'(2594);
			15789: out = 16'(2138);
			15790: out = 16'(2055);
			15791: out = 16'(-4089);
			15792: out = 16'(-4843);
			15793: out = 16'(-440);
			15794: out = 16'(4622);
			15795: out = 16'(5011);
			15796: out = 16'(-10801);
			15797: out = 16'(-6849);
			15798: out = 16'(-2997);
			15799: out = 16'(6973);
			15800: out = 16'(3020);
			15801: out = 16'(-2362);
			15802: out = 16'(-5755);
			15803: out = 16'(-6477);
			15804: out = 16'(-4552);
			15805: out = 16'(2788);
			15806: out = 16'(6638);
			15807: out = 16'(7681);
			15808: out = 16'(2786);
			15809: out = 16'(-1172);
			15810: out = 16'(-3098);
			15811: out = 16'(-3044);
			15812: out = 16'(-1857);
			15813: out = 16'(-2760);
			15814: out = 16'(1805);
			15815: out = 16'(4142);
			15816: out = 16'(4695);
			15817: out = 16'(2643);
			15818: out = 16'(-4);
			15819: out = 16'(-4977);
			15820: out = 16'(-5739);
			15821: out = 16'(-4961);
			15822: out = 16'(1906);
			15823: out = 16'(2826);
			15824: out = 16'(1873);
			15825: out = 16'(-684);
			15826: out = 16'(151);
			15827: out = 16'(4098);
			15828: out = 16'(3590);
			15829: out = 16'(3473);
			15830: out = 16'(2658);
			15831: out = 16'(656);
			15832: out = 16'(-1293);
			15833: out = 16'(-3657);
			15834: out = 16'(-504);
			15835: out = 16'(1462);
			15836: out = 16'(-4432);
			15837: out = 16'(-5549);
			15838: out = 16'(-6219);
			15839: out = 16'(2141);
			15840: out = 16'(3358);
			15841: out = 16'(3742);
			15842: out = 16'(-634);
			15843: out = 16'(-799);
			15844: out = 16'(791);
			15845: out = 16'(563);
			15846: out = 16'(610);
			15847: out = 16'(620);
			15848: out = 16'(-796);
			15849: out = 16'(-1238);
			15850: out = 16'(51);
			15851: out = 16'(998);
			15852: out = 16'(2148);
			15853: out = 16'(1570);
			15854: out = 16'(2034);
			15855: out = 16'(1564);
			15856: out = 16'(2911);
			15857: out = 16'(1041);
			15858: out = 16'(-257);
			15859: out = 16'(-751);
			15860: out = 16'(480);
			15861: out = 16'(1630);
			15862: out = 16'(3354);
			15863: out = 16'(2036);
			15864: out = 16'(-765);
			15865: out = 16'(-825);
			15866: out = 16'(-373);
			15867: out = 16'(-684);
			15868: out = 16'(1878);
			15869: out = 16'(1853);
			15870: out = 16'(774);
			15871: out = 16'(-4311);
			15872: out = 16'(-7278);
			15873: out = 16'(-8309);
			15874: out = 16'(-1890);
			15875: out = 16'(4646);
			15876: out = 16'(5999);
			15877: out = 16'(2317);
			15878: out = 16'(-4684);
			15879: out = 16'(-5836);
			15880: out = 16'(-6543);
			15881: out = 16'(-3735);
			15882: out = 16'(-1525);
			15883: out = 16'(2872);
			15884: out = 16'(8074);
			15885: out = 16'(2300);
			15886: out = 16'(-2109);
			15887: out = 16'(-5412);
			15888: out = 16'(-1748);
			15889: out = 16'(2115);
			15890: out = 16'(2244);
			15891: out = 16'(4306);
			15892: out = 16'(3345);
			15893: out = 16'(-3511);
			15894: out = 16'(-6968);
			15895: out = 16'(-8104);
			15896: out = 16'(2148);
			15897: out = 16'(5639);
			15898: out = 16'(6992);
			15899: out = 16'(2894);
			15900: out = 16'(894);
			15901: out = 16'(-150);
			15902: out = 16'(1220);
			15903: out = 16'(1652);
			15904: out = 16'(571);
			15905: out = 16'(146);
			15906: out = 16'(-1761);
			15907: out = 16'(-5498);
			15908: out = 16'(-6498);
			15909: out = 16'(-5462);
			15910: out = 16'(2680);
			15911: out = 16'(1374);
			15912: out = 16'(-696);
			15913: out = 16'(-3047);
			15914: out = 16'(-777);
			15915: out = 16'(3604);
			15916: out = 16'(803);
			15917: out = 16'(1011);
			15918: out = 16'(-811);
			15919: out = 16'(3550);
			15920: out = 16'(2214);
			15921: out = 16'(257);
			15922: out = 16'(-5998);
			15923: out = 16'(-5508);
			15924: out = 16'(3038);
			15925: out = 16'(5638);
			15926: out = 16'(6380);
			15927: out = 16'(808);
			15928: out = 16'(711);
			15929: out = 16'(158);
			15930: out = 16'(-2538);
			15931: out = 16'(-969);
			15932: out = 16'(690);
			15933: out = 16'(2805);
			15934: out = 16'(-303);
			15935: out = 16'(-4921);
			15936: out = 16'(-3864);
			15937: out = 16'(-398);
			15938: out = 16'(5909);
			15939: out = 16'(4662);
			15940: out = 16'(2947);
			15941: out = 16'(-1781);
			15942: out = 16'(-3558);
			15943: out = 16'(-4228);
			15944: out = 16'(-160);
			15945: out = 16'(-436);
			15946: out = 16'(114);
			15947: out = 16'(-568);
			15948: out = 16'(-192);
			15949: out = 16'(-856);
			15950: out = 16'(-2902);
			15951: out = 16'(-4539);
			15952: out = 16'(-5123);
			15953: out = 16'(-871);
			15954: out = 16'(2725);
			15955: out = 16'(6775);
			15956: out = 16'(869);
			15957: out = 16'(-170);
			15958: out = 16'(715);
			15959: out = 16'(2971);
			15960: out = 16'(2743);
			15961: out = 16'(-1674);
			15962: out = 16'(-407);
			15963: out = 16'(188);
			15964: out = 16'(1861);
			15965: out = 16'(1213);
			15966: out = 16'(640);
			15967: out = 16'(-106);
			15968: out = 16'(-208);
			15969: out = 16'(-38);
			15970: out = 16'(1586);
			15971: out = 16'(927);
			15972: out = 16'(-749);
			15973: out = 16'(-474);
			15974: out = 16'(1202);
			15975: out = 16'(5883);
			15976: out = 16'(-420);
			15977: out = 16'(-2269);
			15978: out = 16'(-5265);
			15979: out = 16'(2147);
			15980: out = 16'(3942);
			15981: out = 16'(1955);
			15982: out = 16'(-4335);
			15983: out = 16'(-8145);
			15984: out = 16'(-5750);
			15985: out = 16'(-2150);
			15986: out = 16'(2153);
			15987: out = 16'(7505);
			15988: out = 16'(4301);
			15989: out = 16'(-1591);
			15990: out = 16'(-5733);
			15991: out = 16'(-4611);
			15992: out = 16'(1745);
			15993: out = 16'(1656);
			15994: out = 16'(4044);
			15995: out = 16'(3980);
			15996: out = 16'(3771);
			15997: out = 16'(317);
			15998: out = 16'(-4434);
			15999: out = 16'(-5055);
			16000: out = 16'(-3556);
			16001: out = 16'(-778);
			16002: out = 16'(1191);
			16003: out = 16'(1773);
			16004: out = 16'(2054);
			16005: out = 16'(519);
			16006: out = 16'(-612);
			16007: out = 16'(-2441);
			16008: out = 16'(-2260);
			16009: out = 16'(-2290);
			16010: out = 16'(6090);
			16011: out = 16'(4901);
			16012: out = 16'(514);
			16013: out = 16'(-3437);
			16014: out = 16'(-2534);
			16015: out = 16'(4114);
			16016: out = 16'(2266);
			16017: out = 16'(429);
			16018: out = 16'(-4547);
			16019: out = 16'(-4649);
			16020: out = 16'(-3452);
			16021: out = 16'(690);
			16022: out = 16'(2232);
			16023: out = 16'(2775);
			16024: out = 16'(3068);
			16025: out = 16'(1546);
			16026: out = 16'(138);
			16027: out = 16'(-9001);
			16028: out = 16'(-7611);
			16029: out = 16'(-2501);
			16030: out = 16'(5246);
			16031: out = 16'(6358);
			16032: out = 16'(2416);
			16033: out = 16'(-3039);
			16034: out = 16'(-4776);
			16035: out = 16'(1366);
			16036: out = 16'(2266);
			16037: out = 16'(4237);
			16038: out = 16'(2358);
			16039: out = 16'(1639);
			16040: out = 16'(-1148);
			16041: out = 16'(-1575);
			16042: out = 16'(-4554);
			16043: out = 16'(-5140);
			16044: out = 16'(-6021);
			16045: out = 16'(-1816);
			16046: out = 16'(2542);
			16047: out = 16'(5253);
			16048: out = 16'(3817);
			16049: out = 16'(-267);
			16050: out = 16'(-104);
			16051: out = 16'(537);
			16052: out = 16'(3014);
			16053: out = 16'(3397);
			16054: out = 16'(2955);
			16055: out = 16'(-176);
			16056: out = 16'(-1457);
			16057: out = 16'(-2423);
			16058: out = 16'(-344);
			16059: out = 16'(1151);
			16060: out = 16'(2992);
			16061: out = 16'(436);
			16062: out = 16'(-88);
			16063: out = 16'(-1394);
			16064: out = 16'(7695);
			16065: out = 16'(7081);
			16066: out = 16'(4653);
			16067: out = 16'(-7153);
			16068: out = 16'(-10506);
			16069: out = 16'(-7265);
			16070: out = 16'(-2222);
			16071: out = 16'(1479);
			16072: out = 16'(-1120);
			16073: out = 16'(2941);
			16074: out = 16'(3270);
			16075: out = 16'(3162);
			16076: out = 16'(580);
			16077: out = 16'(-579);
			16078: out = 16'(-2804);
			16079: out = 16'(352);
			16080: out = 16'(2795);
			16081: out = 16'(3856);
			16082: out = 16'(-728);
			16083: out = 16'(-7343);
			16084: out = 16'(-3123);
			16085: out = 16'(-612);
			16086: out = 16'(3081);
			16087: out = 16'(1047);
			16088: out = 16'(-17);
			16089: out = 16'(-1418);
			16090: out = 16'(-1467);
			16091: out = 16'(-904);
			16092: out = 16'(459);
			16093: out = 16'(1404);
			16094: out = 16'(1946);
			16095: out = 16'(3745);
			16096: out = 16'(749);
			16097: out = 16'(-2034);
			16098: out = 16'(-3552);
			16099: out = 16'(-873);
			16100: out = 16'(3049);
			16101: out = 16'(-264);
			16102: out = 16'(-1581);
			16103: out = 16'(-3725);
			16104: out = 16'(783);
			16105: out = 16'(2234);
			16106: out = 16'(2583);
			16107: out = 16'(1205);
			16108: out = 16'(-161);
			16109: out = 16'(-328);
			16110: out = 16'(-2780);
			16111: out = 16'(-3253);
			16112: out = 16'(-1701);
			16113: out = 16'(567);
			16114: out = 16'(1735);
			16115: out = 16'(822);
			16116: out = 16'(-2615);
			16117: out = 16'(-5613);
			16118: out = 16'(-51);
			16119: out = 16'(3340);
			16120: out = 16'(7539);
			16121: out = 16'(3636);
			16122: out = 16'(3997);
			16123: out = 16'(4003);
			16124: out = 16'(4614);
			16125: out = 16'(1738);
			16126: out = 16'(-4059);
			16127: out = 16'(-4704);
			16128: out = 16'(-3842);
			16129: out = 16'(728);
			16130: out = 16'(1142);
			16131: out = 16'(355);
			16132: out = 16'(-9330);
			16133: out = 16'(-4521);
			16134: out = 16'(1103);
			16135: out = 16'(7740);
			16136: out = 16'(6941);
			16137: out = 16'(3223);
			16138: out = 16'(-441);
			16139: out = 16'(-3563);
			16140: out = 16'(-4778);
			16141: out = 16'(-5824);
			16142: out = 16'(-6234);
			16143: out = 16'(-8089);
			16144: out = 16'(-2061);
			16145: out = 16'(60);
			16146: out = 16'(-266);
			16147: out = 16'(552);
			16148: out = 16'(1969);
			16149: out = 16'(4489);
			16150: out = 16'(4356);
			16151: out = 16'(2950);
			16152: out = 16'(2384);
			16153: out = 16'(-1804);
			16154: out = 16'(-4905);
			16155: out = 16'(-5806);
			16156: out = 16'(-2653);
			16157: out = 16'(1345);
			16158: out = 16'(192);
			16159: out = 16'(-1171);
			16160: out = 16'(-3276);
			16161: out = 16'(-928);
			16162: out = 16'(2552);
			16163: out = 16'(7203);
			16164: out = 16'(7342);
			16165: out = 16'(5284);
			16166: out = 16'(987);
			16167: out = 16'(-4882);
			16168: out = 16'(-7688);
			16169: out = 16'(-2446);
			16170: out = 16'(306);
			16171: out = 16'(3281);
			16172: out = 16'(512);
			16173: out = 16'(2027);
			16174: out = 16'(2556);
			16175: out = 16'(1975);
			16176: out = 16'(739);
			16177: out = 16'(-715);
			16178: out = 16'(-156);
			16179: out = 16'(-216);
			16180: out = 16'(619);
			16181: out = 16'(-4526);
			16182: out = 16'(-4614);
			16183: out = 16'(-204);
			16184: out = 16'(-360);
			16185: out = 16'(-1759);
			16186: out = 16'(-7706);
			16187: out = 16'(-7717);
			16188: out = 16'(-5851);
			16189: out = 16'(3748);
			16190: out = 16'(4481);
			16191: out = 16'(4694);
			16192: out = 16'(169);
			16193: out = 16'(2694);
			16194: out = 16'(5806);
			16195: out = 16'(4059);
			16196: out = 16'(500);
			16197: out = 16'(-6426);
			16198: out = 16'(-1528);
			16199: out = 16'(-1670);
			16200: out = 16'(-712);
			16201: out = 16'(-5589);
			16202: out = 16'(-5650);
			16203: out = 16'(-4611);
			16204: out = 16'(3776);
			16205: out = 16'(8120);
			16206: out = 16'(9084);
			16207: out = 16'(3033);
			16208: out = 16'(-2426);
			16209: out = 16'(-5340);
			16210: out = 16'(-1462);
			16211: out = 16'(3641);
			16212: out = 16'(3659);
			16213: out = 16'(623);
			16214: out = 16'(-5112);
			16215: out = 16'(-3266);
			16216: out = 16'(-2083);
			16217: out = 16'(1273);
			16218: out = 16'(2902);
			16219: out = 16'(4339);
			16220: out = 16'(4523);
			16221: out = 16'(1493);
			16222: out = 16'(-564);
			16223: out = 16'(-251);
			16224: out = 16'(272);
			16225: out = 16'(974);
			16226: out = 16'(852);
			16227: out = 16'(-306);
			16228: out = 16'(-1888);
			16229: out = 16'(-4308);
			16230: out = 16'(-2779);
			16231: out = 16'(607);
			16232: out = 16'(5737);
			16233: out = 16'(8337);
			16234: out = 16'(8951);
			16235: out = 16'(5436);
			16236: out = 16'(2104);
			16237: out = 16'(-2153);
			16238: out = 16'(-137);
			16239: out = 16'(-746);
			16240: out = 16'(-2630);
			16241: out = 16'(-7801);
			16242: out = 16'(-9971);
			16243: out = 16'(-4493);
			16244: out = 16'(-2280);
			16245: out = 16'(994);
			16246: out = 16'(2230);
			16247: out = 16'(2787);
			16248: out = 16'(1495);
			16249: out = 16'(4709);
			16250: out = 16'(3265);
			16251: out = 16'(2444);
			16252: out = 16'(-7512);
			16253: out = 16'(-6877);
			16254: out = 16'(-888);
			16255: out = 16'(40);
			16256: out = 16'(-1431);
			16257: out = 16'(-9488);
			16258: out = 16'(-2675);
			16259: out = 16'(1125);
			16260: out = 16'(3814);
			16261: out = 16'(3378);
			16262: out = 16'(2496);
			16263: out = 16'(869);
			16264: out = 16'(-385);
			16265: out = 16'(-1633);
			16266: out = 16'(-2088);
			16267: out = 16'(-2843);
			16268: out = 16'(-2993);
			16269: out = 16'(506);
			16270: out = 16'(984);
			16271: out = 16'(-57);
			16272: out = 16'(1089);
			16273: out = 16'(953);
			16274: out = 16'(1217);
			16275: out = 16'(150);
			16276: out = 16'(431);
			16277: out = 16'(808);
			16278: out = 16'(3643);
			16279: out = 16'(3636);
			16280: out = 16'(-1203);
			16281: out = 16'(-5047);
			16282: out = 16'(-6900);
			16283: out = 16'(4484);
			16284: out = 16'(4798);
			16285: out = 16'(4862);
			16286: out = 16'(-9022);
			16287: out = 16'(-6998);
			16288: out = 16'(-1320);
			16289: out = 16'(6424);
			16290: out = 16'(6125);
			16291: out = 16'(175);
			16292: out = 16'(541);
			16293: out = 16'(244);
			16294: out = 16'(3210);
			16295: out = 16'(-363);
			16296: out = 16'(-2336);
			16297: out = 16'(-5795);
			16298: out = 16'(-2968);
			16299: out = 16'(-331);
			16300: out = 16'(2755);
			16301: out = 16'(1944);
			16302: out = 16'(1006);
			16303: out = 16'(3683);
			16304: out = 16'(3160);
			16305: out = 16'(2606);
			16306: out = 16'(680);
			16307: out = 16'(478);
			16308: out = 16'(284);
			16309: out = 16'(701);
			16310: out = 16'(-1022);
			16311: out = 16'(-3653);
			16312: out = 16'(-6754);
			16313: out = 16'(-6972);
			16314: out = 16'(-3057);
			16315: out = 16'(-1242);
			16316: out = 16'(780);
			16317: out = 16'(571);
			16318: out = 16'(482);
			16319: out = 16'(174);
			16320: out = 16'(5892);
			16321: out = 16'(2398);
			16322: out = 16'(-767);
			16323: out = 16'(-3228);
			16324: out = 16'(-735);
			16325: out = 16'(3179);
			16326: out = 16'(-1584);
			16327: out = 16'(-3828);
			16328: out = 16'(-6659);
			16329: out = 16'(-685);
			16330: out = 16'(4146);
			16331: out = 16'(10747);
			16332: out = 16'(6725);
			16333: out = 16'(3682);
			16334: out = 16'(-2949);
			16335: out = 16'(549);
			16336: out = 16'(1210);
			16337: out = 16'(48);
			16338: out = 16'(-6605);
			16339: out = 16'(-11446);
			16340: out = 16'(-4686);
			16341: out = 16'(-2065);
			16342: out = 16'(1881);
			16343: out = 16'(3822);
			16344: out = 16'(6561);
			16345: out = 16'(7548);
			16346: out = 16'(1613);
			16347: out = 16'(-824);
			16348: out = 16'(261);
			16349: out = 16'(-2138);
			16350: out = 16'(-3678);
			16351: out = 16'(-9618);
			16352: out = 16'(-2569);
			16353: out = 16'(176);
			16354: out = 16'(1569);
			16355: out = 16'(-3003);
			16356: out = 16'(-5302);
			16357: out = 16'(-5835);
			16358: out = 16'(2012);
			16359: out = 16'(9337);
			16360: out = 16'(10173);
			16361: out = 16'(6376);
			16362: out = 16'(-639);
			16363: out = 16'(-4292);
			16364: out = 16'(-3729);
			16365: out = 16'(2980);
			16366: out = 16'(-2222);
			16367: out = 16'(-1866);
			16368: out = 16'(-2795);
			16369: out = 16'(4976);
			16370: out = 16'(6270);
			16371: out = 16'(1640);
			16372: out = 16'(1110);
			16373: out = 16'(793);
			16374: out = 16'(3721);
			16375: out = 16'(2385);
			16376: out = 16'(1020);
			16377: out = 16'(-3360);
			16378: out = 16'(-3183);
			16379: out = 16'(-2354);
			16380: out = 16'(-357);
			16381: out = 16'(-633);
			16382: out = 16'(-1478);
			16383: out = 16'(-2461);
			16384: out = 16'(-421);
			16385: out = 16'(4046);
			16386: out = 16'(1490);
			16387: out = 16'(-995);
			16388: out = 16'(-7174);
			16389: out = 16'(-2074);
			16390: out = 16'(1981);
			16391: out = 16'(8882);
			16392: out = 16'(4483);
			16393: out = 16'(-156);
			16394: out = 16'(-8570);
			16395: out = 16'(-7478);
			16396: out = 16'(-4362);
			16397: out = 16'(3061);
			16398: out = 16'(2684);
			16399: out = 16'(432);
			16400: out = 16'(-297);
			16401: out = 16'(2662);
			16402: out = 16'(8425);
			16403: out = 16'(2679);
			16404: out = 16'(737);
			16405: out = 16'(-1813);
			16406: out = 16'(-684);
			16407: out = 16'(-618);
			16408: out = 16'(-458);
			16409: out = 16'(-514);
			16410: out = 16'(-1572);
			16411: out = 16'(-7923);
			16412: out = 16'(-5836);
			16413: out = 16'(-3375);
			16414: out = 16'(2764);
			16415: out = 16'(1556);
			16416: out = 16'(52);
			16417: out = 16'(542);
			16418: out = 16'(2883);
			16419: out = 16'(5504);
			16420: out = 16'(1098);
			16421: out = 16'(-3557);
			16422: out = 16'(-10569);
			16423: out = 16'(-8019);
			16424: out = 16'(-5380);
			16425: out = 16'(1725);
			16426: out = 16'(-826);
			16427: out = 16'(-801);
			16428: out = 16'(-3660);
			16429: out = 16'(4539);
			16430: out = 16'(8949);
			16431: out = 16'(9891);
			16432: out = 16'(4425);
			16433: out = 16'(-758);
			16434: out = 16'(101);
			16435: out = 16'(1924);
			16436: out = 16'(4503);
			16437: out = 16'(-2407);
			16438: out = 16'(-6081);
			16439: out = 16'(-10163);
			16440: out = 16'(-1109);
			16441: out = 16'(3092);
			16442: out = 16'(5652);
			16443: out = 16'(6218);
			16444: out = 16'(6058);
			16445: out = 16'(5333);
			16446: out = 16'(2343);
			16447: out = 16'(-490);
			16448: out = 16'(-3548);
			16449: out = 16'(-2603);
			16450: out = 16'(-1336);
			16451: out = 16'(-1612);
			16452: out = 16'(-2434);
			16453: out = 16'(-3423);
			16454: out = 16'(674);
			16455: out = 16'(722);
			16456: out = 16'(744);
			16457: out = 16'(704);
			16458: out = 16'(2273);
			16459: out = 16'(4635);
			16460: out = 16'(1610);
			16461: out = 16'(245);
			16462: out = 16'(-486);
			16463: out = 16'(-1833);
			16464: out = 16'(-3319);
			16465: out = 16'(-5541);
			16466: out = 16'(-4959);
			16467: out = 16'(-3546);
			16468: out = 16'(-425);
			16469: out = 16'(1614);
			16470: out = 16'(3151);
			16471: out = 16'(622);
			16472: out = 16'(1958);
			16473: out = 16'(2929);
			16474: out = 16'(4645);
			16475: out = 16'(1882);
			16476: out = 16'(-2906);
			16477: out = 16'(-586);
			16478: out = 16'(-84);
			16479: out = 16'(1043);
			16480: out = 16'(-1563);
			16481: out = 16'(-3225);
			16482: out = 16'(-5634);
			16483: out = 16'(-1396);
			16484: out = 16'(1243);
			16485: out = 16'(-268);
			16486: out = 16'(1487);
			16487: out = 16'(2171);
			16488: out = 16'(4902);
			16489: out = 16'(1036);
			16490: out = 16'(-2866);
			16491: out = 16'(-2238);
			16492: out = 16'(-1080);
			16493: out = 16'(1235);
			16494: out = 16'(-2799);
			16495: out = 16'(-3282);
			16496: out = 16'(-3220);
			16497: out = 16'(-838);
			16498: out = 16'(317);
			16499: out = 16'(915);
			16500: out = 16'(2821);
			16501: out = 16'(5143);
			16502: out = 16'(8659);
			16503: out = 16'(5129);
			16504: out = 16'(1600);
			16505: out = 16'(1273);
			16506: out = 16'(-422);
			16507: out = 16'(-997);
			16508: out = 16'(-9019);
			16509: out = 16'(-4937);
			16510: out = 16'(277);
			16511: out = 16'(3290);
			16512: out = 16'(1808);
			16513: out = 16'(-1546);
			16514: out = 16'(-929);
			16515: out = 16'(3026);
			16516: out = 16'(10407);
			16517: out = 16'(7075);
			16518: out = 16'(3618);
			16519: out = 16'(-2915);
			16520: out = 16'(-3432);
			16521: out = 16'(-4392);
			16522: out = 16'(-8243);
			16523: out = 16'(-2820);
			16524: out = 16'(1632);
			16525: out = 16'(3555);
			16526: out = 16'(-1331);
			16527: out = 16'(-7000);
			16528: out = 16'(2084);
			16529: out = 16'(4967);
			16530: out = 16'(8895);
			16531: out = 16'(1380);
			16532: out = 16'(1028);
			16533: out = 16'(1161);
			16534: out = 16'(1412);
			16535: out = 16'(-3523);
			16536: out = 16'(-14227);
			16537: out = 16'(-13343);
			16538: out = 16'(-8249);
			16539: out = 16'(8481);
			16540: out = 16'(6662);
			16541: out = 16'(5044);
			16542: out = 16'(-7111);
			16543: out = 16'(-1239);
			16544: out = 16'(3488);
			16545: out = 16'(8822);
			16546: out = 16'(1948);
			16547: out = 16'(-6803);
			16548: out = 16'(-8645);
			16549: out = 16'(-4835);
			16550: out = 16'(3778);
			16551: out = 16'(1141);
			16552: out = 16'(-1927);
			16553: out = 16'(-10797);
			16554: out = 16'(-3357);
			16555: out = 16'(1029);
			16556: out = 16'(6854);
			16557: out = 16'(4630);
			16558: out = 16'(3674);
			16559: out = 16'(3823);
			16560: out = 16'(1439);
			16561: out = 16'(-1345);
			16562: out = 16'(-4143);
			16563: out = 16'(-3288);
			16564: out = 16'(-862);
			16565: out = 16'(-3645);
			16566: out = 16'(-1712);
			16567: out = 16'(67);
			16568: out = 16'(5675);
			16569: out = 16'(5306);
			16570: out = 16'(2519);
			16571: out = 16'(-372);
			16572: out = 16'(-861);
			16573: out = 16'(2155);
			16574: out = 16'(1611);
			16575: out = 16'(948);
			16576: out = 16'(-3906);
			16577: out = 16'(-1406);
			16578: out = 16'(26);
			16579: out = 16'(2952);
			16580: out = 16'(372);
			16581: out = 16'(-2075);
			16582: out = 16'(-5408);
			16583: out = 16'(-4237);
			16584: out = 16'(-1562);
			16585: out = 16'(3747);
			16586: out = 16'(4619);
			16587: out = 16'(3256);
			16588: out = 16'(762);
			16589: out = 16'(-480);
			16590: out = 16'(70);
			16591: out = 16'(-505);
			16592: out = 16'(-119);
			16593: out = 16'(518);
			16594: out = 16'(-81);
			16595: out = 16'(-709);
			16596: out = 16'(-1358);
			16597: out = 16'(-345);
			16598: out = 16'(1235);
			16599: out = 16'(3250);
			16600: out = 16'(4083);
			16601: out = 16'(3958);
			16602: out = 16'(1006);
			16603: out = 16'(27);
			16604: out = 16'(-793);
			16605: out = 16'(-437);
			16606: out = 16'(-2128);
			16607: out = 16'(-4815);
			16608: out = 16'(-3727);
			16609: out = 16'(-2318);
			16610: out = 16'(855);
			16611: out = 16'(332);
			16612: out = 16'(604);
			16613: out = 16'(-747);
			16614: out = 16'(2916);
			16615: out = 16'(4611);
			16616: out = 16'(5301);
			16617: out = 16'(851);
			16618: out = 16'(-3364);
			16619: out = 16'(-2216);
			16620: out = 16'(-2405);
			16621: out = 16'(-1637);
			16622: out = 16'(-9409);
			16623: out = 16'(-7369);
			16624: out = 16'(-2492);
			16625: out = 16'(126);
			16626: out = 16'(923);
			16627: out = 16'(-1496);
			16628: out = 16'(4335);
			16629: out = 16'(5326);
			16630: out = 16'(4611);
			16631: out = 16'(-832);
			16632: out = 16'(-3144);
			16633: out = 16'(1409);
			16634: out = 16'(-185);
			16635: out = 16'(-317);
			16636: out = 16'(-2680);
			16637: out = 16'(1109);
			16638: out = 16'(3935);
			16639: out = 16'(3619);
			16640: out = 16'(2197);
			16641: out = 16'(440);
			16642: out = 16'(2253);
			16643: out = 16'(4719);
			16644: out = 16'(8317);
			16645: out = 16'(309);
			16646: out = 16'(-4145);
			16647: out = 16'(-9234);
			16648: out = 16'(-2580);
			16649: out = 16'(937);
			16650: out = 16'(2528);
			16651: out = 16'(626);
			16652: out = 16'(-161);
			16653: out = 16'(3604);
			16654: out = 16'(3168);
			16655: out = 16'(2722);
			16656: out = 16'(-3547);
			16657: out = 16'(-2959);
			16658: out = 16'(-2356);
			16659: out = 16'(3201);
			16660: out = 16'(1187);
			16661: out = 16'(-1881);
			16662: out = 16'(-6103);
			16663: out = 16'(-4593);
			16664: out = 16'(343);
			16665: out = 16'(1896);
			16666: out = 16'(2334);
			16667: out = 16'(339);
			16668: out = 16'(-1524);
			16669: out = 16'(-1644);
			16670: out = 16'(2870);
			16671: out = 16'(2454);
			16672: out = 16'(2254);
			16673: out = 16'(-543);
			16674: out = 16'(-525);
			16675: out = 16'(-499);
			16676: out = 16'(-386);
			16677: out = 16'(1770);
			16678: out = 16'(4493);
			16679: out = 16'(1691);
			16680: out = 16'(500);
			16681: out = 16'(-2063);
			16682: out = 16'(-258);
			16683: out = 16'(-425);
			16684: out = 16'(1012);
			16685: out = 16'(-3617);
			16686: out = 16'(-4097);
			16687: out = 16'(-2749);
			16688: out = 16'(2193);
			16689: out = 16'(4243);
			16690: out = 16'(2598);
			16691: out = 16'(-1492);
			16692: out = 16'(-5466);
			16693: out = 16'(-6456);
			16694: out = 16'(-3698);
			16695: out = 16'(838);
			16696: out = 16'(97);
			16697: out = 16'(-74);
			16698: out = 16'(-2923);
			16699: out = 16'(809);
			16700: out = 16'(126);
			16701: out = 16'(1190);
			16702: out = 16'(-3891);
			16703: out = 16'(-2426);
			16704: out = 16'(702);
			16705: out = 16'(6846);
			16706: out = 16'(6600);
			16707: out = 16'(-138);
			16708: out = 16'(-5805);
			16709: out = 16'(-7270);
			16710: out = 16'(3318);
			16711: out = 16'(6315);
			16712: out = 16'(7925);
			16713: out = 16'(1285);
			16714: out = 16'(-1742);
			16715: out = 16'(-4911);
			16716: out = 16'(-3547);
			16717: out = 16'(-1838);
			16718: out = 16'(1245);
			16719: out = 16'(1484);
			16720: out = 16'(976);
			16721: out = 16'(-1688);
			16722: out = 16'(-3484);
			16723: out = 16'(-3341);
			16724: out = 16'(2459);
			16725: out = 16'(146);
			16726: out = 16'(123);
			16727: out = 16'(-1831);
			16728: out = 16'(2887);
			16729: out = 16'(5255);
			16730: out = 16'(3726);
			16731: out = 16'(-512);
			16732: out = 16'(-5265);
			16733: out = 16'(-3220);
			16734: out = 16'(-2389);
			16735: out = 16'(481);
			16736: out = 16'(-3323);
			16737: out = 16'(-2851);
			16738: out = 16'(-3485);
			16739: out = 16'(5853);
			16740: out = 16'(7394);
			16741: out = 16'(6201);
			16742: out = 16'(-2862);
			16743: out = 16'(-7243);
			16744: out = 16'(-5198);
			16745: out = 16'(-1190);
			16746: out = 16'(3165);
			16747: out = 16'(4000);
			16748: out = 16'(4340);
			16749: out = 16'(2787);
			16750: out = 16'(-17);
			16751: out = 16'(211);
			16752: out = 16'(2119);
			16753: out = 16'(2138);
			16754: out = 16'(2042);
			16755: out = 16'(-180);
			16756: out = 16'(1089);
			16757: out = 16'(-785);
			16758: out = 16'(-2450);
			16759: out = 16'(-5118);
			16760: out = 16'(-5283);
			16761: out = 16'(-4604);
			16762: out = 16'(-173);
			16763: out = 16'(2651);
			16764: out = 16'(4500);
			16765: out = 16'(1048);
			16766: out = 16'(-1813);
			16767: out = 16'(-248);
			16768: out = 16'(-405);
			16769: out = 16'(-11);
			16770: out = 16'(-161);
			16771: out = 16'(-601);
			16772: out = 16'(-1497);
			16773: out = 16'(-1388);
			16774: out = 16'(-546);
			16775: out = 16'(1081);
			16776: out = 16'(1583);
			16777: out = 16'(567);
			16778: out = 16'(-3794);
			16779: out = 16'(0);
			16780: out = 16'(729);
			16781: out = 16'(37);
			16782: out = 16'(-1575);
			16783: out = 16'(-1501);
			16784: out = 16'(3719);
			16785: out = 16'(2027);
			16786: out = 16'(654);
			16787: out = 16'(650);
			16788: out = 16'(628);
			16789: out = 16'(759);
			16790: out = 16'(-1239);
			16791: out = 16'(-908);
			16792: out = 16'(-32);
			16793: out = 16'(-160);
			16794: out = 16'(-464);
			16795: out = 16'(-1440);
			16796: out = 16'(-433);
			16797: out = 16'(1231);
			16798: out = 16'(5596);
			16799: out = 16'(1202);
			16800: out = 16'(-1153);
			16801: out = 16'(-2504);
			16802: out = 16'(-513);
			16803: out = 16'(1026);
			16804: out = 16'(668);
			16805: out = 16'(682);
			16806: out = 16'(440);
			16807: out = 16'(337);
			16808: out = 16'(1788);
			16809: out = 16'(3419);
			16810: out = 16'(151);
			16811: out = 16'(-1158);
			16812: out = 16'(-2617);
			16813: out = 16'(2922);
			16814: out = 16'(3788);
			16815: out = 16'(1044);
			16816: out = 16'(1058);
			16817: out = 16'(-949);
			16818: out = 16'(-2295);
			16819: out = 16'(-5700);
			16820: out = 16'(-5927);
			16821: out = 16'(-1694);
			16822: out = 16'(-21);
			16823: out = 16'(1358);
			16824: out = 16'(5215);
			16825: out = 16'(2897);
			16826: out = 16'(-16);
			16827: out = 16'(-6055);
			16828: out = 16'(-4268);
			16829: out = 16'(486);
			16830: out = 16'(285);
			16831: out = 16'(-824);
			16832: out = 16'(-4883);
			16833: out = 16'(-685);
			16834: out = 16'(-1196);
			16835: out = 16'(-5661);
			16836: out = 16'(-221);
			16837: out = 16'(3218);
			16838: out = 16'(6293);
			16839: out = 16'(2864);
			16840: out = 16'(-262);
			16841: out = 16'(-2207);
			16842: out = 16'(-902);
			16843: out = 16'(831);
			16844: out = 16'(628);
			16845: out = 16'(-1552);
			16846: out = 16'(-4728);
			16847: out = 16'(-2328);
			16848: out = 16'(-1469);
			16849: out = 16'(449);
			16850: out = 16'(-159);
			16851: out = 16'(295);
			16852: out = 16'(-422);
			16853: out = 16'(753);
			16854: out = 16'(451);
			16855: out = 16'(318);
			16856: out = 16'(-1509);
			16857: out = 16'(-2292);
			16858: out = 16'(-3302);
			16859: out = 16'(-521);
			16860: out = 16'(1602);
			16861: out = 16'(2975);
			16862: out = 16'(963);
			16863: out = 16'(-1178);
			16864: out = 16'(1720);
			16865: out = 16'(3737);
			16866: out = 16'(6428);
			16867: out = 16'(1303);
			16868: out = 16'(180);
			16869: out = 16'(-541);
			16870: out = 16'(722);
			16871: out = 16'(215);
			16872: out = 16'(-1413);
			16873: out = 16'(44);
			16874: out = 16'(1799);
			16875: out = 16'(4264);
			16876: out = 16'(3907);
			16877: out = 16'(2703);
			16878: out = 16'(640);
			16879: out = 16'(-1452);
			16880: out = 16'(-2342);
			16881: out = 16'(1319);
			16882: out = 16'(1581);
			16883: out = 16'(1430);
			16884: out = 16'(752);
			16885: out = 16'(125);
			16886: out = 16'(-473);
			16887: out = 16'(-1425);
			16888: out = 16'(-1142);
			16889: out = 16'(494);
			16890: out = 16'(468);
			16891: out = 16'(29);
			16892: out = 16'(-2952);
			16893: out = 16'(-1600);
			16894: out = 16'(-2178);
			16895: out = 16'(-3061);
			16896: out = 16'(-6893);
			16897: out = 16'(-7204);
			16898: out = 16'(3931);
			16899: out = 16'(6285);
			16900: out = 16'(7007);
			16901: out = 16'(-2496);
			16902: out = 16'(-4057);
			16903: out = 16'(-4323);
			16904: out = 16'(-155);
			16905: out = 16'(773);
			16906: out = 16'(661);
			16907: out = 16'(1673);
			16908: out = 16'(906);
			16909: out = 16'(-2672);
			16910: out = 16'(2150);
			16911: out = 16'(4202);
			16912: out = 16'(6319);
			16913: out = 16'(5);
			16914: out = 16'(-4013);
			16915: out = 16'(-2192);
			16916: out = 16'(-1367);
			16917: out = 16'(242);
			16918: out = 16'(-312);
			16919: out = 16'(-424);
			16920: out = 16'(-1681);
			16921: out = 16'(-1045);
			16922: out = 16'(-1915);
			16923: out = 16'(-2085);
			16924: out = 16'(-2549);
			16925: out = 16'(-183);
			16926: out = 16'(3968);
			16927: out = 16'(1440);
			16928: out = 16'(-155);
			16929: out = 16'(-2361);
			16930: out = 16'(-1503);
			16931: out = 16'(-1349);
			16932: out = 16'(-2151);
			16933: out = 16'(-1636);
			16934: out = 16'(-655);
			16935: out = 16'(886);
			16936: out = 16'(1718);
			16937: out = 16'(1694);
			16938: out = 16'(-662);
			16939: out = 16'(-2199);
			16940: out = 16'(-2920);
			16941: out = 16'(-888);
			16942: out = 16'(2401);
			16943: out = 16'(6567);
			16944: out = 16'(4230);
			16945: out = 16'(2004);
			16946: out = 16'(-2648);
			16947: out = 16'(116);
			16948: out = 16'(1294);
			16949: out = 16'(2825);
			16950: out = 16'(859);
			16951: out = 16'(-433);
			16952: out = 16'(-1333);
			16953: out = 16'(-1368);
			16954: out = 16'(-1032);
			16955: out = 16'(2612);
			16956: out = 16'(1637);
			16957: out = 16'(190);
			16958: out = 16'(-4954);
			16959: out = 16'(-2493);
			16960: out = 16'(3436);
			16961: out = 16'(2447);
			16962: out = 16'(966);
			16963: out = 16'(-5186);
			16964: out = 16'(-118);
			16965: out = 16'(121);
			16966: out = 16'(100);
			16967: out = 16'(-4047);
			16968: out = 16'(-4259);
			16969: out = 16'(433);
			16970: out = 16'(4120);
			16971: out = 16'(6101);
			16972: out = 16'(2793);
			16973: out = 16'(1750);
			16974: out = 16'(510);
			16975: out = 16'(8);
			16976: out = 16'(-1046);
			16977: out = 16'(-2574);
			16978: out = 16'(1422);
			16979: out = 16'(809);
			16980: out = 16'(-341);
			16981: out = 16'(-6280);
			16982: out = 16'(-4950);
			16983: out = 16'(3244);
			16984: out = 16'(5905);
			16985: out = 16'(7450);
			16986: out = 16'(3868);
			16987: out = 16'(2918);
			16988: out = 16'(784);
			16989: out = 16'(912);
			16990: out = 16'(10);
			16991: out = 16'(-70);
			16992: out = 16'(-4737);
			16993: out = 16'(-4171);
			16994: out = 16'(-3525);
			16995: out = 16'(283);
			16996: out = 16'(494);
			16997: out = 16'(410);
			16998: out = 16'(-3035);
			16999: out = 16'(-2638);
			17000: out = 16'(-453);
			17001: out = 16'(-194);
			17002: out = 16'(-158);
			17003: out = 16'(1104);
			17004: out = 16'(-4234);
			17005: out = 16'(-7275);
			17006: out = 16'(-8800);
			17007: out = 16'(-2995);
			17008: out = 16'(1861);
			17009: out = 16'(-64);
			17010: out = 16'(-1113);
			17011: out = 16'(-3222);
			17012: out = 16'(121);
			17013: out = 16'(2322);
			17014: out = 16'(6120);
			17015: out = 16'(1304);
			17016: out = 16'(969);
			17017: out = 16'(-656);
			17018: out = 16'(4058);
			17019: out = 16'(3563);
			17020: out = 16'(2029);
			17021: out = 16'(-2045);
			17022: out = 16'(-3568);
			17023: out = 16'(-4718);
			17024: out = 16'(986);
			17025: out = 16'(4090);
			17026: out = 16'(4766);
			17027: out = 16'(-490);
			17028: out = 16'(-4457);
			17029: out = 16'(222);
			17030: out = 16'(3659);
			17031: out = 16'(7048);
			17032: out = 16'(3803);
			17033: out = 16'(1432);
			17034: out = 16'(-2064);
			17035: out = 16'(-4841);
			17036: out = 16'(-4653);
			17037: out = 16'(-922);
			17038: out = 16'(637);
			17039: out = 16'(2430);
			17040: out = 16'(2388);
			17041: out = 16'(2225);
			17042: out = 16'(1041);
			17043: out = 16'(-448);
			17044: out = 16'(115);
			17045: out = 16'(862);
			17046: out = 16'(578);
			17047: out = 16'(291);
			17048: out = 16'(-837);
			17049: out = 16'(-3988);
			17050: out = 16'(-5683);
			17051: out = 16'(-6298);
			17052: out = 16'(-120);
			17053: out = 16'(1159);
			17054: out = 16'(531);
			17055: out = 16'(234);
			17056: out = 16'(149);
			17057: out = 16'(1088);
			17058: out = 16'(586);
			17059: out = 16'(1481);
			17060: out = 16'(4631);
			17061: out = 16'(1451);
			17062: out = 16'(-1160);
			17063: out = 16'(-4397);
			17064: out = 16'(-2769);
			17065: out = 16'(-1510);
			17066: out = 16'(-5287);
			17067: out = 16'(-5831);
			17068: out = 16'(-5964);
			17069: out = 16'(-374);
			17070: out = 16'(1485);
			17071: out = 16'(3236);
			17072: out = 16'(-1389);
			17073: out = 16'(-1672);
			17074: out = 16'(-1039);
			17075: out = 16'(1033);
			17076: out = 16'(-148);
			17077: out = 16'(-4097);
			17078: out = 16'(-4825);
			17079: out = 16'(-3358);
			17080: out = 16'(3554);
			17081: out = 16'(1780);
			17082: out = 16'(1534);
			17083: out = 16'(3951);
			17084: out = 16'(5707);
			17085: out = 16'(6465);
			17086: out = 16'(-4817);
			17087: out = 16'(-2392);
			17088: out = 16'(1392);
			17089: out = 16'(5215);
			17090: out = 16'(2348);
			17091: out = 16'(-3807);
			17092: out = 16'(-2927);
			17093: out = 16'(-1948);
			17094: out = 16'(1624);
			17095: out = 16'(1538);
			17096: out = 16'(2559);
			17097: out = 16'(2765);
			17098: out = 16'(1854);
			17099: out = 16'(534);
			17100: out = 16'(265);
			17101: out = 16'(-151);
			17102: out = 16'(305);
			17103: out = 16'(476);
			17104: out = 16'(1897);
			17105: out = 16'(2628);
			17106: out = 16'(239);
			17107: out = 16'(-624);
			17108: out = 16'(-1277);
			17109: out = 16'(572);
			17110: out = 16'(1854);
			17111: out = 16'(3765);
			17112: out = 16'(1079);
			17113: out = 16'(255);
			17114: out = 16'(-626);
			17115: out = 16'(2480);
			17116: out = 16'(3187);
			17117: out = 16'(1582);
			17118: out = 16'(468);
			17119: out = 16'(-1162);
			17120: out = 16'(-5598);
			17121: out = 16'(-2890);
			17122: out = 16'(378);
			17123: out = 16'(3140);
			17124: out = 16'(1993);
			17125: out = 16'(-650);
			17126: out = 16'(742);
			17127: out = 16'(-867);
			17128: out = 16'(-2519);
			17129: out = 16'(-527);
			17130: out = 16'(-466);
			17131: out = 16'(-1498);
			17132: out = 16'(-2171);
			17133: out = 16'(-1445);
			17134: out = 16'(2048);
			17135: out = 16'(919);
			17136: out = 16'(-419);
			17137: out = 16'(-5626);
			17138: out = 16'(-3436);
			17139: out = 16'(-2020);
			17140: out = 16'(-1096);
			17141: out = 16'(-2246);
			17142: out = 16'(-2753);
			17143: out = 16'(271);
			17144: out = 16'(2775);
			17145: out = 16'(4621);
			17146: out = 16'(1836);
			17147: out = 16'(-1959);
			17148: out = 16'(-7686);
			17149: out = 16'(-1444);
			17150: out = 16'(2415);
			17151: out = 16'(7414);
			17152: out = 16'(2686);
			17153: out = 16'(67);
			17154: out = 16'(-2256);
			17155: out = 16'(-428);
			17156: out = 16'(1261);
			17157: out = 16'(2741);
			17158: out = 16'(1344);
			17159: out = 16'(-558);
			17160: out = 16'(-1971);
			17161: out = 16'(-1991);
			17162: out = 16'(-1153);
			17163: out = 16'(-3013);
			17164: out = 16'(-4267);
			17165: out = 16'(-6427);
			17166: out = 16'(-756);
			17167: out = 16'(1756);
			17168: out = 16'(5274);
			17169: out = 16'(1464);
			17170: out = 16'(1083);
			17171: out = 16'(362);
			17172: out = 16'(5066);
			17173: out = 16'(5035);
			17174: out = 16'(1159);
			17175: out = 16'(-5129);
			17176: out = 16'(-8257);
			17177: out = 16'(-2658);
			17178: out = 16'(2336);
			17179: out = 16'(7000);
			17180: out = 16'(6818);
			17181: out = 16'(3923);
			17182: out = 16'(-1334);
			17183: out = 16'(-1746);
			17184: out = 16'(-1997);
			17185: out = 16'(378);
			17186: out = 16'(-408);
			17187: out = 16'(-138);
			17188: out = 16'(-1632);
			17189: out = 16'(177);
			17190: out = 16'(1390);
			17191: out = 16'(4692);
			17192: out = 16'(2509);
			17193: out = 16'(1323);
			17194: out = 16'(-330);
			17195: out = 16'(877);
			17196: out = 16'(1555);
			17197: out = 16'(480);
			17198: out = 16'(-112);
			17199: out = 16'(-962);
			17200: out = 16'(-3997);
			17201: out = 16'(-5862);
			17202: out = 16'(-7563);
			17203: out = 16'(-1527);
			17204: out = 16'(665);
			17205: out = 16'(2086);
			17206: out = 16'(-2105);
			17207: out = 16'(-2388);
			17208: out = 16'(931);
			17209: out = 16'(3329);
			17210: out = 16'(4194);
			17211: out = 16'(414);
			17212: out = 16'(-889);
			17213: out = 16'(-2205);
			17214: out = 16'(3149);
			17215: out = 16'(870);
			17216: out = 16'(-299);
			17217: out = 16'(-5412);
			17218: out = 16'(-2959);
			17219: out = 16'(265);
			17220: out = 16'(5539);
			17221: out = 16'(5243);
			17222: out = 16'(3310);
			17223: out = 16'(-3775);
			17224: out = 16'(-4291);
			17225: out = 16'(365);
			17226: out = 16'(4795);
			17227: out = 16'(5839);
			17228: out = 16'(-1195);
			17229: out = 16'(-18);
			17230: out = 16'(-949);
			17231: out = 16'(269);
			17232: out = 16'(-1856);
			17233: out = 16'(-2181);
			17234: out = 16'(-1813);
			17235: out = 16'(-25);
			17236: out = 16'(1064);
			17237: out = 16'(5033);
			17238: out = 16'(3201);
			17239: out = 16'(-15);
			17240: out = 16'(-2006);
			17241: out = 16'(-1966);
			17242: out = 16'(2);
			17243: out = 16'(-1246);
			17244: out = 16'(-1813);
			17245: out = 16'(-2390);
			17246: out = 16'(-3255);
			17247: out = 16'(-1783);
			17248: out = 16'(4601);
			17249: out = 16'(4321);
			17250: out = 16'(3563);
			17251: out = 16'(-2575);
			17252: out = 16'(280);
			17253: out = 16'(2975);
			17254: out = 16'(3226);
			17255: out = 16'(1761);
			17256: out = 16'(-1207);
			17257: out = 16'(716);
			17258: out = 16'(-1508);
			17259: out = 16'(-3586);
			17260: out = 16'(-4666);
			17261: out = 16'(-2954);
			17262: out = 16'(685);
			17263: out = 16'(596);
			17264: out = 16'(2101);
			17265: out = 16'(7160);
			17266: out = 16'(2354);
			17267: out = 16'(317);
			17268: out = 16'(-964);
			17269: out = 16'(2902);
			17270: out = 16'(4348);
			17271: out = 16'(-159);
			17272: out = 16'(-5014);
			17273: out = 16'(-9558);
			17274: out = 16'(-8941);
			17275: out = 16'(-5846);
			17276: out = 16'(-325);
			17277: out = 16'(2499);
			17278: out = 16'(3885);
			17279: out = 16'(2308);
			17280: out = 16'(2296);
			17281: out = 16'(1605);
			17282: out = 16'(2919);
			17283: out = 16'(-430);
			17284: out = 16'(-1855);
			17285: out = 16'(-2522);
			17286: out = 16'(-1223);
			17287: out = 16'(-674);
			17288: out = 16'(-3505);
			17289: out = 16'(-1723);
			17290: out = 16'(389);
			17291: out = 16'(4072);
			17292: out = 16'(4517);
			17293: out = 16'(4021);
			17294: out = 16'(327);
			17295: out = 16'(-483);
			17296: out = 16'(-580);
			17297: out = 16'(302);
			17298: out = 16'(-257);
			17299: out = 16'(-1608);
			17300: out = 16'(-3735);
			17301: out = 16'(-4649);
			17302: out = 16'(-4390);
			17303: out = 16'(-330);
			17304: out = 16'(2660);
			17305: out = 16'(2383);
			17306: out = 16'(2967);
			17307: out = 16'(2718);
			17308: out = 16'(5365);
			17309: out = 16'(3576);
			17310: out = 16'(2207);
			17311: out = 16'(671);
			17312: out = 16'(239);
			17313: out = 16'(-898);
			17314: out = 16'(-1757);
			17315: out = 16'(-6029);
			17316: out = 16'(-11401);
			17317: out = 16'(-9612);
			17318: out = 16'(-4921);
			17319: out = 16'(4448);
			17320: out = 16'(2786);
			17321: out = 16'(3495);
			17322: out = 16'(4377);
			17323: out = 16'(3613);
			17324: out = 16'(1843);
			17325: out = 16'(178);
			17326: out = 16'(-445);
			17327: out = 16'(-373);
			17328: out = 16'(-5649);
			17329: out = 16'(-2269);
			17330: out = 16'(1337);
			17331: out = 16'(2669);
			17332: out = 16'(21);
			17333: out = 16'(-4765);
			17334: out = 16'(-138);
			17335: out = 16'(2005);
			17336: out = 16'(4749);
			17337: out = 16'(5548);
			17338: out = 16'(5162);
			17339: out = 16'(1088);
			17340: out = 16'(558);
			17341: out = 16'(-1158);
			17342: out = 16'(1408);
			17343: out = 16'(-4347);
			17344: out = 16'(-7118);
			17345: out = 16'(-10491);
			17346: out = 16'(-2194);
			17347: out = 16'(5533);
			17348: out = 16'(3333);
			17349: out = 16'(2208);
			17350: out = 16'(-466);
			17351: out = 16'(2513);
			17352: out = 16'(2254);
			17353: out = 16'(1489);
			17354: out = 16'(976);
			17355: out = 16'(-987);
			17356: out = 16'(-3441);
			17357: out = 16'(-6523);
			17358: out = 16'(-6928);
			17359: out = 16'(-4189);
			17360: out = 16'(-999);
			17361: out = 16'(1332);
			17362: out = 16'(1032);
			17363: out = 16'(466);
			17364: out = 16'(113);
			17365: out = 16'(1764);
			17366: out = 16'(4515);
			17367: out = 16'(6872);
			17368: out = 16'(1400);
			17369: out = 16'(300);
			17370: out = 16'(-809);
			17371: out = 16'(-6044);
			17372: out = 16'(-9287);
			17373: out = 16'(-11858);
			17374: out = 16'(-2368);
			17375: out = 16'(2991);
			17376: out = 16'(4554);
			17377: out = 16'(4275);
			17378: out = 16'(4442);
			17379: out = 16'(8722);
			17380: out = 16'(5710);
			17381: out = 16'(3473);
			17382: out = 16'(-345);
			17383: out = 16'(-414);
			17384: out = 16'(-920);
			17385: out = 16'(-2868);
			17386: out = 16'(-4473);
			17387: out = 16'(-4958);
			17388: out = 16'(-2114);
			17389: out = 16'(979);
			17390: out = 16'(3772);
			17391: out = 16'(6209);
			17392: out = 16'(5511);
			17393: out = 16'(2222);
			17394: out = 16'(609);
			17395: out = 16'(-20);
			17396: out = 16'(2736);
			17397: out = 16'(-258);
			17398: out = 16'(-2402);
			17399: out = 16'(-5449);
			17400: out = 16'(-3808);
			17401: out = 16'(-1981);
			17402: out = 16'(-2580);
			17403: out = 16'(-961);
			17404: out = 16'(425);
			17405: out = 16'(4705);
			17406: out = 16'(4513);
			17407: out = 16'(3015);
			17408: out = 16'(-1386);
			17409: out = 16'(-1829);
			17410: out = 16'(788);
			17411: out = 16'(-1115);
			17412: out = 16'(-2560);
			17413: out = 16'(-6813);
			17414: out = 16'(-1744);
			17415: out = 16'(62);
			17416: out = 16'(-1232);
			17417: out = 16'(-1800);
			17418: out = 16'(-1189);
			17419: out = 16'(5313);
			17420: out = 16'(2452);
			17421: out = 16'(-376);
			17422: out = 16'(978);
			17423: out = 16'(2185);
			17424: out = 16'(4283);
			17425: out = 16'(-5288);
			17426: out = 16'(-6017);
			17427: out = 16'(-5103);
			17428: out = 16'(1421);
			17429: out = 16'(2095);
			17430: out = 16'(-307);
			17431: out = 16'(-5258);
			17432: out = 16'(-5966);
			17433: out = 16'(319);
			17434: out = 16'(3230);
			17435: out = 16'(5481);
			17436: out = 16'(209);
			17437: out = 16'(1991);
			17438: out = 16'(1512);
			17439: out = 16'(3233);
			17440: out = 16'(749);
			17441: out = 16'(-569);
			17442: out = 16'(-7163);
			17443: out = 16'(-3867);
			17444: out = 16'(1215);
			17445: out = 16'(4841);
			17446: out = 16'(2256);
			17447: out = 16'(-4714);
			17448: out = 16'(-1948);
			17449: out = 16'(970);
			17450: out = 16'(6270);
			17451: out = 16'(7643);
			17452: out = 16'(6177);
			17453: out = 16'(-2731);
			17454: out = 16'(-2955);
			17455: out = 16'(-2328);
			17456: out = 16'(6723);
			17457: out = 16'(3127);
			17458: out = 16'(170);
			17459: out = 16'(-530);
			17460: out = 16'(587);
			17461: out = 16'(2739);
			17462: out = 16'(1887);
			17463: out = 16'(3763);
			17464: out = 16'(5472);
			17465: out = 16'(4929);
			17466: out = 16'(2718);
			17467: out = 16'(-1406);
			17468: out = 16'(-2216);
			17469: out = 16'(-4210);
			17470: out = 16'(-6944);
			17471: out = 16'(-6352);
			17472: out = 16'(-4597);
			17473: out = 16'(-389);
			17474: out = 16'(161);
			17475: out = 16'(801);
			17476: out = 16'(196);
			17477: out = 16'(250);
			17478: out = 16'(-398);
			17479: out = 16'(3419);
			17480: out = 16'(163);
			17481: out = 16'(-3976);
			17482: out = 16'(-6266);
			17483: out = 16'(-4463);
			17484: out = 16'(359);
			17485: out = 16'(452);
			17486: out = 16'(-64);
			17487: out = 16'(-3620);
			17488: out = 16'(-884);
			17489: out = 16'(816);
			17490: out = 16'(3566);
			17491: out = 16'(2905);
			17492: out = 16'(2181);
			17493: out = 16'(840);
			17494: out = 16'(-984);
			17495: out = 16'(-2607);
			17496: out = 16'(-361);
			17497: out = 16'(-1107);
			17498: out = 16'(-1209);
			17499: out = 16'(-814);
			17500: out = 16'(1282);
			17501: out = 16'(3463);
			17502: out = 16'(469);
			17503: out = 16'(-763);
			17504: out = 16'(-1374);
			17505: out = 16'(-152);
			17506: out = 16'(813);
			17507: out = 16'(510);
			17508: out = 16'(1565);
			17509: out = 16'(1193);
			17510: out = 16'(694);
			17511: out = 16'(-2640);
			17512: out = 16'(-4990);
			17513: out = 16'(-7496);
			17514: out = 16'(-3125);
			17515: out = 16'(1696);
			17516: out = 16'(-303);
			17517: out = 16'(272);
			17518: out = 16'(-483);
			17519: out = 16'(1175);
			17520: out = 16'(-282);
			17521: out = 16'(-2204);
			17522: out = 16'(81);
			17523: out = 16'(780);
			17524: out = 16'(-129);
			17525: out = 16'(249);
			17526: out = 16'(3);
			17527: out = 16'(976);
			17528: out = 16'(-825);
			17529: out = 16'(-536);
			17530: out = 16'(1615);
			17531: out = 16'(3505);
			17532: out = 16'(4191);
			17533: out = 16'(2802);
			17534: out = 16'(1547);
			17535: out = 16'(559);
			17536: out = 16'(-1314);
			17537: out = 16'(-1336);
			17538: out = 16'(-1453);
			17539: out = 16'(3012);
			17540: out = 16'(1982);
			17541: out = 16'(-542);
			17542: out = 16'(-5961);
			17543: out = 16'(-6019);
			17544: out = 16'(-928);
			17545: out = 16'(4107);
			17546: out = 16'(7409);
			17547: out = 16'(6197);
			17548: out = 16'(4404);
			17549: out = 16'(1135);
			17550: out = 16'(-981);
			17551: out = 16'(-3499);
			17552: out = 16'(-4093);
			17553: out = 16'(-4);
			17554: out = 16'(638);
			17555: out = 16'(719);
			17556: out = 16'(409);
			17557: out = 16'(145);
			17558: out = 16'(-621);
			17559: out = 16'(4116);
			17560: out = 16'(4592);
			17561: out = 16'(4085);
			17562: out = 16'(-2498);
			17563: out = 16'(-3688);
			17564: out = 16'(1741);
			17565: out = 16'(3424);
			17566: out = 16'(4132);
			17567: out = 16'(-2130);
			17568: out = 16'(-343);
			17569: out = 16'(-507);
			17570: out = 16'(-3261);
			17571: out = 16'(-4403);
			17572: out = 16'(-3714);
			17573: out = 16'(3737);
			17574: out = 16'(5564);
			17575: out = 16'(5109);
			17576: out = 16'(1484);
			17577: out = 16'(-451);
			17578: out = 16'(-425);
			17579: out = 16'(-4688);
			17580: out = 16'(-6371);
			17581: out = 16'(-7797);
			17582: out = 16'(-4040);
			17583: out = 16'(-1635);
			17584: out = 16'(-92);
			17585: out = 16'(-940);
			17586: out = 16'(-1095);
			17587: out = 16'(-675);
			17588: out = 16'(3195);
			17589: out = 16'(6043);
			17590: out = 16'(3481);
			17591: out = 16'(428);
			17592: out = 16'(-4166);
			17593: out = 16'(-1187);
			17594: out = 16'(-2559);
			17595: out = 16'(-3217);
			17596: out = 16'(-6849);
			17597: out = 16'(-5782);
			17598: out = 16'(-1833);
			17599: out = 16'(760);
			17600: out = 16'(2361);
			17601: out = 16'(1700);
			17602: out = 16'(1388);
			17603: out = 16'(450);
			17604: out = 16'(1243);
			17605: out = 16'(654);
			17606: out = 16'(904);
			17607: out = 16'(-2484);
			17608: out = 16'(-460);
			17609: out = 16'(492);
			17610: out = 16'(1482);
			17611: out = 16'(-2361);
			17612: out = 16'(-6268);
			17613: out = 16'(-4892);
			17614: out = 16'(73);
			17615: out = 16'(7419);
			17616: out = 16'(6768);
			17617: out = 16'(5817);
			17618: out = 16'(3359);
			17619: out = 16'(-588);
			17620: out = 16'(-2780);
			17621: out = 16'(-2319);
			17622: out = 16'(650);
			17623: out = 16'(2969);
			17624: out = 16'(2423);
			17625: out = 16'(510);
			17626: out = 16'(-1924);
			17627: out = 16'(-1306);
			17628: out = 16'(-1021);
			17629: out = 16'(43);
			17630: out = 16'(524);
			17631: out = 16'(377);
			17632: out = 16'(-564);
			17633: out = 16'(-268);
			17634: out = 16'(871);
			17635: out = 16'(3522);
			17636: out = 16'(-887);
			17637: out = 16'(-3163);
			17638: out = 16'(-3046);
			17639: out = 16'(-4358);
			17640: out = 16'(-3640);
			17641: out = 16'(-2648);
			17642: out = 16'(1468);
			17643: out = 16'(4061);
			17644: out = 16'(6122);
			17645: out = 16'(2771);
			17646: out = 16'(-792);
			17647: out = 16'(-3080);
			17648: out = 16'(-1644);
			17649: out = 16'(1244);
			17650: out = 16'(3742);
			17651: out = 16'(3035);
			17652: out = 16'(-33);
			17653: out = 16'(-5546);
			17654: out = 16'(-7479);
			17655: out = 16'(-4827);
			17656: out = 16'(-1338);
			17657: out = 16'(2725);
			17658: out = 16'(4827);
			17659: out = 16'(5096);
			17660: out = 16'(3194);
			17661: out = 16'(230);
			17662: out = 16'(-1108);
			17663: out = 16'(-1148);
			17664: out = 16'(198);
			17665: out = 16'(650);
			17666: out = 16'(-162);
			17667: out = 16'(-5321);
			17668: out = 16'(-7621);
			17669: out = 16'(-7873);
			17670: out = 16'(-1769);
			17671: out = 16'(1588);
			17672: out = 16'(1594);
			17673: out = 16'(5088);
			17674: out = 16'(4364);
			17675: out = 16'(3111);
			17676: out = 16'(-3651);
			17677: out = 16'(-5429);
			17678: out = 16'(748);
			17679: out = 16'(2497);
			17680: out = 16'(2842);
			17681: out = 16'(-3927);
			17682: out = 16'(-4275);
			17683: out = 16'(-3264);
			17684: out = 16'(2826);
			17685: out = 16'(5133);
			17686: out = 16'(5971);
			17687: out = 16'(6294);
			17688: out = 16'(3805);
			17689: out = 16'(440);
			17690: out = 16'(-2624);
			17691: out = 16'(-2197);
			17692: out = 16'(1980);
			17693: out = 16'(785);
			17694: out = 16'(657);
			17695: out = 16'(449);
			17696: out = 16'(-847);
			17697: out = 16'(-1802);
			17698: out = 16'(-3577);
			17699: out = 16'(511);
			17700: out = 16'(3621);
			17701: out = 16'(686);
			17702: out = 16'(-148);
			17703: out = 16'(-1715);
			17704: out = 16'(-424);
			17705: out = 16'(-583);
			17706: out = 16'(-362);
			17707: out = 16'(223);
			17708: out = 16'(563);
			17709: out = 16'(341);
			17710: out = 16'(-1658);
			17711: out = 16'(-2220);
			17712: out = 16'(-132);
			17713: out = 16'(-2618);
			17714: out = 16'(-3139);
			17715: out = 16'(-2319);
			17716: out = 16'(-855);
			17717: out = 16'(371);
			17718: out = 16'(793);
			17719: out = 16'(1517);
			17720: out = 16'(1491);
			17721: out = 16'(-1878);
			17722: out = 16'(-2333);
			17723: out = 16'(-2045);
			17724: out = 16'(-533);
			17725: out = 16'(17);
			17726: out = 16'(116);
			17727: out = 16'(726);
			17728: out = 16'(1838);
			17729: out = 16'(3699);
			17730: out = 16'(2251);
			17731: out = 16'(1260);
			17732: out = 16'(-134);
			17733: out = 16'(-95);
			17734: out = 16'(-3);
			17735: out = 16'(572);
			17736: out = 16'(557);
			17737: out = 16'(-358);
			17738: out = 16'(-6976);
			17739: out = 16'(-7352);
			17740: out = 16'(-6491);
			17741: out = 16'(1205);
			17742: out = 16'(2202);
			17743: out = 16'(1967);
			17744: out = 16'(-1464);
			17745: out = 16'(-1405);
			17746: out = 16'(53);
			17747: out = 16'(2347);
			17748: out = 16'(2696);
			17749: out = 16'(2009);
			17750: out = 16'(-1575);
			17751: out = 16'(-3103);
			17752: out = 16'(-2110);
			17753: out = 16'(3082);
			17754: out = 16'(6194);
			17755: out = 16'(652);
			17756: out = 16'(716);
			17757: out = 16'(-656);
			17758: out = 16'(1393);
			17759: out = 16'(-473);
			17760: out = 16'(-813);
			17761: out = 16'(141);
			17762: out = 16'(3614);
			17763: out = 16'(6662);
			17764: out = 16'(5620);
			17765: out = 16'(3193);
			17766: out = 16'(346);
			17767: out = 16'(-2865);
			17768: out = 16'(-1698);
			17769: out = 16'(4292);
			17770: out = 16'(5155);
			17771: out = 16'(4260);
			17772: out = 16'(-2819);
			17773: out = 16'(-2646);
			17774: out = 16'(-2225);
			17775: out = 16'(1320);
			17776: out = 16'(1391);
			17777: out = 16'(1129);
			17778: out = 16'(-1307);
			17779: out = 16'(-2623);
			17780: out = 16'(-3493);
			17781: out = 16'(-348);
			17782: out = 16'(1229);
			17783: out = 16'(2383);
			17784: out = 16'(779);
			17785: out = 16'(-90);
			17786: out = 16'(-292);
			17787: out = 16'(-672);
			17788: out = 16'(-983);
			17789: out = 16'(-2823);
			17790: out = 16'(-948);
			17791: out = 16'(-88);
			17792: out = 16'(1702);
			17793: out = 16'(656);
			17794: out = 16'(-101);
			17795: out = 16'(-5650);
			17796: out = 16'(-2952);
			17797: out = 16'(-154);
			17798: out = 16'(4035);
			17799: out = 16'(2091);
			17800: out = 16'(-816);
			17801: out = 16'(-7613);
			17802: out = 16'(-5791);
			17803: out = 16'(1116);
			17804: out = 16'(6366);
			17805: out = 16'(7265);
			17806: out = 16'(3048);
			17807: out = 16'(-3706);
			17808: out = 16'(-8317);
			17809: out = 16'(-5960);
			17810: out = 16'(-3794);
			17811: out = 16'(-111);
			17812: out = 16'(114);
			17813: out = 16'(1194);
			17814: out = 16'(-13);
			17815: out = 16'(-2354);
			17816: out = 16'(-4724);
			17817: out = 16'(-5651);
			17818: out = 16'(1560);
			17819: out = 16'(3956);
			17820: out = 16'(4440);
			17821: out = 16'(911);
			17822: out = 16'(-134);
			17823: out = 16'(1275);
			17824: out = 16'(1443);
			17825: out = 16'(1857);
			17826: out = 16'(394);
			17827: out = 16'(1680);
			17828: out = 16'(734);
			17829: out = 16'(-3993);
			17830: out = 16'(-4899);
			17831: out = 16'(-4275);
			17832: out = 16'(2427);
			17833: out = 16'(3257);
			17834: out = 16'(3426);
			17835: out = 16'(-1687);
			17836: out = 16'(-1423);
			17837: out = 16'(73);
			17838: out = 16'(5095);
			17839: out = 16'(5125);
			17840: out = 16'(2226);
			17841: out = 16'(-205);
			17842: out = 16'(-1264);
			17843: out = 16'(1159);
			17844: out = 16'(456);
			17845: out = 16'(816);
			17846: out = 16'(-778);
			17847: out = 16'(1091);
			17848: out = 16'(1412);
			17849: out = 16'(918);
			17850: out = 16'(-94);
			17851: out = 16'(-752);
			17852: out = 16'(-4343);
			17853: out = 16'(-2554);
			17854: out = 16'(-144);
			17855: out = 16'(1592);
			17856: out = 16'(-56);
			17857: out = 16'(-3487);
			17858: out = 16'(-1093);
			17859: out = 16'(2108);
			17860: out = 16'(7722);
			17861: out = 16'(4445);
			17862: out = 16'(808);
			17863: out = 16'(-7919);
			17864: out = 16'(-2362);
			17865: out = 16'(1904);
			17866: out = 16'(5588);
			17867: out = 16'(4111);
			17868: out = 16'(1291);
			17869: out = 16'(-1839);
			17870: out = 16'(-4379);
			17871: out = 16'(-5188);
			17872: out = 16'(-2154);
			17873: out = 16'(495);
			17874: out = 16'(2556);
			17875: out = 16'(419);
			17876: out = 16'(-1679);
			17877: out = 16'(-4467);
			17878: out = 16'(-1097);
			17879: out = 16'(446);
			17880: out = 16'(714);
			17881: out = 16'(166);
			17882: out = 16'(89);
			17883: out = 16'(3843);
			17884: out = 16'(1533);
			17885: out = 16'(-276);
			17886: out = 16'(-8669);
			17887: out = 16'(-4973);
			17888: out = 16'(-1396);
			17889: out = 16'(5930);
			17890: out = 16'(2104);
			17891: out = 16'(-2782);
			17892: out = 16'(-7098);
			17893: out = 16'(-2243);
			17894: out = 16'(6986);
			17895: out = 16'(7746);
			17896: out = 16'(5739);
			17897: out = 16'(-1103);
			17898: out = 16'(-6179);
			17899: out = 16'(-7377);
			17900: out = 16'(1420);
			17901: out = 16'(147);
			17902: out = 16'(1326);
			17903: out = 16'(-629);
			17904: out = 16'(1479);
			17905: out = 16'(1195);
			17906: out = 16'(108);
			17907: out = 16'(-1708);
			17908: out = 16'(-2212);
			17909: out = 16'(-3443);
			17910: out = 16'(-2141);
			17911: out = 16'(-1163);
			17912: out = 16'(1650);
			17913: out = 16'(1698);
			17914: out = 16'(2061);
			17915: out = 16'(-3967);
			17916: out = 16'(-3942);
			17917: out = 16'(-72);
			17918: out = 16'(4434);
			17919: out = 16'(4983);
			17920: out = 16'(-1503);
			17921: out = 16'(-2953);
			17922: out = 16'(-3297);
			17923: out = 16'(4703);
			17924: out = 16'(2786);
			17925: out = 16'(1404);
			17926: out = 16'(-2051);
			17927: out = 16'(-1851);
			17928: out = 16'(-768);
			17929: out = 16'(3616);
			17930: out = 16'(5475);
			17931: out = 16'(6437);
			17932: out = 16'(1906);
			17933: out = 16'(-1248);
			17934: out = 16'(-4621);
			17935: out = 16'(-679);
			17936: out = 16'(2243);
			17937: out = 16'(5915);
			17938: out = 16'(1697);
			17939: out = 16'(-1415);
			17940: out = 16'(-3350);
			17941: out = 16'(-2566);
			17942: out = 16'(-979);
			17943: out = 16'(186);
			17944: out = 16'(-1281);
			17945: out = 16'(-3910);
			17946: out = 16'(-994);
			17947: out = 16'(-2682);
			17948: out = 16'(-2870);
			17949: out = 16'(-3862);
			17950: out = 16'(-474);
			17951: out = 16'(2723);
			17952: out = 16'(5927);
			17953: out = 16'(3328);
			17954: out = 16'(-2405);
			17955: out = 16'(-6993);
			17956: out = 16'(-6747);
			17957: out = 16'(234);
			17958: out = 16'(2953);
			17959: out = 16'(4195);
			17960: out = 16'(1053);
			17961: out = 16'(-1931);
			17962: out = 16'(-4381);
			17963: out = 16'(-3357);
			17964: out = 16'(1747);
			17965: out = 16'(7355);
			17966: out = 16'(1201);
			17967: out = 16'(-472);
			17968: out = 16'(-3453);
			17969: out = 16'(4964);
			17970: out = 16'(4989);
			17971: out = 16'(2255);
			17972: out = 16'(-260);
			17973: out = 16'(-1598);
			17974: out = 16'(316);
			17975: out = 16'(-2773);
			17976: out = 16'(-2752);
			17977: out = 16'(-1712);
			17978: out = 16'(2515);
			17979: out = 16'(3786);
			17980: out = 16'(237);
			17981: out = 16'(-3582);
			17982: out = 16'(-6419);
			17983: out = 16'(-2595);
			17984: out = 16'(136);
			17985: out = 16'(3096);
			17986: out = 16'(820);
			17987: out = 16'(444);
			17988: out = 16'(-60);
			17989: out = 16'(-1716);
			17990: out = 16'(-1917);
			17991: out = 16'(-1019);
			17992: out = 16'(2384);
			17993: out = 16'(3557);
			17994: out = 16'(1615);
			17995: out = 16'(1275);
			17996: out = 16'(197);
			17997: out = 16'(-194);
			17998: out = 16'(60);
			17999: out = 16'(920);
			18000: out = 16'(1643);
			18001: out = 16'(945);
			18002: out = 16'(-364);
			18003: out = 16'(32);
			18004: out = 16'(420);
			18005: out = 16'(1945);
			18006: out = 16'(-2069);
			18007: out = 16'(-839);
			18008: out = 16'(1804);
			18009: out = 16'(2584);
			18010: out = 16'(213);
			18011: out = 16'(-6898);
			18012: out = 16'(-4144);
			18013: out = 16'(-1422);
			18014: out = 16'(5589);
			18015: out = 16'(1649);
			18016: out = 16'(-1833);
			18017: out = 16'(-9476);
			18018: out = 16'(-4592);
			18019: out = 16'(987);
			18020: out = 16'(1405);
			18021: out = 16'(2003);
			18022: out = 16'(607);
			18023: out = 16'(1339);
			18024: out = 16'(-1420);
			18025: out = 16'(-3945);
			18026: out = 16'(-127);
			18027: out = 16'(3288);
			18028: out = 16'(6906);
			18029: out = 16'(3212);
			18030: out = 16'(1111);
			18031: out = 16'(1135);
			18032: out = 16'(-163);
			18033: out = 16'(-1006);
			18034: out = 16'(-5725);
			18035: out = 16'(-393);
			18036: out = 16'(3786);
			18037: out = 16'(8089);
			18038: out = 16'(4429);
			18039: out = 16'(-193);
			18040: out = 16'(-1924);
			18041: out = 16'(-1790);
			18042: out = 16'(350);
			18043: out = 16'(3137);
			18044: out = 16'(5486);
			18045: out = 16'(7004);
			18046: out = 16'(1235);
			18047: out = 16'(-1514);
			18048: out = 16'(-2732);
			18049: out = 16'(-597);
			18050: out = 16'(-1096);
			18051: out = 16'(-6868);
			18052: out = 16'(-7209);
			18053: out = 16'(-6244);
			18054: out = 16'(1661);
			18055: out = 16'(2108);
			18056: out = 16'(1974);
			18057: out = 16'(-6021);
			18058: out = 16'(-5368);
			18059: out = 16'(-3612);
			18060: out = 16'(2793);
			18061: out = 16'(3089);
			18062: out = 16'(1576);
			18063: out = 16'(-2170);
			18064: out = 16'(-2554);
			18065: out = 16'(92);
			18066: out = 16'(-72);
			18067: out = 16'(-1150);
			18068: out = 16'(-6612);
			18069: out = 16'(-1735);
			18070: out = 16'(1446);
			18071: out = 16'(5471);
			18072: out = 16'(2343);
			18073: out = 16'(-709);
			18074: out = 16'(-1635);
			18075: out = 16'(-4857);
			18076: out = 16'(-6847);
			18077: out = 16'(270);
			18078: out = 16'(2143);
			18079: out = 16'(3869);
			18080: out = 16'(-4021);
			18081: out = 16'(-3961);
			18082: out = 16'(-1677);
			18083: out = 16'(3387);
			18084: out = 16'(4875);
			18085: out = 16'(4665);
			18086: out = 16'(-879);
			18087: out = 16'(-2837);
			18088: out = 16'(25);
			18089: out = 16'(2766);
			18090: out = 16'(4296);
			18091: out = 16'(-423);
			18092: out = 16'(196);
			18093: out = 16'(-511);
			18094: out = 16'(-3734);
			18095: out = 16'(-4263);
			18096: out = 16'(-3220);
			18097: out = 16'(5143);
			18098: out = 16'(5518);
			18099: out = 16'(3221);
			18100: out = 16'(1549);
			18101: out = 16'(1506);
			18102: out = 16'(3808);
			18103: out = 16'(3276);
			18104: out = 16'(2623);
			18105: out = 16'(-883);
			18106: out = 16'(-817);
			18107: out = 16'(-1748);
			18108: out = 16'(62);
			18109: out = 16'(-3839);
			18110: out = 16'(-4542);
			18111: out = 16'(62);
			18112: out = 16'(4003);
			18113: out = 16'(6705);
			18114: out = 16'(3633);
			18115: out = 16'(843);
			18116: out = 16'(-2974);
			18117: out = 16'(-283);
			18118: out = 16'(719);
			18119: out = 16'(3632);
			18120: out = 16'(-5625);
			18121: out = 16'(-7475);
			18122: out = 16'(-6354);
			18123: out = 16'(-1146);
			18124: out = 16'(1471);
			18125: out = 16'(735);
			18126: out = 16'(933);
			18127: out = 16'(486);
			18128: out = 16'(12);
			18129: out = 16'(998);
			18130: out = 16'(1846);
			18131: out = 16'(849);
			18132: out = 16'(878);
			18133: out = 16'(353);
			18134: out = 16'(-5626);
			18135: out = 16'(-5314);
			18136: out = 16'(-2537);
			18137: out = 16'(97);
			18138: out = 16'(1488);
			18139: out = 16'(781);
			18140: out = 16'(2671);
			18141: out = 16'(1994);
			18142: out = 16'(0);
			18143: out = 16'(-172);
			18144: out = 16'(-40);
			18145: out = 16'(989);
			18146: out = 16'(901);
			18147: out = 16'(542);
			18148: out = 16'(-2228);
			18149: out = 16'(-1626);
			18150: out = 16'(-1298);
			18151: out = 16'(-2026);
			18152: out = 16'(-1852);
			18153: out = 16'(-610);
			18154: out = 16'(1166);
			18155: out = 16'(3641);
			18156: out = 16'(5145);
			18157: out = 16'(6190);
			18158: out = 16'(3991);
			18159: out = 16'(343);
			18160: out = 16'(-5438);
			18161: out = 16'(-6614);
			18162: out = 16'(-940);
			18163: out = 16'(498);
			18164: out = 16'(1202);
			18165: out = 16'(-5593);
			18166: out = 16'(-3046);
			18167: out = 16'(-1186);
			18168: out = 16'(6005);
			18169: out = 16'(4071);
			18170: out = 16'(2375);
			18171: out = 16'(-1121);
			18172: out = 16'(-520);
			18173: out = 16'(-23);
			18174: out = 16'(6606);
			18175: out = 16'(5062);
			18176: out = 16'(1277);
			18177: out = 16'(-7092);
			18178: out = 16'(-8308);
			18179: out = 16'(-2733);
			18180: out = 16'(780);
			18181: out = 16'(2548);
			18182: out = 16'(-465);
			18183: out = 16'(-2547);
			18184: out = 16'(-3641);
			18185: out = 16'(975);
			18186: out = 16'(3155);
			18187: out = 16'(5038);
			18188: out = 16'(128);
			18189: out = 16'(-1745);
			18190: out = 16'(-4522);
			18191: out = 16'(-1218);
			18192: out = 16'(-622);
			18193: out = 16'(1377);
			18194: out = 16'(-3609);
			18195: out = 16'(-2257);
			18196: out = 16'(1187);
			18197: out = 16'(4829);
			18198: out = 16'(4938);
			18199: out = 16'(246);
			18200: out = 16'(959);
			18201: out = 16'(1401);
			18202: out = 16'(5170);
			18203: out = 16'(3347);
			18204: out = 16'(1231);
			18205: out = 16'(-6094);
			18206: out = 16'(-5395);
			18207: out = 16'(-3226);
			18208: out = 16'(4986);
			18209: out = 16'(5235);
			18210: out = 16'(3644);
			18211: out = 16'(-574);
			18212: out = 16'(-1370);
			18213: out = 16'(-331);
			18214: out = 16'(2408);
			18215: out = 16'(2650);
			18216: out = 16'(287);
			18217: out = 16'(-2676);
			18218: out = 16'(-4966);
			18219: out = 16'(-3942);
			18220: out = 16'(-3358);
			18221: out = 16'(-2516);
			18222: out = 16'(-8741);
			18223: out = 16'(-3157);
			18224: out = 16'(1216);
			18225: out = 16'(6542);
			18226: out = 16'(3837);
			18227: out = 16'(-77);
			18228: out = 16'(-3473);
			18229: out = 16'(-3084);
			18230: out = 16'(-714);
			18231: out = 16'(1301);
			18232: out = 16'(1672);
			18233: out = 16'(557);
			18234: out = 16'(-2067);
			18235: out = 16'(-3198);
			18236: out = 16'(-2935);
			18237: out = 16'(405);
			18238: out = 16'(2437);
			18239: out = 16'(2782);
			18240: out = 16'(452);
			18241: out = 16'(-622);
			18242: out = 16'(4297);
			18243: out = 16'(5072);
			18244: out = 16'(5699);
			18245: out = 16'(3493);
			18246: out = 16'(1224);
			18247: out = 16'(-1952);
			18248: out = 16'(-61);
			18249: out = 16'(-626);
			18250: out = 16'(-378);
			18251: out = 16'(-3801);
			18252: out = 16'(-2775);
			18253: out = 16'(1106);
			18254: out = 16'(637);
			18255: out = 16'(913);
			18256: out = 16'(388);
			18257: out = 16'(645);
			18258: out = 16'(282);
			18259: out = 16'(763);
			18260: out = 16'(-1799);
			18261: out = 16'(-3004);
			18262: out = 16'(-223);
			18263: out = 16'(793);
			18264: out = 16'(1740);
			18265: out = 16'(-83);
			18266: out = 16'(940);
			18267: out = 16'(2662);
			18268: out = 16'(701);
			18269: out = 16'(-375);
			18270: out = 16'(-2630);
			18271: out = 16'(961);
			18272: out = 16'(1915);
			18273: out = 16'(3607);
			18274: out = 16'(-1503);
			18275: out = 16'(-3796);
			18276: out = 16'(-5596);
			18277: out = 16'(260);
			18278: out = 16'(3646);
			18279: out = 16'(2643);
			18280: out = 16'(-1106);
			18281: out = 16'(-4273);
			18282: out = 16'(-467);
			18283: out = 16'(2904);
			18284: out = 16'(6666);
			18285: out = 16'(2824);
			18286: out = 16'(592);
			18287: out = 16'(-2858);
			18288: out = 16'(-3047);
			18289: out = 16'(-2430);
			18290: out = 16'(773);
			18291: out = 16'(-1664);
			18292: out = 16'(-3408);
			18293: out = 16'(-7311);
			18294: out = 16'(-5081);
			18295: out = 16'(-3043);
			18296: out = 16'(88);
			18297: out = 16'(719);
			18298: out = 16'(1135);
			18299: out = 16'(67);
			18300: out = 16'(1127);
			18301: out = 16'(1624);
			18302: out = 16'(-2293);
			18303: out = 16'(-4309);
			18304: out = 16'(-5744);
			18305: out = 16'(-5);
			18306: out = 16'(2860);
			18307: out = 16'(5529);
			18308: out = 16'(1938);
			18309: out = 16'(960);
			18310: out = 16'(956);
			18311: out = 16'(2865);
			18312: out = 16'(3043);
			18313: out = 16'(928);
			18314: out = 16'(-945);
			18315: out = 16'(-2037);
			18316: out = 16'(654);
			18317: out = 16'(2005);
			18318: out = 16'(3609);
			18319: out = 16'(683);
			18320: out = 16'(974);
			18321: out = 16'(310);
			18322: out = 16'(3398);
			18323: out = 16'(1682);
			18324: out = 16'(-207);
			18325: out = 16'(-2991);
			18326: out = 16'(-1454);
			18327: out = 16'(2569);
			18328: out = 16'(2097);
			18329: out = 16'(-1104);
			18330: out = 16'(-9434);
			18331: out = 16'(-9526);
			18332: out = 16'(-6838);
			18333: out = 16'(3502);
			18334: out = 16'(4630);
			18335: out = 16'(4508);
			18336: out = 16'(-1758);
			18337: out = 16'(-3550);
			18338: out = 16'(-4699);
			18339: out = 16'(2916);
			18340: out = 16'(4531);
			18341: out = 16'(5919);
			18342: out = 16'(-2864);
			18343: out = 16'(-2719);
			18344: out = 16'(912);
			18345: out = 16'(194);
			18346: out = 16'(-1347);
			18347: out = 16'(-5250);
			18348: out = 16'(-3060);
			18349: out = 16'(-684);
			18350: out = 16'(2646);
			18351: out = 16'(4899);
			18352: out = 16'(5508);
			18353: out = 16'(1780);
			18354: out = 16'(660);
			18355: out = 16'(-342);
			18356: out = 16'(2445);
			18357: out = 16'(3497);
			18358: out = 16'(4851);
			18359: out = 16'(-918);
			18360: out = 16'(-2158);
			18361: out = 16'(-3569);
			18362: out = 16'(973);
			18363: out = 16'(1411);
			18364: out = 16'(1802);
			18365: out = 16'(-2440);
			18366: out = 16'(-2477);
			18367: out = 16'(-402);
			18368: out = 16'(4094);
			18369: out = 16'(4305);
			18370: out = 16'(-2259);
			18371: out = 16'(-6009);
			18372: out = 16'(-7959);
			18373: out = 16'(-1463);
			18374: out = 16'(-159);
			18375: out = 16'(1084);
			18376: out = 16'(886);
			18377: out = 16'(-1);
			18378: out = 16'(-1370);
			18379: out = 16'(-2198);
			18380: out = 16'(-118);
			18381: out = 16'(3905);
			18382: out = 16'(3945);
			18383: out = 16'(3330);
			18384: out = 16'(97);
			18385: out = 16'(-1226);
			18386: out = 16'(-3015);
			18387: out = 16'(-2886);
			18388: out = 16'(-4705);
			18389: out = 16'(-4700);
			18390: out = 16'(-3209);
			18391: out = 16'(-666);
			18392: out = 16'(1610);
			18393: out = 16'(1576);
			18394: out = 16'(3342);
			18395: out = 16'(4556);
			18396: out = 16'(6454);
			18397: out = 16'(4893);
			18398: out = 16'(1826);
			18399: out = 16'(-1993);
			18400: out = 16'(-4217);
			18401: out = 16'(-3929);
			18402: out = 16'(-5403);
			18403: out = 16'(-3316);
			18404: out = 16'(1014);
			18405: out = 16'(2795);
			18406: out = 16'(2483);
			18407: out = 16'(-3342);
			18408: out = 16'(-1322);
			18409: out = 16'(1004);
			18410: out = 16'(8026);
			18411: out = 16'(5499);
			18412: out = 16'(2093);
			18413: out = 16'(-5590);
			18414: out = 16'(-4479);
			18415: out = 16'(-808);
			18416: out = 16'(-3297);
			18417: out = 16'(-2592);
			18418: out = 16'(-2104);
			18419: out = 16'(1161);
			18420: out = 16'(1693);
			18421: out = 16'(574);
			18422: out = 16'(3294);
			18423: out = 16'(5475);
			18424: out = 16'(8769);
			18425: out = 16'(2804);
			18426: out = 16'(-1360);
			18427: out = 16'(-1051);
			18428: out = 16'(-1932);
			18429: out = 16'(-1978);
			18430: out = 16'(-9756);
			18431: out = 16'(-4595);
			18432: out = 16'(1118);
			18433: out = 16'(6557);
			18434: out = 16'(5476);
			18435: out = 16'(1826);
			18436: out = 16'(373);
			18437: out = 16'(357);
			18438: out = 16'(2707);
			18439: out = 16'(136);
			18440: out = 16'(-851);
			18441: out = 16'(-2581);
			18442: out = 16'(-2295);
			18443: out = 16'(-2110);
			18444: out = 16'(-256);
			18445: out = 16'(-2799);
			18446: out = 16'(-4743);
			18447: out = 16'(-6008);
			18448: out = 16'(-4180);
			18449: out = 16'(-730);
			18450: out = 16'(2705);
			18451: out = 16'(5271);
			18452: out = 16'(5375);
			18453: out = 16'(3561);
			18454: out = 16'(157);
			18455: out = 16'(-2298);
			18456: out = 16'(-8297);
			18457: out = 16'(-7382);
			18458: out = 16'(-2674);
			18459: out = 16'(829);
			18460: out = 16'(1324);
			18461: out = 16'(-1969);
			18462: out = 16'(-3309);
			18463: out = 16'(-2501);
			18464: out = 16'(2786);
			18465: out = 16'(6195);
			18466: out = 16'(8322);
			18467: out = 16'(6748);
			18468: out = 16'(2235);
			18469: out = 16'(-2938);
			18470: out = 16'(125);
			18471: out = 16'(678);
			18472: out = 16'(2714);
			18473: out = 16'(-4262);
			18474: out = 16'(-5554);
			18475: out = 16'(-6102);
			18476: out = 16'(-515);
			18477: out = 16'(1844);
			18478: out = 16'(2727);
			18479: out = 16'(1383);
			18480: out = 16'(422);
			18481: out = 16'(79);
			18482: out = 16'(1121);
			18483: out = 16'(1317);
			18484: out = 16'(-3206);
			18485: out = 16'(-1850);
			18486: out = 16'(-1448);
			18487: out = 16'(-3590);
			18488: out = 16'(-5034);
			18489: out = 16'(-5488);
			18490: out = 16'(-887);
			18491: out = 16'(1604);
			18492: out = 16'(3059);
			18493: out = 16'(4376);
			18494: out = 16'(3970);
			18495: out = 16'(2693);
			18496: out = 16'(862);
			18497: out = 16'(-754);
			18498: out = 16'(-3128);
			18499: out = 16'(-431);
			18500: out = 16'(930);
			18501: out = 16'(811);
			18502: out = 16'(-1425);
			18503: out = 16'(-2773);
			18504: out = 16'(748);
			18505: out = 16'(2112);
			18506: out = 16'(4215);
			18507: out = 16'(5362);
			18508: out = 16'(6439);
			18509: out = 16'(5988);
			18510: out = 16'(4735);
			18511: out = 16'(2003);
			18512: out = 16'(-782);
			18513: out = 16'(-1483);
			18514: out = 16'(-1090);
			18515: out = 16'(280);
			18516: out = 16'(-897);
			18517: out = 16'(-2546);
			18518: out = 16'(-5288);
			18519: out = 16'(-3211);
			18520: out = 16'(375);
			18521: out = 16'(5093);
			18522: out = 16'(6854);
			18523: out = 16'(5987);
			18524: out = 16'(2186);
			18525: out = 16'(-2341);
			18526: out = 16'(-5938);
			18527: out = 16'(-6695);
			18528: out = 16'(-3670);
			18529: out = 16'(1101);
			18530: out = 16'(-1088);
			18531: out = 16'(-2917);
			18532: out = 16'(-6487);
			18533: out = 16'(-1595);
			18534: out = 16'(911);
			18535: out = 16'(1481);
			18536: out = 16'(4785);
			18537: out = 16'(5022);
			18538: out = 16'(1710);
			18539: out = 16'(-1910);
			18540: out = 16'(-4065);
			18541: out = 16'(1741);
			18542: out = 16'(526);
			18543: out = 16'(-458);
			18544: out = 16'(-2975);
			18545: out = 16'(-2920);
			18546: out = 16'(-2140);
			18547: out = 16'(-3997);
			18548: out = 16'(-3320);
			18549: out = 16'(-1828);
			18550: out = 16'(2400);
			18551: out = 16'(3208);
			18552: out = 16'(566);
			18553: out = 16'(611);
			18554: out = 16'(-223);
			18555: out = 16'(1108);
			18556: out = 16'(-4452);
			18557: out = 16'(-6852);
			18558: out = 16'(-2809);
			18559: out = 16'(-1512);
			18560: out = 16'(171);
			18561: out = 16'(-4186);
			18562: out = 16'(164);
			18563: out = 16'(4384);
			18564: out = 16'(5865);
			18565: out = 16'(4234);
			18566: out = 16'(474);
			18567: out = 16'(2104);
			18568: out = 16'(659);
			18569: out = 16'(-1225);
			18570: out = 16'(-1925);
			18571: out = 16'(-1608);
			18572: out = 16'(309);
			18573: out = 16'(-1506);
			18574: out = 16'(-1711);
			18575: out = 16'(-143);
			18576: out = 16'(1099);
			18577: out = 16'(2370);
			18578: out = 16'(3400);
			18579: out = 16'(3527);
			18580: out = 16'(3558);
			18581: out = 16'(4869);
			18582: out = 16'(4593);
			18583: out = 16'(3576);
			18584: out = 16'(254);
			18585: out = 16'(-1677);
			18586: out = 16'(-2466);
			18587: out = 16'(-4939);
			18588: out = 16'(-4757);
			18589: out = 16'(-3130);
			18590: out = 16'(-322);
			18591: out = 16'(1535);
			18592: out = 16'(2547);
			18593: out = 16'(862);
			18594: out = 16'(-232);
			18595: out = 16'(928);
			18596: out = 16'(133);
			18597: out = 16'(5);
			18598: out = 16'(1578);
			18599: out = 16'(1077);
			18600: out = 16'(-134);
			18601: out = 16'(-5609);
			18602: out = 16'(-5295);
			18603: out = 16'(-2522);
			18604: out = 16'(-829);
			18605: out = 16'(1325);
			18606: out = 16'(2556);
			18607: out = 16'(2179);
			18608: out = 16'(771);
			18609: out = 16'(-1264);
			18610: out = 16'(-2010);
			18611: out = 16'(-1675);
			18612: out = 16'(689);
			18613: out = 16'(620);
			18614: out = 16'(46);
			18615: out = 16'(-4106);
			18616: out = 16'(-2498);
			18617: out = 16'(-292);
			18618: out = 16'(3908);
			18619: out = 16'(5163);
			18620: out = 16'(5625);
			18621: out = 16'(526);
			18622: out = 16'(-608);
			18623: out = 16'(-1462);
			18624: out = 16'(2049);
			18625: out = 16'(2069);
			18626: out = 16'(1721);
			18627: out = 16'(-3677);
			18628: out = 16'(-5176);
			18629: out = 16'(-4347);
			18630: out = 16'(2141);
			18631: out = 16'(4669);
			18632: out = 16'(-190);
			18633: out = 16'(-3451);
			18634: out = 16'(-5884);
			18635: out = 16'(1844);
			18636: out = 16'(2321);
			18637: out = 16'(3638);
			18638: out = 16'(-150);
			18639: out = 16'(237);
			18640: out = 16'(-381);
			18641: out = 16'(2580);
			18642: out = 16'(1499);
			18643: out = 16'(604);
			18644: out = 16'(-5162);
			18645: out = 16'(-4969);
			18646: out = 16'(-1070);
			18647: out = 16'(3254);
			18648: out = 16'(5090);
			18649: out = 16'(3173);
			18650: out = 16'(1140);
			18651: out = 16'(-935);
			18652: out = 16'(-218);
			18653: out = 16'(-1146);
			18654: out = 16'(-1177);
			18655: out = 16'(746);
			18656: out = 16'(-650);
			18657: out = 16'(-2742);
			18658: out = 16'(-5788);
			18659: out = 16'(-4010);
			18660: out = 16'(805);
			18661: out = 16'(-486);
			18662: out = 16'(1353);
			18663: out = 16'(2484);
			18664: out = 16'(3027);
			18665: out = 16'(781);
			18666: out = 16'(-4244);
			18667: out = 16'(-2239);
			18668: out = 16'(-667);
			18669: out = 16'(-465);
			18670: out = 16'(1182);
			18671: out = 16'(2038);
			18672: out = 16'(3570);
			18673: out = 16'(1882);
			18674: out = 16'(380);
			18675: out = 16'(-120);
			18676: out = 16'(1390);
			18677: out = 16'(3512);
			18678: out = 16'(1736);
			18679: out = 16'(933);
			18680: out = 16'(-415);
			18681: out = 16'(-175);
			18682: out = 16'(-84);
			18683: out = 16'(772);
			18684: out = 16'(469);
			18685: out = 16'(-410);
			18686: out = 16'(-3506);
			18687: out = 16'(-3222);
			18688: out = 16'(-2354);
			18689: out = 16'(3640);
			18690: out = 16'(1088);
			18691: out = 16'(-500);
			18692: out = 16'(-4446);
			18693: out = 16'(46);
			18694: out = 16'(4477);
			18695: out = 16'(1043);
			18696: out = 16'(-871);
			18697: out = 16'(-3652);
			18698: out = 16'(-3946);
			18699: out = 16'(-3937);
			18700: out = 16'(-2827);
			18701: out = 16'(608);
			18702: out = 16'(2488);
			18703: out = 16'(2544);
			18704: out = 16'(1040);
			18705: out = 16'(-513);
			18706: out = 16'(-988);
			18707: out = 16'(-813);
			18708: out = 16'(392);
			18709: out = 16'(2479);
			18710: out = 16'(2300);
			18711: out = 16'(1262);
			18712: out = 16'(-832);
			18713: out = 16'(-1861);
			18714: out = 16'(-2050);
			18715: out = 16'(-639);
			18716: out = 16'(321);
			18717: out = 16'(972);
			18718: out = 16'(1562);
			18719: out = 16'(1581);
			18720: out = 16'(698);
			18721: out = 16'(945);
			18722: out = 16'(986);
			18723: out = 16'(2843);
			18724: out = 16'(-2544);
			18725: out = 16'(-6151);
			18726: out = 16'(-8016);
			18727: out = 16'(-4380);
			18728: out = 16'(315);
			18729: out = 16'(2135);
			18730: out = 16'(2919);
			18731: out = 16'(1382);
			18732: out = 16'(2399);
			18733: out = 16'(1305);
			18734: out = 16'(2134);
			18735: out = 16'(-4544);
			18736: out = 16'(-3021);
			18737: out = 16'(103);
			18738: out = 16'(6150);
			18739: out = 16'(5343);
			18740: out = 16'(-430);
			18741: out = 16'(-5791);
			18742: out = 16'(-7218);
			18743: out = 16'(-967);
			18744: out = 16'(3472);
			18745: out = 16'(7338);
			18746: out = 16'(5435);
			18747: out = 16'(4411);
			18748: out = 16'(1771);
			18749: out = 16'(2852);
			18750: out = 16'(1099);
			18751: out = 16'(289);
			18752: out = 16'(-1441);
			18753: out = 16'(-1168);
			18754: out = 16'(-592);
			18755: out = 16'(-1295);
			18756: out = 16'(-1286);
			18757: out = 16'(-377);
			18758: out = 16'(-24);
			18759: out = 16'(1203);
			18760: out = 16'(3186);
			18761: out = 16'(3188);
			18762: out = 16'(2502);
			18763: out = 16'(-746);
			18764: out = 16'(-7);
			18765: out = 16'(-708);
			18766: out = 16'(-6890);
			18767: out = 16'(-7151);
			18768: out = 16'(-5645);
			18769: out = 16'(-3007);
			18770: out = 16'(-593);
			18771: out = 16'(710);
			18772: out = 16'(3229);
			18773: out = 16'(3263);
			18774: out = 16'(3529);
			18775: out = 16'(-2656);
			18776: out = 16'(-3609);
			18777: out = 16'(-1176);
			18778: out = 16'(4110);
			18779: out = 16'(6655);
			18780: out = 16'(4614);
			18781: out = 16'(1971);
			18782: out = 16'(-1560);
			18783: out = 16'(-3842);
			18784: out = 16'(-4779);
			18785: out = 16'(-3498);
			18786: out = 16'(975);
			18787: out = 16'(1844);
			18788: out = 16'(1429);
			18789: out = 16'(1610);
			18790: out = 16'(2055);
			18791: out = 16'(3159);
			18792: out = 16'(-1307);
			18793: out = 16'(-4173);
			18794: out = 16'(-7555);
			18795: out = 16'(-3632);
			18796: out = 16'(-1700);
			18797: out = 16'(-1345);
			18798: out = 16'(-551);
			18799: out = 16'(-91);
			18800: out = 16'(666);
			18801: out = 16'(751);
			18802: out = 16'(1125);
			18803: out = 16'(1525);
			18804: out = 16'(3106);
			18805: out = 16'(3975);
			18806: out = 16'(917);
			18807: out = 16'(-1599);
			18808: out = 16'(-4598);
			18809: out = 16'(-678);
			18810: out = 16'(-1146);
			18811: out = 16'(-2177);
			18812: out = 16'(-3197);
			18813: out = 16'(-1188);
			18814: out = 16'(3776);
			18815: out = 16'(2827);
			18816: out = 16'(1471);
			18817: out = 16'(-3444);
			18818: out = 16'(-584);
			18819: out = 16'(1980);
			18820: out = 16'(6364);
			18821: out = 16'(5203);
			18822: out = 16'(2846);
			18823: out = 16'(-4760);
			18824: out = 16'(-4263);
			18825: out = 16'(-1857);
			18826: out = 16'(-924);
			18827: out = 16'(-501);
			18828: out = 16'(-1574);
			18829: out = 16'(464);
			18830: out = 16'(60);
			18831: out = 16'(-224);
			18832: out = 16'(42);
			18833: out = 16'(1362);
			18834: out = 16'(2303);
			18835: out = 16'(3308);
			18836: out = 16'(2655);
			18837: out = 16'(1847);
			18838: out = 16'(-1103);
			18839: out = 16'(-2820);
			18840: out = 16'(-5662);
			18841: out = 16'(-618);
			18842: out = 16'(3718);
			18843: out = 16'(1609);
			18844: out = 16'(650);
			18845: out = 16'(-331);
			18846: out = 16'(3256);
			18847: out = 16'(5196);
			18848: out = 16'(5909);
			18849: out = 16'(6585);
			18850: out = 16'(3212);
			18851: out = 16'(-1926);
			18852: out = 16'(-7901);
			18853: out = 16'(-8427);
			18854: out = 16'(-1365);
			18855: out = 16'(816);
			18856: out = 16'(2197);
			18857: out = 16'(-465);
			18858: out = 16'(-2020);
			18859: out = 16'(-3385);
			18860: out = 16'(-427);
			18861: out = 16'(1744);
			18862: out = 16'(4268);
			18863: out = 16'(2299);
			18864: out = 16'(487);
			18865: out = 16'(-3363);
			18866: out = 16'(-3617);
			18867: out = 16'(-5671);
			18868: out = 16'(-6015);
			18869: out = 16'(-7525);
			18870: out = 16'(-4715);
			18871: out = 16'(845);
			18872: out = 16'(2739);
			18873: out = 16'(3849);
			18874: out = 16'(4336);
			18875: out = 16'(1988);
			18876: out = 16'(284);
			18877: out = 16'(871);
			18878: out = 16'(2021);
			18879: out = 16'(3087);
			18880: out = 16'(-2242);
			18881: out = 16'(-1829);
			18882: out = 16'(-1423);
			18883: out = 16'(-384);
			18884: out = 16'(-1246);
			18885: out = 16'(-2256);
			18886: out = 16'(-1429);
			18887: out = 16'(-1890);
			18888: out = 16'(-4339);
			18889: out = 16'(1777);
			18890: out = 16'(4459);
			18891: out = 16'(6754);
			18892: out = 16'(631);
			18893: out = 16'(-3145);
			18894: out = 16'(-4086);
			18895: out = 16'(-820);
			18896: out = 16'(2246);
			18897: out = 16'(560);
			18898: out = 16'(668);
			18899: out = 16'(-470);
			18900: out = 16'(-825);
			18901: out = 16'(-2259);
			18902: out = 16'(-2931);
			18903: out = 16'(-527);
			18904: out = 16'(827);
			18905: out = 16'(1885);
			18906: out = 16'(837);
			18907: out = 16'(1194);
			18908: out = 16'(2679);
			18909: out = 16'(3791);
			18910: out = 16'(2444);
			18911: out = 16'(-5701);
			18912: out = 16'(-1949);
			18913: out = 16'(303);
			18914: out = 16'(3523);
			18915: out = 16'(1114);
			18916: out = 16'(-166);
			18917: out = 16'(2092);
			18918: out = 16'(4470);
			18919: out = 16'(6017);
			18920: out = 16'(2249);
			18921: out = 16'(-1835);
			18922: out = 16'(-6889);
			18923: out = 16'(-3876);
			18924: out = 16'(-2169);
			18925: out = 16'(692);
			18926: out = 16'(-1705);
			18927: out = 16'(-2608);
			18928: out = 16'(-3183);
			18929: out = 16'(-2579);
			18930: out = 16'(-1459);
			18931: out = 16'(899);
			18932: out = 16'(917);
			18933: out = 16'(1013);
			18934: out = 16'(1776);
			18935: out = 16'(859);
			18936: out = 16'(-269);
			18937: out = 16'(-85);
			18938: out = 16'(-1999);
			18939: out = 16'(-4185);
			18940: out = 16'(115);
			18941: out = 16'(793);
			18942: out = 16'(1013);
			18943: out = 16'(-2301);
			18944: out = 16'(-2265);
			18945: out = 16'(308);
			18946: out = 16'(1225);
			18947: out = 16'(2046);
			18948: out = 16'(1724);
			18949: out = 16'(1306);
			18950: out = 16'(867);
			18951: out = 16'(1835);
			18952: out = 16'(1056);
			18953: out = 16'(286);
			18954: out = 16'(-1175);
			18955: out = 16'(-380);
			18956: out = 16'(1121);
			18957: out = 16'(490);
			18958: out = 16'(1693);
			18959: out = 16'(2272);
			18960: out = 16'(2746);
			18961: out = 16'(399);
			18962: out = 16'(-3391);
			18963: out = 16'(-4767);
			18964: out = 16'(-4004);
			18965: out = 16'(-123);
			18966: out = 16'(927);
			18967: out = 16'(2084);
			18968: out = 16'(2415);
			18969: out = 16'(981);
			18970: out = 16'(-1054);
			18971: out = 16'(-1887);
			18972: out = 16'(-2963);
			18973: out = 16'(-2597);
			18974: out = 16'(207);
			18975: out = 16'(3164);
			18976: out = 16'(5716);
			18977: out = 16'(1368);
			18978: out = 16'(-369);
			18979: out = 16'(-2464);
			18980: out = 16'(2259);
			18981: out = 16'(3240);
			18982: out = 16'(3204);
			18983: out = 16'(-264);
			18984: out = 16'(-1229);
			18985: out = 16'(666);
			18986: out = 16'(1624);
			18987: out = 16'(2093);
			18988: out = 16'(501);
			18989: out = 16'(17);
			18990: out = 16'(-529);
			18991: out = 16'(-1544);
			18992: out = 16'(-496);
			18993: out = 16'(730);
			18994: out = 16'(2178);
			18995: out = 16'(50);
			18996: out = 16'(-3891);
			18997: out = 16'(-3166);
			18998: out = 16'(-2548);
			18999: out = 16'(176);
			19000: out = 16'(-1357);
			19001: out = 16'(-1402);
			19002: out = 16'(-2560);
			19003: out = 16'(-1982);
			19004: out = 16'(-2117);
			19005: out = 16'(431);
			19006: out = 16'(-2284);
			19007: out = 16'(-2728);
			19008: out = 16'(-3644);
			19009: out = 16'(2487);
			19010: out = 16'(6299);
			19011: out = 16'(1556);
			19012: out = 16'(-3207);
			19013: out = 16'(-8191);
			19014: out = 16'(-2040);
			19015: out = 16'(894);
			19016: out = 16'(3674);
			19017: out = 16'(2917);
			19018: out = 16'(1636);
			19019: out = 16'(-223);
			19020: out = 16'(-3910);
			19021: out = 16'(-3337);
			19022: out = 16'(2927);
			19023: out = 16'(4577);
			19024: out = 16'(5257);
			19025: out = 16'(602);
			19026: out = 16'(473);
			19027: out = 16'(-332);
			19028: out = 16'(964);
			19029: out = 16'(-403);
			19030: out = 16'(-1577);
			19031: out = 16'(-3871);
			19032: out = 16'(-2554);
			19033: out = 16'(502);
			19034: out = 16'(-441);
			19035: out = 16'(649);
			19036: out = 16'(214);
			19037: out = 16'(1366);
			19038: out = 16'(-294);
			19039: out = 16'(-592);
			19040: out = 16'(-8658);
			19041: out = 16'(-9883);
			19042: out = 16'(-3959);
			19043: out = 16'(2510);
			19044: out = 16'(6578);
			19045: out = 16'(5130);
			19046: out = 16'(2556);
			19047: out = 16'(-819);
			19048: out = 16'(-5482);
			19049: out = 16'(-2847);
			19050: out = 16'(1996);
			19051: out = 16'(5206);
			19052: out = 16'(3985);
			19053: out = 16'(-568);
			19054: out = 16'(-619);
			19055: out = 16'(-260);
			19056: out = 16'(3107);
			19057: out = 16'(4571);
			19058: out = 16'(5763);
			19059: out = 16'(3517);
			19060: out = 16'(3330);
			19061: out = 16'(898);
			19062: out = 16'(-2012);
			19063: out = 16'(-2843);
			19064: out = 16'(-1689);
			19065: out = 16'(-169);
			19066: out = 16'(1735);
			19067: out = 16'(2383);
			19068: out = 16'(5508);
			19069: out = 16'(3091);
			19070: out = 16'(52);
			19071: out = 16'(-2876);
			19072: out = 16'(-3266);
			19073: out = 16'(-2481);
			19074: out = 16'(-1563);
			19075: out = 16'(-2133);
			19076: out = 16'(-3086);
			19077: out = 16'(-6295);
			19078: out = 16'(-5186);
			19079: out = 16'(1753);
			19080: out = 16'(4341);
			19081: out = 16'(4612);
			19082: out = 16'(-3057);
			19083: out = 16'(-4168);
			19084: out = 16'(-4448);
			19085: out = 16'(2191);
			19086: out = 16'(3336);
			19087: out = 16'(3881);
			19088: out = 16'(-2353);
			19089: out = 16'(-2611);
			19090: out = 16'(-832);
			19091: out = 16'(175);
			19092: out = 16'(1963);
			19093: out = 16'(3182);
			19094: out = 16'(4137);
			19095: out = 16'(2761);
			19096: out = 16'(-520);
			19097: out = 16'(-693);
			19098: out = 16'(280);
			19099: out = 16'(3039);
			19100: out = 16'(1822);
			19101: out = 16'(-202);
			19102: out = 16'(-935);
			19103: out = 16'(-2894);
			19104: out = 16'(-3300);
			19105: out = 16'(-8449);
			19106: out = 16'(-3975);
			19107: out = 16'(1105);
			19108: out = 16'(6050);
			19109: out = 16'(2263);
			19110: out = 16'(-5760);
			19111: out = 16'(-7367);
			19112: out = 16'(-5816);
			19113: out = 16'(627);
			19114: out = 16'(3662);
			19115: out = 16'(3837);
			19116: out = 16'(-3366);
			19117: out = 16'(-3337);
			19118: out = 16'(-2666);
			19119: out = 16'(5363);
			19120: out = 16'(3981);
			19121: out = 16'(3030);
			19122: out = 16'(-1020);
			19123: out = 16'(-551);
			19124: out = 16'(161);
			19125: out = 16'(1578);
			19126: out = 16'(1352);
			19127: out = 16'(478);
			19128: out = 16'(1624);
			19129: out = 16'(1565);
			19130: out = 16'(1686);
			19131: out = 16'(-686);
			19132: out = 16'(-1169);
			19133: out = 16'(-376);
			19134: out = 16'(1021);
			19135: out = 16'(1701);
			19136: out = 16'(1579);
			19137: out = 16'(394);
			19138: out = 16'(-998);
			19139: out = 16'(-3139);
			19140: out = 16'(-1657);
			19141: out = 16'(525);
			19142: out = 16'(2802);
			19143: out = 16'(3423);
			19144: out = 16'(2713);
			19145: out = 16'(-527);
			19146: out = 16'(-3756);
			19147: out = 16'(-7327);
			19148: out = 16'(-588);
			19149: out = 16'(805);
			19150: out = 16'(-135);
			19151: out = 16'(-2859);
			19152: out = 16'(-3449);
			19153: out = 16'(138);
			19154: out = 16'(248);
			19155: out = 16'(2009);
			19156: out = 16'(4730);
			19157: out = 16'(4263);
			19158: out = 16'(2523);
			19159: out = 16'(998);
			19160: out = 16'(-1244);
			19161: out = 16'(-2122);
			19162: out = 16'(-1727);
			19163: out = 16'(1127);
			19164: out = 16'(4197);
			19165: out = 16'(2003);
			19166: out = 16'(-411);
			19167: out = 16'(-4550);
			19168: out = 16'(-889);
			19169: out = 16'(136);
			19170: out = 16'(838);
			19171: out = 16'(-1979);
			19172: out = 16'(-2855);
			19173: out = 16'(-116);
			19174: out = 16'(150);
			19175: out = 16'(1075);
			19176: out = 16'(-461);
			19177: out = 16'(1661);
			19178: out = 16'(2098);
			19179: out = 16'(1108);
			19180: out = 16'(-2833);
			19181: out = 16'(-6057);
			19182: out = 16'(-2963);
			19183: out = 16'(916);
			19184: out = 16'(5239);
			19185: out = 16'(5029);
			19186: out = 16'(2429);
			19187: out = 16'(-3625);
			19188: out = 16'(-3722);
			19189: out = 16'(-3182);
			19190: out = 16'(1227);
			19191: out = 16'(-16);
			19192: out = 16'(10);
			19193: out = 16'(-1468);
			19194: out = 16'(697);
			19195: out = 16'(1566);
			19196: out = 16'(117);
			19197: out = 16'(-1101);
			19198: out = 16'(-1917);
			19199: out = 16'(2159);
			19200: out = 16'(2587);
			19201: out = 16'(2372);
			19202: out = 16'(104);
			19203: out = 16'(-542);
			19204: out = 16'(-339);
			19205: out = 16'(-197);
			19206: out = 16'(-96);
			19207: out = 16'(-139);
			19208: out = 16'(359);
			19209: out = 16'(202);
			19210: out = 16'(-1407);
			19211: out = 16'(-655);
			19212: out = 16'(-342);
			19213: out = 16'(48);
			19214: out = 16'(-815);
			19215: out = 16'(-959);
			19216: out = 16'(462);
			19217: out = 16'(2788);
			19218: out = 16'(4761);
			19219: out = 16'(242);
			19220: out = 16'(-1327);
			19221: out = 16'(-2270);
			19222: out = 16'(-134);
			19223: out = 16'(660);
			19224: out = 16'(272);
			19225: out = 16'(1468);
			19226: out = 16'(1174);
			19227: out = 16'(550);
			19228: out = 16'(-1528);
			19229: out = 16'(-2063);
			19230: out = 16'(-530);
			19231: out = 16'(105);
			19232: out = 16'(746);
			19233: out = 16'(3219);
			19234: out = 16'(1801);
			19235: out = 16'(-31);
			19236: out = 16'(-5596);
			19237: out = 16'(-6321);
			19238: out = 16'(-5776);
			19239: out = 16'(2763);
			19240: out = 16'(3513);
			19241: out = 16'(1428);
			19242: out = 16'(-3606);
			19243: out = 16'(-3902);
			19244: out = 16'(983);
			19245: out = 16'(2968);
			19246: out = 16'(3604);
			19247: out = 16'(-682);
			19248: out = 16'(-1847);
			19249: out = 16'(-3124);
			19250: out = 16'(937);
			19251: out = 16'(-1274);
			19252: out = 16'(-1661);
			19253: out = 16'(1328);
			19254: out = 16'(2271);
			19255: out = 16'(2342);
			19256: out = 16'(1057);
			19257: out = 16'(892);
			19258: out = 16'(1755);
			19259: out = 16'(-98);
			19260: out = 16'(174);
			19261: out = 16'(589);
			19262: out = 16'(1471);
			19263: out = 16'(1093);
			19264: out = 16'(524);
			19265: out = 16'(-2334);
			19266: out = 16'(-2322);
			19267: out = 16'(2383);
			19268: out = 16'(3326);
			19269: out = 16'(3121);
			19270: out = 16'(-3146);
			19271: out = 16'(-3378);
			19272: out = 16'(-2799);
			19273: out = 16'(1908);
			19274: out = 16'(2797);
			19275: out = 16'(3046);
			19276: out = 16'(682);
			19277: out = 16'(310);
			19278: out = 16'(573);
			19279: out = 16'(581);
			19280: out = 16'(-524);
			19281: out = 16'(-3668);
			19282: out = 16'(-601);
			19283: out = 16'(849);
			19284: out = 16'(2435);
			19285: out = 16'(-224);
			19286: out = 16'(-1453);
			19287: out = 16'(335);
			19288: out = 16'(428);
			19289: out = 16'(656);
			19290: out = 16'(1399);
			19291: out = 16'(405);
			19292: out = 16'(-740);
			19293: out = 16'(93);
			19294: out = 16'(1661);
			19295: out = 16'(3923);
			19296: out = 16'(-845);
			19297: out = 16'(-2338);
			19298: out = 16'(-3575);
			19299: out = 16'(-557);
			19300: out = 16'(265);
			19301: out = 16'(-381);
			19302: out = 16'(34);
			19303: out = 16'(910);
			19304: out = 16'(2994);
			19305: out = 16'(2623);
			19306: out = 16'(775);
			19307: out = 16'(-6089);
			19308: out = 16'(-6573);
			19309: out = 16'(-5766);
			19310: out = 16'(-1842);
			19311: out = 16'(-231);
			19312: out = 16'(898);
			19313: out = 16'(-98);
			19314: out = 16'(-26);
			19315: out = 16'(-71);
			19316: out = 16'(3308);
			19317: out = 16'(3932);
			19318: out = 16'(2994);
			19319: out = 16'(1233);
			19320: out = 16'(-433);
			19321: out = 16'(-1421);
			19322: out = 16'(-1549);
			19323: out = 16'(-1716);
			19324: out = 16'(-3347);
			19325: out = 16'(-2686);
			19326: out = 16'(-1561);
			19327: out = 16'(3144);
			19328: out = 16'(1980);
			19329: out = 16'(567);
			19330: out = 16'(1489);
			19331: out = 16'(1830);
			19332: out = 16'(2284);
			19333: out = 16'(-158);
			19334: out = 16'(-276);
			19335: out = 16'(745);
			19336: out = 16'(-1117);
			19337: out = 16'(-1213);
			19338: out = 16'(-517);
			19339: out = 16'(331);
			19340: out = 16'(630);
			19341: out = 16'(384);
			19342: out = 16'(-234);
			19343: out = 16'(-569);
			19344: out = 16'(-592);
			19345: out = 16'(198);
			19346: out = 16'(478);
			19347: out = 16'(-1190);
			19348: out = 16'(-2307);
			19349: out = 16'(-3215);
			19350: out = 16'(-1511);
			19351: out = 16'(-1213);
			19352: out = 16'(-1221);
			19353: out = 16'(235);
			19354: out = 16'(933);
			19355: out = 16'(1803);
			19356: out = 16'(-694);
			19357: out = 16'(-372);
			19358: out = 16'(2573);
			19359: out = 16'(4601);
			19360: out = 16'(3961);
			19361: out = 16'(-5581);
			19362: out = 16'(-2753);
			19363: out = 16'(-191);
			19364: out = 16'(7722);
			19365: out = 16'(3471);
			19366: out = 16'(-1405);
			19367: out = 16'(-6506);
			19368: out = 16'(-4370);
			19369: out = 16'(1441);
			19370: out = 16'(-325);
			19371: out = 16'(2536);
			19372: out = 16'(4607);
			19373: out = 16'(4967);
			19374: out = 16'(3212);
			19375: out = 16'(411);
			19376: out = 16'(367);
			19377: out = 16'(122);
			19378: out = 16'(-1909);
			19379: out = 16'(-256);
			19380: out = 16'(-47);
			19381: out = 16'(-156);
			19382: out = 16'(-1758);
			19383: out = 16'(-3044);
			19384: out = 16'(-9298);
			19385: out = 16'(-5915);
			19386: out = 16'(-1145);
			19387: out = 16'(6796);
			19388: out = 16'(5213);
			19389: out = 16'(-187);
			19390: out = 16'(-4695);
			19391: out = 16'(-4867);
			19392: out = 16'(704);
			19393: out = 16'(-740);
			19394: out = 16'(-810);
			19395: out = 16'(-4579);
			19396: out = 16'(-1134);
			19397: out = 16'(343);
			19398: out = 16'(3737);
			19399: out = 16'(1593);
			19400: out = 16'(601);
			19401: out = 16'(-2398);
			19402: out = 16'(118);
			19403: out = 16'(1869);
			19404: out = 16'(4260);
			19405: out = 16'(1160);
			19406: out = 16'(-2741);
			19407: out = 16'(-6456);
			19408: out = 16'(-4456);
			19409: out = 16'(1364);
			19410: out = 16'(3208);
			19411: out = 16'(3625);
			19412: out = 16'(73);
			19413: out = 16'(792);
			19414: out = 16'(1147);
			19415: out = 16'(5305);
			19416: out = 16'(1843);
			19417: out = 16'(165);
			19418: out = 16'(-2512);
			19419: out = 16'(-697);
			19420: out = 16'(366);
			19421: out = 16'(-111);
			19422: out = 16'(-472);
			19423: out = 16'(-675);
			19424: out = 16'(-4926);
			19425: out = 16'(-3621);
			19426: out = 16'(-774);
			19427: out = 16'(3796);
			19428: out = 16'(4894);
			19429: out = 16'(3785);
			19430: out = 16'(753);
			19431: out = 16'(649);
			19432: out = 16'(5071);
			19433: out = 16'(2763);
			19434: out = 16'(791);
			19435: out = 16'(-5710);
			19436: out = 16'(-2921);
			19437: out = 16'(-1212);
			19438: out = 16'(-303);
			19439: out = 16'(-34);
			19440: out = 16'(233);
			19441: out = 16'(-3340);
			19442: out = 16'(-1531);
			19443: out = 16'(763);
			19444: out = 16'(4299);
			19445: out = 16'(3240);
			19446: out = 16'(115);
			19447: out = 16'(-3208);
			19448: out = 16'(-3882);
			19449: out = 16'(-1029);
			19450: out = 16'(-998);
			19451: out = 16'(-937);
			19452: out = 16'(-4637);
			19453: out = 16'(-98);
			19454: out = 16'(2098);
			19455: out = 16'(3326);
			19456: out = 16'(690);
			19457: out = 16'(-2115);
			19458: out = 16'(-3774);
			19459: out = 16'(-3882);
			19460: out = 16'(-2609);
			19461: out = 16'(-1659);
			19462: out = 16'(-90);
			19463: out = 16'(603);
			19464: out = 16'(1916);
			19465: out = 16'(371);
			19466: out = 16'(-2220);
			19467: out = 16'(-4319);
			19468: out = 16'(-3746);
			19469: out = 16'(630);
			19470: out = 16'(-187);
			19471: out = 16'(1194);
			19472: out = 16'(3302);
			19473: out = 16'(5183);
			19474: out = 16'(4789);
			19475: out = 16'(-1006);
			19476: out = 16'(-2228);
			19477: out = 16'(-3078);
			19478: out = 16'(-184);
			19479: out = 16'(-2042);
			19480: out = 16'(-3839);
			19481: out = 16'(83);
			19482: out = 16'(1962);
			19483: out = 16'(3583);
			19484: out = 16'(2039);
			19485: out = 16'(1700);
			19486: out = 16'(1719);
			19487: out = 16'(2242);
			19488: out = 16'(2389);
			19489: out = 16'(1382);
			19490: out = 16'(2849);
			19491: out = 16'(2130);
			19492: out = 16'(-2228);
			19493: out = 16'(-4090);
			19494: out = 16'(-4099);
			19495: out = 16'(5389);
			19496: out = 16'(5019);
			19497: out = 16'(4303);
			19498: out = 16'(-2054);
			19499: out = 16'(-757);
			19500: out = 16'(1577);
			19501: out = 16'(2224);
			19502: out = 16'(844);
			19503: out = 16'(-1758);
			19504: out = 16'(-3085);
			19505: out = 16'(-2576);
			19506: out = 16'(-212);
			19507: out = 16'(1007);
			19508: out = 16'(518);
			19509: out = 16'(-3365);
			19510: out = 16'(-3985);
			19511: out = 16'(-3042);
			19512: out = 16'(3042);
			19513: out = 16'(4931);
			19514: out = 16'(5686);
			19515: out = 16'(-153);
			19516: out = 16'(-3568);
			19517: out = 16'(-7619);
			19518: out = 16'(-480);
			19519: out = 16'(100);
			19520: out = 16'(2024);
			19521: out = 16'(-7118);
			19522: out = 16'(-5212);
			19523: out = 16'(897);
			19524: out = 16'(6857);
			19525: out = 16'(6789);
			19526: out = 16'(76);
			19527: out = 16'(-1383);
			19528: out = 16'(-1630);
			19529: out = 16'(2378);
			19530: out = 16'(4326);
			19531: out = 16'(4431);
			19532: out = 16'(-2897);
			19533: out = 16'(-6496);
			19534: out = 16'(-8975);
			19535: out = 16'(-200);
			19536: out = 16'(1821);
			19537: out = 16'(3464);
			19538: out = 16'(738);
			19539: out = 16'(289);
			19540: out = 16'(-232);
			19541: out = 16'(1283);
			19542: out = 16'(1130);
			19543: out = 16'(-396);
			19544: out = 16'(-148);
			19545: out = 16'(-1304);
			19546: out = 16'(-3045);
			19547: out = 16'(-3989);
			19548: out = 16'(-3371);
			19549: out = 16'(-480);
			19550: out = 16'(-123);
			19551: out = 16'(52);
			19552: out = 16'(4310);
			19553: out = 16'(2329);
			19554: out = 16'(322);
			19555: out = 16'(-6388);
			19556: out = 16'(-4713);
			19557: out = 16'(-481);
			19558: out = 16'(3919);
			19559: out = 16'(5205);
			19560: out = 16'(4818);
			19561: out = 16'(-1230);
			19562: out = 16'(-3279);
			19563: out = 16'(-2123);
			19564: out = 16'(2663);
			19565: out = 16'(5143);
			19566: out = 16'(3966);
			19567: out = 16'(-247);
			19568: out = 16'(-3712);
			19569: out = 16'(-1138);
			19570: out = 16'(-93);
			19571: out = 16'(2142);
			19572: out = 16'(1955);
			19573: out = 16'(2641);
			19574: out = 16'(1715);
			19575: out = 16'(-2174);
			19576: out = 16'(-5110);
			19577: out = 16'(-7009);
			19578: out = 16'(-1870);
			19579: out = 16'(254);
			19580: out = 16'(-232);
			19581: out = 16'(658);
			19582: out = 16'(2169);
			19583: out = 16'(7449);
			19584: out = 16'(4260);
			19585: out = 16'(2327);
			19586: out = 16'(-1692);
			19587: out = 16'(-48);
			19588: out = 16'(201);
			19589: out = 16'(-18);
			19590: out = 16'(-5124);
			19591: out = 16'(-9367);
			19592: out = 16'(-3917);
			19593: out = 16'(61);
			19594: out = 16'(4789);
			19595: out = 16'(4520);
			19596: out = 16'(4007);
			19597: out = 16'(1047);
			19598: out = 16'(2494);
			19599: out = 16'(2370);
			19600: out = 16'(4258);
			19601: out = 16'(-1991);
			19602: out = 16'(-5241);
			19603: out = 16'(-7231);
			19604: out = 16'(-2534);
			19605: out = 16'(747);
			19606: out = 16'(-3484);
			19607: out = 16'(-1731);
			19608: out = 16'(-1020);
			19609: out = 16'(1841);
			19610: out = 16'(651);
			19611: out = 16'(-187);
			19612: out = 16'(-533);
			19613: out = 16'(740);
			19614: out = 16'(1550);
			19615: out = 16'(1304);
			19616: out = 16'(68);
			19617: out = 16'(-3);
			19618: out = 16'(-6984);
			19619: out = 16'(-8892);
			19620: out = 16'(-7964);
			19621: out = 16'(345);
			19622: out = 16'(5608);
			19623: out = 16'(5789);
			19624: out = 16'(2731);
			19625: out = 16'(155);
			19626: out = 16'(5015);
			19627: out = 16'(5601);
			19628: out = 16'(5830);
			19629: out = 16'(439);
			19630: out = 16'(-3797);
			19631: out = 16'(-8431);
			19632: out = 16'(-3894);
			19633: out = 16'(-247);
			19634: out = 16'(5625);
			19635: out = 16'(674);
			19636: out = 16'(232);
			19637: out = 16'(420);
			19638: out = 16'(3168);
			19639: out = 16'(3990);
			19640: out = 16'(3174);
			19641: out = 16'(1630);
			19642: out = 16'(203);
			19643: out = 16'(-415);
			19644: out = 16'(-635);
			19645: out = 16'(-889);
			19646: out = 16'(-3928);
			19647: out = 16'(-4692);
			19648: out = 16'(-4863);
			19649: out = 16'(-999);
			19650: out = 16'(938);
			19651: out = 16'(2795);
			19652: out = 16'(897);
			19653: out = 16'(1877);
			19654: out = 16'(4157);
			19655: out = 16'(3997);
			19656: out = 16'(3488);
			19657: out = 16'(2210);
			19658: out = 16'(615);
			19659: out = 16'(-1289);
			19660: out = 16'(-4243);
			19661: out = 16'(-3311);
			19662: out = 16'(-2335);
			19663: out = 16'(-4256);
			19664: out = 16'(-3161);
			19665: out = 16'(-1599);
			19666: out = 16'(1904);
			19667: out = 16'(3684);
			19668: out = 16'(4857);
			19669: out = 16'(3415);
			19670: out = 16'(2507);
			19671: out = 16'(1142);
			19672: out = 16'(-1929);
			19673: out = 16'(-4648);
			19674: out = 16'(-5964);
			19675: out = 16'(-6482);
			19676: out = 16'(-4890);
			19677: out = 16'(-2343);
			19678: out = 16'(1164);
			19679: out = 16'(2709);
			19680: out = 16'(1992);
			19681: out = 16'(-827);
			19682: out = 16'(-2748);
			19683: out = 16'(2217);
			19684: out = 16'(4406);
			19685: out = 16'(5906);
			19686: out = 16'(-4447);
			19687: out = 16'(-7647);
			19688: out = 16'(-8857);
			19689: out = 16'(-3596);
			19690: out = 16'(61);
			19691: out = 16'(2869);
			19692: out = 16'(2861);
			19693: out = 16'(2659);
			19694: out = 16'(2813);
			19695: out = 16'(1897);
			19696: out = 16'(2288);
			19697: out = 16'(3970);
			19698: out = 16'(5155);
			19699: out = 16'(4850);
			19700: out = 16'(1026);
			19701: out = 16'(-2400);
			19702: out = 16'(-5758);
			19703: out = 16'(-4039);
			19704: out = 16'(-3992);
			19705: out = 16'(-2808);
			19706: out = 16'(-5120);
			19707: out = 16'(-2673);
			19708: out = 16'(1409);
			19709: out = 16'(3522);
			19710: out = 16'(3659);
			19711: out = 16'(189);
			19712: out = 16'(1812);
			19713: out = 16'(1545);
			19714: out = 16'(2995);
			19715: out = 16'(-2466);
			19716: out = 16'(-5669);
			19717: out = 16'(-6976);
			19718: out = 16'(-3201);
			19719: out = 16'(552);
			19720: out = 16'(-386);
			19721: out = 16'(523);
			19722: out = 16'(1168);
			19723: out = 16'(4591);
			19724: out = 16'(5855);
			19725: out = 16'(6225);
			19726: out = 16'(4080);
			19727: out = 16'(1439);
			19728: out = 16'(-1495);
			19729: out = 16'(-4338);
			19730: out = 16'(-4138);
			19731: out = 16'(292);
			19732: out = 16'(257);
			19733: out = 16'(1102);
			19734: out = 16'(267);
			19735: out = 16'(1869);
			19736: out = 16'(2802);
			19737: out = 16'(4792);
			19738: out = 16'(4245);
			19739: out = 16'(3483);
			19740: out = 16'(-432);
			19741: out = 16'(212);
			19742: out = 16'(1284);
			19743: out = 16'(-227);
			19744: out = 16'(-3099);
			19745: out = 16'(-7497);
			19746: out = 16'(-3863);
			19747: out = 16'(-2332);
			19748: out = 16'(-161);
			19749: out = 16'(-589);
			19750: out = 16'(-123);
			19751: out = 16'(-596);
			19752: out = 16'(1649);
			19753: out = 16'(2884);
			19754: out = 16'(5645);
			19755: out = 16'(2429);
			19756: out = 16'(-998);
			19757: out = 16'(-8708);
			19758: out = 16'(-6302);
			19759: out = 16'(-1942);
			19760: out = 16'(3205);
			19761: out = 16'(3347);
			19762: out = 16'(1042);
			19763: out = 16'(-2904);
			19764: out = 16'(-3462);
			19765: out = 16'(-597);
			19766: out = 16'(1819);
			19767: out = 16'(4634);
			19768: out = 16'(5825);
			19769: out = 16'(4885);
			19770: out = 16'(2383);
			19771: out = 16'(-282);
			19772: out = 16'(-4242);
			19773: out = 16'(-6014);
			19774: out = 16'(-2134);
			19775: out = 16'(-1974);
			19776: out = 16'(-942);
			19777: out = 16'(-2590);
			19778: out = 16'(1053);
			19779: out = 16'(4263);
			19780: out = 16'(4035);
			19781: out = 16'(2187);
			19782: out = 16'(-807);
			19783: out = 16'(-1122);
			19784: out = 16'(-878);
			19785: out = 16'(505);
			19786: out = 16'(539);
			19787: out = 16'(-1111);
			19788: out = 16'(-6166);
			19789: out = 16'(-5868);
			19790: out = 16'(-4612);
			19791: out = 16'(1071);
			19792: out = 16'(3042);
			19793: out = 16'(5332);
			19794: out = 16'(1903);
			19795: out = 16'(4586);
			19796: out = 16'(5064);
			19797: out = 16'(6691);
			19798: out = 16'(1086);
			19799: out = 16'(-4800);
			19800: out = 16'(-8582);
			19801: out = 16'(-5789);
			19802: out = 16'(1301);
			19803: out = 16'(4677);
			19804: out = 16'(5514);
			19805: out = 16'(1761);
			19806: out = 16'(1193);
			19807: out = 16'(306);
			19808: out = 16'(2501);
			19809: out = 16'(1859);
			19810: out = 16'(1917);
			19811: out = 16'(-603);
			19812: out = 16'(-799);
			19813: out = 16'(-1881);
			19814: out = 16'(-300);
			19815: out = 16'(-2602);
			19816: out = 16'(-4328);
			19817: out = 16'(-5195);
			19818: out = 16'(-2857);
			19819: out = 16'(845);
			19820: out = 16'(-1160);
			19821: out = 16'(-1141);
			19822: out = 16'(-1262);
			19823: out = 16'(425);
			19824: out = 16'(427);
			19825: out = 16'(-1357);
			19826: out = 16'(-942);
			19827: out = 16'(-2175);
			19828: out = 16'(-5593);
			19829: out = 16'(-6440);
			19830: out = 16'(-4807);
			19831: out = 16'(5430);
			19832: out = 16'(5878);
			19833: out = 16'(5116);
			19834: out = 16'(-1394);
			19835: out = 16'(-1188);
			19836: out = 16'(462);
			19837: out = 16'(3410);
			19838: out = 16'(4004);
			19839: out = 16'(2959);
			19840: out = 16'(2765);
			19841: out = 16'(1157);
			19842: out = 16'(-1464);
			19843: out = 16'(-468);
			19844: out = 16'(283);
			19845: out = 16'(2527);
			19846: out = 16'(-701);
			19847: out = 16'(-2520);
			19848: out = 16'(-2234);
			19849: out = 16'(-192);
			19850: out = 16'(2126);
			19851: out = 16'(2758);
			19852: out = 16'(3257);
			19853: out = 16'(2674);
			19854: out = 16'(1745);
			19855: out = 16'(80);
			19856: out = 16'(-1678);
			19857: out = 16'(-638);
			19858: out = 16'(-1496);
			19859: out = 16'(-3383);
			19860: out = 16'(-2506);
			19861: out = 16'(-1582);
			19862: out = 16'(578);
			19863: out = 16'(270);
			19864: out = 16'(606);
			19865: out = 16'(545);
			19866: out = 16'(802);
			19867: out = 16'(316);
			19868: out = 16'(-264);
			19869: out = 16'(-1640);
			19870: out = 16'(-2034);
			19871: out = 16'(-594);
			19872: out = 16'(1739);
			19873: out = 16'(3920);
			19874: out = 16'(1020);
			19875: out = 16'(64);
			19876: out = 16'(-514);
			19877: out = 16'(209);
			19878: out = 16'(1385);
			19879: out = 16'(2956);
			19880: out = 16'(2441);
			19881: out = 16'(1501);
			19882: out = 16'(216);
			19883: out = 16'(-1563);
			19884: out = 16'(-3259);
			19885: out = 16'(-6187);
			19886: out = 16'(-5067);
			19887: out = 16'(-3422);
			19888: out = 16'(590);
			19889: out = 16'(-255);
			19890: out = 16'(-1166);
			19891: out = 16'(-729);
			19892: out = 16'(2231);
			19893: out = 16'(5650);
			19894: out = 16'(3516);
			19895: out = 16'(1452);
			19896: out = 16'(-1717);
			19897: out = 16'(-4175);
			19898: out = 16'(-4659);
			19899: out = 16'(-1858);
			19900: out = 16'(-978);
			19901: out = 16'(300);
			19902: out = 16'(-354);
			19903: out = 16'(149);
			19904: out = 16'(142);
			19905: out = 16'(3449);
			19906: out = 16'(1190);
			19907: out = 16'(-139);
			19908: out = 16'(270);
			19909: out = 16'(1424);
			19910: out = 16'(2235);
			19911: out = 16'(942);
			19912: out = 16'(20);
			19913: out = 16'(-466);
			19914: out = 16'(-2172);
			19915: out = 16'(-1384);
			19916: out = 16'(413);
			19917: out = 16'(3060);
			19918: out = 16'(3162);
			19919: out = 16'(489);
			19920: out = 16'(-1872);
			19921: out = 16'(-3137);
			19922: out = 16'(-398);
			19923: out = 16'(524);
			19924: out = 16'(1004);
			19925: out = 16'(-4960);
			19926: out = 16'(-4909);
			19927: out = 16'(-4686);
			19928: out = 16'(555);
			19929: out = 16'(-347);
			19930: out = 16'(-2063);
			19931: out = 16'(-589);
			19932: out = 16'(632);
			19933: out = 16'(1789);
			19934: out = 16'(3005);
			19935: out = 16'(3047);
			19936: out = 16'(2425);
			19937: out = 16'(-1356);
			19938: out = 16'(-3473);
			19939: out = 16'(-2819);
			19940: out = 16'(-964);
			19941: out = 16'(722);
			19942: out = 16'(-2382);
			19943: out = 16'(-1212);
			19944: out = 16'(-676);
			19945: out = 16'(5669);
			19946: out = 16'(3458);
			19947: out = 16'(1412);
			19948: out = 16'(-2891);
			19949: out = 16'(398);
			19950: out = 16'(5892);
			19951: out = 16'(4844);
			19952: out = 16'(1909);
			19953: out = 16'(-4759);
			19954: out = 16'(-1236);
			19955: out = 16'(-631);
			19956: out = 16'(-1505);
			19957: out = 16'(-440);
			19958: out = 16'(-33);
			19959: out = 16'(1843);
			19960: out = 16'(-2565);
			19961: out = 16'(-4608);
			19962: out = 16'(214);
			19963: out = 16'(3104);
			19964: out = 16'(5624);
			19965: out = 16'(3152);
			19966: out = 16'(1576);
			19967: out = 16'(-1009);
			19968: out = 16'(-393);
			19969: out = 16'(-360);
			19970: out = 16'(781);
			19971: out = 16'(-496);
			19972: out = 16'(-528);
			19973: out = 16'(-639);
			19974: out = 16'(324);
			19975: out = 16'(560);
			19976: out = 16'(587);
			19977: out = 16'(-187);
			19978: out = 16'(-367);
			19979: out = 16'(1445);
			19980: out = 16'(881);
			19981: out = 16'(-293);
			19982: out = 16'(-6635);
			19983: out = 16'(-6638);
			19984: out = 16'(-5466);
			19985: out = 16'(-195);
			19986: out = 16'(1169);
			19987: out = 16'(1761);
			19988: out = 16'(-95);
			19989: out = 16'(-434);
			19990: out = 16'(-1359);
			19991: out = 16'(5222);
			19992: out = 16'(7114);
			19993: out = 16'(7557);
			19994: out = 16'(-1142);
			19995: out = 16'(-6968);
			19996: out = 16'(-9984);
			19997: out = 16'(-5568);
			19998: out = 16'(-1119);
			19999: out = 16'(-1525);
			20000: out = 16'(-844);
			20001: out = 16'(-747);
			20002: out = 16'(2256);
			20003: out = 16'(4649);
			20004: out = 16'(7092);
			20005: out = 16'(4333);
			20006: out = 16'(1682);
			20007: out = 16'(-2825);
			20008: out = 16'(197);
			20009: out = 16'(279);
			20010: out = 16'(875);
			20011: out = 16'(-1700);
			20012: out = 16'(-1876);
			20013: out = 16'(-456);
			20014: out = 16'(359);
			20015: out = 16'(689);
			20016: out = 16'(451);
			20017: out = 16'(-137);
			20018: out = 16'(-336);
			20019: out = 16'(619);
			20020: out = 16'(707);
			20021: out = 16'(428);
			20022: out = 16'(-1000);
			20023: out = 16'(-2227);
			20024: out = 16'(-3133);
			20025: out = 16'(-3162);
			20026: out = 16'(-2070);
			20027: out = 16'(-86);
			20028: out = 16'(1163);
			20029: out = 16'(1637);
			20030: out = 16'(660);
			20031: out = 16'(724);
			20032: out = 16'(889);
			20033: out = 16'(3454);
			20034: out = 16'(1458);
			20035: out = 16'(143);
			20036: out = 16'(-3241);
			20037: out = 16'(-1100);
			20038: out = 16'(818);
			20039: out = 16'(2322);
			20040: out = 16'(1413);
			20041: out = 16'(221);
			20042: out = 16'(-2136);
			20043: out = 16'(-170);
			20044: out = 16'(3422);
			20045: out = 16'(1707);
			20046: out = 16'(287);
			20047: out = 16'(-2564);
			20048: out = 16'(-2239);
			20049: out = 16'(-1728);
			20050: out = 16'(614);
			20051: out = 16'(-90);
			20052: out = 16'(4);
			20053: out = 16'(370);
			20054: out = 16'(519);
			20055: out = 16'(-352);
			20056: out = 16'(-5748);
			20057: out = 16'(-4067);
			20058: out = 16'(-1369);
			20059: out = 16'(496);
			20060: out = 16'(667);
			20061: out = 16'(-203);
			20062: out = 16'(3574);
			20063: out = 16'(4573);
			20064: out = 16'(5516);
			20065: out = 16'(1415);
			20066: out = 16'(155);
			20067: out = 16'(392);
			20068: out = 16'(580);
			20069: out = 16'(1);
			20070: out = 16'(-2370);
			20071: out = 16'(-1227);
			20072: out = 16'(390);
			20073: out = 16'(3655);
			20074: out = 16'(3861);
			20075: out = 16'(3377);
			20076: out = 16'(1518);
			20077: out = 16'(667);
			20078: out = 16'(106);
			20079: out = 16'(340);
			20080: out = 16'(1003);
			20081: out = 16'(1984);
			20082: out = 16'(-2451);
			20083: out = 16'(-3677);
			20084: out = 16'(-3212);
			20085: out = 16'(-1405);
			20086: out = 16'(-1090);
			20087: out = 16'(-4655);
			20088: out = 16'(-66);
			20089: out = 16'(1957);
			20090: out = 16'(4090);
			20091: out = 16'(-963);
			20092: out = 16'(-4850);
			20093: out = 16'(-4847);
			20094: out = 16'(-3324);
			20095: out = 16'(-705);
			20096: out = 16'(-1546);
			20097: out = 16'(-217);
			20098: out = 16'(555);
			20099: out = 16'(82);
			20100: out = 16'(477);
			20101: out = 16'(1876);
			20102: out = 16'(2728);
			20103: out = 16'(2687);
			20104: out = 16'(-7);
			20105: out = 16'(428);
			20106: out = 16'(-763);
			20107: out = 16'(165);
			20108: out = 16'(-4998);
			20109: out = 16'(-5728);
			20110: out = 16'(153);
			20111: out = 16'(3922);
			20112: out = 16'(6101);
			20113: out = 16'(3386);
			20114: out = 16'(162);
			20115: out = 16'(-3608);
			20116: out = 16'(-1339);
			20117: out = 16'(-345);
			20118: out = 16'(1891);
			20119: out = 16'(395);
			20120: out = 16'(49);
			20121: out = 16'(-1651);
			20122: out = 16'(-404);
			20123: out = 16'(-369);
			20124: out = 16'(1044);
			20125: out = 16'(-2009);
			20126: out = 16'(-3893);
			20127: out = 16'(-8079);
			20128: out = 16'(-3000);
			20129: out = 16'(1349);
			20130: out = 16'(5462);
			20131: out = 16'(3175);
			20132: out = 16'(-304);
			20133: out = 16'(-4279);
			20134: out = 16'(-2781);
			20135: out = 16'(1385);
			20136: out = 16'(480);
			20137: out = 16'(933);
			20138: out = 16'(-495);
			20139: out = 16'(5187);
			20140: out = 16'(5840);
			20141: out = 16'(4531);
			20142: out = 16'(2364);
			20143: out = 16'(840);
			20144: out = 16'(392);
			20145: out = 16'(-1569);
			20146: out = 16'(-2201);
			20147: out = 16'(393);
			20148: out = 16'(-228);
			20149: out = 16'(7);
			20150: out = 16'(1052);
			20151: out = 16'(2675);
			20152: out = 16'(3650);
			20153: out = 16'(3066);
			20154: out = 16'(1351);
			20155: out = 16'(-809);
			20156: out = 16'(-2156);
			20157: out = 16'(-2397);
			20158: out = 16'(-1511);
			20159: out = 16'(-1577);
			20160: out = 16'(-2198);
			20161: out = 16'(-4398);
			20162: out = 16'(-2342);
			20163: out = 16'(-288);
			20164: out = 16'(3084);
			20165: out = 16'(1616);
			20166: out = 16'(3);
			20167: out = 16'(-1134);
			20168: out = 16'(-2131);
			20169: out = 16'(-2068);
			20170: out = 16'(-1760);
			20171: out = 16'(1222);
			20172: out = 16'(4083);
			20173: out = 16'(2424);
			20174: out = 16'(885);
			20175: out = 16'(-1765);
			20176: out = 16'(339);
			20177: out = 16'(717);
			20178: out = 16'(1480);
			20179: out = 16'(-38);
			20180: out = 16'(-180);
			20181: out = 16'(486);
			20182: out = 16'(503);
			20183: out = 16'(395);
			20184: out = 16'(285);
			20185: out = 16'(-841);
			20186: out = 16'(-1858);
			20187: out = 16'(-3263);
			20188: out = 16'(-1414);
			20189: out = 16'(1087);
			20190: out = 16'(1092);
			20191: out = 16'(594);
			20192: out = 16'(-2051);
			20193: out = 16'(238);
			20194: out = 16'(-2123);
			20195: out = 16'(-3861);
			20196: out = 16'(-7732);
			20197: out = 16'(-4510);
			20198: out = 16'(3585);
			20199: out = 16'(5550);
			20200: out = 16'(4312);
			20201: out = 16'(-3257);
			20202: out = 16'(-5295);
			20203: out = 16'(-6905);
			20204: out = 16'(-4638);
			20205: out = 16'(-2923);
			20206: out = 16'(-114);
			20207: out = 16'(640);
			20208: out = 16'(1403);
			20209: out = 16'(884);
			20210: out = 16'(1986);
			20211: out = 16'(2250);
			20212: out = 16'(3679);
			20213: out = 16'(266);
			20214: out = 16'(518);
			20215: out = 16'(654);
			20216: out = 16'(3062);
			20217: out = 16'(2152);
			20218: out = 16'(-219);
			20219: out = 16'(-3656);
			20220: out = 16'(-4639);
			20221: out = 16'(-3088);
			20222: out = 16'(1904);
			20223: out = 16'(5507);
			20224: out = 16'(4620);
			20225: out = 16'(2466);
			20226: out = 16'(-835);
			20227: out = 16'(131);
			20228: out = 16'(-1583);
			20229: out = 16'(-1972);
			20230: out = 16'(-1631);
			20231: out = 16'(69);
			20232: out = 16'(1693);
			20233: out = 16'(812);
			20234: out = 16'(-88);
			20235: out = 16'(-1274);
			20236: out = 16'(898);
			20237: out = 16'(1426);
			20238: out = 16'(-302);
			20239: out = 16'(450);
			20240: out = 16'(969);
			20241: out = 16'(4231);
			20242: out = 16'(806);
			20243: out = 16'(-1645);
			20244: out = 16'(-1252);
			20245: out = 16'(-503);
			20246: out = 16'(579);
			20247: out = 16'(-452);
			20248: out = 16'(99);
			20249: out = 16'(971);
			20250: out = 16'(3259);
			20251: out = 16'(4106);
			20252: out = 16'(3482);
			20253: out = 16'(3444);
			20254: out = 16'(1592);
			20255: out = 16'(-262);
			20256: out = 16'(-4700);
			20257: out = 16'(-5194);
			20258: out = 16'(469);
			20259: out = 16'(1348);
			20260: out = 16'(1992);
			20261: out = 16'(-1627);
			20262: out = 16'(-801);
			20263: out = 16'(-774);
			20264: out = 16'(-1197);
			20265: out = 16'(-1971);
			20266: out = 16'(-2092);
			20267: out = 16'(-808);
			20268: out = 16'(-237);
			20269: out = 16'(-618);
			20270: out = 16'(519);
			20271: out = 16'(-247);
			20272: out = 16'(-1204);
			20273: out = 16'(-2138);
			20274: out = 16'(-1491);
			20275: out = 16'(-195);
			20276: out = 16'(2252);
			20277: out = 16'(2687);
			20278: out = 16'(-63);
			20279: out = 16'(-1373);
			20280: out = 16'(-1870);
			20281: out = 16'(480);
			20282: out = 16'(3146);
			20283: out = 16'(5318);
			20284: out = 16'(134);
			20285: out = 16'(-1081);
			20286: out = 16'(-2370);
			20287: out = 16'(1056);
			20288: out = 16'(1108);
			20289: out = 16'(277);
			20290: out = 16'(-90);
			20291: out = 16'(-109);
			20292: out = 16'(682);
			20293: out = 16'(-1455);
			20294: out = 16'(-2337);
			20295: out = 16'(-1181);
			20296: out = 16'(-1557);
			20297: out = 16'(-450);
			20298: out = 16'(2889);
			20299: out = 16'(3668);
			20300: out = 16'(3037);
			20301: out = 16'(-2603);
			20302: out = 16'(-4672);
			20303: out = 16'(-6011);
			20304: out = 16'(-2489);
			20305: out = 16'(-2106);
			20306: out = 16'(-1876);
			20307: out = 16'(-1525);
			20308: out = 16'(515);
			20309: out = 16'(3482);
			20310: out = 16'(2673);
			20311: out = 16'(2551);
			20312: out = 16'(3314);
			20313: out = 16'(1293);
			20314: out = 16'(-261);
			20315: out = 16'(-3283);
			20316: out = 16'(193);
			20317: out = 16'(2890);
			20318: out = 16'(3766);
			20319: out = 16'(1849);
			20320: out = 16'(-695);
			20321: out = 16'(541);
			20322: out = 16'(-121);
			20323: out = 16'(-84);
			20324: out = 16'(1664);
			20325: out = 16'(2598);
			20326: out = 16'(2681);
			20327: out = 16'(339);
			20328: out = 16'(-2584);
			20329: out = 16'(-6361);
			20330: out = 16'(-4325);
			20331: out = 16'(-1195);
			20332: out = 16'(5621);
			20333: out = 16'(1685);
			20334: out = 16'(-1451);
			20335: out = 16'(-6059);
			20336: out = 16'(-2603);
			20337: out = 16'(991);
			20338: out = 16'(-423);
			20339: out = 16'(358);
			20340: out = 16'(318);
			20341: out = 16'(1);
			20342: out = 16'(11);
			20343: out = 16'(426);
			20344: out = 16'(-2507);
			20345: out = 16'(-2977);
			20346: out = 16'(-1891);
			20347: out = 16'(-2423);
			20348: out = 16'(-304);
			20349: out = 16'(4178);
			20350: out = 16'(4558);
			20351: out = 16'(3685);
			20352: out = 16'(-1493);
			20353: out = 16'(-679);
			20354: out = 16'(-500);
			20355: out = 16'(-3);
			20356: out = 16'(-1321);
			20357: out = 16'(-2120);
			20358: out = 16'(-646);
			20359: out = 16'(912);
			20360: out = 16'(2471);
			20361: out = 16'(-94);
			20362: out = 16'(-771);
			20363: out = 16'(-1372);
			20364: out = 16'(-224);
			20365: out = 16'(-692);
			20366: out = 16'(-2229);
			20367: out = 16'(-888);
			20368: out = 16'(261);
			20369: out = 16'(1631);
			20370: out = 16'(1091);
			20371: out = 16'(640);
			20372: out = 16'(809);
			20373: out = 16'(647);
			20374: out = 16'(693);
			20375: out = 16'(-497);
			20376: out = 16'(595);
			20377: out = 16'(1614);
			20378: out = 16'(1507);
			20379: out = 16'(793);
			20380: out = 16'(-436);
			20381: out = 16'(-1038);
			20382: out = 16'(-1801);
			20383: out = 16'(-2153);
			20384: out = 16'(-54);
			20385: out = 16'(1170);
			20386: out = 16'(1413);
			20387: out = 16'(1534);
			20388: out = 16'(1986);
			20389: out = 16'(4742);
			20390: out = 16'(3407);
			20391: out = 16'(2291);
			20392: out = 16'(-1632);
			20393: out = 16'(-833);
			20394: out = 16'(-188);
			20395: out = 16'(3619);
			20396: out = 16'(1880);
			20397: out = 16'(-251);
			20398: out = 16'(-3939);
			20399: out = 16'(-3660);
			20400: out = 16'(-2345);
			20401: out = 16'(1480);
			20402: out = 16'(1537);
			20403: out = 16'(281);
			20404: out = 16'(-5338);
			20405: out = 16'(-6013);
			20406: out = 16'(-1234);
			20407: out = 16'(2510);
			20408: out = 16'(5169);
			20409: out = 16'(5252);
			20410: out = 16'(992);
			20411: out = 16'(-3664);
			20412: out = 16'(-5776);
			20413: out = 16'(-3774);
			20414: out = 16'(178);
			20415: out = 16'(-2647);
			20416: out = 16'(-1130);
			20417: out = 16'(-530);
			20418: out = 16'(46);
			20419: out = 16'(-361);
			20420: out = 16'(-256);
			20421: out = 16'(-1161);
			20422: out = 16'(-1611);
			20423: out = 16'(-3248);
			20424: out = 16'(-1516);
			20425: out = 16'(-1010);
			20426: out = 16'(15);
			20427: out = 16'(-2093);
			20428: out = 16'(-2248);
			20429: out = 16'(715);
			20430: out = 16'(3978);
			20431: out = 16'(6197);
			20432: out = 16'(884);
			20433: out = 16'(895);
			20434: out = 16'(806);
			20435: out = 16'(4479);
			20436: out = 16'(3007);
			20437: out = 16'(-115);
			20438: out = 16'(-1560);
			20439: out = 16'(-2928);
			20440: out = 16'(-2935);
			20441: out = 16'(-4073);
			20442: out = 16'(-2885);
			20443: out = 16'(13);
			20444: out = 16'(1646);
			20445: out = 16'(2563);
			20446: out = 16'(1473);
			20447: out = 16'(2136);
			20448: out = 16'(2562);
			20449: out = 16'(3842);
			20450: out = 16'(3084);
			20451: out = 16'(1420);
			20452: out = 16'(-3357);
			20453: out = 16'(-5679);
			20454: out = 16'(-6746);
			20455: out = 16'(-2165);
			20456: out = 16'(-868);
			20457: out = 16'(-1271);
			20458: out = 16'(1208);
			20459: out = 16'(2317);
			20460: out = 16'(4294);
			20461: out = 16'(-595);
			20462: out = 16'(-1603);
			20463: out = 16'(1740);
			20464: out = 16'(2074);
			20465: out = 16'(1210);
			20466: out = 16'(-6058);
			20467: out = 16'(-3826);
			20468: out = 16'(-1298);
			20469: out = 16'(2191);
			20470: out = 16'(1444);
			20471: out = 16'(-228);
			20472: out = 16'(2443);
			20473: out = 16'(1927);
			20474: out = 16'(1585);
			20475: out = 16'(-975);
			20476: out = 16'(-607);
			20477: out = 16'(761);
			20478: out = 16'(1415);
			20479: out = 16'(1153);
			20480: out = 16'(505);
			20481: out = 16'(-2150);
			20482: out = 16'(-2717);
			20483: out = 16'(-450);
			20484: out = 16'(1340);
			20485: out = 16'(2307);
			20486: out = 16'(774);
			20487: out = 16'(-843);
			20488: out = 16'(-2104);
			20489: out = 16'(1300);
			20490: out = 16'(2568);
			20491: out = 16'(3812);
			20492: out = 16'(-788);
			20493: out = 16'(-1547);
			20494: out = 16'(-1357);
			20495: out = 16'(-1379);
			20496: out = 16'(-1777);
			20497: out = 16'(-3301);
			20498: out = 16'(-336);
			20499: out = 16'(204);
			20500: out = 16'(-1260);
			20501: out = 16'(-626);
			20502: out = 16'(1215);
			20503: out = 16'(5908);
			20504: out = 16'(6209);
			20505: out = 16'(5054);
			20506: out = 16'(1031);
			20507: out = 16'(-2510);
			20508: out = 16'(-5366);
			20509: out = 16'(-934);
			20510: out = 16'(-136);
			20511: out = 16'(630);
			20512: out = 16'(-2735);
			20513: out = 16'(-2086);
			20514: out = 16'(727);
			20515: out = 16'(-479);
			20516: out = 16'(-267);
			20517: out = 16'(-618);
			20518: out = 16'(2241);
			20519: out = 16'(2841);
			20520: out = 16'(1465);
			20521: out = 16'(-1248);
			20522: out = 16'(-4155);
			20523: out = 16'(-6520);
			20524: out = 16'(-6068);
			20525: out = 16'(-3917);
			20526: out = 16'(-848);
			20527: out = 16'(1139);
			20528: out = 16'(1839);
			20529: out = 16'(3357);
			20530: out = 16'(2299);
			20531: out = 16'(406);
			20532: out = 16'(-716);
			20533: out = 16'(-1227);
			20534: out = 16'(-1006);
			20535: out = 16'(141);
			20536: out = 16'(403);
			20537: out = 16'(-1235);
			20538: out = 16'(-977);
			20539: out = 16'(-325);
			20540: out = 16'(4305);
			20541: out = 16'(1411);
			20542: out = 16'(-88);
			20543: out = 16'(-483);
			20544: out = 16'(2288);
			20545: out = 16'(4971);
			20546: out = 16'(5100);
			20547: out = 16'(3997);
			20548: out = 16'(1649);
			20549: out = 16'(233);
			20550: out = 16'(-723);
			20551: out = 16'(-492);
			20552: out = 16'(-1405);
			20553: out = 16'(-1411);
			20554: out = 16'(-1450);
			20555: out = 16'(-850);
			20556: out = 16'(96);
			20557: out = 16'(2204);
			20558: out = 16'(2098);
			20559: out = 16'(1887);
			20560: out = 16'(441);
			20561: out = 16'(108);
			20562: out = 16'(-805);
			20563: out = 16'(-1913);
			20564: out = 16'(-4166);
			20565: out = 16'(-5856);
			20566: out = 16'(-2717);
			20567: out = 16'(-591);
			20568: out = 16'(1746);
			20569: out = 16'(82);
			20570: out = 16'(-366);
			20571: out = 16'(-1331);
			20572: out = 16'(945);
			20573: out = 16'(1731);
			20574: out = 16'(2401);
			20575: out = 16'(-685);
			20576: out = 16'(-2059);
			20577: out = 16'(608);
			20578: out = 16'(-203);
			20579: out = 16'(-464);
			20580: out = 16'(-1310);
			20581: out = 16'(-769);
			20582: out = 16'(-332);
			20583: out = 16'(-375);
			20584: out = 16'(-53);
			20585: out = 16'(679);
			20586: out = 16'(1220);
			20587: out = 16'(2175);
			20588: out = 16'(2889);
			20589: out = 16'(1371);
			20590: out = 16'(-925);
			20591: out = 16'(-3989);
			20592: out = 16'(-4742);
			20593: out = 16'(-3353);
			20594: out = 16'(2628);
			20595: out = 16'(765);
			20596: out = 16'(-942);
			20597: out = 16'(-5773);
			20598: out = 16'(-2628);
			20599: out = 16'(557);
			20600: out = 16'(-222);
			20601: out = 16'(-184);
			20602: out = 16'(-1025);
			20603: out = 16'(4381);
			20604: out = 16'(3984);
			20605: out = 16'(2915);
			20606: out = 16'(-4216);
			20607: out = 16'(-5267);
			20608: out = 16'(-2499);
			20609: out = 16'(-510);
			20610: out = 16'(1050);
			20611: out = 16'(374);
			20612: out = 16'(2499);
			20613: out = 16'(3591);
			20614: out = 16'(4567);
			20615: out = 16'(4185);
			20616: out = 16'(3344);
			20617: out = 16'(2367);
			20618: out = 16'(719);
			20619: out = 16'(-443);
			20620: out = 16'(414);
			20621: out = 16'(137);
			20622: out = 16'(-524);
			20623: out = 16'(363);
			20624: out = 16'(-603);
			20625: out = 16'(-1396);
			20626: out = 16'(-2479);
			20627: out = 16'(-618);
			20628: out = 16'(2982);
			20629: out = 16'(4601);
			20630: out = 16'(3845);
			20631: out = 16'(-904);
			20632: out = 16'(-1702);
			20633: out = 16'(-2719);
			20634: out = 16'(-2222);
			20635: out = 16'(-3445);
			20636: out = 16'(-3818);
			20637: out = 16'(-226);
			20638: out = 16'(-1632);
			20639: out = 16'(-3287);
			20640: out = 16'(-4750);
			20641: out = 16'(-3039);
			20642: out = 16'(317);
			20643: out = 16'(2372);
			20644: out = 16'(4192);
			20645: out = 16'(5206);
			20646: out = 16'(-235);
			20647: out = 16'(-2770);
			20648: out = 16'(-1813);
			20649: out = 16'(-2410);
			20650: out = 16'(-2105);
			20651: out = 16'(-4231);
			20652: out = 16'(270);
			20653: out = 16'(2806);
			20654: out = 16'(2347);
			20655: out = 16'(1585);
			20656: out = 16'(917);
			20657: out = 16'(4437);
			20658: out = 16'(4164);
			20659: out = 16'(3232);
			20660: out = 16'(-2186);
			20661: out = 16'(-3807);
			20662: out = 16'(-3932);
			20663: out = 16'(-2588);
			20664: out = 16'(-2195);
			20665: out = 16'(-3078);
			20666: out = 16'(-71);
			20667: out = 16'(1369);
			20668: out = 16'(2429);
			20669: out = 16'(1330);
			20670: out = 16'(456);
			20671: out = 16'(-309);
			20672: out = 16'(-827);
			20673: out = 16'(-1451);
			20674: out = 16'(-1919);
			20675: out = 16'(-1753);
			20676: out = 16'(-893);
			20677: out = 16'(-2217);
			20678: out = 16'(-599);
			20679: out = 16'(724);
			20680: out = 16'(3102);
			20681: out = 16'(2242);
			20682: out = 16'(797);
			20683: out = 16'(-3035);
			20684: out = 16'(-2544);
			20685: out = 16'(1030);
			20686: out = 16'(4150);
			20687: out = 16'(4624);
			20688: out = 16'(258);
			20689: out = 16'(-1068);
			20690: out = 16'(-1773);
			20691: out = 16'(2553);
			20692: out = 16'(1229);
			20693: out = 16'(632);
			20694: out = 16'(453);
			20695: out = 16'(-407);
			20696: out = 16'(-1375);
			20697: out = 16'(-527);
			20698: out = 16'(1234);
			20699: out = 16'(4182);
			20700: out = 16'(1530);
			20701: out = 16'(1311);
			20702: out = 16'(-18);
			20703: out = 16'(3317);
			20704: out = 16'(1991);
			20705: out = 16'(-2351);
			20706: out = 16'(-5444);
			20707: out = 16'(-5755);
			20708: out = 16'(662);
			20709: out = 16'(1332);
			20710: out = 16'(2174);
			20711: out = 16'(-2466);
			20712: out = 16'(83);
			20713: out = 16'(1828);
			20714: out = 16'(5853);
			20715: out = 16'(2549);
			20716: out = 16'(-1934);
			20717: out = 16'(-1262);
			20718: out = 16'(-913);
			20719: out = 16'(451);
			20720: out = 16'(-1140);
			20721: out = 16'(-1112);
			20722: out = 16'(-65);
			20723: out = 16'(-1825);
			20724: out = 16'(-1596);
			20725: out = 16'(357);
			20726: out = 16'(3009);
			20727: out = 16'(5064);
			20728: out = 16'(6339);
			20729: out = 16'(3163);
			20730: out = 16'(-981);
			20731: out = 16'(-4424);
			20732: out = 16'(-5153);
			20733: out = 16'(-3887);
			20734: out = 16'(-7822);
			20735: out = 16'(-5970);
			20736: out = 16'(-3394);
			20737: out = 16'(2098);
			20738: out = 16'(2968);
			20739: out = 16'(1412);
			20740: out = 16'(-1012);
			20741: out = 16'(-1607);
			20742: out = 16'(1202);
			20743: out = 16'(29);
			20744: out = 16'(-639);
			20745: out = 16'(-5074);
			20746: out = 16'(-1155);
			20747: out = 16'(604);
			20748: out = 16'(-849);
			20749: out = 16'(-2473);
			20750: out = 16'(-3317);
			20751: out = 16'(-251);
			20752: out = 16'(2972);
			20753: out = 16'(6587);
			20754: out = 16'(3309);
			20755: out = 16'(3339);
			20756: out = 16'(2815);
			20757: out = 16'(2181);
			20758: out = 16'(-167);
			20759: out = 16'(-3006);
			20760: out = 16'(-3177);
			20761: out = 16'(-2029);
			20762: out = 16'(490);
			20763: out = 16'(300);
			20764: out = 16'(-283);
			20765: out = 16'(-30);
			20766: out = 16'(-1088);
			20767: out = 16'(-444);
			20768: out = 16'(1826);
			20769: out = 16'(4228);
			20770: out = 16'(4958);
			20771: out = 16'(4414);
			20772: out = 16'(176);
			20773: out = 16'(-4431);
			20774: out = 16'(-7353);
			20775: out = 16'(-4956);
			20776: out = 16'(1362);
			20777: out = 16'(1848);
			20778: out = 16'(1694);
			20779: out = 16'(-1397);
			20780: out = 16'(-570);
			20781: out = 16'(323);
			20782: out = 16'(2225);
			20783: out = 16'(4596);
			20784: out = 16'(5574);
			20785: out = 16'(3033);
			20786: out = 16'(135);
			20787: out = 16'(-2791);
			20788: out = 16'(-1349);
			20789: out = 16'(-840);
			20790: out = 16'(522);
			20791: out = 16'(168);
			20792: out = 16'(-532);
			20793: out = 16'(-2482);
			20794: out = 16'(1452);
			20795: out = 16'(2660);
			20796: out = 16'(3712);
			20797: out = 16'(1020);
			20798: out = 16'(243);
			20799: out = 16'(1307);
			20800: out = 16'(578);
			20801: out = 16'(-1420);
			20802: out = 16'(-9010);
			20803: out = 16'(-7190);
			20804: out = 16'(-4996);
			20805: out = 16'(309);
			20806: out = 16'(-1141);
			20807: out = 16'(-3108);
			20808: out = 16'(-2801);
			20809: out = 16'(-1756);
			20810: out = 16'(332);
			20811: out = 16'(3137);
			20812: out = 16'(5690);
			20813: out = 16'(8054);
			20814: out = 16'(2238);
			20815: out = 16'(-2078);
			20816: out = 16'(-8095);
			20817: out = 16'(-1601);
			20818: out = 16'(1087);
			20819: out = 16'(574);
			20820: out = 16'(-3324);
			20821: out = 16'(-5305);
			20822: out = 16'(124);
			20823: out = 16'(2022);
			20824: out = 16'(4205);
			20825: out = 16'(-184);
			20826: out = 16'(1021);
			20827: out = 16'(1566);
			20828: out = 16'(3924);
			20829: out = 16'(1803);
			20830: out = 16'(-1618);
			20831: out = 16'(-2625);
			20832: out = 16'(-2063);
			20833: out = 16'(1150);
			20834: out = 16'(-2176);
			20835: out = 16'(-3305);
			20836: out = 16'(-4902);
			20837: out = 16'(130);
			20838: out = 16'(3797);
			20839: out = 16'(6612);
			20840: out = 16'(4805);
			20841: out = 16'(1613);
			20842: out = 16'(-4246);
			20843: out = 16'(-5613);
			20844: out = 16'(-5133);
			20845: out = 16'(237);
			20846: out = 16'(962);
			20847: out = 16'(450);
			20848: out = 16'(-1591);
			20849: out = 16'(-1303);
			20850: out = 16'(446);
			20851: out = 16'(4598);
			20852: out = 16'(6566);
			20853: out = 16'(5509);
			20854: out = 16'(5294);
			20855: out = 16'(3036);
			20856: out = 16'(795);
			20857: out = 16'(-3194);
			20858: out = 16'(-5394);
			20859: out = 16'(-4927);
			20860: out = 16'(-3552);
			20861: out = 16'(-1470);
			20862: out = 16'(47);
			20863: out = 16'(1607);
			20864: out = 16'(2314);
			20865: out = 16'(1665);
			20866: out = 16'(788);
			20867: out = 16'(-317);
			20868: out = 16'(577);
			20869: out = 16'(253);
			20870: out = 16'(-516);
			20871: out = 16'(-1133);
			20872: out = 16'(-1098);
			20873: out = 16'(-88);
			20874: out = 16'(-854);
			20875: out = 16'(-1981);
			20876: out = 16'(-4849);
			20877: out = 16'(-2714);
			20878: out = 16'(-185);
			20879: out = 16'(2074);
			20880: out = 16'(3091);
			20881: out = 16'(2735);
			20882: out = 16'(1017);
			20883: out = 16'(-1652);
			20884: out = 16'(-3948);
			20885: out = 16'(-1567);
			20886: out = 16'(-301);
			20887: out = 16'(974);
			20888: out = 16'(718);
			20889: out = 16'(1690);
			20890: out = 16'(4100);
			20891: out = 16'(147);
			20892: out = 16'(-2037);
			20893: out = 16'(-3953);
			20894: out = 16'(-840);
			20895: out = 16'(1177);
			20896: out = 16'(638);
			20897: out = 16'(782);
			20898: out = 16'(365);
			20899: out = 16'(104);
			20900: out = 16'(-1026);
			20901: out = 16'(-2042);
			20902: out = 16'(702);
			20903: out = 16'(597);
			20904: out = 16'(495);
			20905: out = 16'(-4911);
			20906: out = 16'(-4244);
			20907: out = 16'(-614);
			20908: out = 16'(2069);
			20909: out = 16'(4531);
			20910: out = 16'(6821);
			20911: out = 16'(2445);
			20912: out = 16'(-524);
			20913: out = 16'(-2080);
			20914: out = 16'(-422);
			20915: out = 16'(813);
			20916: out = 16'(-212);
			20917: out = 16'(-598);
			20918: out = 16'(-1941);
			20919: out = 16'(-7119);
			20920: out = 16'(-6464);
			20921: out = 16'(-3507);
			20922: out = 16'(5280);
			20923: out = 16'(7399);
			20924: out = 16'(6253);
			20925: out = 16'(1476);
			20926: out = 16'(-516);
			20927: out = 16'(846);
			20928: out = 16'(97);
			20929: out = 16'(362);
			20930: out = 16'(-1713);
			20931: out = 16'(1490);
			20932: out = 16'(1733);
			20933: out = 16'(90);
			20934: out = 16'(-3037);
			20935: out = 16'(-4540);
			20936: out = 16'(-220);
			20937: out = 16'(326);
			20938: out = 16'(878);
			20939: out = 16'(496);
			20940: out = 16'(498);
			20941: out = 16'(304);
			20942: out = 16'(-2358);
			20943: out = 16'(-3404);
			20944: out = 16'(-3665);
			20945: out = 16'(-1161);
			20946: out = 16'(1046);
			20947: out = 16'(3343);
			20948: out = 16'(3154);
			20949: out = 16'(2925);
			20950: out = 16'(1352);
			20951: out = 16'(1769);
			20952: out = 16'(723);
			20953: out = 16'(-807);
			20954: out = 16'(-4082);
			20955: out = 16'(-5502);
			20956: out = 16'(-2509);
			20957: out = 16'(351);
			20958: out = 16'(2536);
			20959: out = 16'(1175);
			20960: out = 16'(-706);
			20961: out = 16'(-2873);
			20962: out = 16'(-3041);
			20963: out = 16'(-182);
			20964: out = 16'(5173);
			20965: out = 16'(4681);
			20966: out = 16'(3544);
			20967: out = 16'(-310);
			20968: out = 16'(-669);
			20969: out = 16'(-1393);
			20970: out = 16'(-1075);
			20971: out = 16'(-576);
			20972: out = 16'(209);
			20973: out = 16'(457);
			20974: out = 16'(185);
			20975: out = 16'(-511);
			20976: out = 16'(-967);
			20977: out = 16'(-1573);
			20978: out = 16'(-1877);
			20979: out = 16'(1234);
			20980: out = 16'(1105);
			20981: out = 16'(-410);
			20982: out = 16'(-239);
			20983: out = 16'(259);
			20984: out = 16'(1772);
			20985: out = 16'(804);
			20986: out = 16'(570);
			20987: out = 16'(813);
			20988: out = 16'(1202);
			20989: out = 16'(1297);
			20990: out = 16'(-1367);
			20991: out = 16'(-140);
			20992: out = 16'(690);
			20993: out = 16'(3137);
			20994: out = 16'(1720);
			20995: out = 16'(359);
			20996: out = 16'(-4521);
			20997: out = 16'(-2316);
			20998: out = 16'(2045);
			20999: out = 16'(4616);
			21000: out = 16'(3153);
			21001: out = 16'(-2893);
			21002: out = 16'(-1799);
			21003: out = 16'(-2303);
			21004: out = 16'(-907);
			21005: out = 16'(-1621);
			21006: out = 16'(25);
			21007: out = 16'(3665);
			21008: out = 16'(3084);
			21009: out = 16'(1572);
			21010: out = 16'(93);
			21011: out = 16'(-580);
			21012: out = 16'(-638);
			21013: out = 16'(-4845);
			21014: out = 16'(-2889);
			21015: out = 16'(0);
			21016: out = 16'(1244);
			21017: out = 16'(1040);
			21018: out = 16'(-282);
			21019: out = 16'(-272);
			21020: out = 16'(-303);
			21021: out = 16'(-106);
			21022: out = 16'(1045);
			21023: out = 16'(1543);
			21024: out = 16'(1500);
			21025: out = 16'(-269);
			21026: out = 16'(-1327);
			21027: out = 16'(-98);
			21028: out = 16'(224);
			21029: out = 16'(487);
			21030: out = 16'(-2051);
			21031: out = 16'(-1746);
			21032: out = 16'(-913);
			21033: out = 16'(1119);
			21034: out = 16'(1707);
			21035: out = 16'(1242);
			21036: out = 16'(363);
			21037: out = 16'(-817);
			21038: out = 16'(-1018);
			21039: out = 16'(-2286);
			21040: out = 16'(-895);
			21041: out = 16'(1367);
			21042: out = 16'(2862);
			21043: out = 16'(2158);
			21044: out = 16'(-106);
			21045: out = 16'(-3970);
			21046: out = 16'(-5592);
			21047: out = 16'(-3365);
			21048: out = 16'(1158);
			21049: out = 16'(5024);
			21050: out = 16'(3115);
			21051: out = 16'(1593);
			21052: out = 16'(-1019);
			21053: out = 16'(-4152);
			21054: out = 16'(-4473);
			21055: out = 16'(-2522);
			21056: out = 16'(1116);
			21057: out = 16'(3016);
			21058: out = 16'(2952);
			21059: out = 16'(1302);
			21060: out = 16'(414);
			21061: out = 16'(1615);
			21062: out = 16'(2803);
			21063: out = 16'(3596);
			21064: out = 16'(1149);
			21065: out = 16'(572);
			21066: out = 16'(-682);
			21067: out = 16'(809);
			21068: out = 16'(-1133);
			21069: out = 16'(-2416);
			21070: out = 16'(-3259);
			21071: out = 16'(-1680);
			21072: out = 16'(581);
			21073: out = 16'(-200);
			21074: out = 16'(-191);
			21075: out = 16'(-231);
			21076: out = 16'(-210);
			21077: out = 16'(-205);
			21078: out = 16'(-257);
			21079: out = 16'(-83);
			21080: out = 16'(-977);
			21081: out = 16'(-3965);
			21082: out = 16'(-3424);
			21083: out = 16'(-2015);
			21084: out = 16'(2245);
			21085: out = 16'(2460);
			21086: out = 16'(2085);
			21087: out = 16'(93);
			21088: out = 16'(-641);
			21089: out = 16'(-1309);
			21090: out = 16'(-443);
			21091: out = 16'(13);
			21092: out = 16'(905);
			21093: out = 16'(-326);
			21094: out = 16'(0);
			21095: out = 16'(398);
			21096: out = 16'(3637);
			21097: out = 16'(4301);
			21098: out = 16'(2831);
			21099: out = 16'(1278);
			21100: out = 16'(-498);
			21101: out = 16'(-2259);
			21102: out = 16'(-1179);
			21103: out = 16'(-212);
			21104: out = 16'(-1424);
			21105: out = 16'(-1769);
			21106: out = 16'(-2048);
			21107: out = 16'(1284);
			21108: out = 16'(674);
			21109: out = 16'(-666);
			21110: out = 16'(-1107);
			21111: out = 16'(-889);
			21112: out = 16'(574);
			21113: out = 16'(-4618);
			21114: out = 16'(-5937);
			21115: out = 16'(-5620);
			21116: out = 16'(-443);
			21117: out = 16'(2222);
			21118: out = 16'(561);
			21119: out = 16'(1730);
			21120: out = 16'(1714);
			21121: out = 16'(3528);
			21122: out = 16'(163);
			21123: out = 16'(-2143);
			21124: out = 16'(-7);
			21125: out = 16'(626);
			21126: out = 16'(1699);
			21127: out = 16'(-1962);
			21128: out = 16'(92);
			21129: out = 16'(3585);
			21130: out = 16'(3528);
			21131: out = 16'(3549);
			21132: out = 16'(1884);
			21133: out = 16'(4254);
			21134: out = 16'(2596);
			21135: out = 16'(-2605);
			21136: out = 16'(-575);
			21137: out = 16'(847);
			21138: out = 16'(2870);
			21139: out = 16'(277);
			21140: out = 16'(-1791);
			21141: out = 16'(490);
			21142: out = 16'(-415);
			21143: out = 16'(-563);
			21144: out = 16'(-6035);
			21145: out = 16'(-3181);
			21146: out = 16'(387);
			21147: out = 16'(5833);
			21148: out = 16'(4048);
			21149: out = 16'(-1209);
			21150: out = 16'(-2424);
			21151: out = 16'(-2620);
			21152: out = 16'(101);
			21153: out = 16'(-554);
			21154: out = 16'(-1312);
			21155: out = 16'(-5172);
			21156: out = 16'(-1937);
			21157: out = 16'(943);
			21158: out = 16'(5153);
			21159: out = 16'(4514);
			21160: out = 16'(2921);
			21161: out = 16'(-41);
			21162: out = 16'(-2910);
			21163: out = 16'(-5026);
			21164: out = 16'(-1620);
			21165: out = 16'(-789);
			21166: out = 16'(-19);
			21167: out = 16'(-266);
			21168: out = 16'(223);
			21169: out = 16'(668);
			21170: out = 16'(705);
			21171: out = 16'(406);
			21172: out = 16'(-163);
			21173: out = 16'(-386);
			21174: out = 16'(-31);
			21175: out = 16'(1444);
			21176: out = 16'(2001);
			21177: out = 16'(928);
			21178: out = 16'(-7545);
			21179: out = 16'(-7125);
			21180: out = 16'(-5634);
			21181: out = 16'(2697);
			21182: out = 16'(2916);
			21183: out = 16'(2159);
			21184: out = 16'(-4752);
			21185: out = 16'(-4602);
			21186: out = 16'(-2416);
			21187: out = 16'(3562);
			21188: out = 16'(3812);
			21189: out = 16'(406);
			21190: out = 16'(-3171);
			21191: out = 16'(-3811);
			21192: out = 16'(434);
			21193: out = 16'(3524);
			21194: out = 16'(5329);
			21195: out = 16'(467);
			21196: out = 16'(708);
			21197: out = 16'(71);
			21198: out = 16'(4926);
			21199: out = 16'(2258);
			21200: out = 16'(-19);
			21201: out = 16'(-4496);
			21202: out = 16'(-3025);
			21203: out = 16'(150);
			21204: out = 16'(1098);
			21205: out = 16'(2034);
			21206: out = 16'(2279);
			21207: out = 16'(1772);
			21208: out = 16'(715);
			21209: out = 16'(-1422);
			21210: out = 16'(203);
			21211: out = 16'(782);
			21212: out = 16'(1645);
			21213: out = 16'(-1953);
			21214: out = 16'(-3809);
			21215: out = 16'(-313);
			21216: out = 16'(549);
			21217: out = 16'(1396);
			21218: out = 16'(-2795);
			21219: out = 16'(-3226);
			21220: out = 16'(-3659);
			21221: out = 16'(1954);
			21222: out = 16'(1735);
			21223: out = 16'(454);
			21224: out = 16'(-3076);
			21225: out = 16'(-2271);
			21226: out = 16'(2152);
			21227: out = 16'(635);
			21228: out = 16'(1012);
			21229: out = 16'(1555);
			21230: out = 16'(1733);
			21231: out = 16'(600);
			21232: out = 16'(-3918);
			21233: out = 16'(-1623);
			21234: out = 16'(304);
			21235: out = 16'(-202);
			21236: out = 16'(28);
			21237: out = 16'(-343);
			21238: out = 16'(948);
			21239: out = 16'(-64);
			21240: out = 16'(-1145);
			21241: out = 16'(-446);
			21242: out = 16'(474);
			21243: out = 16'(1733);
			21244: out = 16'(294);
			21245: out = 16'(-129);
			21246: out = 16'(-285);
			21247: out = 16'(495);
			21248: out = 16'(841);
			21249: out = 16'(480);
			21250: out = 16'(231);
			21251: out = 16'(-56);
			21252: out = 16'(884);
			21253: out = 16'(65);
			21254: out = 16'(-186);
			21255: out = 16'(609);
			21256: out = 16'(1552);
			21257: out = 16'(2285);
			21258: out = 16'(675);
			21259: out = 16'(118);
			21260: out = 16'(-148);
			21261: out = 16'(-432);
			21262: out = 16'(-279);
			21263: out = 16'(-139);
			21264: out = 16'(2756);
			21265: out = 16'(3997);
			21266: out = 16'(3487);
			21267: out = 16'(3249);
			21268: out = 16'(2147);
			21269: out = 16'(476);
			21270: out = 16'(-295);
			21271: out = 16'(-855);
			21272: out = 16'(-650);
			21273: out = 16'(-1207);
			21274: out = 16'(-1498);
			21275: out = 16'(-780);
			21276: out = 16'(-268);
			21277: out = 16'(122);
			21278: out = 16'(-1997);
			21279: out = 16'(-2160);
			21280: out = 16'(-1200);
			21281: out = 16'(-34);
			21282: out = 16'(860);
			21283: out = 16'(245);
			21284: out = 16'(2533);
			21285: out = 16'(1981);
			21286: out = 16'(-173);
			21287: out = 16'(-4052);
			21288: out = 16'(-5532);
			21289: out = 16'(-415);
			21290: out = 16'(26);
			21291: out = 16'(782);
			21292: out = 16'(-579);
			21293: out = 16'(38);
			21294: out = 16'(487);
			21295: out = 16'(2090);
			21296: out = 16'(1882);
			21297: out = 16'(1202);
			21298: out = 16'(-69);
			21299: out = 16'(-1542);
			21300: out = 16'(-3211);
			21301: out = 16'(-3128);
			21302: out = 16'(-2224);
			21303: out = 16'(697);
			21304: out = 16'(-372);
			21305: out = 16'(169);
			21306: out = 16'(1284);
			21307: out = 16'(3928);
			21308: out = 16'(4712);
			21309: out = 16'(678);
			21310: out = 16'(-1294);
			21311: out = 16'(-3400);
			21312: out = 16'(-133);
			21313: out = 16'(-950);
			21314: out = 16'(-1398);
			21315: out = 16'(-5549);
			21316: out = 16'(-4168);
			21317: out = 16'(-804);
			21318: out = 16'(1607);
			21319: out = 16'(1946);
			21320: out = 16'(-396);
			21321: out = 16'(1305);
			21322: out = 16'(1069);
			21323: out = 16'(-365);
			21324: out = 16'(-408);
			21325: out = 16'(157);
			21326: out = 16'(3109);
			21327: out = 16'(1007);
			21328: out = 16'(-847);
			21329: out = 16'(-1983);
			21330: out = 16'(-1172);
			21331: out = 16'(82);
			21332: out = 16'(-247);
			21333: out = 16'(198);
			21334: out = 16'(531);
			21335: out = 16'(1262);
			21336: out = 16'(1544);
			21337: out = 16'(1277);
			21338: out = 16'(1542);
			21339: out = 16'(948);
			21340: out = 16'(731);
			21341: out = 16'(-2067);
			21342: out = 16'(-2778);
			21343: out = 16'(-1307);
			21344: out = 16'(386);
			21345: out = 16'(2026);
			21346: out = 16'(4279);
			21347: out = 16'(2753);
			21348: out = 16'(333);
			21349: out = 16'(-5227);
			21350: out = 16'(-5166);
			21351: out = 16'(-3080);
			21352: out = 16'(3233);
			21353: out = 16'(4706);
			21354: out = 16'(3952);
			21355: out = 16'(-1533);
			21356: out = 16'(-2617);
			21357: out = 16'(846);
			21358: out = 16'(-1334);
			21359: out = 16'(-892);
			21360: out = 16'(-720);
			21361: out = 16'(1507);
			21362: out = 16'(1432);
			21363: out = 16'(-2195);
			21364: out = 16'(-611);
			21365: out = 16'(1265);
			21366: out = 16'(3266);
			21367: out = 16'(3370);
			21368: out = 16'(2410);
			21369: out = 16'(3067);
			21370: out = 16'(653);
			21371: out = 16'(-1872);
			21372: out = 16'(-5355);
			21373: out = 16'(-4299);
			21374: out = 16'(-13);
			21375: out = 16'(-668);
			21376: out = 16'(213);
			21377: out = 16'(82);
			21378: out = 16'(2296);
			21379: out = 16'(2459);
			21380: out = 16'(1295);
			21381: out = 16'(-438);
			21382: out = 16'(-1701);
			21383: out = 16'(-1321);
			21384: out = 16'(-1490);
			21385: out = 16'(-1442);
			21386: out = 16'(-2126);
			21387: out = 16'(-3319);
			21388: out = 16'(-4852);
			21389: out = 16'(-1420);
			21390: out = 16'(-263);
			21391: out = 16'(1969);
			21392: out = 16'(-2625);
			21393: out = 16'(-679);
			21394: out = 16'(3127);
			21395: out = 16'(5413);
			21396: out = 16'(3540);
			21397: out = 16'(-3198);
			21398: out = 16'(-4731);
			21399: out = 16'(-5479);
			21400: out = 16'(-3677);
			21401: out = 16'(-1240);
			21402: out = 16'(1402);
			21403: out = 16'(2942);
			21404: out = 16'(2058);
			21405: out = 16'(576);
			21406: out = 16'(1559);
			21407: out = 16'(2404);
			21408: out = 16'(3820);
			21409: out = 16'(724);
			21410: out = 16'(347);
			21411: out = 16'(341);
			21412: out = 16'(7);
			21413: out = 16'(-744);
			21414: out = 16'(-2189);
			21415: out = 16'(-632);
			21416: out = 16'(413);
			21417: out = 16'(2374);
			21418: out = 16'(-58);
			21419: out = 16'(-1791);
			21420: out = 16'(-3853);
			21421: out = 16'(-1671);
			21422: out = 16'(529);
			21423: out = 16'(2835);
			21424: out = 16'(1949);
			21425: out = 16'(290);
			21426: out = 16'(-1634);
			21427: out = 16'(-2446);
			21428: out = 16'(-2798);
			21429: out = 16'(923);
			21430: out = 16'(1539);
			21431: out = 16'(1595);
			21432: out = 16'(-3956);
			21433: out = 16'(-4896);
			21434: out = 16'(-1687);
			21435: out = 16'(2425);
			21436: out = 16'(5026);
			21437: out = 16'(3476);
			21438: out = 16'(2230);
			21439: out = 16'(-7);
			21440: out = 16'(66);
			21441: out = 16'(-1189);
			21442: out = 16'(-790);
			21443: out = 16'(214);
			21444: out = 16'(2237);
			21445: out = 16'(3531);
			21446: out = 16'(919);
			21447: out = 16'(-462);
			21448: out = 16'(-1286);
			21449: out = 16'(-63);
			21450: out = 16'(73);
			21451: out = 16'(-1561);
			21452: out = 16'(877);
			21453: out = 16'(1304);
			21454: out = 16'(1519);
			21455: out = 16'(-1488);
			21456: out = 16'(-3539);
			21457: out = 16'(-4682);
			21458: out = 16'(-3698);
			21459: out = 16'(-2296);
			21460: out = 16'(377);
			21461: out = 16'(682);
			21462: out = 16'(781);
			21463: out = 16'(-2661);
			21464: out = 16'(-836);
			21465: out = 16'(1842);
			21466: out = 16'(3687);
			21467: out = 16'(1410);
			21468: out = 16'(-4108);
			21469: out = 16'(-2329);
			21470: out = 16'(-531);
			21471: out = 16'(3279);
			21472: out = 16'(1659);
			21473: out = 16'(-957);
			21474: out = 16'(-7129);
			21475: out = 16'(-6396);
			21476: out = 16'(-3773);
			21477: out = 16'(1984);
			21478: out = 16'(4769);
			21479: out = 16'(5883);
			21480: out = 16'(5025);
			21481: out = 16'(1549);
			21482: out = 16'(-2250);
			21483: out = 16'(276);
			21484: out = 16'(731);
			21485: out = 16'(682);
			21486: out = 16'(2137);
			21487: out = 16'(2067);
			21488: out = 16'(2478);
			21489: out = 16'(-3048);
			21490: out = 16'(-3907);
			21491: out = 16'(-361);
			21492: out = 16'(3321);
			21493: out = 16'(4654);
			21494: out = 16'(656);
			21495: out = 16'(-2347);
			21496: out = 16'(-5118);
			21497: out = 16'(-2848);
			21498: out = 16'(-1835);
			21499: out = 16'(138);
			21500: out = 16'(467);
			21501: out = 16'(910);
			21502: out = 16'(678);
			21503: out = 16'(1389);
			21504: out = 16'(1787);
			21505: out = 16'(2192);
			21506: out = 16'(2822);
			21507: out = 16'(2373);
			21508: out = 16'(1364);
			21509: out = 16'(-1783);
			21510: out = 16'(-2691);
			21511: out = 16'(436);
			21512: out = 16'(1328);
			21513: out = 16'(1886);
			21514: out = 16'(-1468);
			21515: out = 16'(-806);
			21516: out = 16'(-509);
			21517: out = 16'(325);
			21518: out = 16'(-140);
			21519: out = 16'(-361);
			21520: out = 16'(1726);
			21521: out = 16'(2716);
			21522: out = 16'(3443);
			21523: out = 16'(207);
			21524: out = 16'(-1144);
			21525: out = 16'(-1404);
			21526: out = 16'(-947);
			21527: out = 16'(-480);
			21528: out = 16'(-720);
			21529: out = 16'(58);
			21530: out = 16'(-221);
			21531: out = 16'(-2262);
			21532: out = 16'(-1765);
			21533: out = 16'(-1101);
			21534: out = 16'(-332);
			21535: out = 16'(-239);
			21536: out = 16'(-727);
			21537: out = 16'(-1865);
			21538: out = 16'(-2273);
			21539: out = 16'(-1982);
			21540: out = 16'(-3701);
			21541: out = 16'(-2752);
			21542: out = 16'(-889);
			21543: out = 16'(1023);
			21544: out = 16'(1588);
			21545: out = 16'(675);
			21546: out = 16'(1472);
			21547: out = 16'(1183);
			21548: out = 16'(-355);
			21549: out = 16'(-1267);
			21550: out = 16'(-1873);
			21551: out = 16'(1170);
			21552: out = 16'(-1455);
			21553: out = 16'(-2656);
			21554: out = 16'(-2277);
			21555: out = 16'(783);
			21556: out = 16'(3344);
			21557: out = 16'(3292);
			21558: out = 16'(1312);
			21559: out = 16'(-1282);
			21560: out = 16'(-1317);
			21561: out = 16'(397);
			21562: out = 16'(3177);
			21563: out = 16'(5229);
			21564: out = 16'(4787);
			21565: out = 16'(2073);
			21566: out = 16'(-2019);
			21567: out = 16'(-4066);
			21568: out = 16'(-2079);
			21569: out = 16'(-77);
			21570: out = 16'(1497);
			21571: out = 16'(-203);
			21572: out = 16'(-2034);
			21573: out = 16'(-3856);
			21574: out = 16'(-623);
			21575: out = 16'(2031);
			21576: out = 16'(5528);
			21577: out = 16'(807);
			21578: out = 16'(425);
			21579: out = 16'(-830);
			21580: out = 16'(2713);
			21581: out = 16'(691);
			21582: out = 16'(-4165);
			21583: out = 16'(-5880);
			21584: out = 16'(-5187);
			21585: out = 16'(955);
			21586: out = 16'(-156);
			21587: out = 16'(381);
			21588: out = 16'(251);
			21589: out = 16'(1372);
			21590: out = 16'(1911);
			21591: out = 16'(6624);
			21592: out = 16'(4007);
			21593: out = 16'(1412);
			21594: out = 16'(-6005);
			21595: out = 16'(-4413);
			21596: out = 16'(-617);
			21597: out = 16'(4229);
			21598: out = 16'(3676);
			21599: out = 16'(-29);
			21600: out = 16'(-2229);
			21601: out = 16'(-1595);
			21602: out = 16'(3278);
			21603: out = 16'(4206);
			21604: out = 16'(4146);
			21605: out = 16'(-677);
			21606: out = 16'(-1686);
			21607: out = 16'(-3862);
			21608: out = 16'(-3433);
			21609: out = 16'(-5272);
			21610: out = 16'(-5011);
			21611: out = 16'(-2661);
			21612: out = 16'(1062);
			21613: out = 16'(3951);
			21614: out = 16'(1095);
			21615: out = 16'(6);
			21616: out = 16'(-1228);
			21617: out = 16'(1149);
			21618: out = 16'(1110);
			21619: out = 16'(-280);
			21620: out = 16'(64);
			21621: out = 16'(-668);
			21622: out = 16'(-1919);
			21623: out = 16'(-3256);
			21624: out = 16'(-2534);
			21625: out = 16'(3288);
			21626: out = 16'(1233);
			21627: out = 16'(-915);
			21628: out = 16'(-6052);
			21629: out = 16'(-4228);
			21630: out = 16'(-605);
			21631: out = 16'(4418);
			21632: out = 16'(5834);
			21633: out = 16'(4681);
			21634: out = 16'(3948);
			21635: out = 16'(-392);
			21636: out = 16'(-5896);
			21637: out = 16'(-4210);
			21638: out = 16'(-2124);
			21639: out = 16'(1914);
			21640: out = 16'(191);
			21641: out = 16'(-167);
			21642: out = 16'(13);
			21643: out = 16'(400);
			21644: out = 16'(630);
			21645: out = 16'(519);
			21646: out = 16'(1148);
			21647: out = 16'(1465);
			21648: out = 16'(7);
			21649: out = 16'(-125);
			21650: out = 16'(-337);
			21651: out = 16'(483);
			21652: out = 16'(129);
			21653: out = 16'(-390);
			21654: out = 16'(-2412);
			21655: out = 16'(-2050);
			21656: out = 16'(320);
			21657: out = 16'(401);
			21658: out = 16'(919);
			21659: out = 16'(-321);
			21660: out = 16'(2805);
			21661: out = 16'(3664);
			21662: out = 16'(3102);
			21663: out = 16'(434);
			21664: out = 16'(-1451);
			21665: out = 16'(-351);
			21666: out = 16'(63);
			21667: out = 16'(709);
			21668: out = 16'(-156);
			21669: out = 16'(-246);
			21670: out = 16'(-389);
			21671: out = 16'(-267);
			21672: out = 16'(913);
			21673: out = 16'(3102);
			21674: out = 16'(952);
			21675: out = 16'(480);
			21676: out = 16'(235);
			21677: out = 16'(-722);
			21678: out = 16'(-2440);
			21679: out = 16'(-5739);
			21680: out = 16'(-4068);
			21681: out = 16'(-2092);
			21682: out = 16'(-281);
			21683: out = 16'(605);
			21684: out = 16'(502);
			21685: out = 16'(-813);
			21686: out = 16'(-2424);
			21687: out = 16'(-3306);
			21688: out = 16'(1704);
			21689: out = 16'(3750);
			21690: out = 16'(5135);
			21691: out = 16'(144);
			21692: out = 16'(-3636);
			21693: out = 16'(-8675);
			21694: out = 16'(-2653);
			21695: out = 16'(168);
			21696: out = 16'(2779);
			21697: out = 16'(-2307);
			21698: out = 16'(-4245);
			21699: out = 16'(-1624);
			21700: out = 16'(1681);
			21701: out = 16'(4340);
			21702: out = 16'(569);
			21703: out = 16'(2516);
			21704: out = 16'(3056);
			21705: out = 16'(3395);
			21706: out = 16'(1791);
			21707: out = 16'(506);
			21708: out = 16'(606);
			21709: out = 16'(1391);
			21710: out = 16'(2151);
			21711: out = 16'(408);
			21712: out = 16'(-2215);
			21713: out = 16'(-5629);
			21714: out = 16'(-2621);
			21715: out = 16'(906);
			21716: out = 16'(5071);
			21717: out = 16'(5055);
			21718: out = 16'(2813);
			21719: out = 16'(-2496);
			21720: out = 16'(-5784);
			21721: out = 16'(-6715);
			21722: out = 16'(-472);
			21723: out = 16'(2028);
			21724: out = 16'(3861);
			21725: out = 16'(229);
			21726: out = 16'(-77);
			21727: out = 16'(25);
			21728: out = 16'(1219);
			21729: out = 16'(1656);
			21730: out = 16'(1368);
			21731: out = 16'(3342);
			21732: out = 16'(3011);
			21733: out = 16'(1287);
			21734: out = 16'(-434);
			21735: out = 16'(-1878);
			21736: out = 16'(-2995);
			21737: out = 16'(-2477);
			21738: out = 16'(-1583);
			21739: out = 16'(1585);
			21740: out = 16'(-99);
			21741: out = 16'(-1101);
			21742: out = 16'(-768);
			21743: out = 16'(2951);
			21744: out = 16'(6375);
			21745: out = 16'(618);
			21746: out = 16'(-2134);
			21747: out = 16'(-4900);
			21748: out = 16'(-642);
			21749: out = 16'(607);
			21750: out = 16'(-517);
			21751: out = 16'(896);
			21752: out = 16'(-769);
			21753: out = 16'(-3454);
			21754: out = 16'(-7842);
			21755: out = 16'(-7909);
			21756: out = 16'(-1223);
			21757: out = 16'(4064);
			21758: out = 16'(7320);
			21759: out = 16'(1536);
			21760: out = 16'(1336);
			21761: out = 16'(59);
			21762: out = 16'(-620);
			21763: out = 16'(-3109);
			21764: out = 16'(-5424);
			21765: out = 16'(2062);
			21766: out = 16'(2794);
			21767: out = 16'(1399);
			21768: out = 16'(-3855);
			21769: out = 16'(-4721);
			21770: out = 16'(-422);
			21771: out = 16'(56);
			21772: out = 16'(1299);
			21773: out = 16'(-296);
			21774: out = 16'(2887);
			21775: out = 16'(3729);
			21776: out = 16'(2544);
			21777: out = 16'(887);
			21778: out = 16'(-412);
			21779: out = 16'(550);
			21780: out = 16'(433);
			21781: out = 16'(544);
			21782: out = 16'(-76);
			21783: out = 16'(558);
			21784: out = 16'(1572);
			21785: out = 16'(123);
			21786: out = 16'(-163);
			21787: out = 16'(-97);
			21788: out = 16'(475);
			21789: out = 16'(694);
			21790: out = 16'(383);
			21791: out = 16'(-612);
			21792: out = 16'(-1417);
			21793: out = 16'(-1047);
			21794: out = 16'(-1293);
			21795: out = 16'(-1402);
			21796: out = 16'(-4732);
			21797: out = 16'(-2271);
			21798: out = 16'(670);
			21799: out = 16'(5350);
			21800: out = 16'(5447);
			21801: out = 16'(4011);
			21802: out = 16'(371);
			21803: out = 16'(-399);
			21804: out = 16'(493);
			21805: out = 16'(378);
			21806: out = 16'(-1245);
			21807: out = 16'(-6087);
			21808: out = 16'(-2291);
			21809: out = 16'(-108);
			21810: out = 16'(3257);
			21811: out = 16'(898);
			21812: out = 16'(-344);
			21813: out = 16'(-1206);
			21814: out = 16'(-48);
			21815: out = 16'(894);
			21816: out = 16'(1447);
			21817: out = 16'(1424);
			21818: out = 16'(1458);
			21819: out = 16'(391);
			21820: out = 16'(498);
			21821: out = 16'(142);
			21822: out = 16'(926);
			21823: out = 16'(-850);
			21824: out = 16'(-2910);
			21825: out = 16'(-5325);
			21826: out = 16'(-3840);
			21827: out = 16'(889);
			21828: out = 16'(2473);
			21829: out = 16'(2434);
			21830: out = 16'(-191);
			21831: out = 16'(-3051);
			21832: out = 16'(-4114);
			21833: out = 16'(358);
			21834: out = 16'(2779);
			21835: out = 16'(4280);
			21836: out = 16'(-648);
			21837: out = 16'(-3494);
			21838: out = 16'(-6442);
			21839: out = 16'(-194);
			21840: out = 16'(1947);
			21841: out = 16'(4130);
			21842: out = 16'(1204);
			21843: out = 16'(824);
			21844: out = 16'(664);
			21845: out = 16'(2027);
			21846: out = 16'(1514);
			21847: out = 16'(-1303);
			21848: out = 16'(-1652);
			21849: out = 16'(-2200);
			21850: out = 16'(-1828);
			21851: out = 16'(-2558);
			21852: out = 16'(-2487);
			21853: out = 16'(-1211);
			21854: out = 16'(-124);
			21855: out = 16'(1038);
			21856: out = 16'(3532);
			21857: out = 16'(4547);
			21858: out = 16'(5021);
			21859: out = 16'(-77);
			21860: out = 16'(-2533);
			21861: out = 16'(-4753);
			21862: out = 16'(-280);
			21863: out = 16'(761);
			21864: out = 16'(-47);
			21865: out = 16'(-702);
			21866: out = 16'(-1376);
			21867: out = 16'(-2840);
			21868: out = 16'(-907);
			21869: out = 16'(1036);
			21870: out = 16'(5994);
			21871: out = 16'(3796);
			21872: out = 16'(1711);
			21873: out = 16'(-3664);
			21874: out = 16'(-190);
			21875: out = 16'(4240);
			21876: out = 16'(5652);
			21877: out = 16'(1823);
			21878: out = 16'(-5599);
			21879: out = 16'(-4466);
			21880: out = 16'(-3089);
			21881: out = 16'(2179);
			21882: out = 16'(1054);
			21883: out = 16'(1741);
			21884: out = 16'(235);
			21885: out = 16'(2565);
			21886: out = 16'(2335);
			21887: out = 16'(852);
			21888: out = 16'(-669);
			21889: out = 16'(-1188);
			21890: out = 16'(-641);
			21891: out = 16'(-113);
			21892: out = 16'(-431);
			21893: out = 16'(0);
			21894: out = 16'(-2824);
			21895: out = 16'(-5598);
			21896: out = 16'(-2022);
			21897: out = 16'(677);
			21898: out = 16'(3100);
			21899: out = 16'(3762);
			21900: out = 16'(2497);
			21901: out = 16'(-449);
			21902: out = 16'(-4048);
			21903: out = 16'(-4961);
			21904: out = 16'(41);
			21905: out = 16'(-545);
			21906: out = 16'(-96);
			21907: out = 16'(-1324);
			21908: out = 16'(566);
			21909: out = 16'(1612);
			21910: out = 16'(874);
			21911: out = 16'(377);
			21912: out = 16'(50);
			21913: out = 16'(2030);
			21914: out = 16'(2332);
			21915: out = 16'(2115);
			21916: out = 16'(189);
			21917: out = 16'(-842);
			21918: out = 16'(-1180);
			21919: out = 16'(-652);
			21920: out = 16'(-446);
			21921: out = 16'(-1308);
			21922: out = 16'(-358);
			21923: out = 16'(33);
			21924: out = 16'(555);
			21925: out = 16'(-110);
			21926: out = 16'(33);
			21927: out = 16'(2038);
			21928: out = 16'(3025);
			21929: out = 16'(3451);
			21930: out = 16'(855);
			21931: out = 16'(137);
			21932: out = 16'(-506);
			21933: out = 16'(-3180);
			21934: out = 16'(-4695);
			21935: out = 16'(-5535);
			21936: out = 16'(-2936);
			21937: out = 16'(-854);
			21938: out = 16'(827);
			21939: out = 16'(1944);
			21940: out = 16'(2192);
			21941: out = 16'(563);
			21942: out = 16'(2261);
			21943: out = 16'(2582);
			21944: out = 16'(-108);
			21945: out = 16'(-746);
			21946: out = 16'(-1204);
			21947: out = 16'(619);
			21948: out = 16'(506);
			21949: out = 16'(295);
			21950: out = 16'(-1089);
			21951: out = 16'(-1283);
			21952: out = 16'(-1142);
			21953: out = 16'(237);
			21954: out = 16'(1869);
			21955: out = 16'(4600);
			21956: out = 16'(812);
			21957: out = 16'(-655);
			21958: out = 16'(-1371);
			21959: out = 16'(-539);
			21960: out = 16'(-114);
			21961: out = 16'(668);
			21962: out = 16'(-96);
			21963: out = 16'(-1047);
			21964: out = 16'(-5771);
			21965: out = 16'(-2906);
			21966: out = 16'(359);
			21967: out = 16'(4174);
			21968: out = 16'(2130);
			21969: out = 16'(-1796);
			21970: out = 16'(-2574);
			21971: out = 16'(-1315);
			21972: out = 16'(2839);
			21973: out = 16'(1274);
			21974: out = 16'(1274);
			21975: out = 16'(-589);
			21976: out = 16'(664);
			21977: out = 16'(-812);
			21978: out = 16'(-3660);
			21979: out = 16'(-3520);
			21980: out = 16'(-1768);
			21981: out = 16'(1132);
			21982: out = 16'(3848);
			21983: out = 16'(5307);
			21984: out = 16'(5821);
			21985: out = 16'(3037);
			21986: out = 16'(-431);
			21987: out = 16'(-1852);
			21988: out = 16'(-1415);
			21989: out = 16'(668);
			21990: out = 16'(-5563);
			21991: out = 16'(-7037);
			21992: out = 16'(-7349);
			21993: out = 16'(-2144);
			21994: out = 16'(1439);
			21995: out = 16'(3832);
			21996: out = 16'(3964);
			21997: out = 16'(3123);
			21998: out = 16'(699);
			21999: out = 16'(555);
			22000: out = 16'(601);
			22001: out = 16'(2242);
			22002: out = 16'(1280);
			22003: out = 16'(201);
			22004: out = 16'(-2780);
			22005: out = 16'(-1830);
			22006: out = 16'(225);
			22007: out = 16'(1021);
			22008: out = 16'(1282);
			22009: out = 16'(56);
			22010: out = 16'(864);
			22011: out = 16'(-193);
			22012: out = 16'(-1210);
			22013: out = 16'(-2119);
			22014: out = 16'(-1506);
			22015: out = 16'(-239);
			22016: out = 16'(986);
			22017: out = 16'(1442);
			22018: out = 16'(1497);
			22019: out = 16'(755);
			22020: out = 16'(-296);
			22021: out = 16'(-5706);
			22022: out = 16'(-2995);
			22023: out = 16'(392);
			22024: out = 16'(4039);
			22025: out = 16'(2967);
			22026: out = 16'(298);
			22027: out = 16'(522);
			22028: out = 16'(681);
			22029: out = 16'(1381);
			22030: out = 16'(1472);
			22031: out = 16'(233);
			22032: out = 16'(-2198);
			22033: out = 16'(-4844);
			22034: out = 16'(-4345);
			22035: out = 16'(1660);
			22036: out = 16'(2761);
			22037: out = 16'(3524);
			22038: out = 16'(200);
			22039: out = 16'(623);
			22040: out = 16'(708);
			22041: out = 16'(2757);
			22042: out = 16'(3081);
			22043: out = 16'(3359);
			22044: out = 16'(-4);
			22045: out = 16'(-1095);
			22046: out = 16'(-2632);
			22047: out = 16'(-1868);
			22048: out = 16'(-4110);
			22049: out = 16'(-7596);
			22050: out = 16'(-7643);
			22051: out = 16'(-5008);
			22052: out = 16'(2072);
			22053: out = 16'(2034);
			22054: out = 16'(1888);
			22055: out = 16'(-3083);
			22056: out = 16'(-357);
			22057: out = 16'(722);
			22058: out = 16'(1974);
			22059: out = 16'(67);
			22060: out = 16'(-1242);
			22061: out = 16'(-5324);
			22062: out = 16'(-3220);
			22063: out = 16'(-522);
			22064: out = 16'(3625);
			22065: out = 16'(2505);
			22066: out = 16'(-199);
			22067: out = 16'(-4492);
			22068: out = 16'(-2897);
			22069: out = 16'(3743);
			22070: out = 16'(5661);
			22071: out = 16'(6365);
			22072: out = 16'(4547);
			22073: out = 16'(-615);
			22074: out = 16'(-4414);
			22075: out = 16'(-3504);
			22076: out = 16'(-140);
			22077: out = 16'(3786);
			22078: out = 16'(1157);
			22079: out = 16'(1483);
			22080: out = 16'(109);
			22081: out = 16'(1792);
			22082: out = 16'(1110);
			22083: out = 16'(1749);
			22084: out = 16'(-302);
			22085: out = 16'(878);
			22086: out = 16'(1930);
			22087: out = 16'(1980);
			22088: out = 16'(-391);
			22089: out = 16'(-3652);
			22090: out = 16'(-6651);
			22091: out = 16'(-5919);
			22092: out = 16'(-202);
			22093: out = 16'(3655);
			22094: out = 16'(5471);
			22095: out = 16'(-321);
			22096: out = 16'(-281);
			22097: out = 16'(-342);
			22098: out = 16'(410);
			22099: out = 16'(301);
			22100: out = 16'(-215);
			22101: out = 16'(1518);
			22102: out = 16'(79);
			22103: out = 16'(-2137);
			22104: out = 16'(-3616);
			22105: out = 16'(-1721);
			22106: out = 16'(3400);
			22107: out = 16'(2928);
			22108: out = 16'(2346);
			22109: out = 16'(-559);
			22110: out = 16'(817);
			22111: out = 16'(1536);
			22112: out = 16'(1166);
			22113: out = 16'(1931);
			22114: out = 16'(1808);
			22115: out = 16'(2384);
			22116: out = 16'(-1051);
			22117: out = 16'(-4150);
			22118: out = 16'(-4789);
			22119: out = 16'(-1591);
			22120: out = 16'(3236);
			22121: out = 16'(-1298);
			22122: out = 16'(-3462);
			22123: out = 16'(-6387);
			22124: out = 16'(-1717);
			22125: out = 16'(696);
			22126: out = 16'(1368);
			22127: out = 16'(3284);
			22128: out = 16'(3247);
			22129: out = 16'(2445);
			22130: out = 16'(-2511);
			22131: out = 16'(-5943);
			22132: out = 16'(-4365);
			22133: out = 16'(-2443);
			22134: out = 16'(508);
			22135: out = 16'(144);
			22136: out = 16'(1790);
			22137: out = 16'(2093);
			22138: out = 16'(582);
			22139: out = 16'(-889);
			22140: out = 16'(-1724);
			22141: out = 16'(-1392);
			22142: out = 16'(423);
			22143: out = 16'(3208);
			22144: out = 16'(3528);
			22145: out = 16'(3111);
			22146: out = 16'(435);
			22147: out = 16'(1417);
			22148: out = 16'(673);
			22149: out = 16'(-1815);
			22150: out = 16'(-2228);
			22151: out = 16'(-1415);
			22152: out = 16'(261);
			22153: out = 16'(2730);
			22154: out = 16'(4219);
			22155: out = 16'(2443);
			22156: out = 16'(584);
			22157: out = 16'(-1584);
			22158: out = 16'(-2566);
			22159: out = 16'(-3237);
			22160: out = 16'(-3696);
			22161: out = 16'(-806);
			22162: out = 16'(-9);
			22163: out = 16'(-257);
			22164: out = 16'(-3810);
			22165: out = 16'(-4983);
			22166: out = 16'(-1503);
			22167: out = 16'(-352);
			22168: out = 16'(1762);
			22169: out = 16'(2704);
			22170: out = 16'(3819);
			22171: out = 16'(3196);
			22172: out = 16'(1252);
			22173: out = 16'(-375);
			22174: out = 16'(-1198);
			22175: out = 16'(-4284);
			22176: out = 16'(-2822);
			22177: out = 16'(246);
			22178: out = 16'(3499);
			22179: out = 16'(4327);
			22180: out = 16'(2635);
			22181: out = 16'(3090);
			22182: out = 16'(2777);
			22183: out = 16'(3719);
			22184: out = 16'(810);
			22185: out = 16'(-508);
			22186: out = 16'(-273);
			22187: out = 16'(-334);
			22188: out = 16'(-434);
			22189: out = 16'(-1302);
			22190: out = 16'(-954);
			22191: out = 16'(-552);
			22192: out = 16'(-2031);
			22193: out = 16'(-2375);
			22194: out = 16'(-2686);
			22195: out = 16'(2714);
			22196: out = 16'(3672);
			22197: out = 16'(3325);
			22198: out = 16'(-2084);
			22199: out = 16'(-4747);
			22200: out = 16'(-5348);
			22201: out = 16'(-2134);
			22202: out = 16'(1248);
			22203: out = 16'(4164);
			22204: out = 16'(2746);
			22205: out = 16'(396);
			22206: out = 16'(-1594);
			22207: out = 16'(-3698);
			22208: out = 16'(-4275);
			22209: out = 16'(-2175);
			22210: out = 16'(-849);
			22211: out = 16'(145);
			22212: out = 16'(3);
			22213: out = 16'(-9);
			22214: out = 16'(-228);
			22215: out = 16'(36);
			22216: out = 16'(12);
			22217: out = 16'(85);
			22218: out = 16'(329);
			22219: out = 16'(1628);
			22220: out = 16'(4560);
			22221: out = 16'(3783);
			22222: out = 16'(2804);
			22223: out = 16'(-1515);
			22224: out = 16'(1421);
			22225: out = 16'(2553);
			22226: out = 16'(499);
			22227: out = 16'(-1910);
			22228: out = 16'(-3790);
			22229: out = 16'(169);
			22230: out = 16'(-312);
			22231: out = 16'(-1315);
			22232: out = 16'(297);
			22233: out = 16'(33);
			22234: out = 16'(-450);
			22235: out = 16'(-3040);
			22236: out = 16'(-3749);
			22237: out = 16'(-3569);
			22238: out = 16'(-1012);
			22239: out = 16'(1094);
			22240: out = 16'(3899);
			22241: out = 16'(1194);
			22242: out = 16'(-174);
			22243: out = 16'(-130);
			22244: out = 16'(1729);
			22245: out = 16'(3017);
			22246: out = 16'(3042);
			22247: out = 16'(67);
			22248: out = 16'(-3283);
			22249: out = 16'(-2002);
			22250: out = 16'(-701);
			22251: out = 16'(1904);
			22252: out = 16'(1745);
			22253: out = 16'(2614);
			22254: out = 16'(2616);
			22255: out = 16'(1814);
			22256: out = 16'(806);
			22257: out = 16'(633);
			22258: out = 16'(-239);
			22259: out = 16'(-268);
			22260: out = 16'(-682);
			22261: out = 16'(633);
			22262: out = 16'(1556);
			22263: out = 16'(3427);
			22264: out = 16'(1213);
			22265: out = 16'(-1037);
			22266: out = 16'(-503);
			22267: out = 16'(-462);
			22268: out = 16'(27);
			22269: out = 16'(-4287);
			22270: out = 16'(-4829);
			22271: out = 16'(-4599);
			22272: out = 16'(-1233);
			22273: out = 16'(-95);
			22274: out = 16'(-166);
			22275: out = 16'(-1391);
			22276: out = 16'(-2284);
			22277: out = 16'(-2714);
			22278: out = 16'(-1025);
			22279: out = 16'(842);
			22280: out = 16'(2873);
			22281: out = 16'(2256);
			22282: out = 16'(1099);
			22283: out = 16'(716);
			22284: out = 16'(-158);
			22285: out = 16'(-284);
			22286: out = 16'(-493);
			22287: out = 16'(80);
			22288: out = 16'(483);
			22289: out = 16'(2610);
			22290: out = 16'(2585);
			22291: out = 16'(2037);
			22292: out = 16'(71);
			22293: out = 16'(-811);
			22294: out = 16'(-1369);
			22295: out = 16'(632);
			22296: out = 16'(1351);
			22297: out = 16'(1365);
			22298: out = 16'(-1425);
			22299: out = 16'(-2929);
			22300: out = 16'(-391);
			22301: out = 16'(-25);
			22302: out = 16'(750);
			22303: out = 16'(202);
			22304: out = 16'(400);
			22305: out = 16'(138);
			22306: out = 16'(-298);
			22307: out = 16'(-540);
			22308: out = 16'(-375);
			22309: out = 16'(-471);
			22310: out = 16'(-620);
			22311: out = 16'(-1279);
			22312: out = 16'(228);
			22313: out = 16'(1051);
			22314: out = 16'(2203);
			22315: out = 16'(895);
			22316: out = 16'(218);
			22317: out = 16'(322);
			22318: out = 16'(921);
			22319: out = 16'(1173);
			22320: out = 16'(-274);
			22321: out = 16'(-221);
			22322: out = 16'(-340);
			22323: out = 16'(-223);
			22324: out = 16'(9);
			22325: out = 16'(574);
			22326: out = 16'(-1076);
			22327: out = 16'(-2104);
			22328: out = 16'(-3932);
			22329: out = 16'(519);
			22330: out = 16'(1620);
			22331: out = 16'(2266);
			22332: out = 16'(-1032);
			22333: out = 16'(-1954);
			22334: out = 16'(-1323);
			22335: out = 16'(1079);
			22336: out = 16'(1935);
			22337: out = 16'(772);
			22338: out = 16'(-1881);
			22339: out = 16'(-3967);
			22340: out = 16'(-3731);
			22341: out = 16'(-1663);
			22342: out = 16'(929);
			22343: out = 16'(2103);
			22344: out = 16'(700);
			22345: out = 16'(-2332);
			22346: out = 16'(-3196);
			22347: out = 16'(-2139);
			22348: out = 16'(2117);
			22349: out = 16'(-116);
			22350: out = 16'(141);
			22351: out = 16'(443);
			22352: out = 16'(861);
			22353: out = 16'(663);
			22354: out = 16'(629);
			22355: out = 16'(991);
			22356: out = 16'(1898);
			22357: out = 16'(2683);
			22358: out = 16'(2727);
			22359: out = 16'(1562);
			22360: out = 16'(147);
			22361: out = 16'(-2212);
			22362: out = 16'(-3622);
			22363: out = 16'(-2489);
			22364: out = 16'(-447);
			22365: out = 16'(1523);
			22366: out = 16'(3920);
			22367: out = 16'(2733);
			22368: out = 16'(-1497);
			22369: out = 16'(-2929);
			22370: out = 16'(-3020);
			22371: out = 16'(1005);
			22372: out = 16'(-66);
			22373: out = 16'(-77);
			22374: out = 16'(-1319);
			22375: out = 16'(31);
			22376: out = 16'(881);
			22377: out = 16'(2194);
			22378: out = 16'(1314);
			22379: out = 16'(301);
			22380: out = 16'(598);
			22381: out = 16'(1157);
			22382: out = 16'(2156);
			22383: out = 16'(564);
			22384: out = 16'(99);
			22385: out = 16'(-314);
			22386: out = 16'(-960);
			22387: out = 16'(-1432);
			22388: out = 16'(-1147);
			22389: out = 16'(-161);
			22390: out = 16'(909);
			22391: out = 16'(193);
			22392: out = 16'(2168);
			22393: out = 16'(2438);
			22394: out = 16'(2384);
			22395: out = 16'(-1719);
			22396: out = 16'(-5017);
			22397: out = 16'(-3157);
			22398: out = 16'(-1054);
			22399: out = 16'(1721);
			22400: out = 16'(1151);
			22401: out = 16'(1132);
			22402: out = 16'(394);
			22403: out = 16'(-258);
			22404: out = 16'(-104);
			22405: out = 16'(1430);
			22406: out = 16'(544);
			22407: out = 16'(-859);
			22408: out = 16'(-4932);
			22409: out = 16'(-3463);
			22410: out = 16'(-2375);
			22411: out = 16'(-51);
			22412: out = 16'(-328);
			22413: out = 16'(-78);
			22414: out = 16'(500);
			22415: out = 16'(1551);
			22416: out = 16'(2050);
			22417: out = 16'(670);
			22418: out = 16'(-102);
			22419: out = 16'(-382);
			22420: out = 16'(-1291);
			22421: out = 16'(-223);
			22422: out = 16'(1482);
			22423: out = 16'(2609);
			22424: out = 16'(1558);
			22425: out = 16'(-2378);
			22426: out = 16'(-2000);
			22427: out = 16'(-1485);
			22428: out = 16'(1624);
			22429: out = 16'(588);
			22430: out = 16'(351);
			22431: out = 16'(-597);
			22432: out = 16'(319);
			22433: out = 16'(311);
			22434: out = 16'(-883);
			22435: out = 16'(-2192);
			22436: out = 16'(-2754);
			22437: out = 16'(-3025);
			22438: out = 16'(-1517);
			22439: out = 16'(130);
			22440: out = 16'(3190);
			22441: out = 16'(2311);
			22442: out = 16'(-1452);
			22443: out = 16'(-1632);
			22444: out = 16'(-1508);
			22445: out = 16'(683);
			22446: out = 16'(585);
			22447: out = 16'(652);
			22448: out = 16'(-324);
			22449: out = 16'(-1248);
			22450: out = 16'(-1570);
			22451: out = 16'(2274);
			22452: out = 16'(2471);
			22453: out = 16'(2753);
			22454: out = 16'(-1843);
			22455: out = 16'(-873);
			22456: out = 16'(601);
			22457: out = 16'(2677);
			22458: out = 16'(1756);
			22459: out = 16'(-360);
			22460: out = 16'(-237);
			22461: out = 16'(497);
			22462: out = 16'(2141);
			22463: out = 16'(2615);
			22464: out = 16'(2068);
			22465: out = 16'(-391);
			22466: out = 16'(-371);
			22467: out = 16'(311);
			22468: out = 16'(3298);
			22469: out = 16'(3428);
			22470: out = 16'(2540);
			22471: out = 16'(-1838);
			22472: out = 16'(-4544);
			22473: out = 16'(-6161);
			22474: out = 16'(2442);
			22475: out = 16'(4106);
			22476: out = 16'(4535);
			22477: out = 16'(-1143);
			22478: out = 16'(-2632);
			22479: out = 16'(-2133);
			22480: out = 16'(-926);
			22481: out = 16'(-203);
			22482: out = 16'(-756);
			22483: out = 16'(-452);
			22484: out = 16'(-852);
			22485: out = 16'(-1292);
			22486: out = 16'(-951);
			22487: out = 16'(-445);
			22488: out = 16'(-1504);
			22489: out = 16'(-140);
			22490: out = 16'(688);
			22491: out = 16'(2074);
			22492: out = 16'(946);
			22493: out = 16'(-618);
			22494: out = 16'(-4058);
			22495: out = 16'(-4123);
			22496: out = 16'(-2466);
			22497: out = 16'(1144);
			22498: out = 16'(2077);
			22499: out = 16'(94);
			22500: out = 16'(293);
			22501: out = 16'(85);
			22502: out = 16'(2568);
			22503: out = 16'(-1336);
			22504: out = 16'(-3385);
			22505: out = 16'(-5547);
			22506: out = 16'(-2204);
			22507: out = 16'(464);
			22508: out = 16'(-134);
			22509: out = 16'(85);
			22510: out = 16'(-200);
			22511: out = 16'(831);
			22512: out = 16'(491);
			22513: out = 16'(-10);
			22514: out = 16'(568);
			22515: out = 16'(484);
			22516: out = 16'(584);
			22517: out = 16'(-2734);
			22518: out = 16'(-2611);
			22519: out = 16'(927);
			22520: out = 16'(611);
			22521: out = 16'(871);
			22522: out = 16'(-428);
			22523: out = 16'(1119);
			22524: out = 16'(1314);
			22525: out = 16'(147);
			22526: out = 16'(-1054);
			22527: out = 16'(-1627);
			22528: out = 16'(1447);
			22529: out = 16'(859);
			22530: out = 16'(-84);
			22531: out = 16'(536);
			22532: out = 16'(1117);
			22533: out = 16'(2444);
			22534: out = 16'(-675);
			22535: out = 16'(-736);
			22536: out = 16'(-74);
			22537: out = 16'(3327);
			22538: out = 16'(3464);
			22539: out = 16'(-440);
			22540: out = 16'(353);
			22541: out = 16'(678);
			22542: out = 16'(2950);
			22543: out = 16'(1293);
			22544: out = 16'(-280);
			22545: out = 16'(-2757);
			22546: out = 16'(-2603);
			22547: out = 16'(-1727);
			22548: out = 16'(59);
			22549: out = 16'(673);
			22550: out = 16'(526);
			22551: out = 16'(761);
			22552: out = 16'(-83);
			22553: out = 16'(-1243);
			22554: out = 16'(-646);
			22555: out = 16'(193);
			22556: out = 16'(1414);
			22557: out = 16'(876);
			22558: out = 16'(136);
			22559: out = 16'(-1205);
			22560: out = 16'(-774);
			22561: out = 16'(-510);
			22562: out = 16'(-2163);
			22563: out = 16'(-1008);
			22564: out = 16'(122);
			22565: out = 16'(4192);
			22566: out = 16'(2510);
			22567: out = 16'(177);
			22568: out = 16'(-1715);
			22569: out = 16'(-1429);
			22570: out = 16'(0);
			22571: out = 16'(-257);
			22572: out = 16'(-164);
			22573: out = 16'(-143);
			22574: out = 16'(-898);
			22575: out = 16'(-1915);
			22576: out = 16'(-4854);
			22577: out = 16'(618);
			22578: out = 16'(3681);
			22579: out = 16'(4995);
			22580: out = 16'(1335);
			22581: out = 16'(-1802);
			22582: out = 16'(-1113);
			22583: out = 16'(326);
			22584: out = 16'(2259);
			22585: out = 16'(-350);
			22586: out = 16'(-2086);
			22587: out = 16'(-4922);
			22588: out = 16'(21);
			22589: out = 16'(388);
			22590: out = 16'(903);
			22591: out = 16'(-1704);
			22592: out = 16'(-1160);
			22593: out = 16'(379);
			22594: out = 16'(2417);
			22595: out = 16'(2173);
			22596: out = 16'(-337);
			22597: out = 16'(-1589);
			22598: out = 16'(-1327);
			22599: out = 16'(2010);
			22600: out = 16'(3036);
			22601: out = 16'(3151);
			22602: out = 16'(878);
			22603: out = 16'(-1250);
			22604: out = 16'(-3240);
			22605: out = 16'(-4519);
			22606: out = 16'(-2889);
			22607: out = 16'(383);
			22608: out = 16'(312);
			22609: out = 16'(939);
			22610: out = 16'(519);
			22611: out = 16'(1397);
			22612: out = 16'(953);
			22613: out = 16'(-435);
			22614: out = 16'(-368);
			22615: out = 16'(-118);
			22616: out = 16'(1568);
			22617: out = 16'(-208);
			22618: out = 16'(-1935);
			22619: out = 16'(-6253);
			22620: out = 16'(-3180);
			22621: out = 16'(679);
			22622: out = 16'(3215);
			22623: out = 16'(3324);
			22624: out = 16'(1910);
			22625: out = 16'(2394);
			22626: out = 16'(1454);
			22627: out = 16'(478);
			22628: out = 16'(47);
			22629: out = 16'(-861);
			22630: out = 16'(-2068);
			22631: out = 16'(-3333);
			22632: out = 16'(-3009);
			22633: out = 16'(-175);
			22634: out = 16'(95);
			22635: out = 16'(612);
			22636: out = 16'(-212);
			22637: out = 16'(1312);
			22638: out = 16'(2390);
			22639: out = 16'(2047);
			22640: out = 16'(2249);
			22641: out = 16'(1693);
			22642: out = 16'(-639);
			22643: out = 16'(-2894);
			22644: out = 16'(-4606);
			22645: out = 16'(-3257);
			22646: out = 16'(-960);
			22647: out = 16'(2596);
			22648: out = 16'(1485);
			22649: out = 16'(1403);
			22650: out = 16'(494);
			22651: out = 16'(2374);
			22652: out = 16'(2107);
			22653: out = 16'(-1316);
			22654: out = 16'(-1171);
			22655: out = 16'(-941);
			22656: out = 16'(1521);
			22657: out = 16'(-492);
			22658: out = 16'(-2187);
			22659: out = 16'(-1166);
			22660: out = 16'(-732);
			22661: out = 16'(67);
			22662: out = 16'(-261);
			22663: out = 16'(293);
			22664: out = 16'(648);
			22665: out = 16'(684);
			22666: out = 16'(796);
			22667: out = 16'(1514);
			22668: out = 16'(-614);
			22669: out = 16'(-1038);
			22670: out = 16'(-99);
			22671: out = 16'(1323);
			22672: out = 16'(2067);
			22673: out = 16'(179);
			22674: out = 16'(489);
			22675: out = 16'(158);
			22676: out = 16'(814);
			22677: out = 16'(-928);
			22678: out = 16'(-2182);
			22679: out = 16'(-2145);
			22680: out = 16'(-1181);
			22681: out = 16'(143);
			22682: out = 16'(2315);
			22683: out = 16'(3447);
			22684: out = 16'(4097);
			22685: out = 16'(-689);
			22686: out = 16'(-3010);
			22687: out = 16'(-3693);
			22688: out = 16'(-1350);
			22689: out = 16'(173);
			22690: out = 16'(-636);
			22691: out = 16'(267);
			22692: out = 16'(486);
			22693: out = 16'(1479);
			22694: out = 16'(1656);
			22695: out = 16'(2052);
			22696: out = 16'(-383);
			22697: out = 16'(687);
			22698: out = 16'(1130);
			22699: out = 16'(1550);
			22700: out = 16'(-320);
			22701: out = 16'(-2337);
			22702: out = 16'(-5780);
			22703: out = 16'(-5333);
			22704: out = 16'(-2534);
			22705: out = 16'(989);
			22706: out = 16'(2007);
			22707: out = 16'(-568);
			22708: out = 16'(-197);
			22709: out = 16'(196);
			22710: out = 16'(3068);
			22711: out = 16'(2004);
			22712: out = 16'(510);
			22713: out = 16'(-4291);
			22714: out = 16'(-4652);
			22715: out = 16'(-4018);
			22716: out = 16'(-645);
			22717: out = 16'(134);
			22718: out = 16'(33);
			22719: out = 16'(881);
			22720: out = 16'(430);
			22721: out = 16'(-160);
			22722: out = 16'(-947);
			22723: out = 16'(-425);
			22724: out = 16'(617);
			22725: out = 16'(3033);
			22726: out = 16'(3216);
			22727: out = 16'(622);
			22728: out = 16'(-831);
			22729: out = 16'(-1995);
			22730: out = 16'(-4);
			22731: out = 16'(-957);
			22732: out = 16'(-562);
			22733: out = 16'(1200);
			22734: out = 16'(2771);
			22735: out = 16'(3507);
			22736: out = 16'(1024);
			22737: out = 16'(421);
			22738: out = 16'(470);
			22739: out = 16'(-196);
			22740: out = 16'(407);
			22741: out = 16'(1372);
			22742: out = 16'(692);
			22743: out = 16'(-243);
			22744: out = 16'(-1198);
			22745: out = 16'(-1925);
			22746: out = 16'(-1656);
			22747: out = 16'(-524);
			22748: out = 16'(2144);
			22749: out = 16'(3326);
			22750: out = 16'(-312);
			22751: out = 16'(225);
			22752: out = 16'(309);
			22753: out = 16'(1398);
			22754: out = 16'(440);
			22755: out = 16'(-596);
			22756: out = 16'(-1166);
			22757: out = 16'(-857);
			22758: out = 16'(-44);
			22759: out = 16'(350);
			22760: out = 16'(736);
			22761: out = 16'(473);
			22762: out = 16'(1775);
			22763: out = 16'(1694);
			22764: out = 16'(218);
			22765: out = 16'(290);
			22766: out = 16'(283);
			22767: out = 16'(529);
			22768: out = 16'(-43);
			22769: out = 16'(-880);
			22770: out = 16'(-1939);
			22771: out = 16'(-2624);
			22772: out = 16'(-2718);
			22773: out = 16'(-1530);
			22774: out = 16'(333);
			22775: out = 16'(2350);
			22776: out = 16'(1390);
			22777: out = 16'(1098);
			22778: out = 16'(238);
			22779: out = 16'(1697);
			22780: out = 16'(2750);
			22781: out = 16'(4944);
			22782: out = 16'(985);
			22783: out = 16'(-1937);
			22784: out = 16'(-5795);
			22785: out = 16'(-1924);
			22786: out = 16'(1173);
			22787: out = 16'(935);
			22788: out = 16'(1039);
			22789: out = 16'(-522);
			22790: out = 16'(-3170);
			22791: out = 16'(-4947);
			22792: out = 16'(-5122);
			22793: out = 16'(-2665);
			22794: out = 16'(-778);
			22795: out = 16'(-64);
			22796: out = 16'(2111);
			22797: out = 16'(1610);
			22798: out = 16'(580);
			22799: out = 16'(-2674);
			22800: out = 16'(-2889);
			22801: out = 16'(-134);
			22802: out = 16'(1463);
			22803: out = 16'(2085);
			22804: out = 16'(-79);
			22805: out = 16'(-83);
			22806: out = 16'(-391);
			22807: out = 16'(-1071);
			22808: out = 16'(-611);
			22809: out = 16'(-14);
			22810: out = 16'(2863);
			22811: out = 16'(1585);
			22812: out = 16'(-687);
			22813: out = 16'(-4569);
			22814: out = 16'(-4378);
			22815: out = 16'(-1341);
			22816: out = 16'(1218);
			22817: out = 16'(2799);
			22818: out = 16'(2079);
			22819: out = 16'(1930);
			22820: out = 16'(1722);
			22821: out = 16'(3883);
			22822: out = 16'(2060);
			22823: out = 16'(1180);
			22824: out = 16'(338);
			22825: out = 16'(141);
			22826: out = 16'(-640);
			22827: out = 16'(-2449);
			22828: out = 16'(-4225);
			22829: out = 16'(-5269);
			22830: out = 16'(-2455);
			22831: out = 16'(-83);
			22832: out = 16'(2632);
			22833: out = 16'(896);
			22834: out = 16'(863);
			22835: out = 16'(396);
			22836: out = 16'(2552);
			22837: out = 16'(2208);
			22838: out = 16'(-148);
			22839: out = 16'(-745);
			22840: out = 16'(-1557);
			22841: out = 16'(-2832);
			22842: out = 16'(-1409);
			22843: out = 16'(517);
			22844: out = 16'(4116);
			22845: out = 16'(3689);
			22846: out = 16'(2274);
			22847: out = 16'(-1588);
			22848: out = 16'(-1290);
			22849: out = 16'(750);
			22850: out = 16'(1648);
			22851: out = 16'(1532);
			22852: out = 16'(-693);
			22853: out = 16'(1301);
			22854: out = 16'(542);
			22855: out = 16'(-376);
			22856: out = 16'(-1946);
			22857: out = 16'(-1591);
			22858: out = 16'(-423);
			22859: out = 16'(2663);
			22860: out = 16'(4440);
			22861: out = 16'(4807);
			22862: out = 16'(1894);
			22863: out = 16'(-1248);
			22864: out = 16'(-2725);
			22865: out = 16'(-3335);
			22866: out = 16'(-3015);
			22867: out = 16'(-3805);
			22868: out = 16'(-4129);
			22869: out = 16'(-4547);
			22870: out = 16'(-2501);
			22871: out = 16'(-865);
			22872: out = 16'(906);
			22873: out = 16'(753);
			22874: out = 16'(769);
			22875: out = 16'(784);
			22876: out = 16'(35);
			22877: out = 16'(-201);
			22878: out = 16'(520);
			22879: out = 16'(192);
			22880: out = 16'(-70);
			22881: out = 16'(589);
			22882: out = 16'(-53);
			22883: out = 16'(-530);
			22884: out = 16'(-3576);
			22885: out = 16'(-1925);
			22886: out = 16'(473);
			22887: out = 16'(3865);
			22888: out = 16'(3210);
			22889: out = 16'(325);
			22890: out = 16'(1443);
			22891: out = 16'(1533);
			22892: out = 16'(2229);
			22893: out = 16'(2485);
			22894: out = 16'(3125);
			22895: out = 16'(4102);
			22896: out = 16'(1713);
			22897: out = 16'(-315);
			22898: out = 16'(-1259);
			22899: out = 16'(-2508);
			22900: out = 16'(-3176);
			22901: out = 16'(-3724);
			22902: out = 16'(-2638);
			22903: out = 16'(-683);
			22904: out = 16'(-203);
			22905: out = 16'(1760);
			22906: out = 16'(2504);
			22907: out = 16'(3148);
			22908: out = 16'(-111);
			22909: out = 16'(-4832);
			22910: out = 16'(-5907);
			22911: out = 16'(-4809);
			22912: out = 16'(-815);
			22913: out = 16'(141);
			22914: out = 16'(1199);
			22915: out = 16'(2280);
			22916: out = 16'(99);
			22917: out = 16'(-972);
			22918: out = 16'(346);
			22919: out = 16'(2952);
			22920: out = 16'(4691);
			22921: out = 16'(850);
			22922: out = 16'(-2073);
			22923: out = 16'(-5979);
			22924: out = 16'(-3248);
			22925: out = 16'(-4486);
			22926: out = 16'(-4767);
			22927: out = 16'(-3472);
			22928: out = 16'(454);
			22929: out = 16'(5341);
			22930: out = 16'(4615);
			22931: out = 16'(3394);
			22932: out = 16'(629);
			22933: out = 16'(1252);
			22934: out = 16'(1195);
			22935: out = 16'(-187);
			22936: out = 16'(463);
			22937: out = 16'(547);
			22938: out = 16'(654);
			22939: out = 16'(-2133);
			22940: out = 16'(-4482);
			22941: out = 16'(-1843);
			22942: out = 16'(-1478);
			22943: out = 16'(-755);
			22944: out = 16'(-1038);
			22945: out = 16'(-236);
			22946: out = 16'(742);
			22947: out = 16'(578);
			22948: out = 16'(975);
			22949: out = 16'(1635);
			22950: out = 16'(911);
			22951: out = 16'(296);
			22952: out = 16'(-131);
			22953: out = 16'(-75);
			22954: out = 16'(127);
			22955: out = 16'(-305);
			22956: out = 16'(312);
			22957: out = 16'(796);
			22958: out = 16'(2908);
			22959: out = 16'(2422);
			22960: out = 16'(2027);
			22961: out = 16'(-928);
			22962: out = 16'(-593);
			22963: out = 16'(-74);
			22964: out = 16'(3699);
			22965: out = 16'(2835);
			22966: out = 16'(137);
			22967: out = 16'(-4017);
			22968: out = 16'(-4757);
			22969: out = 16'(-1661);
			22970: out = 16'(288);
			22971: out = 16'(1621);
			22972: out = 16'(561);
			22973: out = 16'(284);
			22974: out = 16'(68);
			22975: out = 16'(1293);
			22976: out = 16'(2546);
			22977: out = 16'(3249);
			22978: out = 16'(707);
			22979: out = 16'(-1530);
			22980: out = 16'(-3812);
			22981: out = 16'(-2171);
			22982: out = 16'(-918);
			22983: out = 16'(888);
			22984: out = 16'(1180);
			22985: out = 16'(1009);
			22986: out = 16'(-519);
			22987: out = 16'(245);
			22988: out = 16'(630);
			22989: out = 16'(1396);
			22990: out = 16'(1280);
			22991: out = 16'(1424);
			22992: out = 16'(2012);
			22993: out = 16'(1040);
			22994: out = 16'(-166);
			22995: out = 16'(-1920);
			22996: out = 16'(-1404);
			22997: out = 16'(-236);
			22998: out = 16'(-364);
			22999: out = 16'(174);
			23000: out = 16'(549);
			23001: out = 16'(545);
			23002: out = 16'(197);
			23003: out = 16'(-466);
			23004: out = 16'(1904);
			23005: out = 16'(3309);
			23006: out = 16'(4582);
			23007: out = 16'(1265);
			23008: out = 16'(-1710);
			23009: out = 16'(-4482);
			23010: out = 16'(-4360);
			23011: out = 16'(-2877);
			23012: out = 16'(-12);
			23013: out = 16'(1380);
			23014: out = 16'(1913);
			23015: out = 16'(413);
			23016: out = 16'(225);
			23017: out = 16'(134);
			23018: out = 16'(-1756);
			23019: out = 16'(-2137);
			23020: out = 16'(-1925);
			23021: out = 16'(-736);
			23022: out = 16'(-711);
			23023: out = 16'(-2115);
			23024: out = 16'(-427);
			23025: out = 16'(-34);
			23026: out = 16'(587);
			23027: out = 16'(-1796);
			23028: out = 16'(-2133);
			23029: out = 16'(1481);
			23030: out = 16'(1717);
			23031: out = 16'(2187);
			23032: out = 16'(1194);
			23033: out = 16'(2153);
			23034: out = 16'(2201);
			23035: out = 16'(-2908);
			23036: out = 16'(-4606);
			23037: out = 16'(-5078);
			23038: out = 16'(-1208);
			23039: out = 16'(317);
			23040: out = 16'(401);
			23041: out = 16'(2550);
			23042: out = 16'(2259);
			23043: out = 16'(603);
			23044: out = 16'(-594);
			23045: out = 16'(-518);
			23046: out = 16'(3072);
			23047: out = 16'(771);
			23048: out = 16'(-499);
			23049: out = 16'(-1998);
			23050: out = 16'(-911);
			23051: out = 16'(-91);
			23052: out = 16'(-1056);
			23053: out = 16'(-1145);
			23054: out = 16'(-948);
			23055: out = 16'(-257);
			23056: out = 16'(273);
			23057: out = 16'(533);
			23058: out = 16'(3038);
			23059: out = 16'(3707);
			23060: out = 16'(4085);
			23061: out = 16'(-1061);
			23062: out = 16'(-3297);
			23063: out = 16'(-2588);
			23064: out = 16'(-1379);
			23065: out = 16'(-270);
			23066: out = 16'(-2251);
			23067: out = 16'(251);
			23068: out = 16'(1861);
			23069: out = 16'(4139);
			23070: out = 16'(2318);
			23071: out = 16'(100);
			23072: out = 16'(-170);
			23073: out = 16'(-690);
			23074: out = 16'(-373);
			23075: out = 16'(-2015);
			23076: out = 16'(-1243);
			23077: out = 16'(-132);
			23078: out = 16'(1106);
			23079: out = 16'(830);
			23080: out = 16'(-480);
			23081: out = 16'(-1575);
			23082: out = 16'(-1659);
			23083: out = 16'(-26);
			23084: out = 16'(136);
			23085: out = 16'(513);
			23086: out = 16'(264);
			23087: out = 16'(1390);
			23088: out = 16'(2021);
			23089: out = 16'(321);
			23090: out = 16'(377);
			23091: out = 16'(294);
			23092: out = 16'(2015);
			23093: out = 16'(881);
			23094: out = 16'(-723);
			23095: out = 16'(-3942);
			23096: out = 16'(-3155);
			23097: out = 16'(824);
			23098: out = 16'(286);
			23099: out = 16'(801);
			23100: out = 16'(139);
			23101: out = 16'(2145);
			23102: out = 16'(2555);
			23103: out = 16'(2022);
			23104: out = 16'(46);
			23105: out = 16'(-1815);
			23106: out = 16'(-1800);
			23107: out = 16'(-3122);
			23108: out = 16'(-3432);
			23109: out = 16'(-2322);
			23110: out = 16'(-14);
			23111: out = 16'(2344);
			23112: out = 16'(668);
			23113: out = 16'(582);
			23114: out = 16'(351);
			23115: out = 16'(2312);
			23116: out = 16'(2570);
			23117: out = 16'(1837);
			23118: out = 16'(423);
			23119: out = 16'(-642);
			23120: out = 16'(-291);
			23121: out = 16'(-2251);
			23122: out = 16'(-2869);
			23123: out = 16'(-2977);
			23124: out = 16'(-354);
			23125: out = 16'(1741);
			23126: out = 16'(1909);
			23127: out = 16'(1406);
			23128: out = 16'(540);
			23129: out = 16'(3181);
			23130: out = 16'(3259);
			23131: out = 16'(3099);
			23132: out = 16'(18);
			23133: out = 16'(-1096);
			23134: out = 16'(-1417);
			23135: out = 16'(-825);
			23136: out = 16'(-915);
			23137: out = 16'(-2343);
			23138: out = 16'(792);
			23139: out = 16'(1818);
			23140: out = 16'(264);
			23141: out = 16'(384);
			23142: out = 16'(55);
			23143: out = 16'(521);
			23144: out = 16'(-217);
			23145: out = 16'(-803);
			23146: out = 16'(-2103);
			23147: out = 16'(-2130);
			23148: out = 16'(-2176);
			23149: out = 16'(-1994);
			23150: out = 16'(-2131);
			23151: out = 16'(-1846);
			23152: out = 16'(-2178);
			23153: out = 16'(-1012);
			23154: out = 16'(424);
			23155: out = 16'(2884);
			23156: out = 16'(2678);
			23157: out = 16'(-281);
			23158: out = 16'(-1833);
			23159: out = 16'(-2213);
			23160: out = 16'(2386);
			23161: out = 16'(527);
			23162: out = 16'(-218);
			23163: out = 16'(-1325);
			23164: out = 16'(1256);
			23165: out = 16'(3393);
			23166: out = 16'(-1759);
			23167: out = 16'(-1331);
			23168: out = 16'(-199);
			23169: out = 16'(2326);
			23170: out = 16'(1766);
			23171: out = 16'(-829);
			23172: out = 16'(-219);
			23173: out = 16'(-919);
			23174: out = 16'(-1061);
			23175: out = 16'(-3123);
			23176: out = 16'(-2887);
			23177: out = 16'(-41);
			23178: out = 16'(393);
			23179: out = 16'(265);
			23180: out = 16'(-2738);
			23181: out = 16'(-1763);
			23182: out = 16'(-747);
			23183: out = 16'(354);
			23184: out = 16'(1031);
			23185: out = 16'(1499);
			23186: out = 16'(760);
			23187: out = 16'(420);
			23188: out = 16'(-175);
			23189: out = 16'(648);
			23190: out = 16'(527);
			23191: out = 16'(476);
			23192: out = 16'(-1389);
			23193: out = 16'(-2146);
			23194: out = 16'(-2747);
			23195: out = 16'(-321);
			23196: out = 16'(1345);
			23197: out = 16'(2914);
			23198: out = 16'(1463);
			23199: out = 16'(1131);
			23200: out = 16'(4635);
			23201: out = 16'(5426);
			23202: out = 16'(5321);
			23203: out = 16'(1014);
			23204: out = 16'(-2605);
			23205: out = 16'(-6568);
			23206: out = 16'(-128);
			23207: out = 16'(691);
			23208: out = 16'(1424);
			23209: out = 16'(-1661);
			23210: out = 16'(-1200);
			23211: out = 16'(480);
			23212: out = 16'(1825);
			23213: out = 16'(463);
			23214: out = 16'(-4535);
			23215: out = 16'(-5588);
			23216: out = 16'(-5337);
			23217: out = 16'(-1085);
			23218: out = 16'(-527);
			23219: out = 16'(-309);
			23220: out = 16'(-1604);
			23221: out = 16'(-2549);
			23222: out = 16'(-3167);
			23223: out = 16'(-1254);
			23224: out = 16'(1421);
			23225: out = 16'(4788);
			23226: out = 16'(2479);
			23227: out = 16'(1625);
			23228: out = 16'(-488);
			23229: out = 16'(2413);
			23230: out = 16'(2959);
			23231: out = 16'(3694);
			23232: out = 16'(-268);
			23233: out = 16'(-2685);
			23234: out = 16'(-4380);
			23235: out = 16'(-1353);
			23236: out = 16'(1637);
			23237: out = 16'(3214);
			23238: out = 16'(3698);
			23239: out = 16'(3152);
			23240: out = 16'(2249);
			23241: out = 16'(1231);
			23242: out = 16'(443);
			23243: out = 16'(1818);
			23244: out = 16'(1265);
			23245: out = 16'(-6);
			23246: out = 16'(-2210);
			23247: out = 16'(-3140);
			23248: out = 16'(-2715);
			23249: out = 16'(-1815);
			23250: out = 16'(-708);
			23251: out = 16'(-255);
			23252: out = 16'(288);
			23253: out = 16'(329);
			23254: out = 16'(407);
			23255: out = 16'(307);
			23256: out = 16'(378);
			23257: out = 16'(291);
			23258: out = 16'(374);
			23259: out = 16'(288);
			23260: out = 16'(632);
			23261: out = 16'(157);
			23262: out = 16'(-250);
			23263: out = 16'(-1087);
			23264: out = 16'(-876);
			23265: out = 16'(-105);
			23266: out = 16'(-371);
			23267: out = 16'(-433);
			23268: out = 16'(-377);
			23269: out = 16'(-266);
			23270: out = 16'(-87);
			23271: out = 16'(-494);
			23272: out = 16'(756);
			23273: out = 16'(1562);
			23274: out = 16'(2766);
			23275: out = 16'(1012);
			23276: out = 16'(-698);
			23277: out = 16'(-203);
			23278: out = 16'(641);
			23279: out = 16'(2107);
			23280: out = 16'(-205);
			23281: out = 16'(56);
			23282: out = 16'(352);
			23283: out = 16'(-112);
			23284: out = 16'(-2073);
			23285: out = 16'(-5594);
			23286: out = 16'(-1781);
			23287: out = 16'(369);
			23288: out = 16'(1220);
			23289: out = 16'(346);
			23290: out = 16'(-761);
			23291: out = 16'(-167);
			23292: out = 16'(-1579);
			23293: out = 16'(-1767);
			23294: out = 16'(-1470);
			23295: out = 16'(978);
			23296: out = 16'(2924);
			23297: out = 16'(2109);
			23298: out = 16'(1354);
			23299: out = 16'(496);
			23300: out = 16'(1671);
			23301: out = 16'(2065);
			23302: out = 16'(1678);
			23303: out = 16'(2145);
			23304: out = 16'(661);
			23305: out = 16'(-1291);
			23306: out = 16'(-5074);
			23307: out = 16'(-5637);
			23308: out = 16'(-2004);
			23309: out = 16'(5);
			23310: out = 16'(1837);
			23311: out = 16'(2597);
			23312: out = 16'(2316);
			23313: out = 16'(1726);
			23314: out = 16'(-385);
			23315: out = 16'(1747);
			23316: out = 16'(4079);
			23317: out = 16'(3395);
			23318: out = 16'(431);
			23319: out = 16'(-4599);
			23320: out = 16'(-4959);
			23321: out = 16'(-5406);
			23322: out = 16'(-3244);
			23323: out = 16'(-4084);
			23324: out = 16'(-2168);
			23325: out = 16'(590);
			23326: out = 16'(1373);
			23327: out = 16'(629);
			23328: out = 16'(-2649);
			23329: out = 16'(-2233);
			23330: out = 16'(-1803);
			23331: out = 16'(-2729);
			23332: out = 16'(-1303);
			23333: out = 16'(392);
			23334: out = 16'(3329);
			23335: out = 16'(3166);
			23336: out = 16'(2061);
			23337: out = 16'(3452);
			23338: out = 16'(3636);
			23339: out = 16'(4065);
			23340: out = 16'(612);
			23341: out = 16'(-1202);
			23342: out = 16'(-3011);
			23343: out = 16'(-1660);
			23344: out = 16'(-822);
			23345: out = 16'(747);
			23346: out = 16'(-244);
			23347: out = 16'(-170);
			23348: out = 16'(84);
			23349: out = 16'(2295);
			23350: out = 16'(3245);
			23351: out = 16'(2191);
			23352: out = 16'(-152);
			23353: out = 16'(-2438);
			23354: out = 16'(-2848);
			23355: out = 16'(-1815);
			23356: out = 16'(175);
			23357: out = 16'(3261);
			23358: out = 16'(4002);
			23359: out = 16'(3017);
			23360: out = 16'(-134);
			23361: out = 16'(-2019);
			23362: out = 16'(-2033);
			23363: out = 16'(-1765);
			23364: out = 16'(-1025);
			23365: out = 16'(-602);
			23366: out = 16'(-494);
			23367: out = 16'(-607);
			23368: out = 16'(-1320);
			23369: out = 16'(-241);
			23370: out = 16'(711);
			23371: out = 16'(1218);
			23372: out = 16'(544);
			23373: out = 16'(-319);
			23374: out = 16'(393);
			23375: out = 16'(800);
			23376: out = 16'(1238);
			23377: out = 16'(2380);
			23378: out = 16'(2323);
			23379: out = 16'(1764);
			23380: out = 16'(-1685);
			23381: out = 16'(-3727);
			23382: out = 16'(-4581);
			23383: out = 16'(-2540);
			23384: out = 16'(-621);
			23385: out = 16'(180);
			23386: out = 16'(157);
			23387: out = 16'(-222);
			23388: out = 16'(646);
			23389: out = 16'(435);
			23390: out = 16'(346);
			23391: out = 16'(361);
			23392: out = 16'(14);
			23393: out = 16'(-646);
			23394: out = 16'(-3088);
			23395: out = 16'(-3203);
			23396: out = 16'(-1578);
			23397: out = 16'(-1469);
			23398: out = 16'(-453);
			23399: out = 16'(-176);
			23400: out = 16'(1263);
			23401: out = 16'(910);
			23402: out = 16'(-966);
			23403: out = 16'(-1154);
			23404: out = 16'(-621);
			23405: out = 16'(303);
			23406: out = 16'(1955);
			23407: out = 16'(3072);
			23408: out = 16'(4192);
			23409: out = 16'(2749);
			23410: out = 16'(1053);
			23411: out = 16'(549);
			23412: out = 16'(1298);
			23413: out = 16'(2720);
			23414: out = 16'(2012);
			23415: out = 16'(1054);
			23416: out = 16'(-791);
			23417: out = 16'(-587);
			23418: out = 16'(-558);
			23419: out = 16'(-359);
			23420: out = 16'(29);
			23421: out = 16'(135);
			23422: out = 16'(241);
			23423: out = 16'(-820);
			23424: out = 16'(-1333);
			23425: out = 16'(-634);
			23426: out = 16'(-104);
			23427: out = 16'(175);
			23428: out = 16'(320);
			23429: out = 16'(-266);
			23430: out = 16'(-670);
			23431: out = 16'(-4966);
			23432: out = 16'(-3693);
			23433: out = 16'(61);
			23434: out = 16'(3025);
			23435: out = 16'(3644);
			23436: out = 16'(771);
			23437: out = 16'(-83);
			23438: out = 16'(-2872);
			23439: out = 16'(-5883);
			23440: out = 16'(-6443);
			23441: out = 16'(-4630);
			23442: out = 16'(482);
			23443: out = 16'(2487);
			23444: out = 16'(3665);
			23445: out = 16'(1321);
			23446: out = 16'(3162);
			23447: out = 16'(4882);
			23448: out = 16'(3518);
			23449: out = 16'(1922);
			23450: out = 16'(-631);
			23451: out = 16'(2366);
			23452: out = 16'(1683);
			23453: out = 16'(56);
			23454: out = 16'(-1688);
			23455: out = 16'(-1653);
			23456: out = 16'(598);
			23457: out = 16'(175);
			23458: out = 16'(-197);
			23459: out = 16'(-2299);
			23460: out = 16'(-1081);
			23461: out = 16'(-500);
			23462: out = 16'(-477);
			23463: out = 16'(-938);
			23464: out = 16'(-1376);
			23465: out = 16'(-1953);
			23466: out = 16'(-2021);
			23467: out = 16'(-1813);
			23468: out = 16'(276);
			23469: out = 16'(947);
			23470: out = 16'(1384);
			23471: out = 16'(-717);
			23472: out = 16'(-804);
			23473: out = 16'(501);
			23474: out = 16'(2462);
			23475: out = 16'(3656);
			23476: out = 16'(3091);
			23477: out = 16'(2584);
			23478: out = 16'(1080);
			23479: out = 16'(-106);
			23480: out = 16'(-2074);
			23481: out = 16'(-2961);
			23482: out = 16'(-2320);
			23483: out = 16'(-808);
			23484: out = 16'(722);
			23485: out = 16'(1045);
			23486: out = 16'(1228);
			23487: out = 16'(1216);
			23488: out = 16'(2891);
			23489: out = 16'(3076);
			23490: out = 16'(2153);
			23491: out = 16'(-202);
			23492: out = 16'(-3301);
			23493: out = 16'(-6196);
			23494: out = 16'(-6198);
			23495: out = 16'(-3629);
			23496: out = 16'(1004);
			23497: out = 16'(3745);
			23498: out = 16'(3847);
			23499: out = 16'(-887);
			23500: out = 16'(-4006);
			23501: out = 16'(-6333);
			23502: out = 16'(-4512);
			23503: out = 16'(-3240);
			23504: out = 16'(-1424);
			23505: out = 16'(-244);
			23506: out = 16'(380);
			23507: out = 16'(646);
			23508: out = 16'(-859);
			23509: out = 16'(705);
			23510: out = 16'(4597);
			23511: out = 16'(3693);
			23512: out = 16'(2635);
			23513: out = 16'(-543);
			23514: out = 16'(192);
			23515: out = 16'(334);
			23516: out = 16'(-241);
			23517: out = 16'(1512);
			23518: out = 16'(2939);
			23519: out = 16'(2604);
			23520: out = 16'(1552);
			23521: out = 16'(-106);
			23522: out = 16'(697);
			23523: out = 16'(-194);
			23524: out = 16'(-587);
			23525: out = 16'(-2705);
			23526: out = 16'(-2005);
			23527: out = 16'(-69);
			23528: out = 16'(-1042);
			23529: out = 16'(-1645);
			23530: out = 16'(-2878);
			23531: out = 16'(-1095);
			23532: out = 16'(83);
			23533: out = 16'(533);
			23534: out = 16'(2060);
			23535: out = 16'(2155);
			23536: out = 16'(-2864);
			23537: out = 16'(-1745);
			23538: out = 16'(-1038);
			23539: out = 16'(848);
			23540: out = 16'(-1771);
			23541: out = 16'(-4500);
			23542: out = 16'(-2145);
			23543: out = 16'(-447);
			23544: out = 16'(1842);
			23545: out = 16'(1303);
			23546: out = 16'(2236);
			23547: out = 16'(3591);
			23548: out = 16'(799);
			23549: out = 16'(-554);
			23550: out = 16'(-1121);
			23551: out = 16'(1031);
			23552: out = 16'(1948);
			23553: out = 16'(-601);
			23554: out = 16'(-101);
			23555: out = 16'(365);
			23556: out = 16'(5433);
			23557: out = 16'(2679);
			23558: out = 16'(164);
			23559: out = 16'(396);
			23560: out = 16'(1862);
			23561: out = 16'(3999);
			23562: out = 16'(-178);
			23563: out = 16'(-1269);
			23564: out = 16'(-2434);
			23565: out = 16'(-155);
			23566: out = 16'(-773);
			23567: out = 16'(-3079);
			23568: out = 16'(-2955);
			23569: out = 16'(-2123);
			23570: out = 16'(647);
			23571: out = 16'(0);
			23572: out = 16'(-487);
			23573: out = 16'(-2009);
			23574: out = 16'(-2005);
			23575: out = 16'(-1758);
			23576: out = 16'(-171);
			23577: out = 16'(225);
			23578: out = 16'(499);
			23579: out = 16'(-3150);
			23580: out = 16'(-3538);
			23581: out = 16'(-3258);
			23582: out = 16'(1344);
			23583: out = 16'(2627);
			23584: out = 16'(2922);
			23585: out = 16'(942);
			23586: out = 16'(1191);
			23587: out = 16'(3610);
			23588: out = 16'(2986);
			23589: out = 16'(1687);
			23590: out = 16'(-2069);
			23591: out = 16'(-2104);
			23592: out = 16'(-1695);
			23593: out = 16'(-335);
			23594: out = 16'(1408);
			23595: out = 16'(2805);
			23596: out = 16'(1305);
			23597: out = 16'(220);
			23598: out = 16'(-1503);
			23599: out = 16'(535);
			23600: out = 16'(273);
			23601: out = 16'(346);
			23602: out = 16'(-2448);
			23603: out = 16'(-2055);
			23604: out = 16'(-33);
			23605: out = 16'(1392);
			23606: out = 16'(1706);
			23607: out = 16'(-470);
			23608: out = 16'(371);
			23609: out = 16'(-269);
			23610: out = 16'(-1869);
			23611: out = 16'(-2607);
			23612: out = 16'(-2425);
			23613: out = 16'(-569);
			23614: out = 16'(143);
			23615: out = 16'(272);
			23616: out = 16'(-874);
			23617: out = 16'(-1225);
			23618: out = 16'(-1030);
			23619: out = 16'(-2529);
			23620: out = 16'(-2512);
			23621: out = 16'(-2559);
			23622: out = 16'(2370);
			23623: out = 16'(4051);
			23624: out = 16'(4251);
			23625: out = 16'(1569);
			23626: out = 16'(217);
			23627: out = 16'(692);
			23628: out = 16'(1418);
			23629: out = 16'(2364);
			23630: out = 16'(3294);
			23631: out = 16'(2968);
			23632: out = 16'(1835);
			23633: out = 16'(-4271);
			23634: out = 16'(-3566);
			23635: out = 16'(-1530);
			23636: out = 16'(3398);
			23637: out = 16'(2512);
			23638: out = 16'(-776);
			23639: out = 16'(-2262);
			23640: out = 16'(-2342);
			23641: out = 16'(138);
			23642: out = 16'(-56);
			23643: out = 16'(328);
			23644: out = 16'(-723);
			23645: out = 16'(-96);
			23646: out = 16'(-276);
			23647: out = 16'(757);
			23648: out = 16'(-1127);
			23649: out = 16'(-2141);
			23650: out = 16'(-2038);
			23651: out = 16'(-1148);
			23652: out = 16'(-179);
			23653: out = 16'(-430);
			23654: out = 16'(77);
			23655: out = 16'(532);
			23656: out = 16'(1287);
			23657: out = 16'(1169);
			23658: out = 16'(507);
			23659: out = 16'(-57);
			23660: out = 16'(-461);
			23661: out = 16'(50);
			23662: out = 16'(-470);
			23663: out = 16'(-102);
			23664: out = 16'(-383);
			23665: out = 16'(2779);
			23666: out = 16'(3809);
			23667: out = 16'(1319);
			23668: out = 16'(-151);
			23669: out = 16'(-1152);
			23670: out = 16'(1884);
			23671: out = 16'(1887);
			23672: out = 16'(1753);
			23673: out = 16'(-103);
			23674: out = 16'(-428);
			23675: out = 16'(-419);
			23676: out = 16'(-2385);
			23677: out = 16'(-3779);
			23678: out = 16'(-5481);
			23679: out = 16'(-1604);
			23680: out = 16'(535);
			23681: out = 16'(2161);
			23682: out = 16'(589);
			23683: out = 16'(-679);
			23684: out = 16'(-2797);
			23685: out = 16'(-1197);
			23686: out = 16'(-267);
			23687: out = 16'(-142);
			23688: out = 16'(-2385);
			23689: out = 16'(-4332);
			23690: out = 16'(-3333);
			23691: out = 16'(-1561);
			23692: out = 16'(1051);
			23693: out = 16'(676);
			23694: out = 16'(1012);
			23695: out = 16'(771);
			23696: out = 16'(881);
			23697: out = 16'(968);
			23698: out = 16'(1552);
			23699: out = 16'(1479);
			23700: out = 16'(1089);
			23701: out = 16'(-257);
			23702: out = 16'(-736);
			23703: out = 16'(-651);
			23704: out = 16'(1479);
			23705: out = 16'(1728);
			23706: out = 16'(2092);
			23707: out = 16'(543);
			23708: out = 16'(1407);
			23709: out = 16'(1900);
			23710: out = 16'(830);
			23711: out = 16'(-219);
			23712: out = 16'(-1137);
			23713: out = 16'(-23);
			23714: out = 16'(1234);
			23715: out = 16'(2651);
			23716: out = 16'(2162);
			23717: out = 16'(844);
			23718: out = 16'(-2176);
			23719: out = 16'(-1439);
			23720: out = 16'(-757);
			23721: out = 16'(1330);
			23722: out = 16'(254);
			23723: out = 16'(-376);
			23724: out = 16'(-1241);
			23725: out = 16'(-250);
			23726: out = 16'(555);
			23727: out = 16'(-345);
			23728: out = 16'(-1112);
			23729: out = 16'(-2012);
			23730: out = 16'(-531);
			23731: out = 16'(-398);
			23732: out = 16'(-356);
			23733: out = 16'(-1007);
			23734: out = 16'(-698);
			23735: out = 16'(506);
			23736: out = 16'(-60);
			23737: out = 16'(-110);
			23738: out = 16'(-207);
			23739: out = 16'(1215);
			23740: out = 16'(2372);
			23741: out = 16'(3168);
			23742: out = 16'(2185);
			23743: out = 16'(539);
			23744: out = 16'(-885);
			23745: out = 16'(-2655);
			23746: out = 16'(-3552);
			23747: out = 16'(-2238);
			23748: out = 16'(-1215);
			23749: out = 16'(-424);
			23750: out = 16'(-2207);
			23751: out = 16'(-3071);
			23752: out = 16'(-3187);
			23753: out = 16'(-459);
			23754: out = 16'(2299);
			23755: out = 16'(4613);
			23756: out = 16'(4525);
			23757: out = 16'(2811);
			23758: out = 16'(39);
			23759: out = 16'(-2899);
			23760: out = 16'(-4645);
			23761: out = 16'(-5211);
			23762: out = 16'(-2153);
			23763: out = 16'(1241);
			23764: out = 16'(1786);
			23765: out = 16'(2365);
			23766: out = 16'(1823);
			23767: out = 16'(983);
			23768: out = 16'(-138);
			23769: out = 16'(-1155);
			23770: out = 16'(-453);
			23771: out = 16'(-157);
			23772: out = 16'(545);
			23773: out = 16'(-870);
			23774: out = 16'(-574);
			23775: out = 16'(599);
			23776: out = 16'(2135);
			23777: out = 16'(2321);
			23778: out = 16'(425);
			23779: out = 16'(-644);
			23780: out = 16'(-835);
			23781: out = 16'(1065);
			23782: out = 16'(2744);
			23783: out = 16'(3910);
			23784: out = 16'(2681);
			23785: out = 16'(1452);
			23786: out = 16'(-256);
			23787: out = 16'(-3809);
			23788: out = 16'(-3884);
			23789: out = 16'(-1655);
			23790: out = 16'(-796);
			23791: out = 16'(75);
			23792: out = 16'(-344);
			23793: out = 16'(1408);
			23794: out = 16'(2469);
			23795: out = 16'(3883);
			23796: out = 16'(3071);
			23797: out = 16'(1192);
			23798: out = 16'(-4393);
			23799: out = 16'(-4567);
			23800: out = 16'(-3982);
			23801: out = 16'(-345);
			23802: out = 16'(-636);
			23803: out = 16'(-1255);
			23804: out = 16'(-2586);
			23805: out = 16'(-1441);
			23806: out = 16'(717);
			23807: out = 16'(-114);
			23808: out = 16'(-36);
			23809: out = 16'(-367);
			23810: out = 16'(516);
			23811: out = 16'(1003);
			23812: out = 16'(2168);
			23813: out = 16'(970);
			23814: out = 16'(408);
			23815: out = 16'(-459);
			23816: out = 16'(89);
			23817: out = 16'(640);
			23818: out = 16'(2769);
			23819: out = 16'(930);
			23820: out = 16'(-921);
			23821: out = 16'(-3375);
			23822: out = 16'(-2193);
			23823: out = 16'(-36);
			23824: out = 16'(-312);
			23825: out = 16'(506);
			23826: out = 16'(1362);
			23827: out = 16'(-672);
			23828: out = 16'(-1385);
			23829: out = 16'(-1939);
			23830: out = 16'(1668);
			23831: out = 16'(2253);
			23832: out = 16'(-293);
			23833: out = 16'(-1172);
			23834: out = 16'(-1788);
			23835: out = 16'(67);
			23836: out = 16'(184);
			23837: out = 16'(794);
			23838: out = 16'(-243);
			23839: out = 16'(459);
			23840: out = 16'(411);
			23841: out = 16'(-692);
			23842: out = 16'(-1869);
			23843: out = 16'(-2544);
			23844: out = 16'(-2588);
			23845: out = 16'(-2361);
			23846: out = 16'(-2474);
			23847: out = 16'(19);
			23848: out = 16'(991);
			23849: out = 16'(1692);
			23850: out = 16'(853);
			23851: out = 16'(1512);
			23852: out = 16'(3389);
			23853: out = 16'(4035);
			23854: out = 16'(3539);
			23855: out = 16'(2321);
			23856: out = 16'(-710);
			23857: out = 16'(-3099);
			23858: out = 16'(-4277);
			23859: out = 16'(-1662);
			23860: out = 16'(1858);
			23861: out = 16'(347);
			23862: out = 16'(286);
			23863: out = 16'(-430);
			23864: out = 16'(-8);
			23865: out = 16'(60);
			23866: out = 16'(501);
			23867: out = 16'(409);
			23868: out = 16'(313);
			23869: out = 16'(-55);
			23870: out = 16'(-172);
			23871: out = 16'(158);
			23872: out = 16'(430);
			23873: out = 16'(2797);
			23874: out = 16'(3279);
			23875: out = 16'(-2382);
			23876: out = 16'(-3990);
			23877: out = 16'(-4711);
			23878: out = 16'(1560);
			23879: out = 16'(2158);
			23880: out = 16'(1983);
			23881: out = 16'(680);
			23882: out = 16'(70);
			23883: out = 16'(-431);
			23884: out = 16'(-289);
			23885: out = 16'(-819);
			23886: out = 16'(-1902);
			23887: out = 16'(-1285);
			23888: out = 16'(-763);
			23889: out = 16'(-31);
			23890: out = 16'(363);
			23891: out = 16'(1114);
			23892: out = 16'(2629);
			23893: out = 16'(2743);
			23894: out = 16'(2514);
			23895: out = 16'(2010);
			23896: out = 16'(1552);
			23897: out = 16'(757);
			23898: out = 16'(-2866);
			23899: out = 16'(-4706);
			23900: out = 16'(-5842);
			23901: out = 16'(-1998);
			23902: out = 16'(-183);
			23903: out = 16'(713);
			23904: out = 16'(196);
			23905: out = 16'(-100);
			23906: out = 16'(60);
			23907: out = 16'(-737);
			23908: out = 16'(-451);
			23909: out = 16'(2225);
			23910: out = 16'(1629);
			23911: out = 16'(835);
			23912: out = 16'(-3379);
			23913: out = 16'(-1748);
			23914: out = 16'(200);
			23915: out = 16'(2573);
			23916: out = 16'(1839);
			23917: out = 16'(52);
			23918: out = 16'(-2814);
			23919: out = 16'(-2274);
			23920: out = 16'(938);
			23921: out = 16'(-1643);
			23922: out = 16'(-983);
			23923: out = 16'(498);
			23924: out = 16'(1255);
			23925: out = 16'(1092);
			23926: out = 16'(-339);
			23927: out = 16'(247);
			23928: out = 16'(118);
			23929: out = 16'(-1803);
			23930: out = 16'(-1725);
			23931: out = 16'(-1641);
			23932: out = 16'(-142);
			23933: out = 16'(-975);
			23934: out = 16'(-1375);
			23935: out = 16'(2324);
			23936: out = 16'(3817);
			23937: out = 16'(4660);
			23938: out = 16'(1381);
			23939: out = 16'(103);
			23940: out = 16'(-299);
			23941: out = 16'(-1018);
			23942: out = 16'(-1058);
			23943: out = 16'(-1130);
			23944: out = 16'(1138);
			23945: out = 16'(2102);
			23946: out = 16'(1228);
			23947: out = 16'(500);
			23948: out = 16'(-42);
			23949: out = 16'(2808);
			23950: out = 16'(972);
			23951: out = 16'(-364);
			23952: out = 16'(-263);
			23953: out = 16'(119);
			23954: out = 16'(443);
			23955: out = 16'(-259);
			23956: out = 16'(-863);
			23957: out = 16'(-1241);
			23958: out = 16'(-3828);
			23959: out = 16'(-3487);
			23960: out = 16'(-780);
			23961: out = 16'(575);
			23962: out = 16'(1413);
			23963: out = 16'(-434);
			23964: out = 16'(1586);
			23965: out = 16'(2036);
			23966: out = 16'(2899);
			23967: out = 16'(359);
			23968: out = 16'(-1629);
			23969: out = 16'(-3441);
			23970: out = 16'(-1978);
			23971: out = 16'(-1);
			23972: out = 16'(234);
			23973: out = 16'(499);
			23974: out = 16'(343);
			23975: out = 16'(-859);
			23976: out = 16'(-758);
			23977: out = 16'(20);
			23978: out = 16'(1610);
			23979: out = 16'(1382);
			23980: out = 16'(-1329);
			23981: out = 16'(-937);
			23982: out = 16'(-1037);
			23983: out = 16'(161);
			23984: out = 16'(-1744);
			23985: out = 16'(-2275);
			23986: out = 16'(-47);
			23987: out = 16'(1037);
			23988: out = 16'(2467);
			23989: out = 16'(1741);
			23990: out = 16'(3515);
			23991: out = 16'(4371);
			23992: out = 16'(2494);
			23993: out = 16'(132);
			23994: out = 16'(-2236);
			23995: out = 16'(-4722);
			23996: out = 16'(-4547);
			23997: out = 16'(-2424);
			23998: out = 16'(-1011);
			23999: out = 16'(180);
			24000: out = 16'(677);
			24001: out = 16'(579);
			24002: out = 16'(264);
			24003: out = 16'(-1206);
			24004: out = 16'(1321);
			24005: out = 16'(3005);
			24006: out = 16'(3396);
			24007: out = 16'(1810);
			24008: out = 16'(-23);
			24009: out = 16'(-1131);
			24010: out = 16'(367);
			24011: out = 16'(2925);
			24012: out = 16'(2406);
			24013: out = 16'(1907);
			24014: out = 16'(83);
			24015: out = 16'(-78);
			24016: out = 16'(-1830);
			24017: out = 16'(-4551);
			24018: out = 16'(-1502);
			24019: out = 16'(521);
			24020: out = 16'(1878);
			24021: out = 16'(56);
			24022: out = 16'(-1457);
			24023: out = 16'(-279);
			24024: out = 16'(-243);
			24025: out = 16'(262);
			24026: out = 16'(-2878);
			24027: out = 16'(-1109);
			24028: out = 16'(405);
			24029: out = 16'(492);
			24030: out = 16'(-919);
			24031: out = 16'(-2703);
			24032: out = 16'(31);
			24033: out = 16'(1081);
			24034: out = 16'(1155);
			24035: out = 16'(1535);
			24036: out = 16'(664);
			24037: out = 16'(32);
			24038: out = 16'(-3692);
			24039: out = 16'(-5266);
			24040: out = 16'(-5167);
			24041: out = 16'(-634);
			24042: out = 16'(2626);
			24043: out = 16'(324);
			24044: out = 16'(738);
			24045: out = 16'(507);
			24046: out = 16'(1480);
			24047: out = 16'(1392);
			24048: out = 16'(1495);
			24049: out = 16'(2536);
			24050: out = 16'(2710);
			24051: out = 16'(2563);
			24052: out = 16'(-375);
			24053: out = 16'(-1405);
			24054: out = 16'(-1111);
			24055: out = 16'(-453);
			24056: out = 16'(0);
			24057: out = 16'(398);
			24058: out = 16'(-233);
			24059: out = 16'(-334);
			24060: out = 16'(-576);
			24061: out = 16'(1438);
			24062: out = 16'(3018);
			24063: out = 16'(5072);
			24064: out = 16'(3069);
			24065: out = 16'(572);
			24066: out = 16'(-1779);
			24067: out = 16'(-1337);
			24068: out = 16'(312);
			24069: out = 16'(-254);
			24070: out = 16'(-988);
			24071: out = 16'(-2098);
			24072: out = 16'(-2860);
			24073: out = 16'(-1258);
			24074: out = 16'(2714);
			24075: out = 16'(4292);
			24076: out = 16'(4215);
			24077: out = 16'(-73);
			24078: out = 16'(-1109);
			24079: out = 16'(-2457);
			24080: out = 16'(-1082);
			24081: out = 16'(-1975);
			24082: out = 16'(-2064);
			24083: out = 16'(-3713);
			24084: out = 16'(-2389);
			24085: out = 16'(-902);
			24086: out = 16'(1041);
			24087: out = 16'(797);
			24088: out = 16'(-282);
			24089: out = 16'(-310);
			24090: out = 16'(-121);
			24091: out = 16'(629);
			24092: out = 16'(589);
			24093: out = 16'(-317);
			24094: out = 16'(-3727);
			24095: out = 16'(-2284);
			24096: out = 16'(-1584);
			24097: out = 16'(138);
			24098: out = 16'(-1625);
			24099: out = 16'(-2390);
			24100: out = 16'(-1166);
			24101: out = 16'(711);
			24102: out = 16'(2278);
			24103: out = 16'(774);
			24104: out = 16'(698);
			24105: out = 16'(704);
			24106: out = 16'(591);
			24107: out = 16'(961);
			24108: out = 16'(1316);
			24109: out = 16'(1434);
			24110: out = 16'(1001);
			24111: out = 16'(683);
			24112: out = 16'(-1713);
			24113: out = 16'(-3051);
			24114: out = 16'(-4300);
			24115: out = 16'(179);
			24116: out = 16'(3710);
			24117: out = 16'(4404);
			24118: out = 16'(3471);
			24119: out = 16'(1519);
			24120: out = 16'(2952);
			24121: out = 16'(945);
			24122: out = 16'(-415);
			24123: out = 16'(-1929);
			24124: out = 16'(-1292);
			24125: out = 16'(-180);
			24126: out = 16'(-306);
			24127: out = 16'(-1668);
			24128: out = 16'(-4527);
			24129: out = 16'(-1885);
			24130: out = 16'(-318);
			24131: out = 16'(1427);
			24132: out = 16'(408);
			24133: out = 16'(-621);
			24134: out = 16'(-2578);
			24135: out = 16'(-2170);
			24136: out = 16'(-1121);
			24137: out = 16'(2695);
			24138: out = 16'(1738);
			24139: out = 16'(322);
			24140: out = 16'(-1548);
			24141: out = 16'(-877);
			24142: out = 16'(1041);
			24143: out = 16'(372);
			24144: out = 16'(1615);
			24145: out = 16'(2665);
			24146: out = 16'(3366);
			24147: out = 16'(1796);
			24148: out = 16'(-2240);
			24149: out = 16'(-1316);
			24150: out = 16'(-589);
			24151: out = 16'(2240);
			24152: out = 16'(-1088);
			24153: out = 16'(-3284);
			24154: out = 16'(-5121);
			24155: out = 16'(-2061);
			24156: out = 16'(686);
			24157: out = 16'(-3484);
			24158: out = 16'(-1644);
			24159: out = 16'(316);
			24160: out = 16'(4274);
			24161: out = 16'(4165);
			24162: out = 16'(2372);
			24163: out = 16'(1116);
			24164: out = 16'(-662);
			24165: out = 16'(-1783);
			24166: out = 16'(-2588);
			24167: out = 16'(-1778);
			24168: out = 16'(519);
			24169: out = 16'(179);
			24170: out = 16'(-279);
			24171: out = 16'(-898);
			24172: out = 16'(-1543);
			24173: out = 16'(-1474);
			24174: out = 16'(-91);
			24175: out = 16'(812);
			24176: out = 16'(1504);
			24177: out = 16'(594);
			24178: out = 16'(277);
			24179: out = 16'(-42);
			24180: out = 16'(-18);
			24181: out = 16'(-69);
			24182: out = 16'(-200);
			24183: out = 16'(1581);
			24184: out = 16'(2736);
			24185: out = 16'(4102);
			24186: out = 16'(1472);
			24187: out = 16'(475);
			24188: out = 16'(1286);
			24189: out = 16'(1650);
			24190: out = 16'(1223);
			24191: out = 16'(-2755);
			24192: out = 16'(-3192);
			24193: out = 16'(-3035);
			24194: out = 16'(2437);
			24195: out = 16'(2206);
			24196: out = 16'(1580);
			24197: out = 16'(-3834);
			24198: out = 16'(-3787);
			24199: out = 16'(-2446);
			24200: out = 16'(1272);
			24201: out = 16'(1657);
			24202: out = 16'(219);
			24203: out = 16'(-1363);
			24204: out = 16'(-1461);
			24205: out = 16'(513);
			24206: out = 16'(360);
			24207: out = 16'(66);
			24208: out = 16'(-1057);
			24209: out = 16'(-2106);
			24210: out = 16'(-2426);
			24211: out = 16'(-1205);
			24212: out = 16'(1029);
			24213: out = 16'(3045);
			24214: out = 16'(2006);
			24215: out = 16'(1425);
			24216: out = 16'(135);
			24217: out = 16'(737);
			24218: out = 16'(354);
			24219: out = 16'(487);
			24220: out = 16'(886);
			24221: out = 16'(2164);
			24222: out = 16'(3925);
			24223: out = 16'(1908);
			24224: out = 16'(353);
			24225: out = 16'(-1318);
			24226: out = 16'(-896);
			24227: out = 16'(-494);
			24228: out = 16'(-599);
			24229: out = 16'(-525);
			24230: out = 16'(-504);
			24231: out = 16'(-289);
			24232: out = 16'(-44);
			24233: out = 16'(387);
			24234: out = 16'(1012);
			24235: out = 16'(949);
			24236: out = 16'(92);
			24237: out = 16'(-1363);
			24238: out = 16'(-3698);
			24239: out = 16'(-6037);
			24240: out = 16'(-4836);
			24241: out = 16'(-2981);
			24242: out = 16'(-113);
			24243: out = 16'(256);
			24244: out = 16'(600);
			24245: out = 16'(499);
			24246: out = 16'(220);
			24247: out = 16'(248);
			24248: out = 16'(2189);
			24249: out = 16'(934);
			24250: out = 16'(-528);
			24251: out = 16'(-2275);
			24252: out = 16'(-2421);
			24253: out = 16'(-1261);
			24254: out = 16'(98);
			24255: out = 16'(3098);
			24256: out = 16'(6107);
			24257: out = 16'(4820);
			24258: out = 16'(4102);
			24259: out = 16'(3073);
			24260: out = 16'(2263);
			24261: out = 16'(663);
			24262: out = 16'(-2325);
			24263: out = 16'(-2087);
			24264: out = 16'(-1564);
			24265: out = 16'(2194);
			24266: out = 16'(-1241);
			24267: out = 16'(-3018);
			24268: out = 16'(-3925);
			24269: out = 16'(785);
			24270: out = 16'(5025);
			24271: out = 16'(3124);
			24272: out = 16'(1364);
			24273: out = 16'(-1880);
			24274: out = 16'(322);
			24275: out = 16'(-645);
			24276: out = 16'(-1304);
			24277: out = 16'(-2674);
			24278: out = 16'(-2199);
			24279: out = 16'(-353);
			24280: out = 16'(-1659);
			24281: out = 16'(-2009);
			24282: out = 16'(-1988);
			24283: out = 16'(-421);
			24284: out = 16'(467);
			24285: out = 16'(-152);
			24286: out = 16'(-632);
			24287: out = 16'(-1049);
			24288: out = 16'(358);
			24289: out = 16'(1146);
			24290: out = 16'(2166);
			24291: out = 16'(477);
			24292: out = 16'(1266);
			24293: out = 16'(1951);
			24294: out = 16'(3179);
			24295: out = 16'(2231);
			24296: out = 16'(259);
			24297: out = 16'(-267);
			24298: out = 16'(-368);
			24299: out = 16'(504);
			24300: out = 16'(359);
			24301: out = 16'(274);
			24302: out = 16'(-381);
			24303: out = 16'(-805);
			24304: out = 16'(-1792);
			24305: out = 16'(-3399);
			24306: out = 16'(-4097);
			24307: out = 16'(-3965);
			24308: out = 16'(-1348);
			24309: out = 16'(-299);
			24310: out = 16'(417);
			24311: out = 16'(-2992);
			24312: out = 16'(-2486);
			24313: out = 16'(-632);
			24314: out = 16'(946);
			24315: out = 16'(1502);
			24316: out = 16'(563);
			24317: out = 16'(786);
			24318: out = 16'(231);
			24319: out = 16'(149);
			24320: out = 16'(-786);
			24321: out = 16'(-661);
			24322: out = 16'(424);
			24323: out = 16'(1125);
			24324: out = 16'(1431);
			24325: out = 16'(1452);
			24326: out = 16'(901);
			24327: out = 16'(259);
			24328: out = 16'(-965);
			24329: out = 16'(-480);
			24330: out = 16'(755);
			24331: out = 16'(3946);
			24332: out = 16'(4397);
			24333: out = 16'(2862);
			24334: out = 16'(780);
			24335: out = 16'(-835);
			24336: out = 16'(109);
			24337: out = 16'(-3558);
			24338: out = 16'(-3555);
			24339: out = 16'(-536);
			24340: out = 16'(1616);
			24341: out = 16'(2220);
			24342: out = 16'(-1110);
			24343: out = 16'(-1642);
			24344: out = 16'(-1786);
			24345: out = 16'(-290);
			24346: out = 16'(173);
			24347: out = 16'(186);
			24348: out = 16'(-1495);
			24349: out = 16'(-2346);
			24350: out = 16'(-2476);
			24351: out = 16'(-3465);
			24352: out = 16'(-2099);
			24353: out = 16'(129);
			24354: out = 16'(2712);
			24355: out = 16'(2833);
			24356: out = 16'(-229);
			24357: out = 16'(424);
			24358: out = 16'(401);
			24359: out = 16'(-123);
			24360: out = 16'(847);
			24361: out = 16'(1294);
			24362: out = 16'(551);
			24363: out = 16'(-128);
			24364: out = 16'(-1);
			24365: out = 16'(1539);
			24366: out = 16'(3624);
			24367: out = 16'(5003);
			24368: out = 16'(4290);
			24369: out = 16'(1725);
			24370: out = 16'(-1503);
			24371: out = 16'(-2778);
			24372: out = 16'(-1316);
			24373: out = 16'(2601);
			24374: out = 16'(4291);
			24375: out = 16'(3939);
			24376: out = 16'(-32);
			24377: out = 16'(-3332);
			24378: out = 16'(-5548);
			24379: out = 16'(-1880);
			24380: out = 16'(-2400);
			24381: out = 16'(-1883);
			24382: out = 16'(-3039);
			24383: out = 16'(-1411);
			24384: out = 16'(7);
			24385: out = 16'(1073);
			24386: out = 16'(990);
			24387: out = 16'(115);
			24388: out = 16'(-186);
			24389: out = 16'(-556);
			24390: out = 16'(-15);
			24391: out = 16'(-2288);
			24392: out = 16'(-2109);
			24393: out = 16'(-384);
			24394: out = 16'(1323);
			24395: out = 16'(1825);
			24396: out = 16'(577);
			24397: out = 16'(-881);
			24398: out = 16'(-2142);
			24399: out = 16'(-1860);
			24400: out = 16'(-782);
			24401: out = 16'(563);
			24402: out = 16'(-1151);
			24403: out = 16'(-643);
			24404: out = 16'(-285);
			24405: out = 16'(379);
			24406: out = 16'(276);
			24407: out = 16'(-59);
			24408: out = 16'(1015);
			24409: out = 16'(1828);
			24410: out = 16'(2716);
			24411: out = 16'(1151);
			24412: out = 16'(34);
			24413: out = 16'(-1192);
			24414: out = 16'(-236);
			24415: out = 16'(387);
			24416: out = 16'(-259);
			24417: out = 16'(-133);
			24418: out = 16'(-180);
			24419: out = 16'(409);
			24420: out = 16'(-787);
			24421: out = 16'(-1973);
			24422: out = 16'(237);
			24423: out = 16'(393);
			24424: out = 16'(643);
			24425: out = 16'(-1646);
			24426: out = 16'(-1135);
			24427: out = 16'(527);
			24428: out = 16'(2652);
			24429: out = 16'(2958);
			24430: out = 16'(1015);
			24431: out = 16'(1271);
			24432: out = 16'(1677);
			24433: out = 16'(4691);
			24434: out = 16'(1297);
			24435: out = 16'(-1574);
			24436: out = 16'(-4298);
			24437: out = 16'(-3421);
			24438: out = 16'(-1824);
			24439: out = 16'(-4622);
			24440: out = 16'(-1898);
			24441: out = 16'(986);
			24442: out = 16'(2398);
			24443: out = 16'(1745);
			24444: out = 16'(-516);
			24445: out = 16'(-64);
			24446: out = 16'(-1501);
			24447: out = 16'(-3515);
			24448: out = 16'(-1285);
			24449: out = 16'(958);
			24450: out = 16'(4123);
			24451: out = 16'(1803);
			24452: out = 16'(-514);
			24453: out = 16'(-4270);
			24454: out = 16'(-1712);
			24455: out = 16'(1139);
			24456: out = 16'(1668);
			24457: out = 16'(1978);
			24458: out = 16'(778);
			24459: out = 16'(208);
			24460: out = 16'(-2386);
			24461: out = 16'(-4250);
			24462: out = 16'(-3077);
			24463: out = 16'(-1420);
			24464: out = 16'(34);
			24465: out = 16'(2813);
			24466: out = 16'(3130);
			24467: out = 16'(2017);
			24468: out = 16'(-197);
			24469: out = 16'(-1087);
			24470: out = 16'(-83);
			24471: out = 16'(1168);
			24472: out = 16'(2050);
			24473: out = 16'(1234);
			24474: out = 16'(503);
			24475: out = 16'(-513);
			24476: out = 16'(-1839);
			24477: out = 16'(-983);
			24478: out = 16'(652);
			24479: out = 16'(1033);
			24480: out = 16'(742);
			24481: out = 16'(-630);
			24482: out = 16'(325);
			24483: out = 16'(64);
			24484: out = 16'(-104);
			24485: out = 16'(-427);
			24486: out = 16'(-104);
			24487: out = 16'(525);
			24488: out = 16'(967);
			24489: out = 16'(1143);
			24490: out = 16'(370);
			24491: out = 16'(1701);
			24492: out = 16'(2410);
			24493: out = 16'(1042);
			24494: out = 16'(710);
			24495: out = 16'(-272);
			24496: out = 16'(-1602);
			24497: out = 16'(-3558);
			24498: out = 16'(-5025);
			24499: out = 16'(-1779);
			24500: out = 16'(171);
			24501: out = 16'(2114);
			24502: out = 16'(1273);
			24503: out = 16'(882);
			24504: out = 16'(-401);
			24505: out = 16'(1932);
			24506: out = 16'(2064);
			24507: out = 16'(392);
			24508: out = 16'(-1016);
			24509: out = 16'(-2615);
			24510: out = 16'(-4042);
			24511: out = 16'(-4769);
			24512: out = 16'(-4311);
			24513: out = 16'(199);
			24514: out = 16'(672);
			24515: out = 16'(621);
			24516: out = 16'(-1502);
			24517: out = 16'(-1620);
			24518: out = 16'(-1570);
			24519: out = 16'(2200);
			24520: out = 16'(2575);
			24521: out = 16'(2061);
			24522: out = 16'(-2065);
			24523: out = 16'(-2879);
			24524: out = 16'(-705);
			24525: out = 16'(1462);
			24526: out = 16'(3470);
			24527: out = 16'(4445);
			24528: out = 16'(3081);
			24529: out = 16'(1196);
			24530: out = 16'(-954);
			24531: out = 16'(-25);
			24532: out = 16'(1561);
			24533: out = 16'(1657);
			24534: out = 16'(989);
			24535: out = 16'(-896);
			24536: out = 16'(-187);
			24537: out = 16'(-691);
			24538: out = 16'(-10);
			24539: out = 16'(-3159);
			24540: out = 16'(-2399);
			24541: out = 16'(-341);
			24542: out = 16'(2854);
			24543: out = 16'(3375);
			24544: out = 16'(975);
			24545: out = 16'(298);
			24546: out = 16'(-331);
			24547: out = 16'(534);
			24548: out = 16'(-33);
			24549: out = 16'(-398);
			24550: out = 16'(-387);
			24551: out = 16'(-1655);
			24552: out = 16'(-2963);
			24553: out = 16'(-4059);
			24554: out = 16'(-3544);
			24555: out = 16'(-2365);
			24556: out = 16'(-2471);
			24557: out = 16'(-3119);
			24558: out = 16'(-4771);
			24559: out = 16'(-1026);
			24560: out = 16'(1079);
			24561: out = 16'(3020);
			24562: out = 16'(2397);
			24563: out = 16'(2328);
			24564: out = 16'(2801);
			24565: out = 16'(2382);
			24566: out = 16'(1639);
			24567: out = 16'(-176);
			24568: out = 16'(-304);
			24569: out = 16'(-87);
			24570: out = 16'(1235);
			24571: out = 16'(1917);
			24572: out = 16'(2600);
			24573: out = 16'(-169);
			24574: out = 16'(-199);
			24575: out = 16'(-209);
			24576: out = 16'(2313);
			24577: out = 16'(1115);
			24578: out = 16'(-2087);
			24579: out = 16'(-2459);
			24580: out = 16'(-1660);
			24581: out = 16'(1459);
			24582: out = 16'(1167);
			24583: out = 16'(1152);
			24584: out = 16'(290);
			24585: out = 16'(-474);
			24586: out = 16'(-1298);
			24587: out = 16'(-981);
			24588: out = 16'(-838);
			24589: out = 16'(11);
			24590: out = 16'(948);
			24591: out = 16'(2000);
			24592: out = 16'(2294);
			24593: out = 16'(-369);
			24594: out = 16'(-2727);
			24595: out = 16'(-5017);
			24596: out = 16'(-1904);
			24597: out = 16'(-264);
			24598: out = 16'(656);
			24599: out = 16'(617);
			24600: out = 16'(271);
			24601: out = 16'(53);
			24602: out = 16'(112);
			24603: out = 16'(1266);
			24604: out = 16'(4327);
			24605: out = 16'(4572);
			24606: out = 16'(3630);
			24607: out = 16'(-747);
			24608: out = 16'(-2125);
			24609: out = 16'(-2512);
			24610: out = 16'(62);
			24611: out = 16'(578);
			24612: out = 16'(75);
			24613: out = 16'(423);
			24614: out = 16'(-160);
			24615: out = 16'(-341);
			24616: out = 16'(-1808);
			24617: out = 16'(-997);
			24618: out = 16'(1150);
			24619: out = 16'(3062);
			24620: out = 16'(3019);
			24621: out = 16'(-298);
			24622: out = 16'(-2107);
			24623: out = 16'(-3846);
			24624: out = 16'(-3233);
			24625: out = 16'(-3548);
			24626: out = 16'(-3079);
			24627: out = 16'(-2699);
			24628: out = 16'(-1104);
			24629: out = 16'(808);
			24630: out = 16'(-78);
			24631: out = 16'(461);
			24632: out = 16'(628);
			24633: out = 16'(2523);
			24634: out = 16'(2003);
			24635: out = 16'(695);
			24636: out = 16'(-1723);
			24637: out = 16'(-2073);
			24638: out = 16'(-273);
			24639: out = 16'(1262);
			24640: out = 16'(2297);
			24641: out = 16'(3383);
			24642: out = 16'(1194);
			24643: out = 16'(-252);
			24644: out = 16'(126);
			24645: out = 16'(2087);
			24646: out = 16'(3653);
			24647: out = 16'(1583);
			24648: out = 16'(-1270);
			24649: out = 16'(-4533);
			24650: out = 16'(-3105);
			24651: out = 16'(-1028);
			24652: out = 16'(2073);
			24653: out = 16'(2894);
			24654: out = 16'(2206);
			24655: out = 16'(-627);
			24656: out = 16'(-3572);
			24657: out = 16'(-5471);
			24658: out = 16'(-4880);
			24659: out = 16'(-2194);
			24660: out = 16'(1046);
			24661: out = 16'(2929);
			24662: out = 16'(2259);
			24663: out = 16'(15);
			24664: out = 16'(947);
			24665: out = 16'(-1677);
			24666: out = 16'(-3423);
			24667: out = 16'(-5544);
			24668: out = 16'(-3563);
			24669: out = 16'(315);
			24670: out = 16'(-107);
			24671: out = 16'(451);
			24672: out = 16'(570);
			24673: out = 16'(1287);
			24674: out = 16'(2108);
			24675: out = 16'(4160);
			24676: out = 16'(3076);
			24677: out = 16'(1999);
			24678: out = 16'(-1156);
			24679: out = 16'(-2);
			24680: out = 16'(888);
			24681: out = 16'(3303);
			24682: out = 16'(980);
			24683: out = 16'(-1537);
			24684: out = 16'(-1776);
			24685: out = 16'(-684);
			24686: out = 16'(1604);
			24687: out = 16'(191);
			24688: out = 16'(807);
			24689: out = 16'(1051);
			24690: out = 16'(884);
			24691: out = 16'(-960);
			24692: out = 16'(-4348);
			24693: out = 16'(-3100);
			24694: out = 16'(-1824);
			24695: out = 16'(489);
			24696: out = 16'(-957);
			24697: out = 16'(-1694);
			24698: out = 16'(-134);
			24699: out = 16'(22);
			24700: out = 16'(780);
			24701: out = 16'(389);
			24702: out = 16'(2443);
			24703: out = 16'(3847);
			24704: out = 16'(1654);
			24705: out = 16'(195);
			24706: out = 16'(-1237);
			24707: out = 16'(-1783);
			24708: out = 16'(-1135);
			24709: out = 16'(487);
			24710: out = 16'(373);
			24711: out = 16'(-148);
			24712: out = 16'(-1930);
			24713: out = 16'(-348);
			24714: out = 16'(1172);
			24715: out = 16'(3179);
			24716: out = 16'(3297);
			24717: out = 16'(2709);
			24718: out = 16'(587);
			24719: out = 16'(250);
			24720: out = 16'(189);
			24721: out = 16'(-339);
			24722: out = 16'(75);
			24723: out = 16'(383);
			24724: out = 16'(475);
			24725: out = 16'(-40);
			24726: out = 16'(-490);
			24727: out = 16'(-1281);
			24728: out = 16'(-422);
			24729: out = 16'(1116);
			24730: out = 16'(1210);
			24731: out = 16'(426);
			24732: out = 16'(-1158);
			24733: out = 16'(-2867);
			24734: out = 16'(-3152);
			24735: out = 16'(-1266);
			24736: out = 16'(298);
			24737: out = 16'(1352);
			24738: out = 16'(1214);
			24739: out = 16'(718);
			24740: out = 16'(-40);
			24741: out = 16'(-3936);
			24742: out = 16'(-2930);
			24743: out = 16'(-628);
			24744: out = 16'(3138);
			24745: out = 16'(3558);
			24746: out = 16'(2333);
			24747: out = 16'(-2010);
			24748: out = 16'(-3154);
			24749: out = 16'(-828);
			24750: out = 16'(905);
			24751: out = 16'(1570);
			24752: out = 16'(-2196);
			24753: out = 16'(-645);
			24754: out = 16'(-551);
			24755: out = 16'(-923);
			24756: out = 16'(-1175);
			24757: out = 16'(-516);
			24758: out = 16'(2291);
			24759: out = 16'(2739);
			24760: out = 16'(2322);
			24761: out = 16'(885);
			24762: out = 16'(251);
			24763: out = 16'(306);
			24764: out = 16'(-1628);
			24765: out = 16'(-1497);
			24766: out = 16'(-326);
			24767: out = 16'(121);
			24768: out = 16'(-257);
			24769: out = 16'(-2802);
			24770: out = 16'(-401);
			24771: out = 16'(1414);
			24772: out = 16'(4491);
			24773: out = 16'(2538);
			24774: out = 16'(208);
			24775: out = 16'(-3858);
			24776: out = 16'(-4383);
			24777: out = 16'(-3509);
			24778: out = 16'(1945);
			24779: out = 16'(3046);
			24780: out = 16'(2890);
			24781: out = 16'(-2941);
			24782: out = 16'(-4720);
			24783: out = 16'(-4661);
			24784: out = 16'(412);
			24785: out = 16'(3046);
			24786: out = 16'(3810);
			24787: out = 16'(1621);
			24788: out = 16'(-310);
			24789: out = 16'(-903);
			24790: out = 16'(-200);
			24791: out = 16'(876);
			24792: out = 16'(336);
			24793: out = 16'(758);
			24794: out = 16'(451);
			24795: out = 16'(2097);
			24796: out = 16'(-17);
			24797: out = 16'(-2027);
			24798: out = 16'(-1239);
			24799: out = 16'(-423);
			24800: out = 16'(644);
			24801: out = 16'(-73);
			24802: out = 16'(-189);
			24803: out = 16'(-149);
			24804: out = 16'(-1351);
			24805: out = 16'(-2434);
			24806: out = 16'(-4191);
			24807: out = 16'(-1465);
			24808: out = 16'(43);
			24809: out = 16'(-306);
			24810: out = 16'(-155);
			24811: out = 16'(185);
			24812: out = 16'(2667);
			24813: out = 16'(2388);
			24814: out = 16'(1807);
			24815: out = 16'(810);
			24816: out = 16'(201);
			24817: out = 16'(-259);
			24818: out = 16'(-2839);
			24819: out = 16'(-2911);
			24820: out = 16'(-1500);
			24821: out = 16'(-1827);
			24822: out = 16'(-1315);
			24823: out = 16'(-911);
			24824: out = 16'(860);
			24825: out = 16'(1480);
			24826: out = 16'(665);
			24827: out = 16'(769);
			24828: out = 16'(1288);
			24829: out = 16'(5233);
			24830: out = 16'(3211);
			24831: out = 16'(1283);
			24832: out = 16'(-2434);
			24833: out = 16'(-1506);
			24834: out = 16'(101);
			24835: out = 16'(1047);
			24836: out = 16'(919);
			24837: out = 16'(209);
			24838: out = 16'(-1578);
			24839: out = 16'(-1213);
			24840: out = 16'(499);
			24841: out = 16'(1010);
			24842: out = 16'(1063);
			24843: out = 16'(272);
			24844: out = 16'(-658);
			24845: out = 16'(-1346);
			24846: out = 16'(-1902);
			24847: out = 16'(-748);
			24848: out = 16'(208);
			24849: out = 16'(2014);
			24850: out = 16'(308);
			24851: out = 16'(-1127);
			24852: out = 16'(-601);
			24853: out = 16'(2096);
			24854: out = 16'(5288);
			24855: out = 16'(3867);
			24856: out = 16'(1492);
			24857: out = 16'(-3387);
			24858: out = 16'(-16);
			24859: out = 16'(7);
			24860: out = 16'(691);
			24861: out = 16'(-3817);
			24862: out = 16'(-4735);
			24863: out = 16'(-2553);
			24864: out = 16'(-1147);
			24865: out = 16'(-576);
			24866: out = 16'(-3435);
			24867: out = 16'(-1196);
			24868: out = 16'(1503);
			24869: out = 16'(5187);
			24870: out = 16'(5914);
			24871: out = 16'(4795);
			24872: out = 16'(1211);
			24873: out = 16'(-2684);
			24874: out = 16'(-5942);
			24875: out = 16'(-3359);
			24876: out = 16'(-848);
			24877: out = 16'(2082);
			24878: out = 16'(1464);
			24879: out = 16'(189);
			24880: out = 16'(-2743);
			24881: out = 16'(-2606);
			24882: out = 16'(-1767);
			24883: out = 16'(1413);
			24884: out = 16'(1646);
			24885: out = 16'(1841);
			24886: out = 16'(-291);
			24887: out = 16'(1108);
			24888: out = 16'(1738);
			24889: out = 16'(62);
			24890: out = 16'(-1655);
			24891: out = 16'(-3486);
			24892: out = 16'(-366);
			24893: out = 16'(47);
			24894: out = 16'(556);
			24895: out = 16'(-449);
			24896: out = 16'(722);
			24897: out = 16'(2625);
			24898: out = 16'(2650);
			24899: out = 16'(1891);
			24900: out = 16'(265);
			24901: out = 16'(-722);
			24902: out = 16'(-1750);
			24903: out = 16'(-4339);
			24904: out = 16'(-2714);
			24905: out = 16'(-1612);
			24906: out = 16'(-119);
			24907: out = 16'(-2318);
			24908: out = 16'(-3824);
			24909: out = 16'(-714);
			24910: out = 16'(1619);
			24911: out = 16'(3473);
			24912: out = 16'(3528);
			24913: out = 16'(1878);
			24914: out = 16'(-517);
			24915: out = 16'(-5228);
			24916: out = 16'(-5697);
			24917: out = 16'(-2079);
			24918: out = 16'(187);
			24919: out = 16'(1754);
			24920: out = 16'(352);
			24921: out = 16'(881);
			24922: out = 16'(809);
			24923: out = 16'(1474);
			24924: out = 16'(1744);
			24925: out = 16'(2286);
			24926: out = 16'(3921);
			24927: out = 16'(2016);
			24928: out = 16'(-483);
			24929: out = 16'(582);
			24930: out = 16'(965);
			24931: out = 16'(1934);
			24932: out = 16'(-622);
			24933: out = 16'(-1976);
			24934: out = 16'(-3518);
			24935: out = 16'(-2727);
			24936: out = 16'(-2314);
			24937: out = 16'(-1680);
			24938: out = 16'(-796);
			24939: out = 16'(189);
			24940: out = 16'(593);
			24941: out = 16'(1601);
			24942: out = 16'(2017);
			24943: out = 16'(1331);
			24944: out = 16'(1318);
			24945: out = 16'(1357);
			24946: out = 16'(2523);
			24947: out = 16'(1614);
			24948: out = 16'(-45);
			24949: out = 16'(-821);
			24950: out = 16'(-903);
			24951: out = 16'(565);
			24952: out = 16'(-3010);
			24953: out = 16'(-2153);
			24954: out = 16'(675);
			24955: out = 16'(2091);
			24956: out = 16'(1723);
			24957: out = 16'(-2061);
			24958: out = 16'(-1282);
			24959: out = 16'(-810);
			24960: out = 16'(628);
			24961: out = 16'(434);
			24962: out = 16'(480);
			24963: out = 16'(1231);
			24964: out = 16'(1179);
			24965: out = 16'(1287);
			24966: out = 16'(976);
			24967: out = 16'(2995);
			24968: out = 16'(5561);
			24969: out = 16'(1668);
			24970: out = 16'(-319);
			24971: out = 16'(-3142);
			24972: out = 16'(-692);
			24973: out = 16'(-871);
			24974: out = 16'(-1994);
			24975: out = 16'(-4665);
			24976: out = 16'(-5802);
			24977: out = 16'(-3935);
			24978: out = 16'(-3406);
			24979: out = 16'(-1278);
			24980: out = 16'(2310);
			24981: out = 16'(4280);
			24982: out = 16'(4599);
			24983: out = 16'(105);
			24984: out = 16'(-852);
			24985: out = 16'(-929);
			24986: out = 16'(918);
			24987: out = 16'(1073);
			24988: out = 16'(92);
			24989: out = 16'(-76);
			24990: out = 16'(-443);
			24991: out = 16'(597);
			24992: out = 16'(-2104);
			24993: out = 16'(-2299);
			24994: out = 16'(-1999);
			24995: out = 16'(1309);
			24996: out = 16'(3140);
			24997: out = 16'(5228);
			24998: out = 16'(877);
			24999: out = 16'(-2647);
			25000: out = 16'(-4159);
			25001: out = 16'(-1543);
			25002: out = 16'(1782);
			25003: out = 16'(1015);
			25004: out = 16'(1018);
			25005: out = 16'(138);
			25006: out = 16'(-287);
			25007: out = 16'(171);
			25008: out = 16'(1362);
			25009: out = 16'(2269);
			25010: out = 16'(1897);
			25011: out = 16'(170);
			25012: out = 16'(-2900);
			25013: out = 16'(-3752);
			25014: out = 16'(155);
			25015: out = 16'(-372);
			25016: out = 16'(-459);
			25017: out = 16'(-4341);
			25018: out = 16'(-1460);
			25019: out = 16'(718);
			25020: out = 16'(349);
			25021: out = 16'(509);
			25022: out = 16'(557);
			25023: out = 16'(2437);
			25024: out = 16'(2141);
			25025: out = 16'(1004);
			25026: out = 16'(-446);
			25027: out = 16'(-2054);
			25028: out = 16'(-3306);
			25029: out = 16'(-3412);
			25030: out = 16'(-2434);
			25031: out = 16'(-82);
			25032: out = 16'(-61);
			25033: out = 16'(137);
			25034: out = 16'(-20);
			25035: out = 16'(500);
			25036: out = 16'(855);
			25037: out = 16'(1402);
			25038: out = 16'(1346);
			25039: out = 16'(1468);
			25040: out = 16'(1858);
			25041: out = 16'(2321);
			25042: out = 16'(2384);
			25043: out = 16'(148);
			25044: out = 16'(-663);
			25045: out = 16'(-240);
			25046: out = 16'(-1719);
			25047: out = 16'(-1894);
			25048: out = 16'(-2763);
			25049: out = 16'(1353);
			25050: out = 16'(2604);
			25051: out = 16'(2012);
			25052: out = 16'(-962);
			25053: out = 16'(-2612);
			25054: out = 16'(-1090);
			25055: out = 16'(1269);
			25056: out = 16'(3516);
			25057: out = 16'(1753);
			25058: out = 16'(1344);
			25059: out = 16'(-252);
			25060: out = 16'(-1309);
			25061: out = 16'(-3392);
			25062: out = 16'(-4815);
			25063: out = 16'(-736);
			25064: out = 16'(1710);
			25065: out = 16'(3209);
			25066: out = 16'(1863);
			25067: out = 16'(826);
			25068: out = 16'(654);
			25069: out = 16'(-670);
			25070: out = 16'(-1284);
			25071: out = 16'(-1945);
			25072: out = 16'(35);
			25073: out = 16'(1384);
			25074: out = 16'(294);
			25075: out = 16'(-320);
			25076: out = 16'(-978);
			25077: out = 16'(3046);
			25078: out = 16'(2760);
			25079: out = 16'(2473);
			25080: out = 16'(458);
			25081: out = 16'(1830);
			25082: out = 16'(4338);
			25083: out = 16'(1687);
			25084: out = 16'(223);
			25085: out = 16'(-606);
			25086: out = 16'(-3964);
			25087: out = 16'(-5930);
			25088: out = 16'(-7625);
			25089: out = 16'(-2967);
			25090: out = 16'(1168);
			25091: out = 16'(3519);
			25092: out = 16'(2174);
			25093: out = 16'(-283);
			25094: out = 16'(910);
			25095: out = 16'(-356);
			25096: out = 16'(-397);
			25097: out = 16'(-4314);
			25098: out = 16'(-1577);
			25099: out = 16'(2145);
			25100: out = 16'(818);
			25101: out = 16'(-806);
			25102: out = 16'(-3555);
			25103: out = 16'(-2247);
			25104: out = 16'(-1087);
			25105: out = 16'(407);
			25106: out = 16'(2432);
			25107: out = 16'(3204);
			25108: out = 16'(1827);
			25109: out = 16'(612);
			25110: out = 16'(-669);
			25111: out = 16'(500);
			25112: out = 16'(-637);
			25113: out = 16'(-1291);
			25114: out = 16'(-2628);
			25115: out = 16'(-1481);
			25116: out = 16'(100);
			25117: out = 16'(-419);
			25118: out = 16'(-476);
			25119: out = 16'(-1115);
			25120: out = 16'(2073);
			25121: out = 16'(2458);
			25122: out = 16'(1913);
			25123: out = 16'(644);
			25124: out = 16'(895);
			25125: out = 16'(3255);
			25126: out = 16'(2222);
			25127: out = 16'(1100);
			25128: out = 16'(-1199);
			25129: out = 16'(-2175);
			25130: out = 16'(-2792);
			25131: out = 16'(-1979);
			25132: out = 16'(-1258);
			25133: out = 16'(-166);
			25134: out = 16'(106);
			25135: out = 16'(266);
			25136: out = 16'(-386);
			25137: out = 16'(-8);
			25138: out = 16'(-438);
			25139: out = 16'(-261);
			25140: out = 16'(-2987);
			25141: out = 16'(-2317);
			25142: out = 16'(537);
			25143: out = 16'(1526);
			25144: out = 16'(1659);
			25145: out = 16'(-253);
			25146: out = 16'(269);
			25147: out = 16'(393);
			25148: out = 16'(506);
			25149: out = 16'(1655);
			25150: out = 16'(2474);
			25151: out = 16'(344);
			25152: out = 16'(-719);
			25153: out = 16'(-2002);
			25154: out = 16'(1719);
			25155: out = 16'(1178);
			25156: out = 16'(393);
			25157: out = 16'(-2221);
			25158: out = 16'(-2470);
			25159: out = 16'(-1884);
			25160: out = 16'(-147);
			25161: out = 16'(195);
			25162: out = 16'(-334);
			25163: out = 16'(-537);
			25164: out = 16'(391);
			25165: out = 16'(2388);
			25166: out = 16'(3863);
			25167: out = 16'(3860);
			25168: out = 16'(1350);
			25169: out = 16'(-671);
			25170: out = 16'(-2506);
			25171: out = 16'(-5730);
			25172: out = 16'(-3517);
			25173: out = 16'(281);
			25174: out = 16'(2614);
			25175: out = 16'(2226);
			25176: out = 16'(-680);
			25177: out = 16'(47);
			25178: out = 16'(-53);
			25179: out = 16'(1473);
			25180: out = 16'(-106);
			25181: out = 16'(7);
			25182: out = 16'(102);
			25183: out = 16'(-15);
			25184: out = 16'(-1223);
			25185: out = 16'(-3204);
			25186: out = 16'(-3624);
			25187: out = 16'(-2816);
			25188: out = 16'(-1459);
			25189: out = 16'(1407);
			25190: out = 16'(3559);
			25191: out = 16'(3915);
			25192: out = 16'(2142);
			25193: out = 16'(-750);
			25194: out = 16'(633);
			25195: out = 16'(297);
			25196: out = 16'(378);
			25197: out = 16'(-1567);
			25198: out = 16'(-932);
			25199: out = 16'(2149);
			25200: out = 16'(761);
			25201: out = 16'(4);
			25202: out = 16'(-2952);
			25203: out = 16'(417);
			25204: out = 16'(1964);
			25205: out = 16'(2089);
			25206: out = 16'(-1908);
			25207: out = 16'(-5053);
			25208: out = 16'(182);
			25209: out = 16'(1003);
			25210: out = 16'(1830);
			25211: out = 16'(-3519);
			25212: out = 16'(-3919);
			25213: out = 16'(-3109);
			25214: out = 16'(-1443);
			25215: out = 16'(-700);
			25216: out = 16'(-980);
			25217: out = 16'(974);
			25218: out = 16'(1520);
			25219: out = 16'(1452);
			25220: out = 16'(810);
			25221: out = 16'(512);
			25222: out = 16'(658);
			25223: out = 16'(1109);
			25224: out = 16'(1209);
			25225: out = 16'(602);
			25226: out = 16'(-1140);
			25227: out = 16'(-2494);
			25228: out = 16'(-504);
			25229: out = 16'(1519);
			25230: out = 16'(4262);
			25231: out = 16'(1379);
			25232: out = 16'(1201);
			25233: out = 16'(296);
			25234: out = 16'(4301);
			25235: out = 16'(3803);
			25236: out = 16'(964);
			25237: out = 16'(-661);
			25238: out = 16'(-646);
			25239: out = 16'(2473);
			25240: out = 16'(2278);
			25241: out = 16'(1738);
			25242: out = 16'(-1316);
			25243: out = 16'(-2188);
			25244: out = 16'(-2782);
			25245: out = 16'(-656);
			25246: out = 16'(-186);
			25247: out = 16'(347);
			25248: out = 16'(-2470);
			25249: out = 16'(-2994);
			25250: out = 16'(-3465);
			25251: out = 16'(-52);
			25252: out = 16'(316);
			25253: out = 16'(-439);
			25254: out = 16'(-3172);
			25255: out = 16'(-3987);
			25256: out = 16'(-2262);
			25257: out = 16'(-2592);
			25258: out = 16'(-1958);
			25259: out = 16'(-957);
			25260: out = 16'(51);
			25261: out = 16'(744);
			25262: out = 16'(503);
			25263: out = 16'(813);
			25264: out = 16'(738);
			25265: out = 16'(1594);
			25266: out = 16'(27);
			25267: out = 16'(-1994);
			25268: out = 16'(-2474);
			25269: out = 16'(-1425);
			25270: out = 16'(1206);
			25271: out = 16'(653);
			25272: out = 16'(809);
			25273: out = 16'(-406);
			25274: out = 16'(2258);
			25275: out = 16'(3120);
			25276: out = 16'(3722);
			25277: out = 16'(1448);
			25278: out = 16'(494);
			25279: out = 16'(2061);
			25280: out = 16'(2436);
			25281: out = 16'(2071);
			25282: out = 16'(-2475);
			25283: out = 16'(-4193);
			25284: out = 16'(-5254);
			25285: out = 16'(-865);
			25286: out = 16'(178);
			25287: out = 16'(763);
			25288: out = 16'(-830);
			25289: out = 16'(-833);
			25290: out = 16'(-205);
			25291: out = 16'(1035);
			25292: out = 16'(1729);
			25293: out = 16'(2141);
			25294: out = 16'(1070);
			25295: out = 16'(-232);
			25296: out = 16'(-1896);
			25297: out = 16'(-1561);
			25298: out = 16'(-527);
			25299: out = 16'(2011);
			25300: out = 16'(2180);
			25301: out = 16'(1809);
			25302: out = 16'(-986);
			25303: out = 16'(-133);
			25304: out = 16'(1794);
			25305: out = 16'(4184);
			25306: out = 16'(3741);
			25307: out = 16'(620);
			25308: out = 16'(3311);
			25309: out = 16'(2417);
			25310: out = 16'(2028);
			25311: out = 16'(-3945);
			25312: out = 16'(-4808);
			25313: out = 16'(-489);
			25314: out = 16'(1831);
			25315: out = 16'(3038);
			25316: out = 16'(-688);
			25317: out = 16'(238);
			25318: out = 16'(59);
			25319: out = 16'(-393);
			25320: out = 16'(-2344);
			25321: out = 16'(-3844);
			25322: out = 16'(-529);
			25323: out = 16'(-438);
			25324: out = 16'(-627);
			25325: out = 16'(-4807);
			25326: out = 16'(-4166);
			25327: out = 16'(-758);
			25328: out = 16'(-147);
			25329: out = 16'(593);
			25330: out = 16'(-317);
			25331: out = 16'(102);
			25332: out = 16'(-440);
			25333: out = 16'(-972);
			25334: out = 16'(-1238);
			25335: out = 16'(-820);
			25336: out = 16'(-462);
			25337: out = 16'(292);
			25338: out = 16'(326);
			25339: out = 16'(-15);
			25340: out = 16'(-1513);
			25341: out = 16'(-2497);
			25342: out = 16'(-513);
			25343: out = 16'(2281);
			25344: out = 16'(5814);
			25345: out = 16'(2638);
			25346: out = 16'(1343);
			25347: out = 16'(-354);
			25348: out = 16'(974);
			25349: out = 16'(1928);
			25350: out = 16'(4253);
			25351: out = 16'(1992);
			25352: out = 16'(643);
			25353: out = 16'(-1489);
			25354: out = 16'(-796);
			25355: out = 16'(-746);
			25356: out = 16'(-290);
			25357: out = 16'(-2800);
			25358: out = 16'(-4800);
			25359: out = 16'(-5502);
			25360: out = 16'(-3034);
			25361: out = 16'(430);
			25362: out = 16'(1121);
			25363: out = 16'(770);
			25364: out = 16'(-1391);
			25365: out = 16'(-1556);
			25366: out = 16'(-1590);
			25367: out = 16'(3);
			25368: out = 16'(-224);
			25369: out = 16'(329);
			25370: out = 16'(449);
			25371: out = 16'(323);
			25372: out = 16'(181);
			25373: out = 16'(2398);
			25374: out = 16'(1115);
			25375: out = 16'(398);
			25376: out = 16'(-417);
			25377: out = 16'(974);
			25378: out = 16'(2137);
			25379: out = 16'(694);
			25380: out = 16'(-924);
			25381: out = 16'(-2803);
			25382: out = 16'(700);
			25383: out = 16'(2246);
			25384: out = 16'(3535);
			25385: out = 16'(2896);
			25386: out = 16'(2267);
			25387: out = 16'(1144);
			25388: out = 16'(667);
			25389: out = 16'(963);
			25390: out = 16'(4129);
			25391: out = 16'(1642);
			25392: out = 16'(-443);
			25393: out = 16'(-3809);
			25394: out = 16'(-2277);
			25395: out = 16'(-440);
			25396: out = 16'(-2208);
			25397: out = 16'(-2373);
			25398: out = 16'(-2901);
			25399: out = 16'(12);
			25400: out = 16'(142);
			25401: out = 16'(-164);
			25402: out = 16'(-433);
			25403: out = 16'(-352);
			25404: out = 16'(-541);
			25405: out = 16'(302);
			25406: out = 16'(-114);
			25407: out = 16'(-1092);
			25408: out = 16'(-2350);
			25409: out = 16'(-2352);
			25410: out = 16'(-423);
			25411: out = 16'(211);
			25412: out = 16'(410);
			25413: out = 16'(589);
			25414: out = 16'(-80);
			25415: out = 16'(-352);
			25416: out = 16'(-2741);
			25417: out = 16'(-1089);
			25418: out = 16'(956);
			25419: out = 16'(4468);
			25420: out = 16'(3375);
			25421: out = 16'(94);
			25422: out = 16'(-3426);
			25423: out = 16'(-3018);
			25424: out = 16'(2655);
			25425: out = 16'(1308);
			25426: out = 16'(1506);
			25427: out = 16'(1243);
			25428: out = 16'(354);
			25429: out = 16'(-760);
			25430: out = 16'(-1141);
			25431: out = 16'(93);
			25432: out = 16'(1310);
			25433: out = 16'(-1932);
			25434: out = 16'(-2251);
			25435: out = 16'(-2788);
			25436: out = 16'(-194);
			25437: out = 16'(-507);
			25438: out = 16'(-1029);
			25439: out = 16'(-1881);
			25440: out = 16'(-726);
			25441: out = 16'(1699);
			25442: out = 16'(1420);
			25443: out = 16'(1303);
			25444: out = 16'(423);
			25445: out = 16'(162);
			25446: out = 16'(75);
			25447: out = 16'(1538);
			25448: out = 16'(837);
			25449: out = 16'(693);
			25450: out = 16'(294);
			25451: out = 16'(972);
			25452: out = 16'(1410);
			25453: out = 16'(2741);
			25454: out = 16'(1392);
			25455: out = 16'(-507);
			25456: out = 16'(-228);
			25457: out = 16'(-53);
			25458: out = 16'(610);
			25459: out = 16'(2658);
			25460: out = 16'(3124);
			25461: out = 16'(1566);
			25462: out = 16'(857);
			25463: out = 16'(-366);
			25464: out = 16'(-96);
			25465: out = 16'(-2225);
			25466: out = 16'(-3474);
			25467: out = 16'(-6456);
			25468: out = 16'(-3766);
			25469: out = 16'(-1385);
			25470: out = 16'(1338);
			25471: out = 16'(-154);
			25472: out = 16'(-2292);
			25473: out = 16'(-4884);
			25474: out = 16'(-3624);
			25475: out = 16'(-429);
			25476: out = 16'(977);
			25477: out = 16'(1851);
			25478: out = 16'(1431);
			25479: out = 16'(350);
			25480: out = 16'(-177);
			25481: out = 16'(707);
			25482: out = 16'(1134);
			25483: out = 16'(1467);
			25484: out = 16'(427);
			25485: out = 16'(274);
			25486: out = 16'(118);
			25487: out = 16'(2244);
			25488: out = 16'(948);
			25489: out = 16'(-512);
			25490: out = 16'(-2325);
			25491: out = 16'(-3213);
			25492: out = 16'(-3235);
			25493: out = 16'(-834);
			25494: out = 16'(949);
			25495: out = 16'(2320);
			25496: out = 16'(1700);
			25497: out = 16'(1147);
			25498: out = 16'(499);
			25499: out = 16'(103);
			25500: out = 16'(-75);
			25501: out = 16'(-69);
			25502: out = 16'(-72);
			25503: out = 16'(453);
			25504: out = 16'(3655);
			25505: out = 16'(1722);
			25506: out = 16'(-239);
			25507: out = 16'(-3393);
			25508: out = 16'(-2460);
			25509: out = 16'(-728);
			25510: out = 16'(451);
			25511: out = 16'(442);
			25512: out = 16'(-442);
			25513: out = 16'(-1576);
			25514: out = 16'(-1203);
			25515: out = 16'(779);
			25516: out = 16'(359);
			25517: out = 16'(561);
			25518: out = 16'(-176);
			25519: out = 16'(1595);
			25520: out = 16'(1989);
			25521: out = 16'(607);
			25522: out = 16'(708);
			25523: out = 16'(757);
			25524: out = 16'(2144);
			25525: out = 16'(1222);
			25526: out = 16'(578);
			25527: out = 16'(1131);
			25528: out = 16'(2230);
			25529: out = 16'(3255);
			25530: out = 16'(199);
			25531: out = 16'(-1363);
			25532: out = 16'(-3080);
			25533: out = 16'(-1530);
			25534: out = 16'(-1469);
			25535: out = 16'(-2070);
			25536: out = 16'(-371);
			25537: out = 16'(823);
			25538: out = 16'(1181);
			25539: out = 16'(1899);
			25540: out = 16'(1669);
			25541: out = 16'(396);
			25542: out = 16'(-1109);
			25543: out = 16'(-2057);
			25544: out = 16'(-208);
			25545: out = 16'(-31);
			25546: out = 16'(468);
			25547: out = 16'(97);
			25548: out = 16'(1087);
			25549: out = 16'(1938);
			25550: out = 16'(1387);
			25551: out = 16'(514);
			25552: out = 16'(-678);
			25553: out = 16'(-1782);
			25554: out = 16'(-2085);
			25555: out = 16'(-1211);
			25556: out = 16'(-1408);
			25557: out = 16'(-708);
			25558: out = 16'(1304);
			25559: out = 16'(690);
			25560: out = 16'(-18);
			25561: out = 16'(-1246);
			25562: out = 16'(-498);
			25563: out = 16'(404);
			25564: out = 16'(-303);
			25565: out = 16'(52);
			25566: out = 16'(205);
			25567: out = 16'(-1055);
			25568: out = 16'(-1331);
			25569: out = 16'(-1164);
			25570: out = 16'(-6);
			25571: out = 16'(249);
			25572: out = 16'(-602);
			25573: out = 16'(300);
			25574: out = 16'(-103);
			25575: out = 16'(-1158);
			25576: out = 16'(-2307);
			25577: out = 16'(-2314);
			25578: out = 16'(512);
			25579: out = 16'(94);
			25580: out = 16'(-253);
			25581: out = 16'(-1891);
			25582: out = 16'(-1105);
			25583: out = 16'(80);
			25584: out = 16'(1903);
			25585: out = 16'(2297);
			25586: out = 16'(1981);
			25587: out = 16'(965);
			25588: out = 16'(-105);
			25589: out = 16'(-1216);
			25590: out = 16'(-365);
			25591: out = 16'(101);
			25592: out = 16'(686);
			25593: out = 16'(457);
			25594: out = 16'(1542);
			25595: out = 16'(4856);
			25596: out = 16'(3874);
			25597: out = 16'(2375);
			25598: out = 16'(-2158);
			25599: out = 16'(-1195);
			25600: out = 16'(58);
			25601: out = 16'(2394);
			25602: out = 16'(1499);
			25603: out = 16'(-120);
			25604: out = 16'(1171);
			25605: out = 16'(622);
			25606: out = 16'(326);
			25607: out = 16'(-1311);
			25608: out = 16'(-254);
			25609: out = 16'(2743);
			25610: out = 16'(558);
			25611: out = 16'(-954);
			25612: out = 16'(-4252);
			25613: out = 16'(-1046);
			25614: out = 16'(569);
			25615: out = 16'(1954);
			25616: out = 16'(-199);
			25617: out = 16'(-1914);
			25618: out = 16'(-3919);
			25619: out = 16'(-1217);
			25620: out = 16'(1736);
			25621: out = 16'(2374);
			25622: out = 16'(1047);
			25623: out = 16'(-2008);
			25624: out = 16'(-1686);
			25625: out = 16'(-2812);
			25626: out = 16'(-2670);
			25627: out = 16'(-3911);
			25628: out = 16'(-2164);
			25629: out = 16'(708);
			25630: out = 16'(1795);
			25631: out = 16'(1419);
			25632: out = 16'(-1315);
			25633: out = 16'(-485);
			25634: out = 16'(267);
			25635: out = 16'(2070);
			25636: out = 16'(1109);
			25637: out = 16'(140);
			25638: out = 16'(694);
			25639: out = 16'(354);
			25640: out = 16'(409);
			25641: out = 16'(-3557);
			25642: out = 16'(-1997);
			25643: out = 16'(643);
			25644: out = 16'(1856);
			25645: out = 16'(774);
			25646: out = 16'(-2347);
			25647: out = 16'(-1926);
			25648: out = 16'(-1183);
			25649: out = 16'(1704);
			25650: out = 16'(-470);
			25651: out = 16'(-1632);
			25652: out = 16'(-3650);
			25653: out = 16'(-1464);
			25654: out = 16'(197);
			25655: out = 16'(608);
			25656: out = 16'(1275);
			25657: out = 16'(1400);
			25658: out = 16'(623);
			25659: out = 16'(55);
			25660: out = 16'(-178);
			25661: out = 16'(1166);
			25662: out = 16'(2279);
			25663: out = 16'(3541);
			25664: out = 16'(1094);
			25665: out = 16'(150);
			25666: out = 16'(-487);
			25667: out = 16'(-197);
			25668: out = 16'(-289);
			25669: out = 16'(-384);
			25670: out = 16'(-1517);
			25671: out = 16'(-1948);
			25672: out = 16'(-1114);
			25673: out = 16'(-597);
			25674: out = 16'(227);
			25675: out = 16'(1257);
			25676: out = 16'(1019);
			25677: out = 16'(199);
			25678: out = 16'(786);
			25679: out = 16'(404);
			25680: out = 16'(681);
			25681: out = 16'(-1829);
			25682: out = 16'(-1098);
			25683: out = 16'(379);
			25684: out = 16'(161);
			25685: out = 16'(-1042);
			25686: out = 16'(-2627);
			25687: out = 16'(-4142);
			25688: out = 16'(-3147);
			25689: out = 16'(746);
			25690: out = 16'(2668);
			25691: out = 16'(3214);
			25692: out = 16'(-229);
			25693: out = 16'(-728);
			25694: out = 16'(-900);
			25695: out = 16'(555);
			25696: out = 16'(1464);
			25697: out = 16'(2189);
			25698: out = 16'(2227);
			25699: out = 16'(1127);
			25700: out = 16'(-261);
			25701: out = 16'(-1105);
			25702: out = 16'(67);
			25703: out = 16'(3019);
			25704: out = 16'(3588);
			25705: out = 16'(4137);
			25706: out = 16'(3854);
			25707: out = 16'(1607);
			25708: out = 16'(-107);
			25709: out = 16'(514);
			25710: out = 16'(-442);
			25711: out = 16'(-795);
			25712: out = 16'(-1553);
			25713: out = 16'(-654);
			25714: out = 16'(26);
			25715: out = 16'(-2129);
			25716: out = 16'(-1867);
			25717: out = 16'(-1317);
			25718: out = 16'(-645);
			25719: out = 16'(-1100);
			25720: out = 16'(-2229);
			25721: out = 16'(-2663);
			25722: out = 16'(-2683);
			25723: out = 16'(-1883);
			25724: out = 16'(-2010);
			25725: out = 16'(-1681);
			25726: out = 16'(-1055);
			25727: out = 16'(-1552);
			25728: out = 16'(-1853);
			25729: out = 16'(-1783);
			25730: out = 16'(-774);
			25731: out = 16'(339);
			25732: out = 16'(-99);
			25733: out = 16'(586);
			25734: out = 16'(823);
			25735: out = 16'(2278);
			25736: out = 16'(933);
			25737: out = 16'(-1230);
			25738: out = 16'(-126);
			25739: out = 16'(624);
			25740: out = 16'(2424);
			25741: out = 16'(-1028);
			25742: out = 16'(-1445);
			25743: out = 16'(678);
			25744: out = 16'(1558);
			25745: out = 16'(2054);
			25746: out = 16'(-434);
			25747: out = 16'(2308);
			25748: out = 16'(3524);
			25749: out = 16'(3576);
			25750: out = 16'(912);
			25751: out = 16'(-1672);
			25752: out = 16'(-1204);
			25753: out = 16'(-295);
			25754: out = 16'(1572);
			25755: out = 16'(181);
			25756: out = 16'(256);
			25757: out = 16'(-481);
			25758: out = 16'(1172);
			25759: out = 16'(370);
			25760: out = 16'(-1306);
			25761: out = 16'(-2578);
			25762: out = 16'(-2206);
			25763: out = 16'(404);
			25764: out = 16'(935);
			25765: out = 16'(1292);
			25766: out = 16'(456);
			25767: out = 16'(193);
			25768: out = 16'(-619);
			25769: out = 16'(-1793);
			25770: out = 16'(-2591);
			25771: out = 16'(-2409);
			25772: out = 16'(833);
			25773: out = 16'(2142);
			25774: out = 16'(2683);
			25775: out = 16'(1585);
			25776: out = 16'(1116);
			25777: out = 16'(1305);
			25778: out = 16'(-169);
			25779: out = 16'(-766);
			25780: out = 16'(-1390);
			25781: out = 16'(-161);
			25782: out = 16'(214);
			25783: out = 16'(-247);
			25784: out = 16'(-385);
			25785: out = 16'(-893);
			25786: out = 16'(-3781);
			25787: out = 16'(-1884);
			25788: out = 16'(-69);
			25789: out = 16'(549);
			25790: out = 16'(189);
			25791: out = 16'(-413);
			25792: out = 16'(-484);
			25793: out = 16'(386);
			25794: out = 16'(1344);
			25795: out = 16'(786);
			25796: out = 16'(-1241);
			25797: out = 16'(-4609);
			25798: out = 16'(-3888);
			25799: out = 16'(-2356);
			25800: out = 16'(855);
			25801: out = 16'(1292);
			25802: out = 16'(1431);
			25803: out = 16'(765);
			25804: out = 16'(584);
			25805: out = 16'(501);
			25806: out = 16'(-147);
			25807: out = 16'(802);
			25808: out = 16'(1388);
			25809: out = 16'(1623);
			25810: out = 16'(-125);
			25811: out = 16'(-2118);
			25812: out = 16'(-3420);
			25813: out = 16'(-2044);
			25814: out = 16'(1103);
			25815: out = 16'(3348);
			25816: out = 16'(4498);
			25817: out = 16'(3978);
			25818: out = 16'(1753);
			25819: out = 16'(-79);
			25820: out = 16'(-332);
			25821: out = 16'(-237);
			25822: out = 16'(576);
			25823: out = 16'(1084);
			25824: out = 16'(898);
			25825: out = 16'(128);
			25826: out = 16'(-1145);
			25827: out = 16'(-766);
			25828: out = 16'(453);
			25829: out = 16'(-673);
			25830: out = 16'(-68);
			25831: out = 16'(121);
			25832: out = 16'(677);
			25833: out = 16'(-706);
			25834: out = 16'(-2987);
			25835: out = 16'(-2344);
			25836: out = 16'(-1351);
			25837: out = 16'(371);
			25838: out = 16'(-90);
			25839: out = 16'(-833);
			25840: out = 16'(-1843);
			25841: out = 16'(-2110);
			25842: out = 16'(-1377);
			25843: out = 16'(384);
			25844: out = 16'(2355);
			25845: out = 16'(3364);
			25846: out = 16'(931);
			25847: out = 16'(-276);
			25848: out = 16'(-1192);
			25849: out = 16'(-358);
			25850: out = 16'(226);
			25851: out = 16'(543);
			25852: out = 16'(1309);
			25853: out = 16'(971);
			25854: out = 16'(685);
			25855: out = 16'(-2655);
			25856: out = 16'(-3011);
			25857: out = 16'(-88);
			25858: out = 16'(2571);
			25859: out = 16'(4161);
			25860: out = 16'(1823);
			25861: out = 16'(893);
			25862: out = 16'(-543);
			25863: out = 16'(1447);
			25864: out = 16'(485);
			25865: out = 16'(267);
			25866: out = 16'(-708);
			25867: out = 16'(-97);
			25868: out = 16'(56);
			25869: out = 16'(644);
			25870: out = 16'(-385);
			25871: out = 16'(-1263);
			25872: out = 16'(-4104);
			25873: out = 16'(-3266);
			25874: out = 16'(743);
			25875: out = 16'(2496);
			25876: out = 16'(2933);
			25877: out = 16'(-731);
			25878: out = 16'(-794);
			25879: out = 16'(-1459);
			25880: out = 16'(-246);
			25881: out = 16'(-1504);
			25882: out = 16'(-1920);
			25883: out = 16'(-1374);
			25884: out = 16'(-711);
			25885: out = 16'(-306);
			25886: out = 16'(1231);
			25887: out = 16'(1568);
			25888: out = 16'(2163);
			25889: out = 16'(-753);
			25890: out = 16'(-686);
			25891: out = 16'(588);
			25892: out = 16'(1231);
			25893: out = 16'(280);
			25894: out = 16'(-2888);
			25895: out = 16'(-4514);
			25896: out = 16'(-4956);
			25897: out = 16'(-1782);
			25898: out = 16'(-639);
			25899: out = 16'(1018);
			25900: out = 16'(459);
			25901: out = 16'(1746);
			25902: out = 16'(2216);
			25903: out = 16'(3670);
			25904: out = 16'(2096);
			25905: out = 16'(72);
			25906: out = 16'(-2341);
			25907: out = 16'(-1885);
			25908: out = 16'(704);
			25909: out = 16'(-383);
			25910: out = 16'(-456);
			25911: out = 16'(-1302);
			25912: out = 16'(798);
			25913: out = 16'(1787);
			25914: out = 16'(2910);
			25915: out = 16'(829);
			25916: out = 16'(-1107);
			25917: out = 16'(-3464);
			25918: out = 16'(-2347);
			25919: out = 16'(-534);
			25920: out = 16'(356);
			25921: out = 16'(1902);
			25922: out = 16'(2786);
			25923: out = 16'(938);
			25924: out = 16'(245);
			25925: out = 16'(-97);
			25926: out = 16'(999);
			25927: out = 16'(2057);
			25928: out = 16'(3455);
			25929: out = 16'(562);
			25930: out = 16'(-1706);
			25931: out = 16'(-4637);
			25932: out = 16'(-715);
			25933: out = 16'(2242);
			25934: out = 16'(3100);
			25935: out = 16'(2880);
			25936: out = 16'(1066);
			25937: out = 16'(-704);
			25938: out = 16'(-4163);
			25939: out = 16'(-5881);
			25940: out = 16'(-837);
			25941: out = 16'(1588);
			25942: out = 16'(3509);
			25943: out = 16'(264);
			25944: out = 16'(-73);
			25945: out = 16'(641);
			25946: out = 16'(-941);
			25947: out = 16'(-1224);
			25948: out = 16'(-1275);
			25949: out = 16'(-327);
			25950: out = 16'(-449);
			25951: out = 16'(-983);
			25952: out = 16'(-3375);
			25953: out = 16'(-3616);
			25954: out = 16'(1412);
			25955: out = 16'(1849);
			25956: out = 16'(1874);
			25957: out = 16'(-1715);
			25958: out = 16'(-1071);
			25959: out = 16'(214);
			25960: out = 16'(260);
			25961: out = 16'(648);
			25962: out = 16'(374);
			25963: out = 16'(3237);
			25964: out = 16'(2717);
			25965: out = 16'(1289);
			25966: out = 16'(-2479);
			25967: out = 16'(-3114);
			25968: out = 16'(-159);
			25969: out = 16'(673);
			25970: out = 16'(1714);
			25971: out = 16'(1965);
			25972: out = 16'(1264);
			25973: out = 16'(126);
			25974: out = 16'(-1075);
			25975: out = 16'(-955);
			25976: out = 16'(-9);
			25977: out = 16'(2323);
			25978: out = 16'(3369);
			25979: out = 16'(3763);
			25980: out = 16'(-1251);
			25981: out = 16'(-2913);
			25982: out = 16'(-3710);
			25983: out = 16'(1320);
			25984: out = 16'(3286);
			25985: out = 16'(3972);
			25986: out = 16'(194);
			25987: out = 16'(-1945);
			25988: out = 16'(-2079);
			25989: out = 16'(-1225);
			25990: out = 16'(-323);
			25991: out = 16'(258);
			25992: out = 16'(-1468);
			25993: out = 16'(-3220);
			25994: out = 16'(-3616);
			25995: out = 16'(-2060);
			25996: out = 16'(268);
			25997: out = 16'(-582);
			25998: out = 16'(-213);
			25999: out = 16'(-407);
			26000: out = 16'(1754);
			26001: out = 16'(2133);
			26002: out = 16'(1983);
			26003: out = 16'(972);
			26004: out = 16'(-91);
			26005: out = 16'(-1260);
			26006: out = 16'(-2941);
			26007: out = 16'(-3713);
			26008: out = 16'(-2675);
			26009: out = 16'(-1468);
			26010: out = 16'(167);
			26011: out = 16'(-471);
			26012: out = 16'(2476);
			26013: out = 16'(4300);
			26014: out = 16'(3619);
			26015: out = 16'(1691);
			26016: out = 16'(-856);
			26017: out = 16'(-82);
			26018: out = 16'(-422);
			26019: out = 16'(-131);
			26020: out = 16'(-1222);
			26021: out = 16'(-752);
			26022: out = 16'(362);
			26023: out = 16'(491);
			26024: out = 16'(542);
			26025: out = 16'(503);
			26026: out = 16'(-2);
			26027: out = 16'(-1311);
			26028: out = 16'(-4478);
			26029: out = 16'(-4098);
			26030: out = 16'(-2915);
			26031: out = 16'(515);
			26032: out = 16'(443);
			26033: out = 16'(-200);
			26034: out = 16'(-833);
			26035: out = 16'(-1131);
			26036: out = 16'(-917);
			26037: out = 16'(-1141);
			26038: out = 16'(-258);
			26039: out = 16'(936);
			26040: out = 16'(1873);
			26041: out = 16'(2399);
			26042: out = 16'(2062);
			26043: out = 16'(2793);
			26044: out = 16'(2090);
			26045: out = 16'(-415);
			26046: out = 16'(-1359);
			26047: out = 16'(-2185);
			26048: out = 16'(-1849);
			26049: out = 16'(-1654);
			26050: out = 16'(-669);
			26051: out = 16'(145);
			26052: out = 16'(1178);
			26053: out = 16'(1551);
			26054: out = 16'(4670);
			26055: out = 16'(4401);
			26056: out = 16'(3867);
			26057: out = 16'(-1211);
			26058: out = 16'(-1439);
			26059: out = 16'(336);
			26060: out = 16'(3999);
			26061: out = 16'(4019);
			26062: out = 16'(-234);
			26063: out = 16'(-1247);
			26064: out = 16'(-2548);
			26065: out = 16'(-1907);
			26066: out = 16'(-3226);
			26067: out = 16'(-3209);
			26068: out = 16'(293);
			26069: out = 16'(-962);
			26070: out = 16'(-2083);
			26071: out = 16'(-2811);
			26072: out = 16'(-241);
			26073: out = 16'(3099);
			26074: out = 16'(1327);
			26075: out = 16'(530);
			26076: out = 16'(-1456);
			26077: out = 16'(215);
			26078: out = 16'(239);
			26079: out = 16'(443);
			26080: out = 16'(170);
			26081: out = 16'(652);
			26082: out = 16'(1177);
			26083: out = 16'(2170);
			26084: out = 16'(2595);
			26085: out = 16'(2516);
			26086: out = 16'(1701);
			26087: out = 16'(718);
			26088: out = 16'(-277);
			26089: out = 16'(-236);
			26090: out = 16'(-3);
			26091: out = 16'(-2805);
			26092: out = 16'(-1977);
			26093: out = 16'(-341);
			26094: out = 16'(209);
			26095: out = 16'(222);
			26096: out = 16'(-674);
			26097: out = 16'(95);
			26098: out = 16'(809);
			26099: out = 16'(2728);
			26100: out = 16'(912);
			26101: out = 16'(-230);
			26102: out = 16'(-3108);
			26103: out = 16'(-773);
			26104: out = 16'(354);
			26105: out = 16'(1406);
			26106: out = 16'(-1976);
			26107: out = 16'(-4688);
			26108: out = 16'(-3638);
			26109: out = 16'(-1311);
			26110: out = 16'(1788);
			26111: out = 16'(406);
			26112: out = 16'(1042);
			26113: out = 16'(1172);
			26114: out = 16'(785);
			26115: out = 16'(176);
			26116: out = 16'(-468);
			26117: out = 16'(163);
			26118: out = 16'(-226);
			26119: out = 16'(-2029);
			26120: out = 16'(-2426);
			26121: out = 16'(-1946);
			26122: out = 16'(2249);
			26123: out = 16'(1008);
			26124: out = 16'(660);
			26125: out = 16'(192);
			26126: out = 16'(1646);
			26127: out = 16'(2539);
			26128: out = 16'(695);
			26129: out = 16'(321);
			26130: out = 16'(269);
			26131: out = 16'(-481);
			26132: out = 16'(-411);
			26133: out = 16'(-574);
			26134: out = 16'(2131);
			26135: out = 16'(1745);
			26136: out = 16'(-397);
			26137: out = 16'(-3186);
			26138: out = 16'(-4384);
			26139: out = 16'(-2558);
			26140: out = 16'(-942);
			26141: out = 16'(629);
			26142: out = 16'(-1440);
			26143: out = 16'(39);
			26144: out = 16'(279);
			26145: out = 16'(982);
			26146: out = 16'(-1443);
			26147: out = 16'(-3434);
			26148: out = 16'(-1379);
			26149: out = 16'(339);
			26150: out = 16'(2325);
			26151: out = 16'(1409);
			26152: out = 16'(1612);
			26153: out = 16'(2060);
			26154: out = 16'(397);
			26155: out = 16'(-342);
			26156: out = 16'(-313);
			26157: out = 16'(-271);
			26158: out = 16'(136);
			26159: out = 16'(1319);
			26160: out = 16'(322);
			26161: out = 16'(-766);
			26162: out = 16'(-1838);
			26163: out = 16'(-1187);
			26164: out = 16'(-170);
			26165: out = 16'(-437);
			26166: out = 16'(-565);
			26167: out = 16'(-1003);
			26168: out = 16'(2856);
			26169: out = 16'(3665);
			26170: out = 16'(3948);
			26171: out = 16'(1713);
			26172: out = 16'(856);
			26173: out = 16'(358);
			26174: out = 16'(985);
			26175: out = 16'(836);
			26176: out = 16'(255);
			26177: out = 16'(-1423);
			26178: out = 16'(-1790);
			26179: out = 16'(350);
			26180: out = 16'(1226);
			26181: out = 16'(1577);
			26182: out = 16'(-1175);
			26183: out = 16'(-1813);
			26184: out = 16'(-1960);
			26185: out = 16'(77);
			26186: out = 16'(1064);
			26187: out = 16'(1790);
			26188: out = 16'(550);
			26189: out = 16'(-945);
			26190: out = 16'(-3038);
			26191: out = 16'(-2249);
			26192: out = 16'(-1652);
			26193: out = 16'(-367);
			26194: out = 16'(-378);
			26195: out = 16'(142);
			26196: out = 16'(1184);
			26197: out = 16'(854);
			26198: out = 16'(123);
			26199: out = 16'(-1030);
			26200: out = 16'(-2148);
			26201: out = 16'(-2437);
			26202: out = 16'(969);
			26203: out = 16'(1647);
			26204: out = 16'(1747);
			26205: out = 16'(-2054);
			26206: out = 16'(-3191);
			26207: out = 16'(-3407);
			26208: out = 16'(-1043);
			26209: out = 16'(225);
			26210: out = 16'(645);
			26211: out = 16'(1175);
			26212: out = 16'(1560);
			26213: out = 16'(2016);
			26214: out = 16'(741);
			26215: out = 16'(-1135);
			26216: out = 16'(-4050);
			26217: out = 16'(-4977);
			26218: out = 16'(-4325);
			26219: out = 16'(-346);
			26220: out = 16'(1590);
			26221: out = 16'(3040);
			26222: out = 16'(2175);
			26223: out = 16'(1626);
			26224: out = 16'(370);
			26225: out = 16'(-503);
			26226: out = 16'(-2084);
			26227: out = 16'(-3292);
			26228: out = 16'(-1111);
			26229: out = 16'(454);
			26230: out = 16'(548);
			26231: out = 16'(1049);
			26232: out = 16'(381);
			26233: out = 16'(969);
			26234: out = 16'(-3246);
			26235: out = 16'(-4404);
			26236: out = 16'(-413);
			26237: out = 16'(2707);
			26238: out = 16'(5151);
			26239: out = 16'(4129);
			26240: out = 16'(2898);
			26241: out = 16'(882);
			26242: out = 16'(-688);
			26243: out = 16'(-921);
			26244: out = 16'(51);
			26245: out = 16'(252);
			26246: out = 16'(-453);
			26247: out = 16'(-2914);
			26248: out = 16'(-826);
			26249: out = 16'(303);
			26250: out = 16'(2234);
			26251: out = 16'(543);
			26252: out = 16'(-242);
			26253: out = 16'(-60);
			26254: out = 16'(-258);
			26255: out = 16'(-501);
			26256: out = 16'(-1910);
			26257: out = 16'(-209);
			26258: out = 16'(1654);
			26259: out = 16'(306);
			26260: out = 16'(538);
			26261: out = 16'(411);
			26262: out = 16'(3728);
			26263: out = 16'(2759);
			26264: out = 16'(229);
			26265: out = 16'(-743);
			26266: out = 16'(-1037);
			26267: out = 16'(495);
			26268: out = 16'(-1497);
			26269: out = 16'(-2027);
			26270: out = 16'(-2016);
			26271: out = 16'(-298);
			26272: out = 16'(684);
			26273: out = 16'(-283);
			26274: out = 16'(290);
			26275: out = 16'(48);
			26276: out = 16'(-1653);
			26277: out = 16'(-2384);
			26278: out = 16'(-2299);
			26279: out = 16'(159);
			26280: out = 16'(2224);
			26281: out = 16'(4165);
			26282: out = 16'(1747);
			26283: out = 16'(906);
			26284: out = 16'(280);
			26285: out = 16'(294);
			26286: out = 16'(519);
			26287: out = 16'(1308);
			26288: out = 16'(527);
			26289: out = 16'(223);
			26290: out = 16'(222);
			26291: out = 16'(286);
			26292: out = 16'(-118);
			26293: out = 16'(-1969);
			26294: out = 16'(-1298);
			26295: out = 16'(-28);
			26296: out = 16'(848);
			26297: out = 16'(2322);
			26298: out = 16'(3091);
			26299: out = 16'(1554);
			26300: out = 16'(40);
			26301: out = 16'(-1486);
			26302: out = 16'(-3902);
			26303: out = 16'(-3954);
			26304: out = 16'(-1713);
			26305: out = 16'(-487);
			26306: out = 16'(605);
			26307: out = 16'(-465);
			26308: out = 16'(1502);
			26309: out = 16'(1669);
			26310: out = 16'(687);
			26311: out = 16'(-986);
			26312: out = 16'(-2012);
			26313: out = 16'(-1211);
			26314: out = 16'(-633);
			26315: out = 16'(-232);
			26316: out = 16'(-2420);
			26317: out = 16'(-2419);
			26318: out = 16'(-1586);
			26319: out = 16'(-661);
			26320: out = 16'(0);
			26321: out = 16'(-380);
			26322: out = 16'(2883);
			26323: out = 16'(3077);
			26324: out = 16'(2102);
			26325: out = 16'(-1766);
			26326: out = 16'(-3988);
			26327: out = 16'(-4158);
			26328: out = 16'(-1274);
			26329: out = 16'(1607);
			26330: out = 16'(2539);
			26331: out = 16'(1973);
			26332: out = 16'(294);
			26333: out = 16'(1709);
			26334: out = 16'(335);
			26335: out = 16'(-317);
			26336: out = 16'(-1884);
			26337: out = 16'(-1036);
			26338: out = 16'(45);
			26339: out = 16'(2864);
			26340: out = 16'(3064);
			26341: out = 16'(1862);
			26342: out = 16'(-240);
			26343: out = 16'(-1790);
			26344: out = 16'(-2672);
			26345: out = 16'(-1220);
			26346: out = 16'(-2);
			26347: out = 16'(334);
			26348: out = 16'(154);
			26349: out = 16'(105);
			26350: out = 16'(1972);
			26351: out = 16'(2351);
			26352: out = 16'(2531);
			26353: out = 16'(675);
			26354: out = 16'(387);
			26355: out = 16'(234);
			26356: out = 16'(205);
			26357: out = 16'(379);
			26358: out = 16'(428);
			26359: out = 16'(1114);
			26360: out = 16'(285);
			26361: out = 16'(-2275);
			26362: out = 16'(-931);
			26363: out = 16'(159);
			26364: out = 16'(2724);
			26365: out = 16'(642);
			26366: out = 16'(-524);
			26367: out = 16'(-513);
			26368: out = 16'(-172);
			26369: out = 16'(279);
			26370: out = 16'(-311);
			26371: out = 16'(-235);
			26372: out = 16'(-457);
			26373: out = 16'(-1648);
			26374: out = 16'(-3042);
			26375: out = 16'(-4388);
			26376: out = 16'(-2324);
			26377: out = 16'(-1023);
			26378: out = 16'(639);
			26379: out = 16'(-223);
			26380: out = 16'(-79);
			26381: out = 16'(-142);
			26382: out = 16'(1572);
			26383: out = 16'(1701);
			26384: out = 16'(-28);
			26385: out = 16'(-1992);
			26386: out = 16'(-3924);
			26387: out = 16'(-4824);
			26388: out = 16'(-3470);
			26389: out = 16'(-897);
			26390: out = 16'(-687);
			26391: out = 16'(1995);
			26392: out = 16'(3628);
			26393: out = 16'(3215);
			26394: out = 16'(1612);
			26395: out = 16'(-241);
			26396: out = 16'(465);
			26397: out = 16'(1296);
			26398: out = 16'(2011);
			26399: out = 16'(2744);
			26400: out = 16'(2061);
			26401: out = 16'(778);
			26402: out = 16'(-2180);
			26403: out = 16'(-3052);
			26404: out = 16'(365);
			26405: out = 16'(2073);
			26406: out = 16'(3411);
			26407: out = 16'(1233);
			26408: out = 16'(917);
			26409: out = 16'(8);
			26410: out = 16'(-191);
			26411: out = 16'(-1483);
			26412: out = 16'(-2744);
			26413: out = 16'(66);
			26414: out = 16'(650);
			26415: out = 16'(525);
			26416: out = 16'(-1883);
			26417: out = 16'(-2516);
			26418: out = 16'(-886);
			26419: out = 16'(-553);
			26420: out = 16'(289);
			26421: out = 16'(475);
			26422: out = 16'(1614);
			26423: out = 16'(1864);
			26424: out = 16'(648);
			26425: out = 16'(197);
			26426: out = 16'(-272);
			26427: out = 16'(-58);
			26428: out = 16'(-953);
			26429: out = 16'(-2026);
			26430: out = 16'(-1805);
			26431: out = 16'(-1878);
			26432: out = 16'(-1726);
			26433: out = 16'(-1240);
			26434: out = 16'(-564);
			26435: out = 16'(40);
			26436: out = 16'(559);
			26437: out = 16'(790);
			26438: out = 16'(716);
			26439: out = 16'(723);
			26440: out = 16'(913);
			26441: out = 16'(2140);
			26442: out = 16'(878);
			26443: out = 16'(-509);
			26444: out = 16'(-1590);
			26445: out = 16'(-2005);
			26446: out = 16'(-1480);
			26447: out = 16'(32);
			26448: out = 16'(1401);
			26449: out = 16'(2026);
			26450: out = 16'(1667);
			26451: out = 16'(415);
			26452: out = 16'(-1098);
			26453: out = 16'(-1838);
			26454: out = 16'(-815);
			26455: out = 16'(2209);
			26456: out = 16'(1996);
			26457: out = 16'(1608);
			26458: out = 16'(-287);
			26459: out = 16'(312);
			26460: out = 16'(450);
			26461: out = 16'(-212);
			26462: out = 16'(-197);
			26463: out = 16'(-122);
			26464: out = 16'(1211);
			26465: out = 16'(775);
			26466: out = 16'(184);
			26467: out = 16'(-1141);
			26468: out = 16'(-309);
			26469: out = 16'(1345);
			26470: out = 16'(41);
			26471: out = 16'(-832);
			26472: out = 16'(-2064);
			26473: out = 16'(-1960);
			26474: out = 16'(-1914);
			26475: out = 16'(-1959);
			26476: out = 16'(-370);
			26477: out = 16'(596);
			26478: out = 16'(349);
			26479: out = 16'(410);
			26480: out = 16'(690);
			26481: out = 16'(2605);
			26482: out = 16'(2395);
			26483: out = 16'(1559);
			26484: out = 16'(-731);
			26485: out = 16'(-2109);
			26486: out = 16'(-2765);
			26487: out = 16'(-4246);
			26488: out = 16'(-3178);
			26489: out = 16'(-758);
			26490: out = 16'(835);
			26491: out = 16'(1296);
			26492: out = 16'(-284);
			26493: out = 16'(691);
			26494: out = 16'(375);
			26495: out = 16'(-121);
			26496: out = 16'(-1878);
			26497: out = 16'(-1846);
			26498: out = 16'(2854);
			26499: out = 16'(2362);
			26500: out = 16'(1805);
			26501: out = 16'(-969);
			26502: out = 16'(-711);
			26503: out = 16'(-299);
			26504: out = 16'(412);
			26505: out = 16'(319);
			26506: out = 16'(507);
			26507: out = 16'(-1050);
			26508: out = 16'(-357);
			26509: out = 16'(622);
			26510: out = 16'(3427);
			26511: out = 16'(3136);
			26512: out = 16'(493);
			26513: out = 16'(-1724);
			26514: out = 16'(-2365);
			26515: out = 16'(389);
			26516: out = 16'(2059);
			26517: out = 16'(3691);
			26518: out = 16'(3729);
			26519: out = 16'(2935);
			26520: out = 16'(1105);
			26521: out = 16'(-1671);
			26522: out = 16'(-2083);
			26523: out = 16'(-1096);
			26524: out = 16'(-897);
			26525: out = 16'(-367);
			26526: out = 16'(-732);
			26527: out = 16'(-381);
			26528: out = 16'(-707);
			26529: out = 16'(-365);
			26530: out = 16'(-1246);
			26531: out = 16'(-786);
			26532: out = 16'(172);
			26533: out = 16'(1004);
			26534: out = 16'(1132);
			26535: out = 16'(1316);
			26536: out = 16'(117);
			26537: out = 16'(-922);
			26538: out = 16'(-3623);
			26539: out = 16'(-2358);
			26540: out = 16'(-1060);
			26541: out = 16'(-39);
			26542: out = 16'(-2262);
			26543: out = 16'(-5452);
			26544: out = 16'(-5084);
			26545: out = 16'(-3189);
			26546: out = 16'(1114);
			26547: out = 16'(-2040);
			26548: out = 16'(-1713);
			26549: out = 16'(40);
			26550: out = 16'(108);
			26551: out = 16'(247);
			26552: out = 16'(-120);
			26553: out = 16'(1504);
			26554: out = 16'(2670);
			26555: out = 16'(3631);
			26556: out = 16'(2013);
			26557: out = 16'(167);
			26558: out = 16'(21);
			26559: out = 16'(-225);
			26560: out = 16'(164);
			26561: out = 16'(-120);
			26562: out = 16'(406);
			26563: out = 16'(710);
			26564: out = 16'(796);
			26565: out = 16'(643);
			26566: out = 16'(776);
			26567: out = 16'(28);
			26568: out = 16'(510);
			26569: out = 16'(2131);
			26570: out = 16'(2056);
			26571: out = 16'(1760);
			26572: out = 16'(318);
			26573: out = 16'(1289);
			26574: out = 16'(2293);
			26575: out = 16'(3083);
			26576: out = 16'(3278);
			26577: out = 16'(2940);
			26578: out = 16'(2634);
			26579: out = 16'(1279);
			26580: out = 16'(-272);
			26581: out = 16'(-2494);
			26582: out = 16'(-3160);
			26583: out = 16'(-2799);
			26584: out = 16'(-1788);
			26585: out = 16'(-838);
			26586: out = 16'(-316);
			26587: out = 16'(130);
			26588: out = 16'(164);
			26589: out = 16'(-315);
			26590: out = 16'(635);
			26591: out = 16'(1148);
			26592: out = 16'(150);
			26593: out = 16'(-6);
			26594: out = 16'(-365);
			26595: out = 16'(472);
			26596: out = 16'(236);
			26597: out = 16'(142);
			26598: out = 16'(-1222);
			26599: out = 16'(-1252);
			26600: out = 16'(-1328);
			26601: out = 16'(-303);
			26602: out = 16'(-397);
			26603: out = 16'(-131);
			26604: out = 16'(-3471);
			26605: out = 16'(-4417);
			26606: out = 16'(-4376);
			26607: out = 16'(1031);
			26608: out = 16'(3393);
			26609: out = 16'(-462);
			26610: out = 16'(216);
			26611: out = 16'(-196);
			26612: out = 16'(1640);
			26613: out = 16'(-485);
			26614: out = 16'(-1873);
			26615: out = 16'(-453);
			26616: out = 16'(-116);
			26617: out = 16'(-112);
			26618: out = 16'(-9);
			26619: out = 16'(-149);
			26620: out = 16'(8);
			26621: out = 16'(-308);
			26622: out = 16'(-398);
			26623: out = 16'(-1213);
			26624: out = 16'(426);
			26625: out = 16'(416);
			26626: out = 16'(139);
			26627: out = 16'(-2320);
			26628: out = 16'(-2960);
			26629: out = 16'(-326);
			26630: out = 16'(1228);
			26631: out = 16'(1971);
			26632: out = 16'(-761);
			26633: out = 16'(-1781);
			26634: out = 16'(-2371);
			26635: out = 16'(-302);
			26636: out = 16'(1308);
			26637: out = 16'(2947);
			26638: out = 16'(1111);
			26639: out = 16'(289);
			26640: out = 16'(-229);
			26641: out = 16'(-453);
			26642: out = 16'(480);
			26643: out = 16'(2054);
			26644: out = 16'(2650);
			26645: out = 16'(2133);
			26646: out = 16'(512);
			26647: out = 16'(-1254);
			26648: out = 16'(-1264);
			26649: out = 16'(2365);
			26650: out = 16'(4444);
			26651: out = 16'(5263);
			26652: out = 16'(178);
			26653: out = 16'(-1939);
			26654: out = 16'(-4013);
			26655: out = 16'(-4193);
			26656: out = 16'(-5035);
			26657: out = 16'(-5759);
			26658: out = 16'(531);
			26659: out = 16'(2754);
			26660: out = 16'(2632);
			26661: out = 16'(659);
			26662: out = 16'(-581);
			26663: out = 16'(126);
			26664: out = 16'(-419);
			26665: out = 16'(-148);
			26666: out = 16'(-211);
			26667: out = 16'(808);
			26668: out = 16'(1152);
			26669: out = 16'(-1034);
			26670: out = 16'(-1077);
			26671: out = 16'(-847);
			26672: out = 16'(2468);
			26673: out = 16'(2137);
			26674: out = 16'(1098);
			26675: out = 16'(-1429);
			26676: out = 16'(-1543);
			26677: out = 16'(-200);
			26678: out = 16'(904);
			26679: out = 16'(1223);
			26680: out = 16'(477);
			26681: out = 16'(-1094);
			26682: out = 16'(-1870);
			26683: out = 16'(-183);
			26684: out = 16'(499);
			26685: out = 16'(1588);
			26686: out = 16'(242);
			26687: out = 16'(1659);
			26688: out = 16'(1718);
			26689: out = 16'(2338);
			26690: out = 16'(-881);
			26691: out = 16'(-3714);
			26692: out = 16'(-2296);
			26693: out = 16'(-259);
			26694: out = 16'(2102);
			26695: out = 16'(151);
			26696: out = 16'(-1793);
			26697: out = 16'(-4439);
			26698: out = 16'(-4283);
			26699: out = 16'(-3895);
			26700: out = 16'(-3365);
			26701: out = 16'(492);
			26702: out = 16'(2809);
			26703: out = 16'(2767);
			26704: out = 16'(1768);
			26705: out = 16'(446);
			26706: out = 16'(702);
			26707: out = 16'(122);
			26708: out = 16'(60);
			26709: out = 16'(614);
			26710: out = 16'(636);
			26711: out = 16'(469);
			26712: out = 16'(591);
			26713: out = 16'(1200);
			26714: out = 16'(2084);
			26715: out = 16'(1462);
			26716: out = 16'(1171);
			26717: out = 16'(1368);
			26718: out = 16'(-591);
			26719: out = 16'(-1093);
			26720: out = 16'(-486);
			26721: out = 16'(1612);
			26722: out = 16'(2333);
			26723: out = 16'(-500);
			26724: out = 16'(-903);
			26725: out = 16'(-760);
			26726: out = 16'(3727);
			26727: out = 16'(3544);
			26728: out = 16'(2786);
			26729: out = 16'(-895);
			26730: out = 16'(-985);
			26731: out = 16'(317);
			26732: out = 16'(-1326);
			26733: out = 16'(-920);
			26734: out = 16'(-385);
			26735: out = 16'(2465);
			26736: out = 16'(2348);
			26737: out = 16'(-664);
			26738: out = 16'(-893);
			26739: out = 16'(-1798);
			26740: out = 16'(-1966);
			26741: out = 16'(-2731);
			26742: out = 16'(-2469);
			26743: out = 16'(-617);
			26744: out = 16'(-262);
			26745: out = 16'(-247);
			26746: out = 16'(-186);
			26747: out = 16'(-334);
			26748: out = 16'(-394);
			26749: out = 16'(-264);
			26750: out = 16'(101);
			26751: out = 16'(528);
			26752: out = 16'(-808);
			26753: out = 16'(-1538);
			26754: out = 16'(-1904);
			26755: out = 16'(-1391);
			26756: out = 16'(-960);
			26757: out = 16'(-1188);
			26758: out = 16'(593);
			26759: out = 16'(1744);
			26760: out = 16'(2729);
			26761: out = 16'(1384);
			26762: out = 16'(138);
			26763: out = 16'(656);
			26764: out = 16'(1125);
			26765: out = 16'(1715);
			26766: out = 16'(-3998);
			26767: out = 16'(-3695);
			26768: out = 16'(-2374);
			26769: out = 16'(1956);
			26770: out = 16'(2188);
			26771: out = 16'(318);
			26772: out = 16'(-1131);
			26773: out = 16'(-2391);
			26774: out = 16'(-2503);
			26775: out = 16'(-1688);
			26776: out = 16'(-386);
			26777: out = 16'(602);
			26778: out = 16'(824);
			26779: out = 16'(580);
			26780: out = 16'(601);
			26781: out = 16'(-55);
			26782: out = 16'(-281);
			26783: out = 16'(-344);
			26784: out = 16'(-90);
			26785: out = 16'(-124);
			26786: out = 16'(-119);
			26787: out = 16'(-978);
			26788: out = 16'(-1727);
			26789: out = 16'(-44);
			26790: out = 16'(1446);
			26791: out = 16'(2799);
			26792: out = 16'(2371);
			26793: out = 16'(1363);
			26794: out = 16'(-105);
			26795: out = 16'(-374);
			26796: out = 16'(-74);
			26797: out = 16'(415);
			26798: out = 16'(3085);
			26799: out = 16'(4500);
			26800: out = 16'(1879);
			26801: out = 16'(726);
			26802: out = 16'(-663);
			26803: out = 16'(2511);
			26804: out = 16'(1402);
			26805: out = 16'(200);
			26806: out = 16'(-1189);
			26807: out = 16'(-1048);
			26808: out = 16'(-306);
			26809: out = 16'(25);
			26810: out = 16'(-75);
			26811: out = 16'(-664);
			26812: out = 16'(-1163);
			26813: out = 16'(-1082);
			26814: out = 16'(242);
			26815: out = 16'(126);
			26816: out = 16'(-129);
			26817: out = 16'(-2187);
			26818: out = 16'(-765);
			26819: out = 16'(861);
			26820: out = 16'(3611);
			26821: out = 16'(3893);
			26822: out = 16'(3481);
			26823: out = 16'(1341);
			26824: out = 16'(294);
			26825: out = 16'(-627);
			26826: out = 16'(84);
			26827: out = 16'(-596);
			26828: out = 16'(-1469);
			26829: out = 16'(-3322);
			26830: out = 16'(-2989);
			26831: out = 16'(-120);
			26832: out = 16'(12);
			26833: out = 16'(475);
			26834: out = 16'(-576);
			26835: out = 16'(1524);
			26836: out = 16'(2374);
			26837: out = 16'(1080);
			26838: out = 16'(220);
			26839: out = 16'(-862);
			26840: out = 16'(-215);
			26841: out = 16'(-1323);
			26842: out = 16'(-2106);
			26843: out = 16'(-1572);
			26844: out = 16'(-309);
			26845: out = 16'(1125);
			26846: out = 16'(-719);
			26847: out = 16'(-2083);
			26848: out = 16'(-3512);
			26849: out = 16'(-2951);
			26850: out = 16'(-2318);
			26851: out = 16'(-1912);
			26852: out = 16'(-732);
			26853: out = 16'(-290);
			26854: out = 16'(-189);
			26855: out = 16'(-1560);
			26856: out = 16'(-2672);
			26857: out = 16'(-3213);
			26858: out = 16'(-1394);
			26859: out = 16'(1082);
			26860: out = 16'(1158);
			26861: out = 16'(1936);
			26862: out = 16'(1943);
			26863: out = 16'(1051);
			26864: out = 16'(491);
			26865: out = 16'(852);
			26866: out = 16'(935);
			26867: out = 16'(2079);
			26868: out = 16'(3108);
			26869: out = 16'(4278);
			26870: out = 16'(3179);
			26871: out = 16'(-1253);
			26872: out = 16'(-1746);
			26873: out = 16'(-1505);
			26874: out = 16'(1833);
			26875: out = 16'(1013);
			26876: out = 16'(386);
			26877: out = 16'(1074);
			26878: out = 16'(1037);
			26879: out = 16'(980);
			26880: out = 16'(-215);
			26881: out = 16'(-148);
			26882: out = 16'(372);
			26883: out = 16'(-979);
			26884: out = 16'(-1609);
			26885: out = 16'(-2033);
			26886: out = 16'(-365);
			26887: out = 16'(-244);
			26888: out = 16'(-3015);
			26889: out = 16'(-996);
			26890: out = 16'(-234);
			26891: out = 16'(1481);
			26892: out = 16'(-1670);
			26893: out = 16'(-3277);
			26894: out = 16'(-1336);
			26895: out = 16'(1167);
			26896: out = 16'(3403);
			26897: out = 16'(1284);
			26898: out = 16'(859);
			26899: out = 16'(74);
			26900: out = 16'(-866);
			26901: out = 16'(-1732);
			26902: out = 16'(-2691);
			26903: out = 16'(-35);
			26904: out = 16'(424);
			26905: out = 16'(-122);
			26906: out = 16'(-1879);
			26907: out = 16'(-2204);
			26908: out = 16'(-266);
			26909: out = 16'(1093);
			26910: out = 16'(2466);
			26911: out = 16'(3760);
			26912: out = 16'(2471);
			26913: out = 16'(284);
			26914: out = 16'(-3764);
			26915: out = 16'(-4159);
			26916: out = 16'(-2956);
			26917: out = 16'(-254);
			26918: out = 16'(731);
			26919: out = 16'(577);
			26920: out = 16'(2804);
			26921: out = 16'(3299);
			26922: out = 16'(3017);
			26923: out = 16'(1249);
			26924: out = 16'(-201);
			26925: out = 16'(-256);
			26926: out = 16'(-3363);
			26927: out = 16'(-3825);
			26928: out = 16'(-1266);
			26929: out = 16'(1079);
			26930: out = 16'(2657);
			26931: out = 16'(1095);
			26932: out = 16'(526);
			26933: out = 16'(-466);
			26934: out = 16'(-188);
			26935: out = 16'(218);
			26936: out = 16'(1480);
			26937: out = 16'(2592);
			26938: out = 16'(3287);
			26939: out = 16'(2668);
			26940: out = 16'(1723);
			26941: out = 16'(-551);
			26942: out = 16'(-2839);
			26943: out = 16'(-4838);
			26944: out = 16'(-4222);
			26945: out = 16'(-440);
			26946: out = 16'(1369);
			26947: out = 16'(2328);
			26948: out = 16'(-761);
			26949: out = 16'(-154);
			26950: out = 16'(-180);
			26951: out = 16'(3275);
			26952: out = 16'(721);
			26953: out = 16'(-1549);
			26954: out = 16'(-2819);
			26955: out = 16'(-619);
			26956: out = 16'(2689);
			26957: out = 16'(21);
			26958: out = 16'(-947);
			26959: out = 16'(-2105);
			26960: out = 16'(-1456);
			26961: out = 16'(-774);
			26962: out = 16'(237);
			26963: out = 16'(465);
			26964: out = 16'(202);
			26965: out = 16'(-358);
			26966: out = 16'(-2377);
			26967: out = 16'(-3622);
			26968: out = 16'(-3416);
			26969: out = 16'(-1825);
			26970: out = 16'(285);
			26971: out = 16'(1716);
			26972: out = 16'(1864);
			26973: out = 16'(1018);
			26974: out = 16'(183);
			26975: out = 16'(-372);
			26976: out = 16'(-249);
			26977: out = 16'(-505);
			26978: out = 16'(243);
			26979: out = 16'(1302);
			26980: out = 16'(195);
			26981: out = 16'(-124);
			26982: out = 16'(438);
			26983: out = 16'(-62);
			26984: out = 16'(-161);
			26985: out = 16'(-420);
			26986: out = 16'(-355);
			26987: out = 16'(-434);
			26988: out = 16'(-310);
			26989: out = 16'(-459);
			26990: out = 16'(-157);
			26991: out = 16'(363);
			26992: out = 16'(1281);
			26993: out = 16'(1861);
			26994: out = 16'(1414);
			26995: out = 16'(733);
			26996: out = 16'(296);
			26997: out = 16'(-1672);
			26998: out = 16'(-1038);
			26999: out = 16'(1288);
			27000: out = 16'(1754);
			27001: out = 16'(557);
			27002: out = 16'(-4437);
			27003: out = 16'(-3742);
			27004: out = 16'(-2429);
			27005: out = 16'(2708);
			27006: out = 16'(1309);
			27007: out = 16'(224);
			27008: out = 16'(376);
			27009: out = 16'(325);
			27010: out = 16'(329);
			27011: out = 16'(343);
			27012: out = 16'(163);
			27013: out = 16'(-197);
			27014: out = 16'(-123);
			27015: out = 16'(-4);
			27016: out = 16'(438);
			27017: out = 16'(-291);
			27018: out = 16'(-170);
			27019: out = 16'(359);
			27020: out = 16'(939);
			27021: out = 16'(1756);
			27022: out = 16'(3861);
			27023: out = 16'(1752);
			27024: out = 16'(-174);
			27025: out = 16'(-1813);
			27026: out = 16'(-1346);
			27027: out = 16'(-179);
			27028: out = 16'(-14);
			27029: out = 16'(794);
			27030: out = 16'(1240);
			27031: out = 16'(3396);
			27032: out = 16'(3451);
			27033: out = 16'(2782);
			27034: out = 16'(259);
			27035: out = 16'(-566);
			27036: out = 16'(203);
			27037: out = 16'(-190);
			27038: out = 16'(382);
			27039: out = 16'(775);
			27040: out = 16'(1035);
			27041: out = 16'(563);
			27042: out = 16'(200);
			27043: out = 16'(-1845);
			27044: out = 16'(-3147);
			27045: out = 16'(-3731);
			27046: out = 16'(-1847);
			27047: out = 16'(709);
			27048: out = 16'(2530);
			27049: out = 16'(2953);
			27050: out = 16'(1915);
			27051: out = 16'(686);
			27052: out = 16'(-1245);
			27053: out = 16'(-2925);
			27054: out = 16'(-1849);
			27055: out = 16'(-811);
			27056: out = 16'(58);
			27057: out = 16'(-298);
			27058: out = 16'(-764);
			27059: out = 16'(-429);
			27060: out = 16'(-1580);
			27061: out = 16'(-2129);
			27062: out = 16'(-2811);
			27063: out = 16'(-1328);
			27064: out = 16'(14);
			27065: out = 16'(209);
			27066: out = 16'(-14);
			27067: out = 16'(-545);
			27068: out = 16'(-1042);
			27069: out = 16'(-897);
			27070: out = 16'(-342);
			27071: out = 16'(199);
			27072: out = 16'(-268);
			27073: out = 16'(-2014);
			27074: out = 16'(-178);
			27075: out = 16'(811);
			27076: out = 16'(1996);
			27077: out = 16'(523);
			27078: out = 16'(-376);
			27079: out = 16'(-311);
			27080: out = 16'(-496);
			27081: out = 16'(-318);
			27082: out = 16'(-509);
			27083: out = 16'(62);
			27084: out = 16'(221);
			27085: out = 16'(-197);
			27086: out = 16'(-1112);
			27087: out = 16'(-1711);
			27088: out = 16'(31);
			27089: out = 16'(2113);
			27090: out = 16'(4601);
			27091: out = 16'(4418);
			27092: out = 16'(3097);
			27093: out = 16'(-688);
			27094: out = 16'(228);
			27095: out = 16'(-185);
			27096: out = 16'(-142);
			27097: out = 16'(-2105);
			27098: out = 16'(-2388);
			27099: out = 16'(226);
			27100: out = 16'(1180);
			27101: out = 16'(1519);
			27102: out = 16'(-1138);
			27103: out = 16'(-1068);
			27104: out = 16'(-386);
			27105: out = 16'(-489);
			27106: out = 16'(33);
			27107: out = 16'(200);
			27108: out = 16'(3640);
			27109: out = 16'(4256);
			27110: out = 16'(4141);
			27111: out = 16'(-2260);
			27112: out = 16'(-4784);
			27113: out = 16'(-2507);
			27114: out = 16'(-1734);
			27115: out = 16'(-11);
			27116: out = 16'(-800);
			27117: out = 16'(1985);
			27118: out = 16'(2635);
			27119: out = 16'(621);
			27120: out = 16'(-1779);
			27121: out = 16'(-3834);
			27122: out = 16'(-2775);
			27123: out = 16'(-2172);
			27124: out = 16'(-1062);
			27125: out = 16'(-2554);
			27126: out = 16'(-2326);
			27127: out = 16'(-1736);
			27128: out = 16'(-171);
			27129: out = 16'(1199);
			27130: out = 16'(2672);
			27131: out = 16'(2566);
			27132: out = 16'(2129);
			27133: out = 16'(92);
			27134: out = 16'(418);
			27135: out = 16'(-14);
			27136: out = 16'(582);
			27137: out = 16'(-2885);
			27138: out = 16'(-5191);
			27139: out = 16'(-3498);
			27140: out = 16'(-1171);
			27141: out = 16'(1777);
			27142: out = 16'(-422);
			27143: out = 16'(209);
			27144: out = 16'(343);
			27145: out = 16'(1922);
			27146: out = 16'(1452);
			27147: out = 16'(587);
			27148: out = 16'(488);
			27149: out = 16'(477);
			27150: out = 16'(-361);
			27151: out = 16'(41);
			27152: out = 16'(-472);
			27153: out = 16'(6);
			27154: out = 16'(-2999);
			27155: out = 16'(-3509);
			27156: out = 16'(14);
			27157: out = 16'(2841);
			27158: out = 16'(4469);
			27159: out = 16'(2910);
			27160: out = 16'(126);
			27161: out = 16'(-2997);
			27162: out = 16'(-3381);
			27163: out = 16'(-1462);
			27164: out = 16'(2422);
			27165: out = 16'(2827);
			27166: out = 16'(2407);
			27167: out = 16'(-857);
			27168: out = 16'(-189);
			27169: out = 16'(-322);
			27170: out = 16'(1490);
			27171: out = 16'(-16);
			27172: out = 16'(-97);
			27173: out = 16'(-715);
			27174: out = 16'(1048);
			27175: out = 16'(1866);
			27176: out = 16'(2635);
			27177: out = 16'(169);
			27178: out = 16'(-2387);
			27179: out = 16'(-2633);
			27180: out = 16'(-1789);
			27181: out = 16'(33);
			27182: out = 16'(-560);
			27183: out = 16'(-563);
			27184: out = 16'(-1292);
			27185: out = 16'(779);
			27186: out = 16'(1070);
			27187: out = 16'(442);
			27188: out = 16'(390);
			27189: out = 16'(121);
			27190: out = 16'(-182);
			27191: out = 16'(-796);
			27192: out = 16'(-1644);
			27193: out = 16'(-4212);
			27194: out = 16'(-2545);
			27195: out = 16'(-836);
			27196: out = 16'(-2605);
			27197: out = 16'(-1677);
			27198: out = 16'(-708);
			27199: out = 16'(1159);
			27200: out = 16'(1495);
			27201: out = 16'(1353);
			27202: out = 16'(206);
			27203: out = 16'(701);
			27204: out = 16'(2915);
			27205: out = 16'(968);
			27206: out = 16'(584);
			27207: out = 16'(266);
			27208: out = 16'(667);
			27209: out = 16'(233);
			27210: out = 16'(-133);
			27211: out = 16'(-2689);
			27212: out = 16'(-4508);
			27213: out = 16'(-5622);
			27214: out = 16'(-3322);
			27215: out = 16'(10);
			27216: out = 16'(2178);
			27217: out = 16'(3968);
			27218: out = 16'(4457);
			27219: out = 16'(2601);
			27220: out = 16'(548);
			27221: out = 16'(-2072);
			27222: out = 16'(-1009);
			27223: out = 16'(-1572);
			27224: out = 16'(-2386);
			27225: out = 16'(-2696);
			27226: out = 16'(-1212);
			27227: out = 16'(2067);
			27228: out = 16'(3805);
			27229: out = 16'(4586);
			27230: out = 16'(3966);
			27231: out = 16'(1917);
			27232: out = 16'(-274);
			27233: out = 16'(-1707);
			27234: out = 16'(-1012);
			27235: out = 16'(495);
			27236: out = 16'(-1150);
			27237: out = 16'(-1041);
			27238: out = 16'(-1065);
			27239: out = 16'(1489);
			27240: out = 16'(1800);
			27241: out = 16'(1122);
			27242: out = 16'(1721);
			27243: out = 16'(2426);
			27244: out = 16'(4542);
			27245: out = 16'(1031);
			27246: out = 16'(-1210);
			27247: out = 16'(-3641);
			27248: out = 16'(-1595);
			27249: out = 16'(-13);
			27250: out = 16'(225);
			27251: out = 16'(-1690);
			27252: out = 16'(-3856);
			27253: out = 16'(-3287);
			27254: out = 16'(-2564);
			27255: out = 16'(-639);
			27256: out = 16'(-1352);
			27257: out = 16'(-183);
			27258: out = 16'(366);
			27259: out = 16'(2471);
			27260: out = 16'(1787);
			27261: out = 16'(-175);
			27262: out = 16'(-814);
			27263: out = 16'(-770);
			27264: out = 16'(410);
			27265: out = 16'(409);
			27266: out = 16'(98);
			27267: out = 16'(-1020);
			27268: out = 16'(-747);
			27269: out = 16'(0);
			27270: out = 16'(347);
			27271: out = 16'(2099);
			27272: out = 16'(3159);
			27273: out = 16'(1510);
			27274: out = 16'(142);
			27275: out = 16'(-1241);
			27276: out = 16'(-1795);
			27277: out = 16'(-1061);
			27278: out = 16'(499);
			27279: out = 16'(610);
			27280: out = 16'(-44);
			27281: out = 16'(-1853);
			27282: out = 16'(-2859);
			27283: out = 16'(-2684);
			27284: out = 16'(123);
			27285: out = 16'(1167);
			27286: out = 16'(2168);
			27287: out = 16'(266);
			27288: out = 16'(675);
			27289: out = 16'(180);
			27290: out = 16'(751);
			27291: out = 16'(-1127);
			27292: out = 16'(-2641);
			27293: out = 16'(-4707);
			27294: out = 16'(-3282);
			27295: out = 16'(-450);
			27296: out = 16'(2089);
			27297: out = 16'(2297);
			27298: out = 16'(-279);
			27299: out = 16'(1343);
			27300: out = 16'(1314);
			27301: out = 16'(1566);
			27302: out = 16'(231);
			27303: out = 16'(-215);
			27304: out = 16'(-39);
			27305: out = 16'(408);
			27306: out = 16'(702);
			27307: out = 16'(501);
			27308: out = 16'(215);
			27309: out = 16'(-32);
			27310: out = 16'(600);
			27311: out = 16'(576);
			27312: out = 16'(504);
			27313: out = 16'(1707);
			27314: out = 16'(2431);
			27315: out = 16'(3222);
			27316: out = 16'(1077);
			27317: out = 16'(278);
			27318: out = 16'(269);
			27319: out = 16'(-718);
			27320: out = 16'(-1780);
			27321: out = 16'(-3361);
			27322: out = 16'(-3925);
			27323: out = 16'(-3587);
			27324: out = 16'(-316);
			27325: out = 16'(-114);
			27326: out = 16'(-116);
			27327: out = 16'(-2359);
			27328: out = 16'(-1377);
			27329: out = 16'(67);
			27330: out = 16'(394);
			27331: out = 16'(364);
			27332: out = 16'(-247);
			27333: out = 16'(503);
			27334: out = 16'(324);
			27335: out = 16'(-188);
			27336: out = 16'(473);
			27337: out = 16'(1275);
			27338: out = 16'(2782);
			27339: out = 16'(1795);
			27340: out = 16'(1104);
			27341: out = 16'(634);
			27342: out = 16'(594);
			27343: out = 16'(573);
			27344: out = 16'(569);
			27345: out = 16'(541);
			27346: out = 16'(509);
			27347: out = 16'(-313);
			27348: out = 16'(-260);
			27349: out = 16'(-163);
			27350: out = 16'(397);
			27351: out = 16'(-684);
			27352: out = 16'(-2678);
			27353: out = 16'(-677);
			27354: out = 16'(892);
			27355: out = 16'(3371);
			27356: out = 16'(1795);
			27357: out = 16'(819);
			27358: out = 16'(-216);
			27359: out = 16'(-280);
			27360: out = 16'(-221);
			27361: out = 16'(301);
			27362: out = 16'(-942);
			27363: out = 16'(-2499);
			27364: out = 16'(-4681);
			27365: out = 16'(-5228);
			27366: out = 16'(-4376);
			27367: out = 16'(-467);
			27368: out = 16'(2042);
			27369: out = 16'(3270);
			27370: out = 16'(1453);
			27371: out = 16'(-1019);
			27372: out = 16'(-4138);
			27373: out = 16'(-1943);
			27374: out = 16'(608);
			27375: out = 16'(4068);
			27376: out = 16'(3654);
			27377: out = 16'(2651);
			27378: out = 16'(480);
			27379: out = 16'(-577);
			27380: out = 16'(-989);
			27381: out = 16'(266);
			27382: out = 16'(1164);
			27383: out = 16'(1966);
			27384: out = 16'(589);
			27385: out = 16'(-118);
			27386: out = 16'(-1248);
			27387: out = 16'(1620);
			27388: out = 16'(1805);
			27389: out = 16'(1825);
			27390: out = 16'(-2409);
			27391: out = 16'(-3520);
			27392: out = 16'(-2493);
			27393: out = 16'(-1159);
			27394: out = 16'(3);
			27395: out = 16'(-284);
			27396: out = 16'(488);
			27397: out = 16'(415);
			27398: out = 16'(-264);
			27399: out = 16'(-256);
			27400: out = 16'(23);
			27401: out = 16'(535);
			27402: out = 16'(-84);
			27403: out = 16'(-1305);
			27404: out = 16'(-188);
			27405: out = 16'(-796);
			27406: out = 16'(-1007);
			27407: out = 16'(-3758);
			27408: out = 16'(-3278);
			27409: out = 16'(-1506);
			27410: out = 16'(1759);
			27411: out = 16'(2884);
			27412: out = 16'(1963);
			27413: out = 16'(714);
			27414: out = 16'(-10);
			27415: out = 16'(1547);
			27416: out = 16'(364);
			27417: out = 16'(-27);
			27418: out = 16'(626);
			27419: out = 16'(530);
			27420: out = 16'(133);
			27421: out = 16'(-2413);
			27422: out = 16'(-1579);
			27423: out = 16'(101);
			27424: out = 16'(1612);
			27425: out = 16'(2409);
			27426: out = 16'(2582);
			27427: out = 16'(2061);
			27428: out = 16'(1858);
			27429: out = 16'(1779);
			27430: out = 16'(343);
			27431: out = 16'(-1861);
			27432: out = 16'(-5052);
			27433: out = 16'(-4692);
			27434: out = 16'(-3233);
			27435: out = 16'(-486);
			27436: out = 16'(1299);
			27437: out = 16'(1858);
			27438: out = 16'(157);
			27439: out = 16'(-1318);
			27440: out = 16'(-2513);
			27441: out = 16'(-1098);
			27442: out = 16'(-440);
			27443: out = 16'(90);
			27444: out = 16'(722);
			27445: out = 16'(133);
			27446: out = 16'(-983);
			27447: out = 16'(-2773);
			27448: out = 16'(-2232);
			27449: out = 16'(900);
			27450: out = 16'(1993);
			27451: out = 16'(3286);
			27452: out = 16'(3183);
			27453: out = 16'(3941);
			27454: out = 16'(3675);
			27455: out = 16'(3388);
			27456: out = 16'(1498);
			27457: out = 16'(-163);
			27458: out = 16'(-1047);
			27459: out = 16'(-878);
			27460: out = 16'(-57);
			27461: out = 16'(-1233);
			27462: out = 16'(-623);
			27463: out = 16'(-141);
			27464: out = 16'(2203);
			27465: out = 16'(1837);
			27466: out = 16'(148);
			27467: out = 16'(-107);
			27468: out = 16'(51);
			27469: out = 16'(1194);
			27470: out = 16'(679);
			27471: out = 16'(162);
			27472: out = 16'(-165);
			27473: out = 16'(-1770);
			27474: out = 16'(-2845);
			27475: out = 16'(-2659);
			27476: out = 16'(-1393);
			27477: out = 16'(268);
			27478: out = 16'(977);
			27479: out = 16'(1417);
			27480: out = 16'(909);
			27481: out = 16'(-1198);
			27482: out = 16'(-2929);
			27483: out = 16'(-4019);
			27484: out = 16'(-475);
			27485: out = 16'(1439);
			27486: out = 16'(1816);
			27487: out = 16'(758);
			27488: out = 16'(-853);
			27489: out = 16'(-1452);
			27490: out = 16'(-4047);
			27491: out = 16'(-4317);
			27492: out = 16'(-1819);
			27493: out = 16'(931);
			27494: out = 16'(3497);
			27495: out = 16'(4883);
			27496: out = 16'(5028);
			27497: out = 16'(3882);
			27498: out = 16'(-293);
			27499: out = 16'(-2612);
			27500: out = 16'(-4296);
			27501: out = 16'(-2085);
			27502: out = 16'(-2244);
			27503: out = 16'(-3256);
			27504: out = 16'(-3322);
			27505: out = 16'(-1829);
			27506: out = 16'(1707);
			27507: out = 16'(1450);
			27508: out = 16'(1393);
			27509: out = 16'(769);
			27510: out = 16'(744);
			27511: out = 16'(707);
			27512: out = 16'(-103);
			27513: out = 16'(1197);
			27514: out = 16'(1985);
			27515: out = 16'(712);
			27516: out = 16'(-955);
			27517: out = 16'(-2621);
			27518: out = 16'(-1800);
			27519: out = 16'(-868);
			27520: out = 16'(739);
			27521: out = 16'(400);
			27522: out = 16'(873);
			27523: out = 16'(1450);
			27524: out = 16'(752);
			27525: out = 16'(140);
			27526: out = 16'(-1092);
			27527: out = 16'(1088);
			27528: out = 16'(2199);
			27529: out = 16'(2021);
			27530: out = 16'(316);
			27531: out = 16'(-1434);
			27532: out = 16'(-1632);
			27533: out = 16'(-870);
			27534: out = 16'(876);
			27535: out = 16'(955);
			27536: out = 16'(2112);
			27537: out = 16'(2479);
			27538: out = 16'(2750);
			27539: out = 16'(1680);
			27540: out = 16'(371);
			27541: out = 16'(-2474);
			27542: out = 16'(-4088);
			27543: out = 16'(-4961);
			27544: out = 16'(-3337);
			27545: out = 16'(-2102);
			27546: out = 16'(-1790);
			27547: out = 16'(-730);
			27548: out = 16'(39);
			27549: out = 16'(-27);
			27550: out = 16'(527);
			27551: out = 16'(1000);
			27552: out = 16'(3383);
			27553: out = 16'(2115);
			27554: out = 16'(462);
			27555: out = 16'(0);
			27556: out = 16'(937);
			27557: out = 16'(2721);
			27558: out = 16'(-280);
			27559: out = 16'(-2619);
			27560: out = 16'(-5852);
			27561: out = 16'(-2718);
			27562: out = 16'(-790);
			27563: out = 16'(791);
			27564: out = 16'(1278);
			27565: out = 16'(1248);
			27566: out = 16'(-196);
			27567: out = 16'(368);
			27568: out = 16'(1309);
			27569: out = 16'(4480);
			27570: out = 16'(3663);
			27571: out = 16'(2101);
			27572: out = 16'(297);
			27573: out = 16'(-1090);
			27574: out = 16'(-1841);
			27575: out = 16'(-1348);
			27576: out = 16'(44);
			27577: out = 16'(2129);
			27578: out = 16'(177);
			27579: out = 16'(6);
			27580: out = 16'(553);
			27581: out = 16'(1509);
			27582: out = 16'(1537);
			27583: out = 16'(-619);
			27584: out = 16'(-119);
			27585: out = 16'(-323);
			27586: out = 16'(757);
			27587: out = 16'(-1820);
			27588: out = 16'(-3459);
			27589: out = 16'(-1970);
			27590: out = 16'(-654);
			27591: out = 16'(860);
			27592: out = 16'(436);
			27593: out = 16'(1452);
			27594: out = 16'(2611);
			27595: out = 16'(166);
			27596: out = 16'(-1618);
			27597: out = 16'(-4495);
			27598: out = 16'(-435);
			27599: out = 16'(-122);
			27600: out = 16'(-1693);
			27601: out = 16'(-4468);
			27602: out = 16'(-4603);
			27603: out = 16'(692);
			27604: out = 16'(1512);
			27605: out = 16'(2121);
			27606: out = 16'(-17);
			27607: out = 16'(451);
			27608: out = 16'(390);
			27609: out = 16'(-770);
			27610: out = 16'(-639);
			27611: out = 16'(159);
			27612: out = 16'(3431);
			27613: out = 16'(3739);
			27614: out = 16'(2316);
			27615: out = 16'(11);
			27616: out = 16'(-2129);
			27617: out = 16'(-3139);
			27618: out = 16'(-2450);
			27619: out = 16'(-662);
			27620: out = 16'(1244);
			27621: out = 16'(3247);
			27622: out = 16'(3399);
			27623: out = 16'(-131);
			27624: out = 16'(292);
			27625: out = 16'(916);
			27626: out = 16'(3105);
			27627: out = 16'(2269);
			27628: out = 16'(849);
			27629: out = 16'(557);
			27630: out = 16'(-580);
			27631: out = 16'(-1189);
			27632: out = 16'(-1367);
			27633: out = 16'(-524);
			27634: out = 16'(465);
			27635: out = 16'(1079);
			27636: out = 16'(497);
			27637: out = 16'(-1177);
			27638: out = 16'(-2147);
			27639: out = 16'(-2355);
			27640: out = 16'(-992);
			27641: out = 16'(-1071);
			27642: out = 16'(-1081);
			27643: out = 16'(-1744);
			27644: out = 16'(-508);
			27645: out = 16'(1178);
			27646: out = 16'(2109);
			27647: out = 16'(3411);
			27648: out = 16'(3472);
			27649: out = 16'(4641);
			27650: out = 16'(1071);
			27651: out = 16'(-3838);
			27652: out = 16'(-5229);
			27653: out = 16'(-4122);
			27654: out = 16'(327);
			27655: out = 16'(128);
			27656: out = 16'(630);
			27657: out = 16'(-526);
			27658: out = 16'(-629);
			27659: out = 16'(-942);
			27660: out = 16'(843);
			27661: out = 16'(-13);
			27662: out = 16'(-283);
			27663: out = 16'(-3335);
			27664: out = 16'(-1203);
			27665: out = 16'(678);
			27666: out = 16'(1357);
			27667: out = 16'(26);
			27668: out = 16'(-1811);
			27669: out = 16'(-1090);
			27670: out = 16'(335);
			27671: out = 16'(2858);
			27672: out = 16'(1467);
			27673: out = 16'(1078);
			27674: out = 16'(278);
			27675: out = 16'(-491);
			27676: out = 16'(-1498);
			27677: out = 16'(-2344);
			27678: out = 16'(-1225);
			27679: out = 16'(481);
			27680: out = 16'(1698);
			27681: out = 16'(2506);
			27682: out = 16'(2327);
			27683: out = 16'(2081);
			27684: out = 16'(1326);
			27685: out = 16'(1184);
			27686: out = 16'(-448);
			27687: out = 16'(92);
			27688: out = 16'(449);
			27689: out = 16'(4246);
			27690: out = 16'(3637);
			27691: out = 16'(1515);
			27692: out = 16'(-2309);
			27693: out = 16'(-3168);
			27694: out = 16'(-1154);
			27695: out = 16'(773);
			27696: out = 16'(1321);
			27697: out = 16'(-1271);
			27698: out = 16'(-2097);
			27699: out = 16'(-2354);
			27700: out = 16'(135);
			27701: out = 16'(421);
			27702: out = 16'(614);
			27703: out = 16'(3617);
			27704: out = 16'(1703);
			27705: out = 16'(-736);
			27706: out = 16'(-5089);
			27707: out = 16'(-3835);
			27708: out = 16'(263);
			27709: out = 16'(1330);
			27710: out = 16'(766);
			27711: out = 16'(-2934);
			27712: out = 16'(-2877);
			27713: out = 16'(-2956);
			27714: out = 16'(-743);
			27715: out = 16'(-1173);
			27716: out = 16'(-422);
			27717: out = 16'(1266);
			27718: out = 16'(909);
			27719: out = 16'(-62);
			27720: out = 16'(-3025);
			27721: out = 16'(-1497);
			27722: out = 16'(1183);
			27723: out = 16'(3246);
			27724: out = 16'(4374);
			27725: out = 16'(3925);
			27726: out = 16'(766);
			27727: out = 16'(-2463);
			27728: out = 16'(-5472);
			27729: out = 16'(-1162);
			27730: out = 16'(2098);
			27731: out = 16'(4819);
			27732: out = 16'(4209);
			27733: out = 16'(2513);
			27734: out = 16'(-1165);
			27735: out = 16'(-359);
			27736: out = 16'(564);
			27737: out = 16'(1646);
			27738: out = 16'(998);
			27739: out = 16'(-134);
			27740: out = 16'(-326);
			27741: out = 16'(-401);
			27742: out = 16'(415);
			27743: out = 16'(-547);
			27744: out = 16'(886);
			27745: out = 16'(2211);
			27746: out = 16'(2044);
			27747: out = 16'(-106);
			27748: out = 16'(-3566);
			27749: out = 16'(-4631);
			27750: out = 16'(-4085);
			27751: out = 16'(-992);
			27752: out = 16'(-638);
			27753: out = 16'(-510);
			27754: out = 16'(-1718);
			27755: out = 16'(-1771);
			27756: out = 16'(-1306);
			27757: out = 16'(369);
			27758: out = 16'(2031);
			27759: out = 16'(2994);
			27760: out = 16'(326);
			27761: out = 16'(-1497);
			27762: out = 16'(-3223);
			27763: out = 16'(-824);
			27764: out = 16'(647);
			27765: out = 16'(1949);
			27766: out = 16'(1523);
			27767: out = 16'(342);
			27768: out = 16'(-1770);
			27769: out = 16'(-3243);
			27770: out = 16'(-3892);
			27771: out = 16'(-3026);
			27772: out = 16'(-1420);
			27773: out = 16'(859);
			27774: out = 16'(3585);
			27775: out = 16'(4658);
			27776: out = 16'(4262);
			27777: out = 16'(-1150);
			27778: out = 16'(-2510);
			27779: out = 16'(-2897);
			27780: out = 16'(2999);
			27781: out = 16'(3215);
			27782: out = 16'(1631);
			27783: out = 16'(-417);
			27784: out = 16'(-791);
			27785: out = 16'(741);
			27786: out = 16'(-101);
			27787: out = 16'(-136);
			27788: out = 16'(-177);
			27789: out = 16'(269);
			27790: out = 16'(395);
			27791: out = 16'(-1196);
			27792: out = 16'(-355);
			27793: out = 16'(-232);
			27794: out = 16'(841);
			27795: out = 16'(-1841);
			27796: out = 16'(-3939);
			27797: out = 16'(-2142);
			27798: out = 16'(777);
			27799: out = 16'(4131);
			27800: out = 16'(4222);
			27801: out = 16'(3240);
			27802: out = 16'(865);
			27803: out = 16'(-1615);
			27804: out = 16'(-2274);
			27805: out = 16'(100);
			27806: out = 16'(485);
			27807: out = 16'(1295);
			27808: out = 16'(137);
			27809: out = 16'(1073);
			27810: out = 16'(296);
			27811: out = 16'(-3155);
			27812: out = 16'(-3185);
			27813: out = 16'(-1911);
			27814: out = 16'(1308);
			27815: out = 16'(2057);
			27816: out = 16'(1497);
			27817: out = 16'(841);
			27818: out = 16'(-123);
			27819: out = 16'(-169);
			27820: out = 16'(-4288);
			27821: out = 16'(-3420);
			27822: out = 16'(618);
			27823: out = 16'(951);
			27824: out = 16'(30);
			27825: out = 16'(-5233);
			27826: out = 16'(-1641);
			27827: out = 16'(216);
			27828: out = 16'(1312);
			27829: out = 16'(882);
			27830: out = 16'(598);
			27831: out = 16'(580);
			27832: out = 16'(556);
			27833: out = 16'(388);
			27834: out = 16'(1906);
			27835: out = 16'(934);
			27836: out = 16'(-473);
			27837: out = 16'(-4117);
			27838: out = 16'(-3765);
			27839: out = 16'(-421);
			27840: out = 16'(453);
			27841: out = 16'(1975);
			27842: out = 16'(1582);
			27843: out = 16'(3178);
			27844: out = 16'(2643);
			27845: out = 16'(2828);
			27846: out = 16'(-621);
			27847: out = 16'(-2072);
			27848: out = 16'(-3694);
			27849: out = 16'(548);
			27850: out = 16'(3264);
			27851: out = 16'(3313);
			27852: out = 16'(-497);
			27853: out = 16'(-4517);
			27854: out = 16'(-3503);
			27855: out = 16'(-674);
			27856: out = 16'(3596);
			27857: out = 16'(3506);
			27858: out = 16'(2438);
			27859: out = 16'(-881);
			27860: out = 16'(-3017);
			27861: out = 16'(-4471);
			27862: out = 16'(-3856);
			27863: out = 16'(-2119);
			27864: out = 16'(-599);
			27865: out = 16'(-1120);
			27866: out = 16'(-1193);
			27867: out = 16'(-1539);
			27868: out = 16'(142);
			27869: out = 16'(298);
			27870: out = 16'(877);
			27871: out = 16'(-96);
			27872: out = 16'(1028);
			27873: out = 16'(2061);
			27874: out = 16'(656);
			27875: out = 16'(161);
			27876: out = 16'(-329);
			27877: out = 16'(424);
			27878: out = 16'(-233);
			27879: out = 16'(-1751);
			27880: out = 16'(-652);
			27881: out = 16'(153);
			27882: out = 16'(607);
			27883: out = 16'(1185);
			27884: out = 16'(1256);
			27885: out = 16'(1423);
			27886: out = 16'(-74);
			27887: out = 16'(-1269);
			27888: out = 16'(-2408);
			27889: out = 16'(-1221);
			27890: out = 16'(454);
			27891: out = 16'(2890);
			27892: out = 16'(2538);
			27893: out = 16'(946);
			27894: out = 16'(73);
			27895: out = 16'(-303);
			27896: out = 16'(598);
			27897: out = 16'(1317);
			27898: out = 16'(2590);
			27899: out = 16'(3548);
			27900: out = 16'(2035);
			27901: out = 16'(67);
			27902: out = 16'(-1718);
			27903: out = 16'(-3042);
			27904: out = 16'(-3079);
			27905: out = 16'(-2013);
			27906: out = 16'(-402);
			27907: out = 16'(806);
			27908: out = 16'(1823);
			27909: out = 16'(937);
			27910: out = 16'(-390);
			27911: out = 16'(-876);
			27912: out = 16'(-876);
			27913: out = 16'(-187);
			27914: out = 16'(344);
			27915: out = 16'(647);
			27916: out = 16'(478);
			27917: out = 16'(542);
			27918: out = 16'(657);
			27919: out = 16'(1209);
			27920: out = 16'(-241);
			27921: out = 16'(-2006);
			27922: out = 16'(-4714);
			27923: out = 16'(-3545);
			27924: out = 16'(-1650);
			27925: out = 16'(-420);
			27926: out = 16'(1951);
			27927: out = 16'(3180);
			27928: out = 16'(2245);
			27929: out = 16'(-10);
			27930: out = 16'(-2638);
			27931: out = 16'(-490);
			27932: out = 16'(83);
			27933: out = 16'(712);
			27934: out = 16'(463);
			27935: out = 16'(281);
			27936: out = 16'(-50);
			27937: out = 16'(-132);
			27938: out = 16'(259);
			27939: out = 16'(1240);
			27940: out = 16'(2090);
			27941: out = 16'(2257);
			27942: out = 16'(467);
			27943: out = 16'(477);
			27944: out = 16'(-43);
			27945: out = 16'(-1627);
			27946: out = 16'(-2556);
			27947: out = 16'(-3165);
			27948: out = 16'(-576);
			27949: out = 16'(-30);
			27950: out = 16'(563);
			27951: out = 16'(-409);
			27952: out = 16'(1001);
			27953: out = 16'(3257);
			27954: out = 16'(4059);
			27955: out = 16'(3474);
			27956: out = 16'(894);
			27957: out = 16'(610);
			27958: out = 16'(-498);
			27959: out = 16'(-2665);
			27960: out = 16'(-2197);
			27961: out = 16'(-1686);
			27962: out = 16'(-339);
			27963: out = 16'(-1601);
			27964: out = 16'(-2300);
			27965: out = 16'(-9);
			27966: out = 16'(1708);
			27967: out = 16'(3254);
			27968: out = 16'(3600);
			27969: out = 16'(2683);
			27970: out = 16'(728);
			27971: out = 16'(-1697);
			27972: out = 16'(-3409);
			27973: out = 16'(-4008);
			27974: out = 16'(-3124);
			27975: out = 16'(-1670);
			27976: out = 16'(372);
			27977: out = 16'(931);
			27978: out = 16'(1298);
			27979: out = 16'(364);
			27980: out = 16'(1769);
			27981: out = 16'(2664);
			27982: out = 16'(4859);
			27983: out = 16'(2169);
			27984: out = 16'(-847);
			27985: out = 16'(-2350);
			27986: out = 16'(-1961);
			27987: out = 16'(-241);
			27988: out = 16'(-20);
			27989: out = 16'(140);
			27990: out = 16'(-322);
			27991: out = 16'(-1516);
			27992: out = 16'(-1411);
			27993: out = 16'(352);
			27994: out = 16'(2877);
			27995: out = 16'(4197);
			27996: out = 16'(1965);
			27997: out = 16'(1268);
			27998: out = 16'(-654);
			27999: out = 16'(-82);
			28000: out = 16'(-3345);
			28001: out = 16'(-5116);
			28002: out = 16'(-5887);
			28003: out = 16'(-3040);
			28004: out = 16'(334);
			28005: out = 16'(950);
			28006: out = 16'(1045);
			28007: out = 16'(281);
			28008: out = 16'(474);
			28009: out = 16'(1322);
			28010: out = 16'(3150);
			28011: out = 16'(2617);
			28012: out = 16'(1461);
			28013: out = 16'(-1272);
			28014: out = 16'(-2593);
			28015: out = 16'(-3455);
			28016: out = 16'(-2438);
			28017: out = 16'(-2202);
			28018: out = 16'(-1580);
			28019: out = 16'(-1854);
			28020: out = 16'(-1255);
			28021: out = 16'(-757);
			28022: out = 16'(485);
			28023: out = 16'(1492);
			28024: out = 16'(2677);
			28025: out = 16'(231);
			28026: out = 16'(-370);
			28027: out = 16'(-1094);
			28028: out = 16'(372);
			28029: out = 16'(721);
			28030: out = 16'(1409);
			28031: out = 16'(-1433);
			28032: out = 16'(-2586);
			28033: out = 16'(-2429);
			28034: out = 16'(-466);
			28035: out = 16'(999);
			28036: out = 16'(1271);
			28037: out = 16'(885);
			28038: out = 16'(368);
			28039: out = 16'(-131);
			28040: out = 16'(1749);
			28041: out = 16'(3814);
			28042: out = 16'(286);
			28043: out = 16'(-1611);
			28044: out = 16'(-4240);
			28045: out = 16'(-41);
			28046: out = 16'(854);
			28047: out = 16'(1363);
			28048: out = 16'(512);
			28049: out = 16'(653);
			28050: out = 16'(1168);
			28051: out = 16'(2470);
			28052: out = 16'(3466);
			28053: out = 16'(4722);
			28054: out = 16'(3288);
			28055: out = 16'(1382);
			28056: out = 16'(-2542);
			28057: out = 16'(-2119);
			28058: out = 16'(-1404);
			28059: out = 16'(-3956);
			28060: out = 16'(-4831);
			28061: out = 16'(-5429);
			28062: out = 16'(-1124);
			28063: out = 16'(290);
			28064: out = 16'(621);
			28065: out = 16'(1697);
			28066: out = 16'(1946);
			28067: out = 16'(1868);
			28068: out = 16'(403);
			28069: out = 16'(-58);
			28070: out = 16'(1297);
			28071: out = 16'(178);
			28072: out = 16'(-1215);
			28073: out = 16'(-4771);
			28074: out = 16'(-4386);
			28075: out = 16'(-3364);
			28076: out = 16'(246);
			28077: out = 16'(365);
			28078: out = 16'(-18);
			28079: out = 16'(-821);
			28080: out = 16'(33);
			28081: out = 16'(1531);
			28082: out = 16'(163);
			28083: out = 16'(-227);
			28084: out = 16'(-967);
			28085: out = 16'(907);
			28086: out = 16'(1434);
			28087: out = 16'(1328);
			28088: out = 16'(308);
			28089: out = 16'(-243);
			28090: out = 16'(822);
			28091: out = 16'(31);
			28092: out = 16'(418);
			28093: out = 16'(2317);
			28094: out = 16'(3617);
			28095: out = 16'(3937);
			28096: out = 16'(857);
			28097: out = 16'(-1325);
			28098: out = 16'(-3584);
			28099: out = 16'(-1250);
			28100: out = 16'(-702);
			28101: out = 16'(494);
			28102: out = 16'(-3447);
			28103: out = 16'(-2920);
			28104: out = 16'(-59);
			28105: out = 16'(1750);
			28106: out = 16'(2543);
			28107: out = 16'(1018);
			28108: out = 16'(1377);
			28109: out = 16'(1010);
			28110: out = 16'(1368);
			28111: out = 16'(-257);
			28112: out = 16'(-1148);
			28113: out = 16'(-437);
			28114: out = 16'(67);
			28115: out = 16'(482);
			28116: out = 16'(-982);
			28117: out = 16'(-815);
			28118: out = 16'(-317);
			28119: out = 16'(-395);
			28120: out = 16'(-345);
			28121: out = 16'(-343);
			28122: out = 16'(-173);
			28123: out = 16'(61);
			28124: out = 16'(603);
			28125: out = 16'(1418);
			28126: out = 16'(1849);
			28127: out = 16'(1001);
			28128: out = 16'(491);
			28129: out = 16'(-613);
			28130: out = 16'(-22);
			28131: out = 16'(-3103);
			28132: out = 16'(-4959);
			28133: out = 16'(-4947);
			28134: out = 16'(-2149);
			28135: out = 16'(1252);
			28136: out = 16'(1710);
			28137: out = 16'(1646);
			28138: out = 16'(156);
			28139: out = 16'(100);
			28140: out = 16'(-850);
			28141: out = 16'(-1609);
			28142: out = 16'(-147);
			28143: out = 16'(759);
			28144: out = 16'(568);
			28145: out = 16'(242);
			28146: out = 16'(-688);
			28147: out = 16'(-1499);
			28148: out = 16'(-992);
			28149: out = 16'(467);
			28150: out = 16'(1649);
			28151: out = 16'(2918);
			28152: out = 16'(3034);
			28153: out = 16'(3447);
			28154: out = 16'(1454);
			28155: out = 16'(-497);
			28156: out = 16'(-4909);
			28157: out = 16'(-4094);
			28158: out = 16'(-503);
			28159: out = 16'(1183);
			28160: out = 16'(1898);
			28161: out = 16'(342);
			28162: out = 16'(2132);
			28163: out = 16'(2658);
			28164: out = 16'(3084);
			28165: out = 16'(2631);
			28166: out = 16'(2115);
			28167: out = 16'(1792);
			28168: out = 16'(0);
			28169: out = 16'(-1695);
			28170: out = 16'(-2563);
			28171: out = 16'(-2076);
			28172: out = 16'(-1145);
			28173: out = 16'(-3889);
			28174: out = 16'(-3123);
			28175: out = 16'(-1337);
			28176: out = 16'(624);
			28177: out = 16'(1634);
			28178: out = 16'(1006);
			28179: out = 16'(2541);
			28180: out = 16'(1731);
			28181: out = 16'(750);
			28182: out = 16'(-3314);
			28183: out = 16'(-4244);
			28184: out = 16'(-989);
			28185: out = 16'(1568);
			28186: out = 16'(3093);
			28187: out = 16'(-152);
			28188: out = 16'(-762);
			28189: out = 16'(-1970);
			28190: out = 16'(-779);
			28191: out = 16'(-1454);
			28192: out = 16'(-1392);
			28193: out = 16'(-41);
			28194: out = 16'(1718);
			28195: out = 16'(3157);
			28196: out = 16'(61);
			28197: out = 16'(-2359);
			28198: out = 16'(-4676);
			28199: out = 16'(-2574);
			28200: out = 16'(-680);
			28201: out = 16'(637);
			28202: out = 16'(2075);
			28203: out = 16'(3064);
			28204: out = 16'(4426);
			28205: out = 16'(3672);
			28206: out = 16'(2546);
			28207: out = 16'(-905);
			28208: out = 16'(-482);
			28209: out = 16'(488);
			28210: out = 16'(1666);
			28211: out = 16'(937);
			28212: out = 16'(-709);
			28213: out = 16'(-1537);
			28214: out = 16'(-1540);
			28215: out = 16'(-166);
			28216: out = 16'(-71);
			28217: out = 16'(738);
			28218: out = 16'(1018);
			28219: out = 16'(2140);
			28220: out = 16'(1843);
			28221: out = 16'(-281);
			28222: out = 16'(-365);
			28223: out = 16'(-613);
			28224: out = 16'(-1141);
			28225: out = 16'(-829);
			28226: out = 16'(-317);
			28227: out = 16'(-277);
			28228: out = 16'(-216);
			28229: out = 16'(-513);
			28230: out = 16'(-77);
			28231: out = 16'(-626);
			28232: out = 16'(-1089);
			28233: out = 16'(-3523);
			28234: out = 16'(-3051);
			28235: out = 16'(28);
			28236: out = 16'(-271);
			28237: out = 16'(257);
			28238: out = 16'(299);
			28239: out = 16'(601);
			28240: out = 16'(-84);
			28241: out = 16'(-1486);
			28242: out = 16'(-2641);
			28243: out = 16'(-2498);
			28244: out = 16'(1678);
			28245: out = 16'(3003);
			28246: out = 16'(3655);
			28247: out = 16'(86);
			28248: out = 16'(-375);
			28249: out = 16'(-306);
			28250: out = 16'(365);
			28251: out = 16'(-726);
			28252: out = 16'(-3412);
			28253: out = 16'(-150);
			28254: out = 16'(1217);
			28255: out = 16'(2687);
			28256: out = 16'(-399);
			28257: out = 16'(-2200);
			28258: out = 16'(-2337);
			28259: out = 16'(-1724);
			28260: out = 16'(-290);
			28261: out = 16'(1709);
			28262: out = 16'(2716);
			28263: out = 16'(3006);
			28264: out = 16'(1354);
			28265: out = 16'(583);
			28266: out = 16'(-546);
			28267: out = 16'(-1939);
			28268: out = 16'(-3891);
			28269: out = 16'(-5430);
			28270: out = 16'(-3849);
			28271: out = 16'(-1441);
			28272: out = 16'(1545);
			28273: out = 16'(3713);
			28274: out = 16'(4253);
			28275: out = 16'(2408);
			28276: out = 16'(1803);
			28277: out = 16'(1175);
			28278: out = 16'(2645);
			28279: out = 16'(1060);
			28280: out = 16'(-37);
			28281: out = 16'(-1106);
			28282: out = 16'(-863);
			28283: out = 16'(-367);
			28284: out = 16'(-503);
			28285: out = 16'(-279);
			28286: out = 16'(-103);
			28287: out = 16'(1395);
			28288: out = 16'(2700);
			28289: out = 16'(4271);
			28290: out = 16'(1674);
			28291: out = 16'(99);
			28292: out = 16'(-2229);
			28293: out = 16'(-673);
			28294: out = 16'(-454);
			28295: out = 16'(-141);
			28296: out = 16'(-2392);
			28297: out = 16'(-3581);
			28298: out = 16'(-4267);
			28299: out = 16'(-1494);
			28300: out = 16'(1104);
			28301: out = 16'(2293);
			28302: out = 16'(1930);
			28303: out = 16'(922);
			28304: out = 16'(-863);
			28305: out = 16'(-862);
			28306: out = 16'(-503);
			28307: out = 16'(-133);
			28308: out = 16'(-2188);
			28309: out = 16'(-5651);
			28310: out = 16'(-6247);
			28311: out = 16'(-4627);
			28312: out = 16'(74);
			28313: out = 16'(2225);
			28314: out = 16'(3767);
			28315: out = 16'(3867);
			28316: out = 16'(2004);
			28317: out = 16'(541);
			28318: out = 16'(1917);
			28319: out = 16'(3677);
			28320: out = 16'(5225);
			28321: out = 16'(72);
			28322: out = 16'(-1834);
			28323: out = 16'(-4514);
			28324: out = 16'(-476);
			28325: out = 16'(-1405);
			28326: out = 16'(-2359);
			28327: out = 16'(-3406);
			28328: out = 16'(-1433);
			28329: out = 16'(2093);
			28330: out = 16'(2953);
			28331: out = 16'(2695);
			28332: out = 16'(1281);
			28333: out = 16'(-769);
			28334: out = 16'(-1835);
			28335: out = 16'(-1080);
			28336: out = 16'(303);
			28337: out = 16'(1205);
			28338: out = 16'(-175);
			28339: out = 16'(-2131);
			28340: out = 16'(-4130);
			28341: out = 16'(-1801);
			28342: out = 16'(-976);
			28343: out = 16'(263);
			28344: out = 16'(494);
			28345: out = 16'(586);
			28346: out = 16'(-367);
			28347: out = 16'(466);
			28348: out = 16'(480);
			28349: out = 16'(797);
			28350: out = 16'(-915);
			28351: out = 16'(-2451);
			28352: out = 16'(-5457);
			28353: out = 16'(-2533);
			28354: out = 16'(-15);
			28355: out = 16'(1367);
			28356: out = 16'(928);
			28357: out = 16'(242);
			28358: out = 16'(2741);
			28359: out = 16'(3185);
			28360: out = 16'(3971);
			28361: out = 16'(51);
			28362: out = 16'(275);
			28363: out = 16'(622);
			28364: out = 16'(3965);
			28365: out = 16'(3133);
			28366: out = 16'(377);
			28367: out = 16'(-3837);
			28368: out = 16'(-5558);
			28369: out = 16'(-3614);
			28370: out = 16'(-1110);
			28371: out = 16'(1962);
			28372: out = 16'(3483);
			28373: out = 16'(4528);
			28374: out = 16'(3728);
			28375: out = 16'(1601);
			28376: out = 16'(-460);
			28377: out = 16'(-2117);
			28378: out = 16'(-2994);
			28379: out = 16'(-3633);
			28380: out = 16'(-3736);
			28381: out = 16'(-1460);
			28382: out = 16'(118);
			28383: out = 16'(1486);
			28384: out = 16'(333);
			28385: out = 16'(-57);
			28386: out = 16'(-106);
			28387: out = 16'(388);
			28388: out = 16'(1233);
			28389: out = 16'(2580);
			28390: out = 16'(2259);
			28391: out = 16'(1694);
			28392: out = 16'(1343);
			28393: out = 16'(772);
			28394: out = 16'(360);
			28395: out = 16'(-1007);
			28396: out = 16'(-1029);
			28397: out = 16'(-1038);
			28398: out = 16'(279);
			28399: out = 16'(2);
			28400: out = 16'(-300);
			28401: out = 16'(-1641);
			28402: out = 16'(-909);
			28403: out = 16'(652);
			28404: out = 16'(1671);
			28405: out = 16'(1347);
			28406: out = 16'(-321);
			28407: out = 16'(-2761);
			28408: out = 16'(-4059);
			28409: out = 16'(-3044);
			28410: out = 16'(-1473);
			28411: out = 16'(207);
			28412: out = 16'(-306);
			28413: out = 16'(-644);
			28414: out = 16'(-1642);
			28415: out = 16'(882);
			28416: out = 16'(321);
			28417: out = 16'(80);
			28418: out = 16'(-4058);
			28419: out = 16'(-3228);
			28420: out = 16'(-385);
			28421: out = 16'(333);
			28422: out = 16'(497);
			28423: out = 16'(-806);
			28424: out = 16'(556);
			28425: out = 16'(1334);
			28426: out = 16'(2806);
			28427: out = 16'(1876);
			28428: out = 16'(1153);
			28429: out = 16'(133);
			28430: out = 16'(752);
			28431: out = 16'(1808);
			28432: out = 16'(3467);
			28433: out = 16'(4101);
			28434: out = 16'(3790);
			28435: out = 16'(485);
			28436: out = 16'(-1017);
			28437: out = 16'(-1649);
			28438: out = 16'(-565);
			28439: out = 16'(676);
			28440: out = 16'(1730);
			28441: out = 16'(1925);
			28442: out = 16'(578);
			28443: out = 16'(-2598);
			28444: out = 16'(-2978);
			28445: out = 16'(-2546);
			28446: out = 16'(702);
			28447: out = 16'(305);
			28448: out = 16'(538);
			28449: out = 16'(312);
			28450: out = 16'(2273);
			28451: out = 16'(3375);
			28452: out = 16'(-109);
			28453: out = 16'(-1078);
			28454: out = 16'(-1760);
			28455: out = 16'(832);
			28456: out = 16'(861);
			28457: out = 16'(182);
			28458: out = 16'(258);
			28459: out = 16'(219);
			28460: out = 16'(234);
			28461: out = 16'(-752);
			28462: out = 16'(-725);
			28463: out = 16'(1292);
			28464: out = 16'(112);
			28465: out = 16'(-848);
			28466: out = 16'(-4907);
			28467: out = 16'(-1553);
			28468: out = 16'(1104);
			28469: out = 16'(2943);
			28470: out = 16'(1049);
			28471: out = 16'(-1376);
			28472: out = 16'(-1005);
			28473: out = 16'(304);
			28474: out = 16'(2613);
			28475: out = 16'(696);
			28476: out = 16'(-900);
			28477: out = 16'(-4342);
			28478: out = 16'(-2470);
			28479: out = 16'(-2047);
			28480: out = 16'(168);
			28481: out = 16'(-2536);
			28482: out = 16'(-2379);
			28483: out = 16'(-1116);
			28484: out = 16'(1601);
			28485: out = 16'(2254);
			28486: out = 16'(838);
			28487: out = 16'(-2391);
			28488: out = 16'(-4355);
			28489: out = 16'(-1855);
			28490: out = 16'(890);
			28491: out = 16'(3378);
			28492: out = 16'(1707);
			28493: out = 16'(-352);
			28494: out = 16'(-3154);
			28495: out = 16'(-3595);
			28496: out = 16'(-1858);
			28497: out = 16'(2512);
			28498: out = 16'(2804);
			28499: out = 16'(2878);
			28500: out = 16'(423);
			28501: out = 16'(911);
			28502: out = 16'(388);
			28503: out = 16'(141);
			28504: out = 16'(176);
			28505: out = 16'(437);
			28506: out = 16'(-1001);
			28507: out = 16'(10);
			28508: out = 16'(810);
			28509: out = 16'(1837);
			28510: out = 16'(1374);
			28511: out = 16'(485);
			28512: out = 16'(1199);
			28513: out = 16'(948);
			28514: out = 16'(507);
			28515: out = 16'(410);
			28516: out = 16'(110);
			28517: out = 16'(-401);
			28518: out = 16'(-1250);
			28519: out = 16'(-1850);
			28520: out = 16'(-1538);
			28521: out = 16'(-938);
			28522: out = 16'(181);
			28523: out = 16'(81);
			28524: out = 16'(2175);
			28525: out = 16'(2986);
			28526: out = 16'(3304);
			28527: out = 16'(-46);
			28528: out = 16'(-3539);
			28529: out = 16'(-1797);
			28530: out = 16'(-867);
			28531: out = 16'(792);
			28532: out = 16'(271);
			28533: out = 16'(299);
			28534: out = 16'(-210);
			28535: out = 16'(-41);
			28536: out = 16'(-207);
			28537: out = 16'(-278);
			28538: out = 16'(-170);
			28539: out = 16'(-96);
			28540: out = 16'(-79);
			28541: out = 16'(-254);
			28542: out = 16'(-44);
			28543: out = 16'(1084);
			28544: out = 16'(1860);
			28545: out = 16'(2283);
			28546: out = 16'(436);
			28547: out = 16'(-80);
			28548: out = 16'(-477);
			28549: out = 16'(-355);
			28550: out = 16'(-666);
			28551: out = 16'(-1086);
			28552: out = 16'(-528);
			28553: out = 16'(109);
			28554: out = 16'(1260);
			28555: out = 16'(149);
			28556: out = 16'(-796);
			28557: out = 16'(-3365);
			28558: out = 16'(-1026);
			28559: out = 16'(491);
			28560: out = 16'(3206);
			28561: out = 16'(232);
			28562: out = 16'(-2323);
			28563: out = 16'(-4500);
			28564: out = 16'(-2401);
			28565: out = 16'(731);
			28566: out = 16'(3111);
			28567: out = 16'(3678);
			28568: out = 16'(2673);
			28569: out = 16'(940);
			28570: out = 16'(-416);
			28571: out = 16'(-1055);
			28572: out = 16'(-539);
			28573: out = 16'(-539);
			28574: out = 16'(-1057);
			28575: out = 16'(-2952);
			28576: out = 16'(-4302);
			28577: out = 16'(-5154);
			28578: out = 16'(-2635);
			28579: out = 16'(361);
			28580: out = 16'(2919);
			28581: out = 16'(3137);
			28582: out = 16'(2137);
			28583: out = 16'(993);
			28584: out = 16'(132);
			28585: out = 16'(22);
			28586: out = 16'(-929);
			28587: out = 16'(-584);
			28588: out = 16'(-160);
			28589: out = 16'(2090);
			28590: out = 16'(2167);
			28591: out = 16'(1115);
			28592: out = 16'(-345);
			28593: out = 16'(-976);
			28594: out = 16'(96);
			28595: out = 16'(-321);
			28596: out = 16'(-517);
			28597: out = 16'(-2545);
			28598: out = 16'(266);
			28599: out = 16'(2238);
			28600: out = 16'(2339);
			28601: out = 16'(1527);
			28602: out = 16'(-136);
			28603: out = 16'(-629);
			28604: out = 16'(-1591);
			28605: out = 16'(-1499);
			28606: out = 16'(-1939);
			28607: out = 16'(-581);
			28608: out = 16'(636);
			28609: out = 16'(3127);
			28610: out = 16'(3292);
			28611: out = 16'(2359);
			28612: out = 16'(370);
			28613: out = 16'(-974);
			28614: out = 16'(-2635);
			28615: out = 16'(-828);
			28616: out = 16'(-155);
			28617: out = 16'(644);
			28618: out = 16'(-3462);
			28619: out = 16'(-6100);
			28620: out = 16'(-3267);
			28621: out = 16'(-188);
			28622: out = 16'(3216);
			28623: out = 16'(3999);
			28624: out = 16'(3521);
			28625: out = 16'(1464);
			28626: out = 16'(473);
			28627: out = 16'(-770);
			28628: out = 16'(-1658);
			28629: out = 16'(-566);
			28630: out = 16'(-205);
			28631: out = 16'(109);
			28632: out = 16'(-2690);
			28633: out = 16'(-3048);
			28634: out = 16'(511);
			28635: out = 16'(2463);
			28636: out = 16'(3399);
			28637: out = 16'(-939);
			28638: out = 16'(-489);
			28639: out = 16'(-55);
			28640: out = 16'(1772);
			28641: out = 16'(1079);
			28642: out = 16'(-285);
			28643: out = 16'(1294);
			28644: out = 16'(497);
			28645: out = 16'(-74);
			28646: out = 16'(-4386);
			28647: out = 16'(-4105);
			28648: out = 16'(-588);
			28649: out = 16'(1913);
			28650: out = 16'(3457);
			28651: out = 16'(2890);
			28652: out = 16'(1636);
			28653: out = 16'(-245);
			28654: out = 16'(-2162);
			28655: out = 16'(-2482);
			28656: out = 16'(-1851);
			28657: out = 16'(1057);
			28658: out = 16'(982);
			28659: out = 16'(427);
			28660: out = 16'(-1343);
			28661: out = 16'(-1875);
			28662: out = 16'(-2189);
			28663: out = 16'(1834);
			28664: out = 16'(2729);
			28665: out = 16'(3177);
			28666: out = 16'(-1218);
			28667: out = 16'(-1760);
			28668: out = 16'(429);
			28669: out = 16'(3078);
			28670: out = 16'(3692);
			28671: out = 16'(1189);
			28672: out = 16'(-2664);
			28673: out = 16'(-5619);
			28674: out = 16'(-2898);
			28675: out = 16'(-1376);
			28676: out = 16'(1278);
			28677: out = 16'(20);
			28678: out = 16'(1464);
			28679: out = 16'(1779);
			28680: out = 16'(3655);
			28681: out = 16'(2521);
			28682: out = 16'(1064);
			28683: out = 16'(-31);
			28684: out = 16'(165);
			28685: out = 16'(1033);
			28686: out = 16'(624);
			28687: out = 16'(-725);
			28688: out = 16'(-3148);
			28689: out = 16'(-2843);
			28690: out = 16'(-2055);
			28691: out = 16'(-1949);
			28692: out = 16'(184);
			28693: out = 16'(1438);
			28694: out = 16'(3178);
			28695: out = 16'(636);
			28696: out = 16'(-2030);
			28697: out = 16'(-3078);
			28698: out = 16'(-621);
			28699: out = 16'(3467);
			28700: out = 16'(1355);
			28701: out = 16'(122);
			28702: out = 16'(-2680);
			28703: out = 16'(-1149);
			28704: out = 16'(-696);
			28705: out = 16'(475);
			28706: out = 16'(-30);
			28707: out = 16'(-97);
			28708: out = 16'(-138);
			28709: out = 16'(-600);
			28710: out = 16'(-970);
			28711: out = 16'(-44);
			28712: out = 16'(-143);
			28713: out = 16'(-292);
			28714: out = 16'(-2868);
			28715: out = 16'(-2791);
			28716: out = 16'(-1992);
			28717: out = 16'(167);
			28718: out = 16'(1763);
			28719: out = 16'(3210);
			28720: out = 16'(1623);
			28721: out = 16'(558);
			28722: out = 16'(-1128);
			28723: out = 16'(-144);
			28724: out = 16'(-208);
			28725: out = 16'(116);
			28726: out = 16'(-2147);
			28727: out = 16'(-2887);
			28728: out = 16'(-1664);
			28729: out = 16'(510);
			28730: out = 16'(2092);
			28731: out = 16'(445);
			28732: out = 16'(-113);
			28733: out = 16'(-983);
			28734: out = 16'(703);
			28735: out = 16'(301);
			28736: out = 16'(52);
			28737: out = 16'(320);
			28738: out = 16'(800);
			28739: out = 16'(1291);
			28740: out = 16'(1260);
			28741: out = 16'(1053);
			28742: out = 16'(520);
			28743: out = 16'(1032);
			28744: out = 16'(1051);
			28745: out = 16'(502);
			28746: out = 16'(25);
			28747: out = 16'(-590);
			28748: out = 16'(-949);
			28749: out = 16'(-1120);
			28750: out = 16'(-843);
			28751: out = 16'(-488);
			28752: out = 16'(485);
			28753: out = 16'(1353);
			28754: out = 16'(2254);
			28755: out = 16'(1938);
			28756: out = 16'(952);
			28757: out = 16'(1145);
			28758: out = 16'(1159);
			28759: out = 16'(1759);
			28760: out = 16'(560);
			28761: out = 16'(500);
			28762: out = 16'(924);
			28763: out = 16'(1010);
			28764: out = 16'(489);
			28765: out = 16'(-1222);
			28766: out = 16'(-1304);
			28767: out = 16'(-1062);
			28768: out = 16'(-387);
			28769: out = 16'(-259);
			28770: out = 16'(-390);
			28771: out = 16'(-339);
			28772: out = 16'(-1468);
			28773: out = 16'(-2563);
			28774: out = 16'(-696);
			28775: out = 16'(-229);
			28776: out = 16'(-216);
			28777: out = 16'(237);
			28778: out = 16'(214);
			28779: out = 16'(313);
			28780: out = 16'(-1754);
			28781: out = 16'(-2577);
			28782: out = 16'(-2392);
			28783: out = 16'(-925);
			28784: out = 16'(147);
			28785: out = 16'(-189);
			28786: out = 16'(-64);
			28787: out = 16'(-249);
			28788: out = 16'(652);
			28789: out = 16'(534);
			28790: out = 16'(527);
			28791: out = 16'(-858);
			28792: out = 16'(-959);
			28793: out = 16'(-855);
			28794: out = 16'(1464);
			28795: out = 16'(1926);
			28796: out = 16'(1749);
			28797: out = 16'(-339);
			28798: out = 16'(-896);
			28799: out = 16'(544);
			28800: out = 16'(126);
			28801: out = 16'(506);
			28802: out = 16'(85);
			28803: out = 16'(1806);
			28804: out = 16'(2013);
			28805: out = 16'(466);
			28806: out = 16'(-1695);
			28807: out = 16'(-3124);
			28808: out = 16'(-204);
			28809: out = 16'(-160);
			28810: out = 16'(-3);
			28811: out = 16'(238);
			28812: out = 16'(715);
			28813: out = 16'(1212);
			28814: out = 16'(466);
			28815: out = 16'(180);
			28816: out = 16'(-202);
			28817: out = 16'(858);
			28818: out = 16'(953);
			28819: out = 16'(256);
			28820: out = 16'(-1043);
			28821: out = 16'(-1936);
			28822: out = 16'(-1623);
			28823: out = 16'(-1393);
			28824: out = 16'(-817);
			28825: out = 16'(-1087);
			28826: out = 16'(-188);
			28827: out = 16'(588);
			28828: out = 16'(1754);
			28829: out = 16'(1576);
			28830: out = 16'(1115);
			28831: out = 16'(1121);
			28832: out = 16'(1742);
			28833: out = 16'(2989);
			28834: out = 16'(402);
			28835: out = 16'(-984);
			28836: out = 16'(-2601);
			28837: out = 16'(-836);
			28838: out = 16'(292);
			28839: out = 16'(1781);
			28840: out = 16'(332);
			28841: out = 16'(-658);
			28842: out = 16'(-1105);
			28843: out = 16'(103);
			28844: out = 16'(1214);
			28845: out = 16'(362);
			28846: out = 16'(418);
			28847: out = 16'(147);
			28848: out = 16'(479);
			28849: out = 16'(101);
			28850: out = 16'(-277);
			28851: out = 16'(156);
			28852: out = 16'(-14);
			28853: out = 16'(-529);
			28854: out = 16'(-938);
			28855: out = 16'(-1022);
			28856: out = 16'(-324);
			28857: out = 16'(-371);
			28858: out = 16'(123);
			28859: out = 16'(1014);
			28860: out = 16'(1144);
			28861: out = 16'(881);
			28862: out = 16'(317);
			28863: out = 16'(-247);
			28864: out = 16'(-518);
			28865: out = 16'(-1189);
			28866: out = 16'(-406);
			28867: out = 16'(566);
			28868: out = 16'(1503);
			28869: out = 16'(1190);
			28870: out = 16'(16);
			28871: out = 16'(-124);
			28872: out = 16'(-36);
			28873: out = 16'(1152);
			28874: out = 16'(277);
			28875: out = 16'(16);
			28876: out = 16'(-644);
			28877: out = 16'(-417);
			28878: out = 16'(-677);
			28879: out = 16'(-316);
			28880: out = 16'(-2168);
			28881: out = 16'(-3428);
			28882: out = 16'(-3967);
			28883: out = 16'(-1889);
			28884: out = 16'(784);
			28885: out = 16'(124);
			28886: out = 16'(418);
			28887: out = 16'(-329);
			28888: out = 16'(145);
			28889: out = 16'(-579);
			28890: out = 16'(-820);
			28891: out = 16'(-2261);
			28892: out = 16'(-1524);
			28893: out = 16'(382);
			28894: out = 16'(1546);
			28895: out = 16'(1575);
			28896: out = 16'(703);
			28897: out = 16'(-1707);
			28898: out = 16'(-3109);
			28899: out = 16'(-1621);
			28900: out = 16'(188);
			28901: out = 16'(2422);
			28902: out = 16'(2132);
			28903: out = 16'(2980);
			28904: out = 16'(2789);
			28905: out = 16'(3195);
			28906: out = 16'(1552);
			28907: out = 16'(-418);
			28908: out = 16'(-402);
			28909: out = 16'(-506);
			28910: out = 16'(-486);
			28911: out = 16'(-318);
			28912: out = 16'(160);
			28913: out = 16'(1816);
			28914: out = 16'(605);
			28915: out = 16'(-169);
			28916: out = 16'(-2048);
			28917: out = 16'(628);
			28918: out = 16'(2422);
			28919: out = 16'(1621);
			28920: out = 16'(-33);
			28921: out = 16'(-2233);
			28922: out = 16'(-402);
			28923: out = 16'(-712);
			28924: out = 16'(-331);
			28925: out = 16'(-1244);
			28926: out = 16'(-993);
			28927: out = 16'(-1239);
			28928: out = 16'(1229);
			28929: out = 16'(2084);
			28930: out = 16'(3694);
			28931: out = 16'(-1431);
			28932: out = 16'(-3912);
			28933: out = 16'(-4806);
			28934: out = 16'(-1616);
			28935: out = 16'(798);
			28936: out = 16'(1073);
			28937: out = 16'(39);
			28938: out = 16'(-1255);
			28939: out = 16'(-997);
			28940: out = 16'(-431);
			28941: out = 16'(587);
			28942: out = 16'(2114);
			28943: out = 16'(2386);
			28944: out = 16'(2230);
			28945: out = 16'(-1137);
			28946: out = 16'(-1701);
			28947: out = 16'(-1066);
			28948: out = 16'(2477);
			28949: out = 16'(2850);
			28950: out = 16'(29);
			28951: out = 16'(-2568);
			28952: out = 16'(-3658);
			28953: out = 16'(543);
			28954: out = 16'(144);
			28955: out = 16'(606);
			28956: out = 16'(-596);
			28957: out = 16'(106);
			28958: out = 16'(278);
			28959: out = 16'(1749);
			28960: out = 16'(1301);
			28961: out = 16'(1099);
			28962: out = 16'(144);
			28963: out = 16'(804);
			28964: out = 16'(1599);
			28965: out = 16'(1218);
			28966: out = 16'(172);
			28967: out = 16'(-1215);
			28968: out = 16'(-1853);
			28969: out = 16'(-1301);
			28970: out = 16'(307);
			28971: out = 16'(1641);
			28972: out = 16'(1927);
			28973: out = 16'(202);
			28974: out = 16'(-1459);
			28975: out = 16'(-2488);
			28976: out = 16'(263);
			28977: out = 16'(611);
			28978: out = 16'(1019);
			28979: out = 16'(158);
			28980: out = 16'(92);
			28981: out = 16'(24);
			28982: out = 16'(-1600);
			28983: out = 16'(-1560);
			28984: out = 16'(-317);
			28985: out = 16'(48);
			28986: out = 16'(534);
			28987: out = 16'(231);
			28988: out = 16'(935);
			28989: out = 16'(643);
			28990: out = 16'(-251);
			28991: out = 16'(-1698);
			28992: out = 16'(-2679);
			28993: out = 16'(-1717);
			28994: out = 16'(-1934);
			28995: out = 16'(-1553);
			28996: out = 16'(-1283);
			28997: out = 16'(134);
			28998: out = 16'(1216);
			28999: out = 16'(641);
			29000: out = 16'(-97);
			29001: out = 16'(-1065);
			29002: out = 16'(10);
			29003: out = 16'(521);
			29004: out = 16'(400);
			29005: out = 16'(1135);
			29006: out = 16'(358);
			29007: out = 16'(-1725);
			29008: out = 16'(-2751);
			29009: out = 16'(-2634);
			29010: out = 16'(-51);
			29011: out = 16'(237);
			29012: out = 16'(911);
			29013: out = 16'(2346);
			29014: out = 16'(1843);
			29015: out = 16'(878);
			29016: out = 16'(-145);
			29017: out = 16'(-235);
			29018: out = 16'(381);
			29019: out = 16'(-406);
			29020: out = 16'(-232);
			29021: out = 16'(-209);
			29022: out = 16'(866);
			29023: out = 16'(985);
			29024: out = 16'(402);
			29025: out = 16'(349);
			29026: out = 16'(159);
			29027: out = 16'(291);
			29028: out = 16'(-129);
			29029: out = 16'(227);
			29030: out = 16'(2881);
			29031: out = 16'(1867);
			29032: out = 16'(577);
			29033: out = 16'(-975);
			29034: out = 16'(-756);
			29035: out = 16'(322);
			29036: out = 16'(-1276);
			29037: out = 16'(-748);
			29038: out = 16'(-533);
			29039: out = 16'(2502);
			29040: out = 16'(1982);
			29041: out = 16'(233);
			29042: out = 16'(-3014);
			29043: out = 16'(-3455);
			29044: out = 16'(-206);
			29045: out = 16'(-567);
			29046: out = 16'(-817);
			29047: out = 16'(-3358);
			29048: out = 16'(-2241);
			29049: out = 16'(-1538);
			29050: out = 16'(-1036);
			29051: out = 16'(-263);
			29052: out = 16'(609);
			29053: out = 16'(1119);
			29054: out = 16'(754);
			29055: out = 16'(-312);
			29056: out = 16'(63);
			29057: out = 16'(-103);
			29058: out = 16'(506);
			29059: out = 16'(-2602);
			29060: out = 16'(-2474);
			29061: out = 16'(-838);
			29062: out = 16'(1109);
			29063: out = 16'(2073);
			29064: out = 16'(1812);
			29065: out = 16'(948);
			29066: out = 16'(238);
			29067: out = 16'(580);
			29068: out = 16'(1159);
			29069: out = 16'(1816);
			29070: out = 16'(269);
			29071: out = 16'(392);
			29072: out = 16'(217);
			29073: out = 16'(581);
			29074: out = 16'(125);
			29075: out = 16'(-215);
			29076: out = 16'(-1459);
			29077: out = 16'(-1975);
			29078: out = 16'(-2345);
			29079: out = 16'(328);
			29080: out = 16'(1886);
			29081: out = 16'(3004);
			29082: out = 16'(877);
			29083: out = 16'(-502);
			29084: out = 16'(-192);
			29085: out = 16'(-913);
			29086: out = 16'(-1068);
			29087: out = 16'(-1790);
			29088: out = 16'(-1248);
			29089: out = 16'(-789);
			29090: out = 16'(1162);
			29091: out = 16'(589);
			29092: out = 16'(-232);
			29093: out = 16'(-2111);
			29094: out = 16'(-1304);
			29095: out = 16'(945);
			29096: out = 16'(1869);
			29097: out = 16'(2865);
			29098: out = 16'(2780);
			29099: out = 16'(2695);
			29100: out = 16'(1335);
			29101: out = 16'(-1121);
			29102: out = 16'(-787);
			29103: out = 16'(-169);
			29104: out = 16'(304);
			29105: out = 16'(837);
			29106: out = 16'(1115);
			29107: out = 16'(2278);
			29108: out = 16'(1243);
			29109: out = 16'(134);
			29110: out = 16'(-453);
			29111: out = 16'(-226);
			29112: out = 16'(387);
			29113: out = 16'(132);
			29114: out = 16'(-124);
			29115: out = 16'(-640);
			29116: out = 16'(-1500);
			29117: out = 16'(-2358);
			29118: out = 16'(-3257);
			29119: out = 16'(-1819);
			29120: out = 16'(-599);
			29121: out = 16'(216);
			29122: out = 16'(287);
			29123: out = 16'(557);
			29124: out = 16'(2301);
			29125: out = 16'(2277);
			29126: out = 16'(1892);
			29127: out = 16'(-1549);
			29128: out = 16'(-2186);
			29129: out = 16'(-2542);
			29130: out = 16'(-1130);
			29131: out = 16'(-1841);
			29132: out = 16'(-3238);
			29133: out = 16'(-3053);
			29134: out = 16'(-2619);
			29135: out = 16'(-1426);
			29136: out = 16'(-671);
			29137: out = 16'(549);
			29138: out = 16'(1917);
			29139: out = 16'(3491);
			29140: out = 16'(3950);
			29141: out = 16'(1016);
			29142: out = 16'(1037);
			29143: out = 16'(234);
			29144: out = 16'(2215);
			29145: out = 16'(-1646);
			29146: out = 16'(-4893);
			29147: out = 16'(-5434);
			29148: out = 16'(-1789);
			29149: out = 16'(3749);
			29150: out = 16'(1849);
			29151: out = 16'(945);
			29152: out = 16'(-2034);
			29153: out = 16'(367);
			29154: out = 16'(386);
			29155: out = 16'(518);
			29156: out = 16'(-1668);
			29157: out = 16'(-2090);
			29158: out = 16'(-205);
			29159: out = 16'(-714);
			29160: out = 16'(-1030);
			29161: out = 16'(-1638);
			29162: out = 16'(-421);
			29163: out = 16'(1054);
			29164: out = 16'(1618);
			29165: out = 16'(2607);
			29166: out = 16'(2912);
			29167: out = 16'(2096);
			29168: out = 16'(833);
			29169: out = 16'(-458);
			29170: out = 16'(28);
			29171: out = 16'(1119);
			29172: out = 16'(3038);
			29173: out = 16'(1953);
			29174: out = 16'(933);
			29175: out = 16'(-1340);
			29176: out = 16'(-688);
			29177: out = 16'(-403);
			29178: out = 16'(459);
			29179: out = 16'(133);
			29180: out = 16'(253);
			29181: out = 16'(-539);
			29182: out = 16'(1682);
			29183: out = 16'(3491);
			29184: out = 16'(2245);
			29185: out = 16'(960);
			29186: out = 16'(-976);
			29187: out = 16'(-1091);
			29188: out = 16'(-1265);
			29189: out = 16'(-487);
			29190: out = 16'(-2273);
			29191: out = 16'(-3236);
			29192: out = 16'(-4984);
			29193: out = 16'(-2124);
			29194: out = 16'(-406);
			29195: out = 16'(1198);
			29196: out = 16'(255);
			29197: out = 16'(-116);
			29198: out = 16'(221);
			29199: out = 16'(1140);
			29200: out = 16'(1852);
			29201: out = 16'(2323);
			29202: out = 16'(1004);
			29203: out = 16'(-1028);
			29204: out = 16'(-3429);
			29205: out = 16'(-4246);
			29206: out = 16'(-3558);
			29207: out = 16'(-1043);
			29208: out = 16'(1457);
			29209: out = 16'(3637);
			29210: out = 16'(1822);
			29211: out = 16'(708);
			29212: out = 16'(358);
			29213: out = 16'(690);
			29214: out = 16'(1102);
			29215: out = 16'(189);
			29216: out = 16'(959);
			29217: out = 16'(702);
			29218: out = 16'(500);
			29219: out = 16'(-2124);
			29220: out = 16'(-3791);
			29221: out = 16'(-1341);
			29222: out = 16'(282);
			29223: out = 16'(1877);
			29224: out = 16'(1623);
			29225: out = 16'(1228);
			29226: out = 16'(207);
			29227: out = 16'(-662);
			29228: out = 16'(-1622);
			29229: out = 16'(-2392);
			29230: out = 16'(-968);
			29231: out = 16'(-73);
			29232: out = 16'(229);
			29233: out = 16'(304);
			29234: out = 16'(170);
			29235: out = 16'(-408);
			29236: out = 16'(146);
			29237: out = 16'(832);
			29238: out = 16'(3337);
			29239: out = 16'(2444);
			29240: out = 16'(1330);
			29241: out = 16'(-335);
			29242: out = 16'(-145);
			29243: out = 16'(306);
			29244: out = 16'(1006);
			29245: out = 16'(-550);
			29246: out = 16'(-3419);
			29247: out = 16'(-3737);
			29248: out = 16'(-2723);
			29249: out = 16'(773);
			29250: out = 16'(1130);
			29251: out = 16'(1840);
			29252: out = 16'(774);
			29253: out = 16'(1662);
			29254: out = 16'(1036);
			29255: out = 16'(-803);
			29256: out = 16'(-2018);
			29257: out = 16'(-1881);
			29258: out = 16'(1260);
			29259: out = 16'(2886);
			29260: out = 16'(3643);
			29261: out = 16'(148);
			29262: out = 16'(-1953);
			29263: out = 16'(-4064);
			29264: out = 16'(-3078);
			29265: out = 16'(-3299);
			29266: out = 16'(-3591);
			29267: out = 16'(-1281);
			29268: out = 16'(1088);
			29269: out = 16'(3484);
			29270: out = 16'(2832);
			29271: out = 16'(1852);
			29272: out = 16'(1306);
			29273: out = 16'(-675);
			29274: out = 16'(-1736);
			29275: out = 16'(-1074);
			29276: out = 16'(101);
			29277: out = 16'(1223);
			29278: out = 16'(285);
			29279: out = 16'(149);
			29280: out = 16'(-221);
			29281: out = 16'(408);
			29282: out = 16'(451);
			29283: out = 16'(418);
			29284: out = 16'(-125);
			29285: out = 16'(-1180);
			29286: out = 16'(-3164);
			29287: out = 16'(-1492);
			29288: out = 16'(-857);
			29289: out = 16'(-915);
			29290: out = 16'(-2132);
			29291: out = 16'(-2783);
			29292: out = 16'(-645);
			29293: out = 16'(-982);
			29294: out = 16'(-727);
			29295: out = 16'(-3001);
			29296: out = 16'(-569);
			29297: out = 16'(1734);
			29298: out = 16'(4053);
			29299: out = 16'(2483);
			29300: out = 16'(-569);
			29301: out = 16'(-1708);
			29302: out = 16'(-1602);
			29303: out = 16'(290);
			29304: out = 16'(-15);
			29305: out = 16'(-545);
			29306: out = 16'(-2968);
			29307: out = 16'(-1387);
			29308: out = 16'(254);
			29309: out = 16'(3718);
			29310: out = 16'(3584);
			29311: out = 16'(3415);
			29312: out = 16'(1728);
			29313: out = 16'(2416);
			29314: out = 16'(2719);
			29315: out = 16'(1233);
			29316: out = 16'(368);
			29317: out = 16'(-547);
			29318: out = 16'(-153);
			29319: out = 16'(-366);
			29320: out = 16'(-329);
			29321: out = 16'(-575);
			29322: out = 16'(622);
			29323: out = 16'(2903);
			29324: out = 16'(2293);
			29325: out = 16'(1818);
			29326: out = 16'(891);
			29327: out = 16'(126);
			29328: out = 16'(-535);
			29329: out = 16'(-449);
			29330: out = 16'(-301);
			29331: out = 16'(102);
			29332: out = 16'(-1281);
			29333: out = 16'(-735);
			29334: out = 16'(-415);
			29335: out = 16'(2030);
			29336: out = 16'(1263);
			29337: out = 16'(195);
			29338: out = 16'(-1600);
			29339: out = 16'(-1134);
			29340: out = 16'(368);
			29341: out = 16'(1683);
			29342: out = 16'(1590);
			29343: out = 16'(-20);
			29344: out = 16'(-1771);
			29345: out = 16'(-2375);
			29346: out = 16'(-494);
			29347: out = 16'(646);
			29348: out = 16'(1821);
			29349: out = 16'(1952);
			29350: out = 16'(911);
			29351: out = 16'(-1044);
			29352: out = 16'(-2769);
			29353: out = 16'(-3842);
			29354: out = 16'(-3696);
			29355: out = 16'(-4074);
			29356: out = 16'(-2333);
			29357: out = 16'(-144);
			29358: out = 16'(-352);
			29359: out = 16'(-231);
			29360: out = 16'(-289);
			29361: out = 16'(-692);
			29362: out = 16'(-1241);
			29363: out = 16'(-2239);
			29364: out = 16'(-1331);
			29365: out = 16'(-568);
			29366: out = 16'(-220);
			29367: out = 16'(14);
			29368: out = 16'(244);
			29369: out = 16'(1890);
			29370: out = 16'(950);
			29371: out = 16'(-76);
			29372: out = 16'(1184);
			29373: out = 16'(1410);
			29374: out = 16'(1770);
			29375: out = 16'(-1123);
			29376: out = 16'(-1663);
			29377: out = 16'(-1516);
			29378: out = 16'(112);
			29379: out = 16'(866);
			29380: out = 16'(1226);
			29381: out = 16'(703);
			29382: out = 16'(575);
			29383: out = 16'(438);
			29384: out = 16'(2078);
			29385: out = 16'(2880);
			29386: out = 16'(2265);
			29387: out = 16'(804);
			29388: out = 16'(-705);
			29389: out = 16'(-90);
			29390: out = 16'(-376);
			29391: out = 16'(-185);
			29392: out = 16'(-1059);
			29393: out = 16'(-1049);
			29394: out = 16'(-1115);
			29395: out = 16'(-1512);
			29396: out = 16'(-1753);
			29397: out = 16'(-1534);
			29398: out = 16'(-582);
			29399: out = 16'(304);
			29400: out = 16'(382);
			29401: out = 16'(1148);
			29402: out = 16'(765);
			29403: out = 16'(95);
			29404: out = 16'(-1926);
			29405: out = 16'(-2891);
			29406: out = 16'(-1708);
			29407: out = 16'(209);
			29408: out = 16'(2133);
			29409: out = 16'(1680);
			29410: out = 16'(1368);
			29411: out = 16'(295);
			29412: out = 16'(590);
			29413: out = 16'(-316);
			29414: out = 16'(-919);
			29415: out = 16'(-396);
			29416: out = 16'(536);
			29417: out = 16'(1749);
			29418: out = 16'(1732);
			29419: out = 16'(1381);
			29420: out = 16'(400);
			29421: out = 16'(330);
			29422: out = 16'(219);
			29423: out = 16'(440);
			29424: out = 16'(274);
			29425: out = 16'(-77);
			29426: out = 16'(-2367);
			29427: out = 16'(-1490);
			29428: out = 16'(-215);
			29429: out = 16'(-514);
			29430: out = 16'(-60);
			29431: out = 16'(315);
			29432: out = 16'(972);
			29433: out = 16'(860);
			29434: out = 16'(124);
			29435: out = 16'(-164);
			29436: out = 16'(-419);
			29437: out = 16'(452);
			29438: out = 16'(-2188);
			29439: out = 16'(-2787);
			29440: out = 16'(-966);
			29441: out = 16'(648);
			29442: out = 16'(1957);
			29443: out = 16'(898);
			29444: out = 16'(1861);
			29445: out = 16'(1962);
			29446: out = 16'(71);
			29447: out = 16'(-1260);
			29448: out = 16'(-2373);
			29449: out = 16'(666);
			29450: out = 16'(1311);
			29451: out = 16'(1604);
			29452: out = 16'(-1601);
			29453: out = 16'(-2584);
			29454: out = 16'(-2279);
			29455: out = 16'(-797);
			29456: out = 16'(332);
			29457: out = 16'(1115);
			29458: out = 16'(660);
			29459: out = 16'(873);
			29460: out = 16'(2808);
			29461: out = 16'(2536);
			29462: out = 16'(1244);
			29463: out = 16'(-4153);
			29464: out = 16'(-4755);
			29465: out = 16'(-4107);
			29466: out = 16'(-2092);
			29467: out = 16'(-529);
			29468: out = 16'(478);
			29469: out = 16'(1815);
			29470: out = 16'(454);
			29471: out = 16'(-2483);
			29472: out = 16'(-2687);
			29473: out = 16'(-1881);
			29474: out = 16'(1714);
			29475: out = 16'(80);
			29476: out = 16'(745);
			29477: out = 16'(2269);
			29478: out = 16'(3325);
			29479: out = 16'(2906);
			29480: out = 16'(602);
			29481: out = 16'(-1631);
			29482: out = 16'(-2858);
			29483: out = 16'(138);
			29484: out = 16'(1055);
			29485: out = 16'(1798);
			29486: out = 16'(630);
			29487: out = 16'(236);
			29488: out = 16'(-206);
			29489: out = 16'(-130);
			29490: out = 16'(-23);
			29491: out = 16'(336);
			29492: out = 16'(266);
			29493: out = 16'(140);
			29494: out = 16'(-403);
			29495: out = 16'(-340);
			29496: out = 16'(-258);
			29497: out = 16'(309);
			29498: out = 16'(414);
			29499: out = 16'(266);
			29500: out = 16'(-1633);
			29501: out = 16'(-1644);
			29502: out = 16'(-1397);
			29503: out = 16'(1615);
			29504: out = 16'(925);
			29505: out = 16'(-284);
			29506: out = 16'(-1398);
			29507: out = 16'(-1020);
			29508: out = 16'(549);
			29509: out = 16'(-268);
			29510: out = 16'(-237);
			29511: out = 16'(-358);
			29512: out = 16'(-676);
			29513: out = 16'(-1143);
			29514: out = 16'(-1534);
			29515: out = 16'(-782);
			29516: out = 16'(77);
			29517: out = 16'(282);
			29518: out = 16'(1019);
			29519: out = 16'(1499);
			29520: out = 16'(3484);
			29521: out = 16'(2920);
			29522: out = 16'(1871);
			29523: out = 16'(-2388);
			29524: out = 16'(-2887);
			29525: out = 16'(-2061);
			29526: out = 16'(-618);
			29527: out = 16'(-686);
			29528: out = 16'(-2377);
			29529: out = 16'(-520);
			29530: out = 16'(64);
			29531: out = 16'(791);
			29532: out = 16'(507);
			29533: out = 16'(1234);
			29534: out = 16'(2876);
			29535: out = 16'(3374);
			29536: out = 16'(2888);
			29537: out = 16'(29);
			29538: out = 16'(-981);
			29539: out = 16'(-1736);
			29540: out = 16'(-974);
			29541: out = 16'(-765);
			29542: out = 16'(-140);
			29543: out = 16'(-469);
			29544: out = 16'(380);
			29545: out = 16'(1210);
			29546: out = 16'(3410);
			29547: out = 16'(3864);
			29548: out = 16'(3174);
			29549: out = 16'(1293);
			29550: out = 16'(-606);
			29551: out = 16'(-2410);
			29552: out = 16'(-2149);
			29553: out = 16'(-1386);
			29554: out = 16'(-334);
			29555: out = 16'(93);
			29556: out = 16'(237);
			29557: out = 16'(184);
			29558: out = 16'(618);
			29559: out = 16'(1050);
			29560: out = 16'(971);
			29561: out = 16'(502);
			29562: out = 16'(-475);
			29563: out = 16'(-847);
			29564: out = 16'(-1094);
			29565: out = 16'(-234);
			29566: out = 16'(-678);
			29567: out = 16'(-45);
			29568: out = 16'(-39);
			29569: out = 16'(1824);
			29570: out = 16'(1645);
			29571: out = 16'(419);
			29572: out = 16'(-2859);
			29573: out = 16'(-4311);
			29574: out = 16'(-1237);
			29575: out = 16'(1300);
			29576: out = 16'(3615);
			29577: out = 16'(1543);
			29578: out = 16'(1440);
			29579: out = 16'(713);
			29580: out = 16'(571);
			29581: out = 16'(-318);
			29582: out = 16'(-1213);
			29583: out = 16'(-1116);
			29584: out = 16'(-1194);
			29585: out = 16'(-1015);
			29586: out = 16'(-1712);
			29587: out = 16'(-813);
			29588: out = 16'(2270);
			29589: out = 16'(2182);
			29590: out = 16'(1645);
			29591: out = 16'(-1120);
			29592: out = 16'(-652);
			29593: out = 16'(-72);
			29594: out = 16'(836);
			29595: out = 16'(446);
			29596: out = 16'(-499);
			29597: out = 16'(374);
			29598: out = 16'(-1069);
			29599: out = 16'(-2566);
			29600: out = 16'(-4234);
			29601: out = 16'(-3848);
			29602: out = 16'(-2164);
			29603: out = 16'(-374);
			29604: out = 16'(534);
			29605: out = 16'(253);
			29606: out = 16'(71);
			29607: out = 16'(200);
			29608: out = 16'(1769);
			29609: out = 16'(1358);
			29610: out = 16'(717);
			29611: out = 16'(-867);
			29612: out = 16'(-1464);
			29613: out = 16'(-1725);
			29614: out = 16'(-2352);
			29615: out = 16'(-1650);
			29616: out = 16'(-539);
			29617: out = 16'(3396);
			29618: out = 16'(4160);
			29619: out = 16'(3821);
			29620: out = 16'(1089);
			29621: out = 16'(530);
			29622: out = 16'(1670);
			29623: out = 16'(174);
			29624: out = 16'(-689);
			29625: out = 16'(-1005);
			29626: out = 16'(-2631);
			29627: out = 16'(-2936);
			29628: out = 16'(-1877);
			29629: out = 16'(364);
			29630: out = 16'(1718);
			29631: out = 16'(358);
			29632: out = 16'(-1398);
			29633: out = 16'(-3135);
			29634: out = 16'(-284);
			29635: out = 16'(102);
			29636: out = 16'(601);
			29637: out = 16'(310);
			29638: out = 16'(177);
			29639: out = 16'(-217);
			29640: out = 16'(-1208);
			29641: out = 16'(-2115);
			29642: out = 16'(-2986);
			29643: out = 16'(-674);
			29644: out = 16'(1140);
			29645: out = 16'(2297);
			29646: out = 16'(1749);
			29647: out = 16'(654);
			29648: out = 16'(-803);
			29649: out = 16'(-1084);
			29650: out = 16'(-626);
			29651: out = 16'(936);
			29652: out = 16'(1785);
			29653: out = 16'(2236);
			29654: out = 16'(534);
			29655: out = 16'(-272);
			29656: out = 16'(-1064);
			29657: out = 16'(1299);
			29658: out = 16'(1518);
			29659: out = 16'(996);
			29660: out = 16'(-62);
			29661: out = 16'(-305);
			29662: out = 16'(478);
			29663: out = 16'(743);
			29664: out = 16'(1182);
			29665: out = 16'(1557);
			29666: out = 16'(427);
			29667: out = 16'(-1109);
			29668: out = 16'(-2966);
			29669: out = 16'(-2603);
			29670: out = 16'(-1449);
			29671: out = 16'(-1969);
			29672: out = 16'(-774);
			29673: out = 16'(-135);
			29674: out = 16'(580);
			29675: out = 16'(-119);
			29676: out = 16'(-917);
			29677: out = 16'(-1155);
			29678: out = 16'(170);
			29679: out = 16'(2397);
			29680: out = 16'(2824);
			29681: out = 16'(1942);
			29682: out = 16'(-1141);
			29683: out = 16'(-1482);
			29684: out = 16'(-1516);
			29685: out = 16'(-119);
			29686: out = 16'(-202);
			29687: out = 16'(67);
			29688: out = 16'(1667);
			29689: out = 16'(1079);
			29690: out = 16'(170);
			29691: out = 16'(-2121);
			29692: out = 16'(-1518);
			29693: out = 16'(204);
			29694: out = 16'(2291);
			29695: out = 16'(2295);
			29696: out = 16'(48);
			29697: out = 16'(1657);
			29698: out = 16'(1215);
			29699: out = 16'(1150);
			29700: out = 16'(-2065);
			29701: out = 16'(-2925);
			29702: out = 16'(-996);
			29703: out = 16'(-310);
			29704: out = 16'(271);
			29705: out = 16'(-1137);
			29706: out = 16'(-213);
			29707: out = 16'(419);
			29708: out = 16'(1083);
			29709: out = 16'(734);
			29710: out = 16'(44);
			29711: out = 16'(-1341);
			29712: out = 16'(-2549);
			29713: out = 16'(-3673);
			29714: out = 16'(-397);
			29715: out = 16'(1361);
			29716: out = 16'(3032);
			29717: out = 16'(601);
			29718: out = 16'(-286);
			29719: out = 16'(-299);
			29720: out = 16'(101);
			29721: out = 16'(273);
			29722: out = 16'(-124);
			29723: out = 16'(-224);
			29724: out = 16'(-618);
			29725: out = 16'(-3009);
			29726: out = 16'(-1259);
			29727: out = 16'(868);
			29728: out = 16'(2040);
			29729: out = 16'(2482);
			29730: out = 16'(2058);
			29731: out = 16'(154);
			29732: out = 16'(-1005);
			29733: out = 16'(-1648);
			29734: out = 16'(-133);
			29735: out = 16'(242);
			29736: out = 16'(-430);
			29737: out = 16'(-135);
			29738: out = 16'(220);
			29739: out = 16'(1828);
			29740: out = 16'(773);
			29741: out = 16'(-189);
			29742: out = 16'(-2362);
			29743: out = 16'(-1228);
			29744: out = 16'(-218);
			29745: out = 16'(-1013);
			29746: out = 16'(-882);
			29747: out = 16'(-892);
			29748: out = 16'(286);
			29749: out = 16'(113);
			29750: out = 16'(-312);
			29751: out = 16'(-812);
			29752: out = 16'(-636);
			29753: out = 16'(59);
			29754: out = 16'(337);
			29755: out = 16'(995);
			29756: out = 16'(1763);
			29757: out = 16'(1004);
			29758: out = 16'(-29);
			29759: out = 16'(-1536);
			29760: out = 16'(-1684);
			29761: out = 16'(-1342);
			29762: out = 16'(-325);
			29763: out = 16'(-202);
			29764: out = 16'(-67);
			29765: out = 16'(1721);
			29766: out = 16'(1776);
			29767: out = 16'(1754);
			29768: out = 16'(466);
			29769: out = 16'(400);
			29770: out = 16'(489);
			29771: out = 16'(1968);
			29772: out = 16'(2088);
			29773: out = 16'(1606);
			29774: out = 16'(133);
			29775: out = 16'(-837);
			29776: out = 16'(-1834);
			29777: out = 16'(88);
			29778: out = 16'(1138);
			29779: out = 16'(1027);
			29780: out = 16'(-525);
			29781: out = 16'(-1795);
			29782: out = 16'(210);
			29783: out = 16'(534);
			29784: out = 16'(1050);
			29785: out = 16'(-352);
			29786: out = 16'(-680);
			29787: out = 16'(-1103);
			29788: out = 16'(159);
			29789: out = 16'(957);
			29790: out = 16'(2296);
			29791: out = 16'(146);
			29792: out = 16'(-353);
			29793: out = 16'(-373);
			29794: out = 16'(617);
			29795: out = 16'(799);
			29796: out = 16'(176);
			29797: out = 16'(-1495);
			29798: out = 16'(-2346);
			29799: out = 16'(251);
			29800: out = 16'(51);
			29801: out = 16'(20);
			29802: out = 16'(-3078);
			29803: out = 16'(-1864);
			29804: out = 16'(-56);
			29805: out = 16'(1344);
			29806: out = 16'(1755);
			29807: out = 16'(1498);
			29808: out = 16'(-1005);
			29809: out = 16'(-2164);
			29810: out = 16'(-2249);
			29811: out = 16'(-921);
			29812: out = 16'(811);
			29813: out = 16'(2802);
			29814: out = 16'(2871);
			29815: out = 16'(2306);
			29816: out = 16'(322);
			29817: out = 16'(310);
			29818: out = 16'(-256);
			29819: out = 16'(-1587);
			29820: out = 16'(-2950);
			29821: out = 16'(-3801);
			29822: out = 16'(-2563);
			29823: out = 16'(-1100);
			29824: out = 16'(752);
			29825: out = 16'(-263);
			29826: out = 16'(-649);
			29827: out = 16'(-1763);
			29828: out = 16'(726);
			29829: out = 16'(1184);
			29830: out = 16'(1190);
			29831: out = 16'(-319);
			29832: out = 16'(-1457);
			29833: out = 16'(-3059);
			29834: out = 16'(-1611);
			29835: out = 16'(-558);
			29836: out = 16'(428);
			29837: out = 16'(379);
			29838: out = 16'(558);
			29839: out = 16'(240);
			29840: out = 16'(1261);
			29841: out = 16'(1856);
			29842: out = 16'(4038);
			29843: out = 16'(2238);
			29844: out = 16'(-390);
			29845: out = 16'(-1513);
			29846: out = 16'(-617);
			29847: out = 16'(1828);
			29848: out = 16'(2585);
			29849: out = 16'(1963);
			29850: out = 16'(-490);
			29851: out = 16'(-2798);
			29852: out = 16'(-3227);
			29853: out = 16'(493);
			29854: out = 16'(2106);
			29855: out = 16'(3301);
			29856: out = 16'(258);
			29857: out = 16'(439);
			29858: out = 16'(-132);
			29859: out = 16'(-903);
			29860: out = 16'(-1260);
			29861: out = 16'(-982);
			29862: out = 16'(-610);
			29863: out = 16'(-542);
			29864: out = 16'(-1188);
			29865: out = 16'(-250);
			29866: out = 16'(-128);
			29867: out = 16'(378);
			29868: out = 16'(-1263);
			29869: out = 16'(-1457);
			29870: out = 16'(-323);
			29871: out = 16'(54);
			29872: out = 16'(364);
			29873: out = 16'(238);
			29874: out = 16'(460);
			29875: out = 16'(237);
			29876: out = 16'(-1570);
			29877: out = 16'(-1394);
			29878: out = 16'(-787);
			29879: out = 16'(364);
			29880: out = 16'(317);
			29881: out = 16'(-158);
			29882: out = 16'(413);
			29883: out = 16'(1088);
			29884: out = 16'(2435);
			29885: out = 16'(1249);
			29886: out = 16'(919);
			29887: out = 16'(292);
			29888: out = 16'(1734);
			29889: out = 16'(1844);
			29890: out = 16'(301);
			29891: out = 16'(-466);
			29892: out = 16'(-1745);
			29893: out = 16'(-3646);
			29894: out = 16'(-3983);
			29895: out = 16'(-3082);
			29896: out = 16'(1216);
			29897: out = 16'(2459);
			29898: out = 16'(2687);
			29899: out = 16'(258);
			29900: out = 16'(-351);
			29901: out = 16'(-121);
			29902: out = 16'(-951);
			29903: out = 16'(-643);
			29904: out = 16'(321);
			29905: out = 16'(440);
			29906: out = 16'(13);
			29907: out = 16'(-1835);
			29908: out = 16'(-714);
			29909: out = 16'(-242);
			29910: out = 16'(410);
			29911: out = 16'(-892);
			29912: out = 16'(-1647);
			29913: out = 16'(-993);
			29914: out = 16'(112);
			29915: out = 16'(1474);
			29916: out = 16'(2099);
			29917: out = 16'(2184);
			29918: out = 16'(1437);
			29919: out = 16'(656);
			29920: out = 16'(-440);
			29921: out = 16'(-957);
			29922: out = 16'(-253);
			29923: out = 16'(1169);
			29924: out = 16'(2733);
			29925: out = 16'(2859);
			29926: out = 16'(2030);
			29927: out = 16'(144);
			29928: out = 16'(-1202);
			29929: out = 16'(-1906);
			29930: out = 16'(-1158);
			29931: out = 16'(-846);
			29932: out = 16'(-411);
			29933: out = 16'(-508);
			29934: out = 16'(-719);
			29935: out = 16'(-1334);
			29936: out = 16'(-2780);
			29937: out = 16'(-3195);
			29938: out = 16'(-2824);
			29939: out = 16'(-1435);
			29940: out = 16'(-293);
			29941: out = 16'(372);
			29942: out = 16'(638);
			29943: out = 16'(525);
			29944: out = 16'(651);
			29945: out = 16'(-440);
			29946: out = 16'(-1094);
			29947: out = 16'(-1571);
			29948: out = 16'(-757);
			29949: out = 16'(-64);
			29950: out = 16'(-9);
			29951: out = 16'(-395);
			29952: out = 16'(-835);
			29953: out = 16'(-7);
			29954: out = 16'(523);
			29955: out = 16'(1362);
			29956: out = 16'(-135);
			29957: out = 16'(368);
			29958: out = 16'(1322);
			29959: out = 16'(2125);
			29960: out = 16'(2096);
			29961: out = 16'(971);
			29962: out = 16'(1647);
			29963: out = 16'(1331);
			29964: out = 16'(244);
			29965: out = 16'(-199);
			29966: out = 16'(-365);
			29967: out = 16'(514);
			29968: out = 16'(-812);
			29969: out = 16'(-1783);
			29970: out = 16'(-344);
			29971: out = 16'(-360);
			29972: out = 16'(-132);
			29973: out = 16'(-1681);
			29974: out = 16'(-681);
			29975: out = 16'(720);
			29976: out = 16'(2533);
			29977: out = 16'(2021);
			29978: out = 16'(-491);
			29979: out = 16'(-2);
			29980: out = 16'(-1244);
			29981: out = 16'(-2927);
			29982: out = 16'(-2667);
			29983: out = 16'(-1035);
			29984: out = 16'(2980);
			29985: out = 16'(2248);
			29986: out = 16'(1434);
			29987: out = 16'(438);
			29988: out = 16'(40);
			29989: out = 16'(-161);
			29990: out = 16'(-155);
			29991: out = 16'(-200);
			29992: out = 16'(-302);
			29993: out = 16'(395);
			29994: out = 16'(693);
			29995: out = 16'(1144);
			29996: out = 16'(370);
			29997: out = 16'(343);
			29998: out = 16'(407);
			29999: out = 16'(484);
			30000: out = 16'(170);
			30001: out = 16'(-350);
			30002: out = 16'(-829);
			30003: out = 16'(-1177);
			30004: out = 16'(-2337);
			30005: out = 16'(-1093);
			30006: out = 16'(-206);
			30007: out = 16'(-16);
			30008: out = 16'(-1120);
			30009: out = 16'(-2221);
			30010: out = 16'(-1613);
			30011: out = 16'(-361);
			30012: out = 16'(1363);
			30013: out = 16'(51);
			30014: out = 16'(125);
			30015: out = 16'(440);
			30016: out = 16'(-9);
			30017: out = 16'(434);
			30018: out = 16'(1744);
			30019: out = 16'(2068);
			30020: out = 16'(1893);
			30021: out = 16'(417);
			30022: out = 16'(1);
			30023: out = 16'(-416);
			30024: out = 16'(-112);
			30025: out = 16'(72);
			30026: out = 16'(539);
			30027: out = 16'(189);
			30028: out = 16'(313);
			30029: out = 16'(172);
			30030: out = 16'(472);
			30031: out = 16'(268);
			30032: out = 16'(269);
			30033: out = 16'(-880);
			30034: out = 16'(-573);
			30035: out = 16'(486);
			30036: out = 16'(1196);
			30037: out = 16'(1761);
			30038: out = 16'(2002);
			30039: out = 16'(1402);
			30040: out = 16'(106);
			30041: out = 16'(-2972);
			30042: out = 16'(-2692);
			30043: out = 16'(-2047);
			30044: out = 16'(-445);
			30045: out = 16'(-976);
			30046: out = 16'(-1596);
			30047: out = 16'(-474);
			30048: out = 16'(512);
			30049: out = 16'(1736);
			30050: out = 16'(68);
			30051: out = 16'(-401);
			30052: out = 16'(-1041);
			30053: out = 16'(-879);
			30054: out = 16'(-1018);
			30055: out = 16'(-812);
			30056: out = 16'(-1016);
			30057: out = 16'(-474);
			30058: out = 16'(445);
			30059: out = 16'(1598);
			30060: out = 16'(2200);
			30061: out = 16'(1606);
			30062: out = 16'(1272);
			30063: out = 16'(760);
			30064: out = 16'(-254);
			30065: out = 16'(-1303);
			30066: out = 16'(-2483);
			30067: out = 16'(-1009);
			30068: out = 16'(-1365);
			30069: out = 16'(-1509);
			30070: out = 16'(-2854);
			30071: out = 16'(-1882);
			30072: out = 16'(8);
			30073: out = 16'(2523);
			30074: out = 16'(3101);
			30075: out = 16'(1593);
			30076: out = 16'(-417);
			30077: out = 16'(-1913);
			30078: out = 16'(-1513);
			30079: out = 16'(-465);
			30080: out = 16'(759);
			30081: out = 16'(189);
			30082: out = 16'(-192);
			30083: out = 16'(-937);
			30084: out = 16'(1610);
			30085: out = 16'(1320);
			30086: out = 16'(1058);
			30087: out = 16'(-121);
			30088: out = 16'(633);
			30089: out = 16'(2252);
			30090: out = 16'(718);
			30091: out = 16'(105);
			30092: out = 16'(-463);
			30093: out = 16'(977);
			30094: out = 16'(1427);
			30095: out = 16'(190);
			30096: out = 16'(-20);
			30097: out = 16'(-513);
			30098: out = 16'(1190);
			30099: out = 16'(-752);
			30100: out = 16'(-1804);
			30101: out = 16'(-2554);
			30102: out = 16'(-91);
			30103: out = 16'(2209);
			30104: out = 16'(-75);
			30105: out = 16'(-2041);
			30106: out = 16'(-4514);
			30107: out = 16'(-1529);
			30108: out = 16'(-141);
			30109: out = 16'(1143);
			30110: out = 16'(160);
			30111: out = 16'(-1411);
			30112: out = 16'(-4313);
			30113: out = 16'(-3806);
			30114: out = 16'(-2295);
			30115: out = 16'(1870);
			30116: out = 16'(2455);
			30117: out = 16'(2694);
			30118: out = 16'(-268);
			30119: out = 16'(228);
			30120: out = 16'(344);
			30121: out = 16'(1306);
			30122: out = 16'(107);
			30123: out = 16'(-871);
			30124: out = 16'(-1070);
			30125: out = 16'(806);
			30126: out = 16'(3554);
			30127: out = 16'(2424);
			30128: out = 16'(1238);
			30129: out = 16'(-1152);
			30130: out = 16'(-361);
			30131: out = 16'(490);
			30132: out = 16'(2816);
			30133: out = 16'(2585);
			30134: out = 16'(2322);
			30135: out = 16'(189);
			30136: out = 16'(49);
			30137: out = 16'(-368);
			30138: out = 16'(1661);
			30139: out = 16'(-22);
			30140: out = 16'(-1425);
			30141: out = 16'(-4332);
			30142: out = 16'(-2785);
			30143: out = 16'(-54);
			30144: out = 16'(1246);
			30145: out = 16'(829);
			30146: out = 16'(-1258);
			30147: out = 16'(-520);
			30148: out = 16'(251);
			30149: out = 16'(2283);
			30150: out = 16'(859);
			30151: out = 16'(-296);
			30152: out = 16'(-2347);
			30153: out = 16'(-2366);
			30154: out = 16'(-1900);
			30155: out = 16'(197);
			30156: out = 16'(381);
			30157: out = 16'(711);
			30158: out = 16'(2578);
			30159: out = 16'(2443);
			30160: out = 16'(1764);
			30161: out = 16'(-1760);
			30162: out = 16'(-2259);
			30163: out = 16'(-1463);
			30164: out = 16'(-537);
			30165: out = 16'(126);
			30166: out = 16'(196);
			30167: out = 16'(317);
			30168: out = 16'(77);
			30169: out = 16'(-389);
			30170: out = 16'(-337);
			30171: out = 16'(-375);
			30172: out = 16'(-300);
			30173: out = 16'(-58);
			30174: out = 16'(451);
			30175: out = 16'(290);
			30176: out = 16'(1183);
			30177: out = 16'(1446);
			30178: out = 16'(1248);
			30179: out = 16'(-552);
			30180: out = 16'(-2513);
			30181: out = 16'(-3488);
			30182: out = 16'(-2275);
			30183: out = 16'(678);
			30184: out = 16'(775);
			30185: out = 16'(956);
			30186: out = 16'(-343);
			30187: out = 16'(486);
			30188: out = 16'(234);
			30189: out = 16'(-28);
			30190: out = 16'(-276);
			30191: out = 16'(355);
			30192: out = 16'(2004);
			30193: out = 16'(2861);
			30194: out = 16'(2934);
			30195: out = 16'(1088);
			30196: out = 16'(477);
			30197: out = 16'(46);
			30198: out = 16'(-284);
			30199: out = 16'(-104);
			30200: out = 16'(365);
			30201: out = 16'(679);
			30202: out = 16'(1260);
			30203: out = 16'(1967);
			30204: out = 16'(104);
			30205: out = 16'(-1386);
			30206: out = 16'(-3182);
			30207: out = 16'(-959);
			30208: out = 16'(372);
			30209: out = 16'(-57);
			30210: out = 16'(250);
			30211: out = 16'(-70);
			30212: out = 16'(-116);
			30213: out = 16'(-1151);
			30214: out = 16'(-1824);
			30215: out = 16'(-2352);
			30216: out = 16'(-1472);
			30217: out = 16'(-202);
			30218: out = 16'(-464);
			30219: out = 16'(-302);
			30220: out = 16'(-392);
			30221: out = 16'(-333);
			30222: out = 16'(-296);
			30223: out = 16'(-102);
			30224: out = 16'(185);
			30225: out = 16'(-340);
			30226: out = 16'(-3091);
			30227: out = 16'(-751);
			30228: out = 16'(896);
			30229: out = 16'(2774);
			30230: out = 16'(1780);
			30231: out = 16'(706);
			30232: out = 16'(-896);
			30233: out = 16'(-443);
			30234: out = 16'(609);
			30235: out = 16'(3372);
			30236: out = 16'(3150);
			30237: out = 16'(1640);
			30238: out = 16'(-937);
			30239: out = 16'(-2300);
			30240: out = 16'(-2181);
			30241: out = 16'(-1583);
			30242: out = 16'(-409);
			30243: out = 16'(258);
			30244: out = 16'(1710);
			30245: out = 16'(1759);
			30246: out = 16'(286);
			30247: out = 16'(232);
			30248: out = 16'(-21);
			30249: out = 16'(-479);
			30250: out = 16'(-831);
			30251: out = 16'(-1234);
			30252: out = 16'(-1677);
			30253: out = 16'(-954);
			30254: out = 16'(485);
			30255: out = 16'(-448);
			30256: out = 16'(675);
			30257: out = 16'(1513);
			30258: out = 16'(3855);
			30259: out = 16'(2899);
			30260: out = 16'(38);
			30261: out = 16'(-3145);
			30262: out = 16'(-4441);
			30263: out = 16'(-2039);
			30264: out = 16'(-2198);
			30265: out = 16'(-1106);
			30266: out = 16'(-630);
			30267: out = 16'(972);
			30268: out = 16'(1837);
			30269: out = 16'(3239);
			30270: out = 16'(2316);
			30271: out = 16'(1194);
			30272: out = 16'(-875);
			30273: out = 16'(-695);
			30274: out = 16'(206);
			30275: out = 16'(171);
			30276: out = 16'(-1349);
			30277: out = 16'(-4793);
			30278: out = 16'(-1536);
			30279: out = 16'(-665);
			30280: out = 16'(730);
			30281: out = 16'(-1689);
			30282: out = 16'(-1758);
			30283: out = 16'(-443);
			30284: out = 16'(2099);
			30285: out = 16'(3436);
			30286: out = 16'(3270);
			30287: out = 16'(1550);
			30288: out = 16'(-408);
			30289: out = 16'(-2837);
			30290: out = 16'(-1878);
			30291: out = 16'(-46);
			30292: out = 16'(1303);
			30293: out = 16'(942);
			30294: out = 16'(-386);
			30295: out = 16'(-261);
			30296: out = 16'(658);
			30297: out = 16'(2771);
			30298: out = 16'(1768);
			30299: out = 16'(600);
			30300: out = 16'(-1879);
			30301: out = 16'(-2205);
			30302: out = 16'(-1982);
			30303: out = 16'(226);
			30304: out = 16'(127);
			30305: out = 16'(125);
			30306: out = 16'(-433);
			30307: out = 16'(-447);
			30308: out = 16'(-373);
			30309: out = 16'(-303);
			30310: out = 16'(343);
			30311: out = 16'(1015);
			30312: out = 16'(981);
			30313: out = 16'(428);
			30314: out = 16'(-549);
			30315: out = 16'(-944);
			30316: out = 16'(-750);
			30317: out = 16'(248);
			30318: out = 16'(-277);
			30319: out = 16'(-723);
			30320: out = 16'(-1692);
			30321: out = 16'(-1668);
			30322: out = 16'(-1506);
			30323: out = 16'(-968);
			30324: out = 16'(-278);
			30325: out = 16'(700);
			30326: out = 16'(1987);
			30327: out = 16'(2783);
			30328: out = 16'(3085);
			30329: out = 16'(1174);
			30330: out = 16'(565);
			30331: out = 16'(22);
			30332: out = 16'(348);
			30333: out = 16'(-15);
			30334: out = 16'(-328);
			30335: out = 16'(-1471);
			30336: out = 16'(-1800);
			30337: out = 16'(-1737);
			30338: out = 16'(-394);
			30339: out = 16'(235);
			30340: out = 16'(-254);
			30341: out = 16'(-223);
			30342: out = 16'(-177);
			30343: out = 16'(-316);
			30344: out = 16'(777);
			30345: out = 16'(1646);
			30346: out = 16'(1562);
			30347: out = 16'(362);
			30348: out = 16'(-1554);
			30349: out = 16'(-3818);
			30350: out = 16'(-4135);
			30351: out = 16'(-2477);
			30352: out = 16'(-1636);
			30353: out = 16'(187);
			30354: out = 16'(992);
			30355: out = 16'(3732);
			30356: out = 16'(4030);
			30357: out = 16'(3306);
			30358: out = 16'(741);
			30359: out = 16'(-696);
			30360: out = 16'(-414);
			30361: out = 16'(-338);
			30362: out = 16'(-183);
			30363: out = 16'(1032);
			30364: out = 16'(-186);
			30365: out = 16'(-1088);
			30366: out = 16'(-1310);
			30367: out = 16'(1105);
			30368: out = 16'(3974);
			30369: out = 16'(4024);
			30370: out = 16'(2725);
			30371: out = 16'(-201);
			30372: out = 16'(-245);
			30373: out = 16'(-1328);
			30374: out = 16'(-2587);
			30375: out = 16'(-1987);
			30376: out = 16'(-2004);
			30377: out = 16'(-2285);
			30378: out = 16'(-4166);
			30379: out = 16'(-4590);
			30380: out = 16'(-1650);
			30381: out = 16'(-412);
			30382: out = 16'(858);
			30383: out = 16'(1587);
			30384: out = 16'(1178);
			30385: out = 16'(309);
			30386: out = 16'(-168);
			30387: out = 16'(-274);
			30388: out = 16'(-127);
			30389: out = 16'(-41);
			30390: out = 16'(-834);
			30391: out = 16'(-2269);
			30392: out = 16'(-3252);
			30393: out = 16'(-2652);
			30394: out = 16'(233);
			30395: out = 16'(1050);
			30396: out = 16'(2392);
			30397: out = 16'(3216);
			30398: out = 16'(3493);
			30399: out = 16'(2680);
			30400: out = 16'(-15);
			30401: out = 16'(-60);
			30402: out = 16'(262);
			30403: out = 16'(-251);
			30404: out = 16'(-173);
			30405: out = 16'(-256);
			30406: out = 16'(243);
			30407: out = 16'(-277);
			30408: out = 16'(-1123);
			30409: out = 16'(-963);
			30410: out = 16'(-1032);
			30411: out = 16'(-941);
			30412: out = 16'(-1015);
			30413: out = 16'(-695);
			30414: out = 16'(-105);
			30415: out = 16'(-196);
			30416: out = 16'(-531);
			30417: out = 16'(-1565);
			30418: out = 16'(-1174);
			30419: out = 16'(-1075);
			30420: out = 16'(-3444);
			30421: out = 16'(-2484);
			30422: out = 16'(-901);
			30423: out = 16'(1930);
			30424: out = 16'(2798);
			30425: out = 16'(2723);
			30426: out = 16'(517);
			30427: out = 16'(-240);
			30428: out = 16'(-66);
			30429: out = 16'(161);
			30430: out = 16'(618);
			30431: out = 16'(473);
			30432: out = 16'(1097);
			30433: out = 16'(964);
			30434: out = 16'(636);
			30435: out = 16'(-35);
			30436: out = 16'(-140);
			30437: out = 16'(200);
			30438: out = 16'(1987);
			30439: out = 16'(3432);
			30440: out = 16'(2040);
			30441: out = 16'(2420);
			30442: out = 16'(2588);
			30443: out = 16'(3108);
			30444: out = 16'(1934);
			30445: out = 16'(-317);
			30446: out = 16'(279);
			30447: out = 16'(-991);
			30448: out = 16'(-2459);
			30449: out = 16'(-4976);
			30450: out = 16'(-5625);
			30451: out = 16'(-4224);
			30452: out = 16'(-1798);
			30453: out = 16'(288);
			30454: out = 16'(-386);
			30455: out = 16'(1827);
			30456: out = 16'(2735);
			30457: out = 16'(1737);
			30458: out = 16'(700);
			30459: out = 16'(-700);
			30460: out = 16'(-1239);
			30461: out = 16'(-2836);
			30462: out = 16'(-4104);
			30463: out = 16'(-459);
			30464: out = 16'(1680);
			30465: out = 16'(3405);
			30466: out = 16'(2101);
			30467: out = 16'(1043);
			30468: out = 16'(-173);
			30469: out = 16'(-174);
			30470: out = 16'(-56);
			30471: out = 16'(279);
			30472: out = 16'(231);
			30473: out = 16'(250);
			30474: out = 16'(251);
			30475: out = 16'(50);
			30476: out = 16'(-229);
			30477: out = 16'(-172);
			30478: out = 16'(60);
			30479: out = 16'(534);
			30480: out = 16'(859);
			30481: out = 16'(865);
			30482: out = 16'(208);
			30483: out = 16'(44);
			30484: out = 16'(-472);
			30485: out = 16'(-269);
			30486: out = 16'(-3370);
			30487: out = 16'(-4402);
			30488: out = 16'(-4235);
			30489: out = 16'(-1605);
			30490: out = 16'(180);
			30491: out = 16'(-311);
			30492: out = 16'(-48);
			30493: out = 16'(-41);
			30494: out = 16'(1249);
			30495: out = 16'(894);
			30496: out = 16'(589);
			30497: out = 16'(461);
			30498: out = 16'(459);
			30499: out = 16'(675);
			30500: out = 16'(904);
			30501: out = 16'(1992);
			30502: out = 16'(3335);
			30503: out = 16'(3361);
			30504: out = 16'(1766);
			30505: out = 16'(-2604);
			30506: out = 16'(-464);
			30507: out = 16'(637);
			30508: out = 16'(2151);
			30509: out = 16'(474);
			30510: out = 16'(-868);
			30511: out = 16'(-1672);
			30512: out = 16'(-1056);
			30513: out = 16'(238);
			30514: out = 16'(2212);
			30515: out = 16'(3038);
			30516: out = 16'(2746);
			30517: out = 16'(803);
			30518: out = 16'(-1295);
			30519: out = 16'(-3306);
			30520: out = 16'(-3124);
			30521: out = 16'(-3074);
			30522: out = 16'(-3049);
			30523: out = 16'(-1990);
			30524: out = 16'(-1420);
			30525: out = 16'(-874);
			30526: out = 16'(-1838);
			30527: out = 16'(-1822);
			30528: out = 16'(-25);
			30529: out = 16'(253);
			30530: out = 16'(42);
			30531: out = 16'(-2711);
			30532: out = 16'(-1838);
			30533: out = 16'(-438);
			30534: out = 16'(-235);
			30535: out = 16'(997);
			30536: out = 16'(1874);
			30537: out = 16'(2865);
			30538: out = 16'(1798);
			30539: out = 16'(-259);
			30540: out = 16'(-634);
			30541: out = 16'(-733);
			30542: out = 16'(33);
			30543: out = 16'(344);
			30544: out = 16'(329);
			30545: out = 16'(-959);
			30546: out = 16'(-1211);
			30547: out = 16'(-1326);
			30548: out = 16'(516);
			30549: out = 16'(-70);
			30550: out = 16'(-98);
			30551: out = 16'(-421);
			30552: out = 16'(1623);
			30553: out = 16'(3607);
			30554: out = 16'(2754);
			30555: out = 16'(1947);
			30556: out = 16'(47);
			30557: out = 16'(204);
			30558: out = 16'(-965);
			30559: out = 16'(-1524);
			30560: out = 16'(-4317);
			30561: out = 16'(-4431);
			30562: out = 16'(-2745);
			30563: out = 16'(-881);
			30564: out = 16'(812);
			30565: out = 16'(2982);
			30566: out = 16'(1513);
			30567: out = 16'(22);
			30568: out = 16'(-2755);
			30569: out = 16'(-951);
			30570: out = 16'(1097);
			30571: out = 16'(2708);
			30572: out = 16'(1908);
			30573: out = 16'(305);
			30574: out = 16'(50);
			30575: out = 16'(305);
			30576: out = 16'(1250);
			30577: out = 16'(1993);
			30578: out = 16'(1884);
			30579: out = 16'(918);
			30580: out = 16'(-836);
			30581: out = 16'(-2146);
			30582: out = 16'(-2913);
			30583: out = 16'(-1614);
			30584: out = 16'(-647);
			30585: out = 16'(-245);
			30586: out = 16'(-1323);
			30587: out = 16'(-2022);
			30588: out = 16'(-294);
			30589: out = 16'(1077);
			30590: out = 16'(2556);
			30591: out = 16'(1650);
			30592: out = 16'(1800);
			30593: out = 16'(1608);
			30594: out = 16'(2679);
			30595: out = 16'(2112);
			30596: out = 16'(787);
			30597: out = 16'(-6);
			30598: out = 16'(-542);
			30599: out = 16'(405);
			30600: out = 16'(-3208);
			30601: out = 16'(-4512);
			30602: out = 16'(-4331);
			30603: out = 16'(-893);
			30604: out = 16'(1927);
			30605: out = 16'(2570);
			30606: out = 16'(2422);
			30607: out = 16'(1171);
			30608: out = 16'(228);
			30609: out = 16'(-1283);
			30610: out = 16'(-2072);
			30611: out = 16'(-40);
			30612: out = 16'(994);
			30613: out = 16'(1676);
			30614: out = 16'(186);
			30615: out = 16'(-230);
			30616: out = 16'(-294);
			30617: out = 16'(-162);
			30618: out = 16'(-137);
			30619: out = 16'(-299);
			30620: out = 16'(-731);
			30621: out = 16'(-788);
			30622: out = 16'(-49);
			30623: out = 16'(-83);
			30624: out = 16'(-271);
			30625: out = 16'(-1419);
			30626: out = 16'(-2504);
			30627: out = 16'(-3311);
			30628: out = 16'(262);
			30629: out = 16'(734);
			30630: out = 16'(1346);
			30631: out = 16'(-1288);
			30632: out = 16'(-528);
			30633: out = 16'(660);
			30634: out = 16'(2643);
			30635: out = 16'(1777);
			30636: out = 16'(-934);
			30637: out = 16'(-2802);
			30638: out = 16'(-2703);
			30639: out = 16'(623);
			30640: out = 16'(923);
			30641: out = 16'(1116);
			30642: out = 16'(26);
			30643: out = 16'(-392);
			30644: out = 16'(-966);
			30645: out = 16'(-2034);
			30646: out = 16'(-701);
			30647: out = 16'(1064);
			30648: out = 16'(2637);
			30649: out = 16'(2353);
			30650: out = 16'(918);
			30651: out = 16'(293);
			30652: out = 16'(-30);
			30653: out = 16'(449);
			30654: out = 16'(-1123);
			30655: out = 16'(-1418);
			30656: out = 16'(-706);
			30657: out = 16'(-1744);
			30658: out = 16'(-2167);
			30659: out = 16'(-2814);
			30660: out = 16'(-525);
			30661: out = 16'(1182);
			30662: out = 16'(2394);
			30663: out = 16'(1183);
			30664: out = 16'(36);
			30665: out = 16'(1699);
			30666: out = 16'(2528);
			30667: out = 16'(3324);
			30668: out = 16'(899);
			30669: out = 16'(-319);
			30670: out = 16'(-1652);
			30671: out = 16'(-526);
			30672: out = 16'(24);
			30673: out = 16'(577);
			30674: out = 16'(1314);
			30675: out = 16'(2000);
			30676: out = 16'(2729);
			30677: out = 16'(1246);
			30678: out = 16'(25);
			30679: out = 16'(-74);
			30680: out = 16'(-747);
			30681: out = 16'(-1162);
			30682: out = 16'(-2273);
			30683: out = 16'(-1635);
			30684: out = 16'(-839);
			30685: out = 16'(-1590);
			30686: out = 16'(-969);
			30687: out = 16'(-144);
			30688: out = 16'(-121);
			30689: out = 16'(137);
			30690: out = 16'(408);
			30691: out = 16'(526);
			30692: out = 16'(397);
			30693: out = 16'(-142);
			30694: out = 16'(-126);
			30695: out = 16'(-398);
			30696: out = 16'(-166);
			30697: out = 16'(-1511);
			30698: out = 16'(-2342);
			30699: out = 16'(-2817);
			30700: out = 16'(-1429);
			30701: out = 16'(468);
			30702: out = 16'(2582);
			30703: out = 16'(3062);
			30704: out = 16'(2593);
			30705: out = 16'(1490);
			30706: out = 16'(180);
			30707: out = 16'(-977);
			30708: out = 16'(233);
			30709: out = 16'(711);
			30710: out = 16'(1067);
			30711: out = 16'(145);
			30712: out = 16'(-241);
			30713: out = 16'(-116);
			30714: out = 16'(117);
			30715: out = 16'(97);
			30716: out = 16'(-1033);
			30717: out = 16'(-532);
			30718: out = 16'(-319);
			30719: out = 16'(-300);
			30720: out = 16'(-337);
			30721: out = 16'(-193);
			30722: out = 16'(427);
			30723: out = 16'(284);
			30724: out = 16'(-251);
			30725: out = 16'(-104);
			30726: out = 16'(-882);
			30727: out = 16'(-1532);
			30728: out = 16'(-2136);
			30729: out = 16'(-1386);
			30730: out = 16'(514);
			30731: out = 16'(541);
			30732: out = 16'(468);
			30733: out = 16'(-56);
			30734: out = 16'(698);
			30735: out = 16'(1130);
			30736: out = 16'(-243);
			30737: out = 16'(763);
			30738: out = 16'(920);
			30739: out = 16'(824);
			30740: out = 16'(-1572);
			30741: out = 16'(-3604);
			30742: out = 16'(-2424);
			30743: out = 16'(-2);
			30744: out = 16'(3189);
			30745: out = 16'(1343);
			30746: out = 16'(711);
			30747: out = 16'(-352);
			30748: out = 16'(-86);
			30749: out = 16'(100);
			30750: out = 16'(506);
			30751: out = 16'(1754);
			30752: out = 16'(1838);
			30753: out = 16'(-173);
			30754: out = 16'(-1679);
			30755: out = 16'(-3062);
			30756: out = 16'(-1271);
			30757: out = 16'(-2401);
			30758: out = 16'(-2528);
			30759: out = 16'(-1714);
			30760: out = 16'(-15);
			30761: out = 16'(1305);
			30762: out = 16'(310);
			30763: out = 16'(-737);
			30764: out = 16'(-2082);
			30765: out = 16'(-1502);
			30766: out = 16'(-830);
			30767: out = 16'(226);
			30768: out = 16'(497);
			30769: out = 16'(-76);
			30770: out = 16'(-2784);
			30771: out = 16'(-715);
			30772: out = 16'(829);
			30773: out = 16'(3046);
			30774: out = 16'(2067);
			30775: out = 16'(1013);
			30776: out = 16'(7);
			30777: out = 16'(120);
			30778: out = 16'(554);
			30779: out = 16'(39);
			30780: out = 16'(6);
			30781: out = 16'(-184);
			30782: out = 16'(-142);
			30783: out = 16'(100);
			30784: out = 16'(758);
			30785: out = 16'(57);
			30786: out = 16'(246);
			30787: out = 16'(591);
			30788: out = 16'(1104);
			30789: out = 16'(945);
			30790: out = 16'(-13);
			30791: out = 16'(-40);
			30792: out = 16'(104);
			30793: out = 16'(523);
			30794: out = 16'(305);
			30795: out = 16'(-139);
			30796: out = 16'(715);
			30797: out = 16'(-474);
			30798: out = 16'(-1522);
			30799: out = 16'(-2647);
			30800: out = 16'(-1104);
			30801: out = 16'(1479);
			30802: out = 16'(1081);
			30803: out = 16'(851);
			30804: out = 16'(-309);
			30805: out = 16'(72);
			30806: out = 16'(35);
			30807: out = 16'(494);
			30808: out = 16'(-73);
			30809: out = 16'(-43);
			30810: out = 16'(593);
			30811: out = 16'(194);
			30812: out = 16'(15);
			30813: out = 16'(376);
			30814: out = 16'(484);
			30815: out = 16'(386);
			30816: out = 16'(-1191);
			30817: out = 16'(-2024);
			30818: out = 16'(-2557);
			30819: out = 16'(10);
			30820: out = 16'(658);
			30821: out = 16'(595);
			30822: out = 16'(529);
			30823: out = 16'(366);
			30824: out = 16'(473);
			30825: out = 16'(357);
			30826: out = 16'(395);
			30827: out = 16'(-85);
			30828: out = 16'(792);
			30829: out = 16'(1054);
			30830: out = 16'(591);
			30831: out = 16'(111);
			30832: out = 16'(-422);
			30833: out = 16'(-1370);
			30834: out = 16'(-1400);
			30835: out = 16'(-1360);
			30836: out = 16'(-194);
			30837: out = 16'(-451);
			30838: out = 16'(-666);
			30839: out = 16'(-900);
			30840: out = 16'(261);
			30841: out = 16'(1823);
			30842: out = 16'(3001);
			30843: out = 16'(2842);
			30844: out = 16'(1611);
			30845: out = 16'(-521);
			30846: out = 16'(-1474);
			30847: out = 16'(-195);
			30848: out = 16'(1125);
			30849: out = 16'(2251);
			30850: out = 16'(859);
			30851: out = 16'(769);
			30852: out = 16'(78);
			30853: out = 16'(1139);
			30854: out = 16'(-27);
			30855: out = 16'(-1174);
			30856: out = 16'(-3120);
			30857: out = 16'(-3287);
			30858: out = 16'(-2562);
			30859: out = 16'(-1788);
			30860: out = 16'(-634);
			30861: out = 16'(692);
			30862: out = 16'(940);
			30863: out = 16'(1519);
			30864: out = 16'(2137);
			30865: out = 16'(2631);
			30866: out = 16'(1830);
			30867: out = 16'(-2140);
			30868: out = 16'(-2124);
			30869: out = 16'(-1678);
			30870: out = 16'(1579);
			30871: out = 16'(1042);
			30872: out = 16'(286);
			30873: out = 16'(-1785);
			30874: out = 16'(-2027);
			30875: out = 16'(-1856);
			30876: out = 16'(749);
			30877: out = 16'(1214);
			30878: out = 16'(1101);
			30879: out = 16'(-2755);
			30880: out = 16'(-3972);
			30881: out = 16'(-2989);
			30882: out = 16'(-238);
			30883: out = 16'(2226);
			30884: out = 16'(3137);
			30885: out = 16'(2951);
			30886: out = 16'(1652);
			30887: out = 16'(759);
			30888: out = 16'(-1423);
			30889: out = 16'(-2740);
			30890: out = 16'(-2599);
			30891: out = 16'(-1977);
			30892: out = 16'(-1096);
			30893: out = 16'(-765);
			30894: out = 16'(-334);
			30895: out = 16'(62);
			30896: out = 16'(564);
			30897: out = 16'(1281);
			30898: out = 16'(2420);
			30899: out = 16'(1901);
			30900: out = 16'(1614);
			30901: out = 16'(1127);
			30902: out = 16'(1542);
			30903: out = 16'(1493);
			30904: out = 16'(505);
			30905: out = 16'(455);
			30906: out = 16'(224);
			30907: out = 16'(19);
			30908: out = 16'(-496);
			30909: out = 16'(-801);
			30910: out = 16'(-159);
			30911: out = 16'(419);
			30912: out = 16'(1106);
			30913: out = 16'(-608);
			30914: out = 16'(-518);
			30915: out = 16'(455);
			30916: out = 16'(-21);
			30917: out = 16'(-203);
			30918: out = 16'(-964);
			30919: out = 16'(222);
			30920: out = 16'(401);
			30921: out = 16'(-13);
			30922: out = 16'(-953);
			30923: out = 16'(-1245);
			30924: out = 16'(343);
			30925: out = 16'(356);
			30926: out = 16'(319);
			30927: out = 16'(29);
			30928: out = 16'(-103);
			30929: out = 16'(-122);
			30930: out = 16'(-1774);
			30931: out = 16'(-2236);
			30932: out = 16'(-2640);
			30933: out = 16'(-490);
			30934: out = 16'(-259);
			30935: out = 16'(-621);
			30936: out = 16'(-1276);
			30937: out = 16'(-306);
			30938: out = 16'(2368);
			30939: out = 16'(3359);
			30940: out = 16'(3495);
			30941: out = 16'(1647);
			30942: out = 16'(923);
			30943: out = 16'(173);
			30944: out = 16'(347);
			30945: out = 16'(391);
			30946: out = 16'(388);
			30947: out = 16'(-123);
			30948: out = 16'(-1127);
			30949: out = 16'(-2155);
			30950: out = 16'(-2111);
			30951: out = 16'(-1285);
			30952: out = 16'(161);
			30953: out = 16'(2039);
			30954: out = 16'(2900);
			30955: out = 16'(2533);
			30956: out = 16'(1556);
			30957: out = 16'(615);
			30958: out = 16'(465);
			30959: out = 16'(157);
			30960: out = 16'(190);
			30961: out = 16'(76);
			30962: out = 16'(218);
			30963: out = 16'(-310);
			30964: out = 16'(-3206);
			30965: out = 16'(-3938);
			30966: out = 16'(-3809);
			30967: out = 16'(-137);
			30968: out = 16'(1314);
			30969: out = 16'(2159);
			30970: out = 16'(276);
			30971: out = 16'(-188);
			30972: out = 16'(-113);
			30973: out = 16'(1156);
			30974: out = 16'(1509);
			30975: out = 16'(926);
			30976: out = 16'(138);
			30977: out = 16'(-628);
			30978: out = 16'(-899);
			30979: out = 16'(-217);
			30980: out = 16'(742);
			30981: out = 16'(1346);
			30982: out = 16'(1352);
			30983: out = 16'(773);
			30984: out = 16'(1607);
			30985: out = 16'(738);
			30986: out = 16'(-94);
			30987: out = 16'(-3648);
			30988: out = 16'(-4312);
			30989: out = 16'(-4036);
			30990: out = 16'(-1106);
			30991: out = 16'(179);
			30992: out = 16'(529);
			30993: out = 16'(56);
			30994: out = 16'(76);
			30995: out = 16'(279);
			30996: out = 16'(1240);
			30997: out = 16'(1681);
			30998: out = 16'(2232);
			30999: out = 16'(640);
			31000: out = 16'(-743);
			31001: out = 16'(-2769);
			31002: out = 16'(-1558);
			31003: out = 16'(-137);
			31004: out = 16'(359);
			31005: out = 16'(-1233);
			31006: out = 16'(-3570);
			31007: out = 16'(-3405);
			31008: out = 16'(-1575);
			31009: out = 16'(2148);
			31010: out = 16'(1997);
			31011: out = 16'(1949);
			31012: out = 16'(198);
			31013: out = 16'(596);
			31014: out = 16'(1082);
			31015: out = 16'(3880);
			31016: out = 16'(2912);
			31017: out = 16'(2026);
			31018: out = 16'(-1664);
			31019: out = 16'(-844);
			31020: out = 16'(-368);
			31021: out = 16'(547);
			31022: out = 16'(-1185);
			31023: out = 16'(-2923);
			31024: out = 16'(-2294);
			31025: out = 16'(-659);
			31026: out = 16'(1896);
			31027: out = 16'(54);
			31028: out = 16'(-69);
			31029: out = 16'(-168);
			31030: out = 16'(-122);
			31031: out = 16'(-787);
			31032: out = 16'(-2135);
			31033: out = 16'(-716);
			31034: out = 16'(143);
			31035: out = 16'(-176);
			31036: out = 16'(329);
			31037: out = 16'(334);
			31038: out = 16'(632);
			31039: out = 16'(84);
			31040: out = 16'(-283);
			31041: out = 16'(-881);
			31042: out = 16'(-176);
			31043: out = 16'(606);
			31044: out = 16'(574);
			31045: out = 16'(41);
			31046: out = 16'(-893);
			31047: out = 16'(-218);
			31048: out = 16'(481);
			31049: out = 16'(1731);
			31050: out = 16'(1199);
			31051: out = 16'(789);
			31052: out = 16'(-173);
			31053: out = 16'(288);
			31054: out = 16'(368);
			31055: out = 16'(-136);
			31056: out = 16'(-118);
			31057: out = 16'(-141);
			31058: out = 16'(-224);
			31059: out = 16'(-594);
			31060: out = 16'(-793);
			31061: out = 16'(386);
			31062: out = 16'(490);
			31063: out = 16'(273);
			31064: out = 16'(337);
			31065: out = 16'(494);
			31066: out = 16'(1131);
			31067: out = 16'(28);
			31068: out = 16'(-78);
			31069: out = 16'(-226);
			31070: out = 16'(2167);
			31071: out = 16'(3148);
			31072: out = 16'(2458);
			31073: out = 16'(1172);
			31074: out = 16'(-439);
			31075: out = 16'(-1449);
			31076: out = 16'(-1854);
			31077: out = 16'(-1346);
			31078: out = 16'(-464);
			31079: out = 16'(426);
			31080: out = 16'(888);
			31081: out = 16'(349);
			31082: out = 16'(-134);
			31083: out = 16'(-424);
			31084: out = 16'(-879);
			31085: out = 16'(-1331);
			31086: out = 16'(-2262);
			31087: out = 16'(-376);
			31088: out = 16'(779);
			31089: out = 16'(2159);
			31090: out = 16'(526);
			31091: out = 16'(-213);
			31092: out = 16'(187);
			31093: out = 16'(976);
			31094: out = 16'(1345);
			31095: out = 16'(-151);
			31096: out = 16'(-902);
			31097: out = 16'(-1701);
			31098: out = 16'(-991);
			31099: out = 16'(-762);
			31100: out = 16'(-298);
			31101: out = 16'(-1425);
			31102: out = 16'(-1343);
			31103: out = 16'(-818);
			31104: out = 16'(-25);
			31105: out = 16'(445);
			31106: out = 16'(195);
			31107: out = 16'(1628);
			31108: out = 16'(2220);
			31109: out = 16'(2612);
			31110: out = 16'(1100);
			31111: out = 16'(-209);
			31112: out = 16'(-941);
			31113: out = 16'(-647);
			31114: out = 16'(-146);
			31115: out = 16'(-272);
			31116: out = 16'(-251);
			31117: out = 16'(-502);
			31118: out = 16'(-1428);
			31119: out = 16'(-1409);
			31120: out = 16'(-788);
			31121: out = 16'(116);
			31122: out = 16'(577);
			31123: out = 16'(293);
			31124: out = 16'(-389);
			31125: out = 16'(-1463);
			31126: out = 16'(-1930);
			31127: out = 16'(-3132);
			31128: out = 16'(-2710);
			31129: out = 16'(-309);
			31130: out = 16'(1617);
			31131: out = 16'(2662);
			31132: out = 16'(-87);
			31133: out = 16'(329);
			31134: out = 16'(588);
			31135: out = 16'(2099);
			31136: out = 16'(1404);
			31137: out = 16'(285);
			31138: out = 16'(-117);
			31139: out = 16'(-815);
			31140: out = 16'(-1551);
			31141: out = 16'(-576);
			31142: out = 16'(115);
			31143: out = 16'(1117);
			31144: out = 16'(519);
			31145: out = 16'(474);
			31146: out = 16'(119);
			31147: out = 16'(1782);
			31148: out = 16'(2734);
			31149: out = 16'(3049);
			31150: out = 16'(1204);
			31151: out = 16'(-673);
			31152: out = 16'(-270);
			31153: out = 16'(-957);
			31154: out = 16'(-859);
			31155: out = 16'(512);
			31156: out = 16'(1412);
			31157: out = 16'(1752);
			31158: out = 16'(-899);
			31159: out = 16'(-2802);
			31160: out = 16'(-4232);
			31161: out = 16'(-3291);
			31162: out = 16'(-2168);
			31163: out = 16'(-904);
			31164: out = 16'(451);
			31165: out = 16'(1289);
			31166: out = 16'(1534);
			31167: out = 16'(563);
			31168: out = 16'(-545);
			31169: out = 16'(496);
			31170: out = 16'(-564);
			31171: out = 16'(-904);
			31172: out = 16'(-2318);
			31173: out = 16'(128);
			31174: out = 16'(3026);
			31175: out = 16'(3834);
			31176: out = 16'(2805);
			31177: out = 16'(-38);
			31178: out = 16'(1387);
			31179: out = 16'(1559);
			31180: out = 16'(2588);
			31181: out = 16'(258);
			31182: out = 16'(-626);
			31183: out = 16'(-1196);
			31184: out = 16'(-1071);
			31185: out = 16'(-1425);
			31186: out = 16'(-2194);
			31187: out = 16'(-2455);
			31188: out = 16'(-1703);
			31189: out = 16'(558);
			31190: out = 16'(2140);
			31191: out = 16'(3015);
			31192: out = 16'(2623);
			31193: out = 16'(1165);
			31194: out = 16'(-864);
			31195: out = 16'(-2461);
			31196: out = 16'(-3165);
			31197: out = 16'(-2768);
			31198: out = 16'(-1559);
			31199: out = 16'(-739);
			31200: out = 16'(-1107);
			31201: out = 16'(4);
			31202: out = 16'(176);
			31203: out = 16'(-87);
			31204: out = 16'(-297);
			31205: out = 16'(-241);
			31206: out = 16'(-200);
			31207: out = 16'(504);
			31208: out = 16'(974);
			31209: out = 16'(-129);
			31210: out = 16'(34);
			31211: out = 16'(260);
			31212: out = 16'(196);
			31213: out = 16'(337);
			31214: out = 16'(390);
			31215: out = 16'(871);
			31216: out = 16'(623);
			31217: out = 16'(-328);
			31218: out = 16'(280);
			31219: out = 16'(191);
			31220: out = 16'(-214);
			31221: out = 16'(-760);
			31222: out = 16'(-701);
			31223: out = 16'(997);
			31224: out = 16'(560);
			31225: out = 16'(105);
			31226: out = 16'(-1557);
			31227: out = 16'(-1297);
			31228: out = 16'(-961);
			31229: out = 16'(-934);
			31230: out = 16'(-1236);
			31231: out = 16'(-1445);
			31232: out = 16'(-30);
			31233: out = 16'(504);
			31234: out = 16'(344);
			31235: out = 16'(109);
			31236: out = 16'(-1338);
			31237: out = 16'(-3354);
			31238: out = 16'(-4355);
			31239: out = 16'(-3510);
			31240: out = 16'(619);
			31241: out = 16'(1242);
			31242: out = 16'(1659);
			31243: out = 16'(-877);
			31244: out = 16'(196);
			31245: out = 16'(998);
			31246: out = 16'(4166);
			31247: out = 16'(3422);
			31248: out = 16'(2552);
			31249: out = 16'(1050);
			31250: out = 16'(1682);
			31251: out = 16'(2538);
			31252: out = 16'(3503);
			31253: out = 16'(2294);
			31254: out = 16'(-143);
			31255: out = 16'(-3207);
			31256: out = 16'(-4118);
			31257: out = 16'(-2022);
			31258: out = 16'(-1197);
			31259: out = 16'(39);
			31260: out = 16'(42);
			31261: out = 16'(463);
			31262: out = 16'(523);
			31263: out = 16'(2042);
			31264: out = 16'(2207);
			31265: out = 16'(2351);
			31266: out = 16'(-216);
			31267: out = 16'(-298);
			31268: out = 16'(-607);
			31269: out = 16'(391);
			31270: out = 16'(-574);
			31271: out = 16'(-1708);
			31272: out = 16'(-2805);
			31273: out = 16'(-1883);
			31274: out = 16'(524);
			31275: out = 16'(783);
			31276: out = 16'(678);
			31277: out = 16'(-415);
			31278: out = 16'(-1181);
			31279: out = 16'(-1378);
			31280: out = 16'(250);
			31281: out = 16'(224);
			31282: out = 16'(23);
			31283: out = 16'(-1472);
			31284: out = 16'(-1313);
			31285: out = 16'(-598);
			31286: out = 16'(611);
			31287: out = 16'(2283);
			31288: out = 16'(3641);
			31289: out = 16'(3220);
			31290: out = 16'(1767);
			31291: out = 16'(-726);
			31292: out = 16'(-296);
			31293: out = 16'(-96);
			31294: out = 16'(908);
			31295: out = 16'(-503);
			31296: out = 16'(-1747);
			31297: out = 16'(-3569);
			31298: out = 16'(-3221);
			31299: out = 16'(-2359);
			31300: out = 16'(-450);
			31301: out = 16'(-154);
			31302: out = 16'(75);
			31303: out = 16'(2004);
			31304: out = 16'(1840);
			31305: out = 16'(1425);
			31306: out = 16'(468);
			31307: out = 16'(376);
			31308: out = 16'(239);
			31309: out = 16'(-68);
			31310: out = 16'(-1540);
			31311: out = 16'(-3544);
			31312: out = 16'(-3099);
			31313: out = 16'(-1957);
			31314: out = 16'(-107);
			31315: out = 16'(1149);
			31316: out = 16'(1363);
			31317: out = 16'(-65);
			31318: out = 16'(-584);
			31319: out = 16'(-683);
			31320: out = 16'(336);
			31321: out = 16'(1691);
			31322: out = 16'(2662);
			31323: out = 16'(1730);
			31324: out = 16'(196);
			31325: out = 16'(-1735);
			31326: out = 16'(-992);
			31327: out = 16'(102);
			31328: out = 16'(2346);
			31329: out = 16'(616);
			31330: out = 16'(102);
			31331: out = 16'(-1119);
			31332: out = 16'(-228);
			31333: out = 16'(-298);
			31334: out = 16'(-154);
			31335: out = 16'(-2377);
			31336: out = 16'(-3257);
			31337: out = 16'(-1431);
			31338: out = 16'(-683);
			31339: out = 16'(182);
			31340: out = 16'(-302);
			31341: out = 16'(291);
			31342: out = 16'(641);
			31343: out = 16'(1563);
			31344: out = 16'(1648);
			31345: out = 16'(1572);
			31346: out = 16'(707);
			31347: out = 16'(-329);
			31348: out = 16'(-2293);
			31349: out = 16'(-594);
			31350: out = 16'(-118);
			31351: out = 16'(714);
			31352: out = 16'(-2186);
			31353: out = 16'(-3225);
			31354: out = 16'(-1993);
			31355: out = 16'(-99);
			31356: out = 16'(1330);
			31357: out = 16'(-67);
			31358: out = 16'(344);
			31359: out = 16'(420);
			31360: out = 16'(5);
			31361: out = 16'(932);
			31362: out = 16'(2404);
			31363: out = 16'(2095);
			31364: out = 16'(1610);
			31365: out = 16'(22);
			31366: out = 16'(40);
			31367: out = 16'(-727);
			31368: out = 16'(-688);
			31369: out = 16'(-2383);
			31370: out = 16'(-2131);
			31371: out = 16'(-240);
			31372: out = 16'(665);
			31373: out = 16'(1403);
			31374: out = 16'(2742);
			31375: out = 16'(1408);
			31376: out = 16'(321);
			31377: out = 16'(247);
			31378: out = 16'(1361);
			31379: out = 16'(2663);
			31380: out = 16'(1070);
			31381: out = 16'(181);
			31382: out = 16'(-1153);
			31383: out = 16'(221);
			31384: out = 16'(477);
			31385: out = 16'(976);
			31386: out = 16'(-46);
			31387: out = 16'(-141);
			31388: out = 16'(346);
			31389: out = 16'(-82);
			31390: out = 16'(-245);
			31391: out = 16'(237);
			31392: out = 16'(-590);
			31393: out = 16'(-1391);
			31394: out = 16'(-3417);
			31395: out = 16'(-2550);
			31396: out = 16'(-1143);
			31397: out = 16'(5);
			31398: out = 16'(540);
			31399: out = 16'(498);
			31400: out = 16'(2371);
			31401: out = 16'(2596);
			31402: out = 16'(2488);
			31403: out = 16'(805);
			31404: out = 16'(121);
			31405: out = 16'(135);
			31406: out = 16'(-1194);
			31407: out = 16'(-1863);
			31408: out = 16'(-1560);
			31409: out = 16'(-1404);
			31410: out = 16'(-780);
			31411: out = 16'(-1249);
			31412: out = 16'(864);
			31413: out = 16'(2243);
			31414: out = 16'(3059);
			31415: out = 16'(1662);
			31416: out = 16'(-14);
			31417: out = 16'(-912);
			31418: out = 16'(-827);
			31419: out = 16'(-230);
			31420: out = 16'(690);
			31421: out = 16'(234);
			31422: out = 16'(-1209);
			31423: out = 16'(-2039);
			31424: out = 16'(-1700);
			31425: out = 16'(529);
			31426: out = 16'(232);
			31427: out = 16'(292);
			31428: out = 16'(-542);
			31429: out = 16'(12);
			31430: out = 16'(-166);
			31431: out = 16'(-2182);
			31432: out = 16'(-2204);
			31433: out = 16'(-2009);
			31434: out = 16'(186);
			31435: out = 16'(-297);
			31436: out = 16'(-1054);
			31437: out = 16'(-3134);
			31438: out = 16'(-2690);
			31439: out = 16'(-1179);
			31440: out = 16'(584);
			31441: out = 16'(1632);
			31442: out = 16'(2228);
			31443: out = 16'(987);
			31444: out = 16'(-95);
			31445: out = 16'(-2258);
			31446: out = 16'(152);
			31447: out = 16'(1509);
			31448: out = 16'(3406);
			31449: out = 16'(1);
			31450: out = 16'(-2488);
			31451: out = 16'(-2794);
			31452: out = 16'(-3);
			31453: out = 16'(3270);
			31454: out = 16'(3423);
			31455: out = 16'(2464);
			31456: out = 16'(-68);
			31457: out = 16'(121);
			31458: out = 16'(-70);
			31459: out = 16'(1164);
			31460: out = 16'(-173);
			31461: out = 16'(-469);
			31462: out = 16'(-1858);
			31463: out = 16'(-1786);
			31464: out = 16'(-2377);
			31465: out = 16'(-1153);
			31466: out = 16'(-3436);
			31467: out = 16'(-3552);
			31468: out = 16'(-2356);
			31469: out = 16'(924);
			31470: out = 16'(3002);
			31471: out = 16'(2891);
			31472: out = 16'(991);
			31473: out = 16'(-1030);
			31474: out = 16'(-910);
			31475: out = 16'(422);
			31476: out = 16'(2307);
			31477: out = 16'(1798);
			31478: out = 16'(330);
			31479: out = 16'(-2267);
			31480: out = 16'(-2175);
			31481: out = 16'(-1065);
			31482: out = 16'(1748);
			31483: out = 16'(3051);
			31484: out = 16'(3494);
			31485: out = 16'(2024);
			31486: out = 16'(251);
			31487: out = 16'(-1118);
			31488: out = 16'(466);
			31489: out = 16'(1077);
			31490: out = 16'(2042);
			31491: out = 16'(-481);
			31492: out = 16'(-91);
			31493: out = 16'(63);
			31494: out = 16'(421);
			31495: out = 16'(-80);
			31496: out = 16'(-399);
			31497: out = 16'(-426);
			31498: out = 16'(335);
			31499: out = 16'(1424);
			31500: out = 16'(1470);
			31501: out = 16'(867);
			31502: out = 16'(-501);
			31503: out = 16'(-2517);
			31504: out = 16'(-3606);
			31505: out = 16'(-1397);
			31506: out = 16'(-2473);
			31507: out = 16'(-2864);
			31508: out = 16'(-4776);
			31509: out = 16'(-2640);
			31510: out = 16'(-127);
			31511: out = 16'(2866);
			31512: out = 16'(3013);
			31513: out = 16'(1930);
			31514: out = 16'(766);
			31515: out = 16'(-46);
			31516: out = 16'(-172);
			31517: out = 16'(1097);
			31518: out = 16'(2001);
			31519: out = 16'(2571);
			31520: out = 16'(1013);
			31521: out = 16'(-414);
			31522: out = 16'(-1537);
			31523: out = 16'(-925);
			31524: out = 16'(-51);
			31525: out = 16'(274);
			31526: out = 16'(769);
			31527: out = 16'(1052);
			31528: out = 16'(1958);
			31529: out = 16'(1735);
			31530: out = 16'(1275);
			31531: out = 16'(362);
			31532: out = 16'(-857);
			31533: out = 16'(-2486);
			31534: out = 16'(-1076);
			31535: out = 16'(-1831);
			31536: out = 16'(-3554);
			31537: out = 16'(-3021);
			31538: out = 16'(-1611);
			31539: out = 16'(1824);
			31540: out = 16'(300);
			31541: out = 16'(-523);
			31542: out = 16'(-1495);
			31543: out = 16'(-598);
			31544: out = 16'(52);
			31545: out = 16'(-236);
			31546: out = 16'(-455);
			31547: out = 16'(-955);
			31548: out = 16'(-1276);
			31549: out = 16'(-1481);
			31550: out = 16'(-1090);
			31551: out = 16'(638);
			31552: out = 16'(2316);
			31553: out = 16'(3788);
			31554: out = 16'(2546);
			31555: out = 16'(1667);
			31556: out = 16'(1020);
			31557: out = 16'(910);
			31558: out = 16'(1011);
			31559: out = 16'(812);
			31560: out = 16'(1386);
			31561: out = 16'(1159);
			31562: out = 16'(308);
			31563: out = 16'(-999);
			31564: out = 16'(-1568);
			31565: out = 16'(-575);
			31566: out = 16'(306);
			31567: out = 16'(850);
			31568: out = 16'(-36);
			31569: out = 16'(-668);
			31570: out = 16'(-909);
			31571: out = 16'(-1221);
			31572: out = 16'(27);
			31573: out = 16'(1449);
			31574: out = 16'(3283);
			31575: out = 16'(2138);
			31576: out = 16'(-1772);
			31577: out = 16'(-3829);
			31578: out = 16'(-4155);
			31579: out = 16'(408);
			31580: out = 16'(90);
			31581: out = 16'(53);
			31582: out = 16'(-2087);
			31583: out = 16'(-1428);
			31584: out = 16'(-509);
			31585: out = 16'(1247);
			31586: out = 16'(2094);
			31587: out = 16'(2402);
			31588: out = 16'(1233);
			31589: out = 16'(291);
			31590: out = 16'(-377);
			31591: out = 16'(-962);
			31592: out = 16'(-734);
			31593: out = 16'(-462);
			31594: out = 16'(1382);
			31595: out = 16'(1925);
			31596: out = 16'(1978);
			31597: out = 16'(-72);
			31598: out = 16'(-1161);
			31599: out = 16'(-1084);
			31600: out = 16'(382);
			31601: out = 16'(1576);
			31602: out = 16'(2435);
			31603: out = 16'(127);
			31604: out = 16'(-2780);
			31605: out = 16'(-3761);
			31606: out = 16'(-3489);
			31607: out = 16'(-1686);
			31608: out = 16'(-388);
			31609: out = 16'(959);
			31610: out = 16'(1421);
			31611: out = 16'(1165);
			31612: out = 16'(664);
			31613: out = 16'(210);
			31614: out = 16'(-75);
			31615: out = 16'(-182);
			31616: out = 16'(300);
			31617: out = 16'(-1291);
			31618: out = 16'(-2081);
			31619: out = 16'(-926);
			31620: out = 16'(-303);
			31621: out = 16'(376);
			31622: out = 16'(215);
			31623: out = 16'(119);
			31624: out = 16'(-151);
			31625: out = 16'(206);
			31626: out = 16'(515);
			31627: out = 16'(1089);
			31628: out = 16'(2501);
			31629: out = 16'(3076);
			31630: out = 16'(2699);
			31631: out = 16'(1002);
			31632: out = 16'(-871);
			31633: out = 16'(-2096);
			31634: out = 16'(-2421);
			31635: out = 16'(-1903);
			31636: out = 16'(-1791);
			31637: out = 16'(-541);
			31638: out = 16'(-167);
			31639: out = 16'(1169);
			31640: out = 16'(-1360);
			31641: out = 16'(-3513);
			31642: out = 16'(-3411);
			31643: out = 16'(-1156);
			31644: out = 16'(1957);
			31645: out = 16'(409);
			31646: out = 16'(-215);
			31647: out = 16'(-1522);
			31648: out = 16'(178);
			31649: out = 16'(994);
			31650: out = 16'(2151);
			31651: out = 16'(1692);
			31652: out = 16'(1215);
			31653: out = 16'(215);
			31654: out = 16'(-115);
			31655: out = 16'(-350);
			31656: out = 16'(-142);
			31657: out = 16'(140);
			31658: out = 16'(258);
			31659: out = 16'(-1409);
			31660: out = 16'(-1502);
			31661: out = 16'(-1272);
			31662: out = 16'(734);
			31663: out = 16'(865);
			31664: out = 16'(320);
			31665: out = 16'(39);
			31666: out = 16'(95);
			31667: out = 16'(1171);
			31668: out = 16'(223);
			31669: out = 16'(710);
			31670: out = 16'(1321);
			31671: out = 16'(2335);
			31672: out = 16'(1757);
			31673: out = 16'(-262);
			31674: out = 16'(-2336);
			31675: out = 16'(-3519);
			31676: out = 16'(-3461);
			31677: out = 16'(-1417);
			31678: out = 16'(554);
			31679: out = 16'(250);
			31680: out = 16'(-660);
			31681: out = 16'(-2172);
			31682: out = 16'(-897);
			31683: out = 16'(-117);
			31684: out = 16'(1255);
			31685: out = 16'(408);
			31686: out = 16'(234);
			31687: out = 16'(-305);
			31688: out = 16'(748);
			31689: out = 16'(1091);
			31690: out = 16'(965);
			31691: out = 16'(1046);
			31692: out = 16'(800);
			31693: out = 16'(345);
			31694: out = 16'(-798);
			31695: out = 16'(-1523);
			31696: out = 16'(-866);
			31697: out = 16'(-609);
			31698: out = 16'(-157);
			31699: out = 16'(208);
			31700: out = 16'(337);
			31701: out = 16'(218);
			31702: out = 16'(-1186);
			31703: out = 16'(-942);
			31704: out = 16'(577);
			31705: out = 16'(1070);
			31706: out = 16'(2189);
			31707: out = 16'(2878);
			31708: out = 16'(2845);
			31709: out = 16'(1385);
			31710: out = 16'(-1449);
			31711: out = 16'(-2838);
			31712: out = 16'(-2917);
			31713: out = 16'(129);
			31714: out = 16'(686);
			31715: out = 16'(761);
			31716: out = 16'(-1287);
			31717: out = 16'(-2081);
			31718: out = 16'(-2543);
			31719: out = 16'(128);
			31720: out = 16'(969);
			31721: out = 16'(1610);
			31722: out = 16'(595);
			31723: out = 16'(444);
			31724: out = 16'(424);
			31725: out = 16'(1576);
			31726: out = 16'(2188);
			31727: out = 16'(2406);
			31728: out = 16'(1761);
			31729: out = 16'(918);
			31730: out = 16'(-445);
			31731: out = 16'(-198);
			31732: out = 16'(236);
			31733: out = 16'(754);
			31734: out = 16'(235);
			31735: out = 16'(-464);
			31736: out = 16'(-259);
			31737: out = 16'(-161);
			31738: out = 16'(318);
			31739: out = 16'(-449);
			31740: out = 16'(-819);
			31741: out = 16'(-1816);
			31742: out = 16'(-89);
			31743: out = 16'(17);
			31744: out = 16'(269);
			31745: out = 16'(-2132);
			31746: out = 16'(-2652);
			31747: out = 16'(-2239);
			31748: out = 16'(644);
			31749: out = 16'(2007);
			31750: out = 16'(988);
			31751: out = 16'(-1746);
			31752: out = 16'(-4358);
			31753: out = 16'(-2454);
			31754: out = 16'(-2257);
			31755: out = 16'(-1119);
			31756: out = 16'(-3293);
			31757: out = 16'(-1735);
			31758: out = 16'(120);
			31759: out = 16'(1887);
			31760: out = 16'(1978);
			31761: out = 16'(1036);
			31762: out = 16'(1916);
			31763: out = 16'(2412);
			31764: out = 16'(3097);
			31765: out = 16'(1653);
			31766: out = 16'(480);
			31767: out = 16'(-219);
			31768: out = 16'(-1498);
			31769: out = 16'(-2080);
			31770: out = 16'(-1413);
			31771: out = 16'(-1093);
			31772: out = 16'(-700);
			31773: out = 16'(-815);
			31774: out = 16'(-371);
			31775: out = 16'(113);
			31776: out = 16'(390);
			31777: out = 16'(1201);
			31778: out = 16'(2162);
			31779: out = 16'(1721);
			31780: out = 16'(688);
			31781: out = 16'(-1631);
			31782: out = 16'(-27);
			31783: out = 16'(217);
			31784: out = 16'(-20);
			31785: out = 16'(-964);
			31786: out = 16'(-1365);
			31787: out = 16'(-786);
			31788: out = 16'(-333);
			31789: out = 16'(-29);
			31790: out = 16'(-756);
			31791: out = 16'(-464);
			31792: out = 16'(-116);
			31793: out = 16'(-168);
			31794: out = 16'(-794);
			31795: out = 16'(-1978);
			31796: out = 16'(1281);
			31797: out = 16'(1603);
			31798: out = 16'(1721);
			31799: out = 16'(-2185);
			31800: out = 16'(-2538);
			31801: out = 16'(45);
			31802: out = 16'(1710);
			31803: out = 16'(2851);
			31804: out = 16'(1893);
			31805: out = 16'(2521);
			31806: out = 16'(2250);
			31807: out = 16'(1010);
			31808: out = 16'(632);
			31809: out = 16'(218);
			31810: out = 16'(567);
			31811: out = 16'(-1362);
			31812: out = 16'(-3589);
			31813: out = 16'(-3242);
			31814: out = 16'(-2417);
			31815: out = 16'(-483);
			31816: out = 16'(-484);
			31817: out = 16'(93);
			31818: out = 16'(-127);
			31819: out = 16'(934);
			31820: out = 16'(923);
			31821: out = 16'(392);
			31822: out = 16'(433);
			31823: out = 16'(491);
			31824: out = 16'(-124);
			31825: out = 16'(259);
			31826: out = 16'(341);
			31827: out = 16'(1133);
			31828: out = 16'(320);
			31829: out = 16'(-341);
			31830: out = 16'(-1421);
			31831: out = 16'(-553);
			31832: out = 16'(607);
			31833: out = 16'(1441);
			31834: out = 16'(977);
			31835: out = 16'(-183);
			31836: out = 16'(-674);
			31837: out = 16'(-637);
			31838: out = 16'(-107);
			31839: out = 16'(1087);
			31840: out = 16'(1225);
			31841: out = 16'(-78);
			31842: out = 16'(-1305);
			31843: out = 16'(-1829);
			31844: out = 16'(248);
			31845: out = 16'(949);
			31846: out = 16'(1712);
			31847: out = 16'(2456);
			31848: out = 16'(1579);
			31849: out = 16'(80);
			31850: out = 16'(-148);
			31851: out = 16'(-415);
			31852: out = 16'(-141);
			31853: out = 16'(-786);
			31854: out = 16'(-1519);
			31855: out = 16'(-2846);
			31856: out = 16'(-2236);
			31857: out = 16'(-1626);
			31858: out = 16'(-204);
			31859: out = 16'(82);
			31860: out = 16'(67);
			31861: out = 16'(-2141);
			31862: out = 16'(-769);
			31863: out = 16'(276);
			31864: out = 16'(2114);
			31865: out = 16'(672);
			31866: out = 16'(-1035);
			31867: out = 16'(-219);
			31868: out = 16'(231);
			31869: out = 16'(1145);
			31870: out = 16'(-623);
			31871: out = 16'(-1021);
			31872: out = 16'(-1464);
			31873: out = 16'(564);
			31874: out = 16'(1277);
			31875: out = 16'(1590);
			31876: out = 16'(357);
			31877: out = 16'(-99);
			31878: out = 16'(312);
			31879: out = 16'(698);
			31880: out = 16'(1097);
			31881: out = 16'(1494);
			31882: out = 16'(596);
			31883: out = 16'(-342);
			31884: out = 16'(320);
			31885: out = 16'(-416);
			31886: out = 16'(-951);
			31887: out = 16'(-435);
			31888: out = 16'(-231);
			31889: out = 16'(-156);
			31890: out = 16'(-314);
			31891: out = 16'(-87);
			31892: out = 16'(454);
			31893: out = 16'(1);
			31894: out = 16'(-750);
			31895: out = 16'(-2830);
			31896: out = 16'(-1372);
			31897: out = 16'(-445);
			31898: out = 16'(1147);
			31899: out = 16'(-463);
			31900: out = 16'(-1593);
			31901: out = 16'(-1972);
			31902: out = 16'(-785);
			31903: out = 16'(653);
			31904: out = 16'(424);
			31905: out = 16'(868);
			31906: out = 16'(1039);
			31907: out = 16'(496);
			31908: out = 16'(-94);
			31909: out = 16'(-917);
			31910: out = 16'(-199);
			31911: out = 16'(-794);
			31912: out = 16'(-1940);
			31913: out = 16'(-2077);
			31914: out = 16'(-765);
			31915: out = 16'(2801);
			31916: out = 16'(2663);
			31917: out = 16'(2284);
			31918: out = 16'(497);
			31919: out = 16'(93);
			31920: out = 16'(-277);
			31921: out = 16'(483);
			31922: out = 16'(654);
			31923: out = 16'(1090);
			31924: out = 16'(882);
			31925: out = 16'(812);
			31926: out = 16'(262);
			31927: out = 16'(994);
			31928: out = 16'(423);
			31929: out = 16'(-212);
			31930: out = 16'(-2165);
			31931: out = 16'(-2813);
			31932: out = 16'(-2655);
			31933: out = 16'(-473);
			31934: out = 16'(771);
			31935: out = 16'(360);
			31936: out = 16'(244);
			31937: out = 16'(-60);
			31938: out = 16'(1140);
			31939: out = 16'(343);
			31940: out = 16'(-250);
			31941: out = 16'(-1364);
			31942: out = 16'(-1144);
			31943: out = 16'(-740);
			31944: out = 16'(-311);
			31945: out = 16'(0);
			31946: out = 16'(408);
			31947: out = 16'(-185);
			31948: out = 16'(-104);
			31949: out = 16'(-91);
			31950: out = 16'(79);
			31951: out = 16'(-593);
			31952: out = 16'(-1907);
			31953: out = 16'(-2435);
			31954: out = 16'(-1970);
			31955: out = 16'(39);
			31956: out = 16'(1645);
			31957: out = 16'(3004);
			31958: out = 16'(2495);
			31959: out = 16'(2779);
			31960: out = 16'(2333);
			31961: out = 16'(1769);
			31962: out = 16'(816);
			31963: out = 16'(150);
			31964: out = 16'(-772);
			31965: out = 16'(-1110);
			31966: out = 16'(-1532);
			31967: out = 16'(-481);
			31968: out = 16'(-156);
			31969: out = 16'(388);
			31970: out = 16'(-2280);
			31971: out = 16'(-3413);
			31972: out = 16'(-3114);
			31973: out = 16'(-1198);
			31974: out = 16'(618);
			31975: out = 16'(914);
			31976: out = 16'(1641);
			31977: out = 16'(1419);
			31978: out = 16'(793);
			31979: out = 16'(-433);
			31980: out = 16'(-1378);
			31981: out = 16'(-273);
			31982: out = 16'(-51);
			31983: out = 16'(49);
			31984: out = 16'(341);
			31985: out = 16'(485);
			31986: out = 16'(552);
			31987: out = 16'(136);
			31988: out = 16'(-226);
			31989: out = 16'(-750);
			31990: out = 16'(-52);
			31991: out = 16'(953);
			31992: out = 16'(2590);
			31993: out = 16'(2606);
			31994: out = 16'(2217);
			31995: out = 16'(298);
			31996: out = 16'(222);
			31997: out = 16'(236);
			31998: out = 16'(963);
			31999: out = 16'(291);
			32000: out = 16'(-419);
			32001: out = 16'(-448);
			32002: out = 16'(515);
			32003: out = 16'(2040);
			32004: out = 16'(174);
			32005: out = 16'(-847);
			32006: out = 16'(-2235);
			32007: out = 16'(-1610);
			32008: out = 16'(-1749);
			32009: out = 16'(-2688);
			32010: out = 16'(-1486);
			32011: out = 16'(-473);
			32012: out = 16'(-134);
			32013: out = 16'(293);
			32014: out = 16'(297);
			32015: out = 16'(46);
			32016: out = 16'(-163);
			32017: out = 16'(-314);
			32018: out = 16'(-2437);
			32019: out = 16'(-1588);
			32020: out = 16'(65);
			32021: out = 16'(267);
			32022: out = 16'(-25);
			32023: out = 16'(-1489);
			32024: out = 16'(185);
			32025: out = 16'(305);
			32026: out = 16'(134);
			32027: out = 16'(-943);
			32028: out = 16'(-1001);
			32029: out = 16'(76);
			32030: out = 16'(1035);
			32031: out = 16'(1796);
			32032: out = 16'(1015);
			32033: out = 16'(1481);
			32034: out = 16'(1558);
			32035: out = 16'(1658);
			32036: out = 16'(782);
			32037: out = 16'(-245);
			32038: out = 16'(-149);
			32039: out = 16'(-568);
			32040: out = 16'(-844);
			32041: out = 16'(-1395);
			32042: out = 16'(-896);
			32043: out = 16'(443);
			32044: out = 16'(-2);
			32045: out = 16'(-186);
			32046: out = 16'(-872);
			32047: out = 16'(1);
			32048: out = 16'(350);
			32049: out = 16'(-38);
			32050: out = 16'(-114);
			32051: out = 16'(-179);
			32052: out = 16'(-58);
			32053: out = 16'(483);
			32054: out = 16'(1240);
			32055: out = 16'(1415);
			32056: out = 16'(1640);
			32057: out = 16'(1366);
			32058: out = 16'(1169);
			32059: out = 16'(176);
			32060: out = 16'(-990);
			32061: out = 16'(-1854);
			32062: out = 16'(-1801);
			32063: out = 16'(-753);
			32064: out = 16'(-128);
			32065: out = 16'(607);
			32066: out = 16'(945);
			32067: out = 16'(1349);
			32068: out = 16'(1677);
			32069: out = 16'(2446);
			32070: out = 16'(2459);
			32071: out = 16'(2092);
			32072: out = 16'(-152);
			32073: out = 16'(-337);
			32074: out = 16'(-206);
			32075: out = 16'(1150);
			32076: out = 16'(1165);
			32077: out = 16'(591);
			32078: out = 16'(-610);
			32079: out = 16'(-2003);
			32080: out = 16'(-3521);
			32081: out = 16'(-2509);
			32082: out = 16'(-1646);
			32083: out = 16'(-260);
			32084: out = 16'(-47);
			32085: out = 16'(413);
			32086: out = 16'(30);
			32087: out = 16'(1456);
			32088: out = 16'(1707);
			32089: out = 16'(566);
			32090: out = 16'(-1341);
			32091: out = 16'(-2844);
			32092: out = 16'(-1589);
			32093: out = 16'(-731);
			32094: out = 16'(406);
			32095: out = 16'(-141);
			32096: out = 16'(53);
			32097: out = 16'(249);
			32098: out = 16'(-1136);
			32099: out = 16'(-1198);
			32100: out = 16'(-162);
			32101: out = 16'(219);
			32102: out = 16'(535);
			32103: out = 16'(256);
			32104: out = 16'(-415);
			32105: out = 16'(-885);
			32106: out = 16'(-183);
			32107: out = 16'(-32);
			32108: out = 16'(319);
			32109: out = 16'(-917);
			32110: out = 16'(-328);
			32111: out = 16'(81);
			32112: out = 16'(2409);
			32113: out = 16'(1905);
			32114: out = 16'(719);
			32115: out = 16'(-1987);
			32116: out = 16'(-3054);
			32117: out = 16'(-3196);
			32118: out = 16'(-1797);
			32119: out = 16'(-1496);
			32120: out = 16'(-2580);
			32121: out = 16'(-1253);
			32122: out = 16'(413);
			32123: out = 16'(3750);
			32124: out = 16'(3693);
			32125: out = 16'(3115);
			32126: out = 16'(-43);
			32127: out = 16'(-51);
			32128: out = 16'(-44);
			32129: out = 16'(1538);
			32130: out = 16'(891);
			32131: out = 16'(118);
			32132: out = 16'(-1317);
			32133: out = 16'(-1056);
			32134: out = 16'(-202);
			32135: out = 16'(-93);
			32136: out = 16'(-491);
			32137: out = 16'(-1475);
			32138: out = 16'(-1875);
			32139: out = 16'(-1368);
			32140: out = 16'(674);
			32141: out = 16'(1480);
			32142: out = 16'(2167);
			32143: out = 16'(816);
			32144: out = 16'(1512);
			32145: out = 16'(1398);
			32146: out = 16'(2200);
			32147: out = 16'(895);
			32148: out = 16'(-9);
			32149: out = 16'(-2694);
			32150: out = 16'(-1403);
			32151: out = 16'(467);
			32152: out = 16'(2264);
			32153: out = 16'(1528);
			32154: out = 16'(-372);
			32155: out = 16'(-1719);
			32156: out = 16'(-1554);
			32157: out = 16'(354);
			32158: out = 16'(740);
			32159: out = 16'(571);
			32160: out = 16'(-916);
			32161: out = 16'(-1731);
			32162: out = 16'(-1596);
			32163: out = 16'(874);
			32164: out = 16'(2161);
			32165: out = 16'(2813);
			32166: out = 16'(359);
			32167: out = 16'(-700);
			32168: out = 16'(-1596);
			32169: out = 16'(-345);
			32170: out = 16'(499);
			32171: out = 16'(1470);
			32172: out = 16'(93);
			32173: out = 16'(-895);
			32174: out = 16'(-2220);
			32175: out = 16'(-2077);
			32176: out = 16'(-2054);
			32177: out = 16'(-2034);
			32178: out = 16'(-806);
			32179: out = 16'(152);
			32180: out = 16'(1091);
			32181: out = 16'(323);
			32182: out = 16'(76);
			32183: out = 16'(931);
			32184: out = 16'(2123);
			32185: out = 16'(2969);
			32186: out = 16'(1046);
			32187: out = 16'(380);
			32188: out = 16'(-626);
			32189: out = 16'(-1214);
			32190: out = 16'(-2314);
			32191: out = 16'(-3279);
			32192: out = 16'(-757);
			32193: out = 16'(441);
			32194: out = 16'(998);
			32195: out = 16'(141);
			32196: out = 16'(-345);
			32197: out = 16'(31);
			32198: out = 16'(-187);
			32199: out = 16'(11);
			32200: out = 16'(-218);
			32201: out = 16'(940);
			32202: out = 16'(1414);
			32203: out = 16'(-81);
			32204: out = 16'(-136);
			32205: out = 16'(-10);
			32206: out = 16'(1350);
			32207: out = 16'(1106);
			32208: out = 16'(171);
			32209: out = 16'(-34);
			32210: out = 16'(-1147);
			32211: out = 16'(-2059);
			32212: out = 16'(-2689);
			32213: out = 16'(-1881);
			32214: out = 16'(13);
			32215: out = 16'(367);
			32216: out = 16'(153);
			32217: out = 16'(-1408);
			32218: out = 16'(-1366);
			32219: out = 16'(-1013);
			32220: out = 16'(369);
			32221: out = 16'(860);
			32222: out = 16'(1178);
			32223: out = 16'(1134);
			32224: out = 16'(771);
			32225: out = 16'(352);
			32226: out = 16'(468);
			32227: out = 16'(1316);
			32228: out = 16'(2668);
			32229: out = 16'(803);
			32230: out = 16'(-170);
			32231: out = 16'(-1551);
			32232: out = 16'(24);
			32233: out = 16'(624);
			32234: out = 16'(1020);
			32235: out = 16'(-253);
			32236: out = 16'(-864);
			32237: out = 16'(-23);
			32238: out = 16'(106);
			32239: out = 16'(449);
			32240: out = 16'(-973);
			32241: out = 16'(-62);
			32242: out = 16'(465);
			32243: out = 16'(1050);
			32244: out = 16'(114);
			32245: out = 16'(-1017);
			32246: out = 16'(-2412);
			32247: out = 16'(-2055);
			32248: out = 16'(-632);
			32249: out = 16'(-386);
			32250: out = 16'(-146);
			32251: out = 16'(-185);
			32252: out = 16'(-635);
			32253: out = 16'(-475);
			32254: out = 16'(339);
			32255: out = 16'(1239);
			32256: out = 16'(1214);
			32257: out = 16'(-1263);
			32258: out = 16'(-2022);
			32259: out = 16'(-2310);
			32260: out = 16'(258);
			32261: out = 16'(799);
			32262: out = 16'(1243);
			32263: out = 16'(1532);
			32264: out = 16'(1468);
			32265: out = 16'(935);
			32266: out = 16'(555);
			32267: out = 16'(251);
			32268: out = 16'(590);
			32269: out = 16'(254);
			32270: out = 16'(306);
			32271: out = 16'(-248);
			32272: out = 16'(1440);
			32273: out = 16'(1669);
			32274: out = 16'(-144);
			32275: out = 16'(-902);
			32276: out = 16'(-1422);
			32277: out = 16'(-108);
			32278: out = 16'(87);
			32279: out = 16'(382);
			32280: out = 16'(-1913);
			32281: out = 16'(-1511);
			32282: out = 16'(-660);
			32283: out = 16'(783);
			32284: out = 16'(724);
			32285: out = 16'(-220);
			32286: out = 16'(-73);
			32287: out = 16'(-643);
			32288: out = 16'(-1387);
			32289: out = 16'(-988);
			32290: out = 16'(-438);
			32291: out = 16'(555);
			32292: out = 16'(176);
			32293: out = 16'(-63);
			32294: out = 16'(-8);
			32295: out = 16'(255);
			32296: out = 16'(600);
			32297: out = 16'(423);
			32298: out = 16'(1050);
			32299: out = 16'(1573);
			32300: out = 16'(1050);
			32301: out = 16'(720);
			32302: out = 16'(216);
			32303: out = 16'(1666);
			32304: out = 16'(1960);
			32305: out = 16'(1836);
			32306: out = 16'(290);
			32307: out = 16'(-497);
			32308: out = 16'(-183);
			32309: out = 16'(-411);
			32310: out = 16'(-95);
			32311: out = 16'(163);
			32312: out = 16'(314);
			32313: out = 16'(-437);
			32314: out = 16'(-2562);
			32315: out = 16'(-3303);
			32316: out = 16'(-3180);
			32317: out = 16'(-3018);
			32318: out = 16'(-458);
			32319: out = 16'(2377);
			32320: out = 16'(1977);
			32321: out = 16'(1118);
			32322: out = 16'(-1192);
			32323: out = 16'(1227);
			32324: out = 16'(1383);
			32325: out = 16'(1547);
			32326: out = 16'(-1201);
			32327: out = 16'(-2194);
			32328: out = 16'(-1433);
			32329: out = 16'(-1169);
			32330: out = 16'(-773);
			32331: out = 16'(-917);
			32332: out = 16'(-377);
			32333: out = 16'(5);
			32334: out = 16'(-158);
			32335: out = 16'(492);
			32336: out = 16'(1073);
			32337: out = 16'(1013);
			32338: out = 16'(501);
			32339: out = 16'(-418);
			32340: out = 16'(-116);
			32341: out = 16'(349);
			32342: out = 16'(1692);
			32343: out = 16'(381);
			32344: out = 16'(274);
			32345: out = 16'(81);
			32346: out = 16'(1250);
			32347: out = 16'(901);
			32348: out = 16'(-883);
			32349: out = 16'(-2507);
			32350: out = 16'(-3242);
			32351: out = 16'(-1469);
			32352: out = 16'(-569);
			32353: out = 16'(477);
			32354: out = 16'(-369);
			32355: out = 16'(-19);
			32356: out = 16'(-183);
			32357: out = 16'(85);
			32358: out = 16'(-872);
			32359: out = 16'(-1972);
			32360: out = 16'(-427);
			32361: out = 16'(450);
			32362: out = 16'(1090);
			32363: out = 16'(1441);
			32364: out = 16'(2040);
			32365: out = 16'(3665);
			32366: out = 16'(1279);
			32367: out = 16'(-398);
			32368: out = 16'(-2052);
			32369: out = 16'(-731);
			32370: out = 16'(291);
			32371: out = 16'(-937);
			32372: out = 16'(-509);
			32373: out = 16'(-293);
			32374: out = 16'(-284);
			32375: out = 16'(-55);
			32376: out = 16'(414);
			32377: out = 16'(1609);
			32378: out = 16'(2336);
			32379: out = 16'(2803);
			32380: out = 16'(1987);
			32381: out = 16'(1831);
			32382: out = 16'(2219);
			32383: out = 16'(443);
			32384: out = 16'(-1253);
			32385: out = 16'(-3329);
			32386: out = 16'(-3087);
			32387: out = 16'(-2079);
			32388: out = 16'(22);
			32389: out = 16'(367);
			32390: out = 16'(122);
			32391: out = 16'(-715);
			32392: out = 16'(-1563);
			32393: out = 16'(-1953);
			32394: out = 16'(-1575);
			32395: out = 16'(-561);
			32396: out = 16'(580);
			32397: out = 16'(1286);
			32398: out = 16'(1114);
			32399: out = 16'(131);
			32400: out = 16'(-15);
			32401: out = 16'(63);
			32402: out = 16'(987);
			32403: out = 16'(835);
			32404: out = 16'(731);
			32405: out = 16'(-249);
			32406: out = 16'(-97);
			32407: out = 16'(-259);
			32408: out = 16'(-49);
			32409: out = 16'(-895);
			32410: out = 16'(-1567);
			32411: out = 16'(-2496);
			32412: out = 16'(-1740);
			32413: out = 16'(-619);
			32414: out = 16'(-1335);
			32415: out = 16'(-1009);
			32416: out = 16'(-670);
			32417: out = 16'(-684);
			32418: out = 16'(-661);
			32419: out = 16'(-623);
			32420: out = 16'(1016);
			32421: out = 16'(1574);
			32422: out = 16'(333);
			32423: out = 16'(411);
			32424: out = 16'(-296);
			32425: out = 16'(362);
			32426: out = 16'(-2307);
			32427: out = 16'(-3646);
			32428: out = 16'(-3713);
			32429: out = 16'(-1067);
			32430: out = 16'(1823);
			32431: out = 16'(3596);
			32432: out = 16'(3928);
			32433: out = 16'(3249);
			32434: out = 16'(1013);
			32435: out = 16'(310);
			32436: out = 16'(339);
			32437: out = 16'(2362);
			32438: out = 16'(2684);
			32439: out = 16'(1805);
			32440: out = 16'(-64);
			32441: out = 16'(-1117);
			32442: out = 16'(-850);
			32443: out = 16'(-438);
			32444: out = 16'(-198);
			32445: out = 16'(-211);
			32446: out = 16'(-1626);
			32447: out = 16'(-2506);
			32448: out = 16'(-1555);
			32449: out = 16'(273);
			32450: out = 16'(2236);
			32451: out = 16'(2784);
			32452: out = 16'(1747);
			32453: out = 16'(-497);
			32454: out = 16'(-1064);
			32455: out = 16'(-1286);
			32456: out = 16'(-105);
			32457: out = 16'(-305);
			32458: out = 16'(-28);
			32459: out = 16'(-227);
			32460: out = 16'(-79);
			32461: out = 16'(0);
			32462: out = 16'(993);
			32463: out = 16'(229);
			32464: out = 16'(-222);
			32465: out = 16'(-272);
			32466: out = 16'(-600);
			32467: out = 16'(-968);
			32468: out = 16'(-1847);
			32469: out = 16'(-1520);
			32470: out = 16'(-494);
			32471: out = 16'(556);
			32472: out = 16'(1858);
			32473: out = 16'(2896);
			32474: out = 16'(2908);
			32475: out = 16'(2337);
			32476: out = 16'(1249);
			32477: out = 16'(507);
			32478: out = 16'(-127);
			32479: out = 16'(-193);
			32480: out = 16'(-766);
			32481: out = 16'(-1170);
			32482: out = 16'(-2080);
			32483: out = 16'(-1704);
			32484: out = 16'(-1496);
			32485: out = 16'(-1943);
			32486: out = 16'(-1964);
			32487: out = 16'(-1756);
			32488: out = 16'(-474);
			32489: out = 16'(78);
			32490: out = 16'(291);
			32491: out = 16'(345);
			32492: out = 16'(248);
			32493: out = 16'(329);
			32494: out = 16'(-1004);
			32495: out = 16'(-1255);
			32496: out = 16'(-705);
			32497: out = 16'(-57);
			32498: out = 16'(501);
			32499: out = 16'(446);
			32500: out = 16'(271);
			32501: out = 16'(-467);
			32502: out = 16'(-2284);
			32503: out = 16'(-2537);
			32504: out = 16'(-1877);
			32505: out = 16'(1664);
			32506: out = 16'(2656);
			32507: out = 16'(2853);
			32508: out = 16'(391);
			32509: out = 16'(-177);
			32510: out = 16'(21);
			32511: out = 16'(312);
			32512: out = 16'(391);
			32513: out = 16'(-168);
			32514: out = 16'(296);
			32515: out = 16'(262);
			32516: out = 16'(557);
			32517: out = 16'(4);
			32518: out = 16'(-65);
			32519: out = 16'(-336);
			32520: out = 16'(-28);
			32521: out = 16'(-237);
			32522: out = 16'(137);
			32523: out = 16'(-1385);
			32524: out = 16'(-2532);
			32525: out = 16'(-2560);
			32526: out = 16'(-1387);
			32527: out = 16'(69);
			32528: out = 16'(1374);
			32529: out = 16'(1264);
			32530: out = 16'(536);
			32531: out = 16'(-522);
			32532: out = 16'(66);
			32533: out = 16'(2089);
			32534: out = 16'(3067);
			32535: out = 16'(2689);
			32536: out = 16'(-356);
			32537: out = 16'(-967);
			32538: out = 16'(-1232);
			32539: out = 16'(401);
			32540: out = 16'(1416);
			32541: out = 16'(2727);
			32542: out = 16'(3059);
			32543: out = 16'(3148);
			32544: out = 16'(2355);
			32545: out = 16'(641);
			32546: out = 16'(-258);
			32547: out = 16'(-249);
			32548: out = 16'(-197);
			32549: out = 16'(343);
			32550: out = 16'(594);
			32551: out = 16'(437);
			32552: out = 16'(-576);
			32553: out = 16'(-2156);
			32554: out = 16'(-3052);
			32555: out = 16'(-2843);
			32556: out = 16'(-378);
			32557: out = 16'(-394);
			32558: out = 16'(-640);
			32559: out = 16'(-2558);
			32560: out = 16'(-2288);
			32561: out = 16'(-1679);
			32562: out = 16'(212);
			32563: out = 16'(749);
			32564: out = 16'(846);
			32565: out = 16'(-954);
			32566: out = 16'(-2068);
			32567: out = 16'(-3093);
			32568: out = 16'(-641);
			32569: out = 16'(575);
			32570: out = 16'(1602);
			32571: out = 16'(-55);
			32572: out = 16'(-1120);
			32573: out = 16'(-1824);
			32574: out = 16'(-834);
			32575: out = 16'(246);
			32576: out = 16'(977);
			32577: out = 16'(837);
			32578: out = 16'(351);
			32579: out = 16'(-41);
			32580: out = 16'(-526);
			32581: out = 16'(-521);
			32582: out = 16'(1248);
			32583: out = 16'(2185);
			32584: out = 16'(2960);
			32585: out = 16'(1211);
			32586: out = 16'(1032);
			32587: out = 16'(1412);
			32588: out = 16'(1404);
			32589: out = 16'(903);
			32590: out = 16'(-492);
			32591: out = 16'(-688);
			32592: out = 16'(-1164);
			32593: out = 16'(-1367);
			32594: out = 16'(-2204);
			32595: out = 16'(-2376);
			32596: out = 16'(-844);
			32597: out = 16'(-247);
			32598: out = 16'(386);
			32599: out = 16'(-871);
			32600: out = 16'(-87);
			32601: out = 16'(590);
			32602: out = 16'(2282);
			32603: out = 16'(1883);
			32604: out = 16'(775);
			32605: out = 16'(-466);
			32606: out = 16'(-972);
			32607: out = 16'(-800);
			32608: out = 16'(66);
			32609: out = 16'(587);
			32610: out = 16'(943);
			32611: out = 16'(170);
			32612: out = 16'(0);
			32613: out = 16'(822);
			32614: out = 16'(1782);
			32615: out = 16'(2196);
			32616: out = 16'(928);
			32617: out = 16'(-628);
			32618: out = 16'(-2247);
			32619: out = 16'(-406);
			32620: out = 16'(-391);
			32621: out = 16'(-87);
			32622: out = 16'(-434);
			32623: out = 16'(-208);
			32624: out = 16'(-268);
			32625: out = 16'(-66);
			32626: out = 16'(-603);
			32627: out = 16'(-1407);
			32628: out = 16'(-1514);
			32629: out = 16'(-1081);
			32630: out = 16'(-316);
			32631: out = 16'(254);
			32632: out = 16'(339);
			32633: out = 16'(-18);
			32634: out = 16'(-824);
			32635: out = 16'(-1351);
			32636: out = 16'(-861);
			32637: out = 16'(96);
			32638: out = 16'(1102);
			32639: out = 16'(380);
			32640: out = 16'(-324);
			32641: out = 16'(-1418);
			32642: out = 16'(640);
			32643: out = 16'(1471);
			32644: out = 16'(2555);
			32645: out = 16'(706);
			32646: out = 16'(39);
			32647: out = 16'(-381);
			32648: out = 16'(1231);
			32649: out = 16'(1702);
			32650: out = 16'(95);
			32651: out = 16'(-109);
			32652: out = 16'(-419);
			32653: out = 16'(228);
			32654: out = 16'(70);
			32655: out = 16'(229);
			32656: out = 16'(-292);
			32657: out = 16'(330);
			32658: out = 16'(898);
			32659: out = 16'(2148);
			32660: out = 16'(1903);
			32661: out = 16'(1084);
			32662: out = 16'(-1872);
			32663: out = 16'(-3009);
			32664: out = 16'(-2532);
			32665: out = 16'(-2336);
			32666: out = 16'(-1827);
			32667: out = 16'(-2039);
			32668: out = 16'(-603);
			32669: out = 16'(52);
			32670: out = 16'(-60);
			32671: out = 16'(-8);
			32672: out = 16'(119);
			32673: out = 16'(1504);
			32674: out = 16'(692);
			32675: out = 16'(-397);
			32676: out = 16'(-143);
			32677: out = 16'(-33);
			32678: out = 16'(538);
			32679: out = 16'(-1635);
			32680: out = 16'(-1484);
			32681: out = 16'(-661);
			32682: out = 16'(1007);
			32683: out = 16'(1639);
			32684: out = 16'(1440);
			32685: out = 16'(447);
			32686: out = 16'(-141);
			32687: out = 16'(538);
			32688: out = 16'(270);
			32689: out = 16'(159);
			32690: out = 16'(-877);
			32691: out = 16'(-200);
			32692: out = 16'(328);
			32693: out = 16'(237);
			32694: out = 16'(277);
			32695: out = 16'(227);
			32696: out = 16'(273);
			32697: out = 16'(31);
			32698: out = 16'(-301);
			32699: out = 16'(-148);
			32700: out = 16'(37);
			32701: out = 16'(447);
			32702: out = 16'(-13);
			32703: out = 16'(-56);
			32704: out = 16'(270);
			32705: out = 16'(215);
			32706: out = 16'(202);
			32707: out = 16'(-158);
			32708: out = 16'(-111);
			32709: out = 16'(-128);
			32710: out = 16'(443);
			32711: out = 16'(11);
			32712: out = 16'(-321);
			32713: out = 16'(-370);
			32714: out = 16'(242);
			32715: out = 16'(983);
			32716: out = 16'(1286);
			32717: out = 16'(1219);
			32718: out = 16'(747);
			32719: out = 16'(20);
			32720: out = 16'(-1082);
			32721: out = 16'(-2683);
			32722: out = 16'(-1400);
			32723: out = 16'(-582);
			32724: out = 16'(-151);
			32725: out = 16'(115);
			32726: out = 16'(268);
			32727: out = 16'(-190);
			32728: out = 16'(497);
			32729: out = 16'(802);
			32730: out = 16'(-112);
			32731: out = 16'(-1372);
			32732: out = 16'(-2596);
			32733: out = 16'(-1504);
			32734: out = 16'(-800);
			32735: out = 16'(56);
			32736: out = 16'(-63);
			32737: out = 16'(-191);
			32738: out = 16'(-756);
			32739: out = 16'(31);
			32740: out = 16'(821);
			32741: out = 16'(2002);
			32742: out = 16'(2291);
			32743: out = 16'(2105);
			32744: out = 16'(345);
			32745: out = 16'(421);
			32746: out = 16'(225);
			32747: out = 16'(-74);
			32748: out = 16'(-558);
			32749: out = 16'(-838);
			32750: out = 16'(-242);
			32751: out = 16'(45);
			32752: out = 16'(335);
			32753: out = 16'(-203);
			32754: out = 16'(-929);
			32755: out = 16'(-2113);
			32756: out = 16'(-702);
			32757: out = 16'(76);
			32758: out = 16'(999);
			32759: out = 16'(379);
			32760: out = 16'(123);
			32761: out = 16'(-427);
			32762: out = 16'(513);
			32763: out = 16'(933);
			32764: out = 16'(1475);
			32765: out = 16'(82);
			32766: out = 16'(-1161);
			32767: out = 16'(-2025);
			32768: out = 16'(-708);
			32769: out = 16'(1193);
			32770: out = 16'(1216);
			32771: out = 16'(915);
			32772: out = 16'(-463);
			32773: out = 16'(335);
			32774: out = 16'(-337);
			32775: out = 16'(-852);
			32776: out = 16'(-1855);
			32777: out = 16'(-1602);
			32778: out = 16'(-267);
			32779: out = 16'(178);
			32780: out = 16'(398);
			32781: out = 16'(-220);
			32782: out = 16'(787);
			32783: out = 16'(1737);
			32784: out = 16'(2697);
			32785: out = 16'(2394);
			32786: out = 16'(1470);
			32787: out = 16'(1042);
			32788: out = 16'(-202);
			32789: out = 16'(-1127);
			32790: out = 16'(-2610);
			32791: out = 16'(-1726);
			32792: out = 16'(325);
			32793: out = 16'(-231);
			32794: out = 16'(-376);
			32795: out = 16'(-1013);
			32796: out = 16'(-475);
			32797: out = 16'(-586);
			32798: out = 16'(-1544);
			32799: out = 16'(-362);
			32800: out = 16'(360);
			32801: out = 16'(350);
			32802: out = 16'(34);
			32803: out = 16'(-600);
			32804: out = 16'(-1877);
			32805: out = 16'(-1750);
			32806: out = 16'(-1163);
			32807: out = 16'(41);
			32808: out = 16'(678);
			32809: out = 16'(976);
			32810: out = 16'(390);
			32811: out = 16'(242);
			32812: out = 16'(266);
			32813: out = 16'(395);
			32814: out = 16'(527);
			32815: out = 16'(973);
			32816: out = 16'(381);
			32817: out = 16'(25);
			32818: out = 16'(-1008);
			32819: out = 16'(624);
			32820: out = 16'(1626);
			32821: out = 16'(2369);
			32822: out = 16'(928);
			32823: out = 16'(-454);
			32824: out = 16'(-190);
			32825: out = 16'(-48);
			32826: out = 16'(277);
			32827: out = 16'(-135);
			32828: out = 16'(-974);
			32829: out = 16'(-2204);
			32830: out = 16'(-2522);
			32831: out = 16'(-1972);
			32832: out = 16'(-54);
			32833: out = 16'(-294);
			32834: out = 16'(35);
			32835: out = 16'(-252);
			32836: out = 16'(737);
			32837: out = 16'(709);
			32838: out = 16'(-55);
			32839: out = 16'(-591);
			32840: out = 16'(-742);
			32841: out = 16'(-154);
			32842: out = 16'(185);
			32843: out = 16'(407);
			32844: out = 16'(-59);
			32845: out = 16'(18);
			32846: out = 16'(278);
			32847: out = 16'(-756);
			32848: out = 16'(-415);
			32849: out = 16'(287);
			32850: out = 16'(57);
			32851: out = 16'(-530);
			32852: out = 16'(-1311);
			32853: out = 16'(-1438);
			32854: out = 16'(-583);
			32855: out = 16'(1547);
			32856: out = 16'(2147);
			32857: out = 16'(2273);
			32858: out = 16'(918);
			32859: out = 16'(642);
			32860: out = 16'(370);
			32861: out = 16'(867);
			32862: out = 16'(859);
			32863: out = 16'(684);
			32864: out = 16'(-1141);
			32865: out = 16'(-2241);
			32866: out = 16'(-3193);
			32867: out = 16'(-1693);
			32868: out = 16'(-847);
			32869: out = 16'(47);
			32870: out = 16'(218);
			32871: out = 16'(119);
			32872: out = 16'(-889);
			32873: out = 16'(99);
			32874: out = 16'(310);
			32875: out = 16'(401);
			32876: out = 16'(-411);
			32877: out = 16'(-643);
			32878: out = 16'(-135);
			32879: out = 16'(1059);
			32880: out = 16'(2087);
			32881: out = 16'(1485);
			32882: out = 16'(812);
			32883: out = 16'(-376);
			32884: out = 16'(-55);
			32885: out = 16'(-1218);
			32886: out = 16'(-2585);
			32887: out = 16'(-1587);
			32888: out = 16'(-795);
			32889: out = 16'(459);
			32890: out = 16'(-168);
			32891: out = 16'(173);
			32892: out = 16'(981);
			32893: out = 16'(2278);
			32894: out = 16'(2878);
			32895: out = 16'(1837);
			32896: out = 16'(1374);
			32897: out = 16'(609);
			32898: out = 16'(322);
			32899: out = 16'(-235);
			32900: out = 16'(-263);
			32901: out = 16'(628);
			32902: out = 16'(909);
			32903: out = 16'(659);
			32904: out = 16'(496);
			32905: out = 16'(-296);
			32906: out = 16'(-953);
			32907: out = 16'(-2363);
			32908: out = 16'(-2222);
			32909: out = 16'(-811);
			32910: out = 16'(-402);
			32911: out = 16'(-109);
			32912: out = 16'(-311);
			32913: out = 16'(-958);
			32914: out = 16'(-1422);
			32915: out = 16'(-764);
			32916: out = 16'(-303);
			32917: out = 16'(460);
			32918: out = 16'(-205);
			32919: out = 16'(503);
			32920: out = 16'(951);
			32921: out = 16'(1487);
			32922: out = 16'(793);
			32923: out = 16'(-250);
			32924: out = 16'(-1124);
			32925: out = 16'(-1333);
			32926: out = 16'(-742);
			32927: out = 16'(-857);
			32928: out = 16'(-743);
			32929: out = 16'(-793);
			32930: out = 16'(-68);
			32931: out = 16'(482);
			32932: out = 16'(366);
			32933: out = 16'(1401);
			32934: out = 16'(1905);
			32935: out = 16'(963);
			32936: out = 16'(395);
			32937: out = 16'(-216);
			32938: out = 16'(851);
			32939: out = 16'(611);
			32940: out = 16'(303);
			32941: out = 16'(182);
			32942: out = 16'(138);
			32943: out = 16'(131);
			32944: out = 16'(-282);
			32945: out = 16'(-89);
			32946: out = 16'(932);
			32947: out = 16'(50);
			32948: out = 16'(-682);
			32949: out = 16'(-2780);
			32950: out = 16'(-807);
			32951: out = 16'(392);
			32952: out = 16'(375);
			32953: out = 16'(-277);
			32954: out = 16'(-928);
			32955: out = 16'(-312);
			32956: out = 16'(-77);
			32957: out = 16'(210);
			32958: out = 16'(-735);
			32959: out = 16'(-877);
			32960: out = 16'(-738);
			32961: out = 16'(-24);
			32962: out = 16'(627);
			32963: out = 16'(875);
			32964: out = 16'(1787);
			32965: out = 16'(1203);
			32966: out = 16'(-929);
			32967: out = 16'(-1640);
			32968: out = 16'(-1411);
			32969: out = 16'(2068);
			32970: out = 16'(891);
			32971: out = 16'(270);
			32972: out = 16'(-353);
			32973: out = 16'(52);
			32974: out = 16'(369);
			32975: out = 16'(382);
			32976: out = 16'(48);
			32977: out = 16'(-396);
			32978: out = 16'(119);
			32979: out = 16'(87);
			32980: out = 16'(-215);
			32981: out = 16'(661);
			32982: out = 16'(847);
			32983: out = 16'(842);
			32984: out = 16'(-401);
			32985: out = 16'(-1191);
			32986: out = 16'(-1455);
			32987: out = 16'(-806);
			32988: out = 16'(-178);
			32989: out = 16'(-230);
			32990: out = 16'(-110);
			32991: out = 16'(-139);
			32992: out = 16'(250);
			32993: out = 16'(22);
			32994: out = 16'(-157);
			32995: out = 16'(-311);
			32996: out = 16'(-103);
			32997: out = 16'(249);
			32998: out = 16'(-68);
			32999: out = 16'(-369);
			33000: out = 16'(-909);
			33001: out = 16'(-822);
			33002: out = 16'(-740);
			33003: out = 16'(-176);
			33004: out = 16'(-387);
			33005: out = 16'(100);
			33006: out = 16'(839);
			33007: out = 16'(2178);
			33008: out = 16'(2857);
			33009: out = 16'(2364);
			33010: out = 16'(997);
			33011: out = 16'(-488);
			33012: out = 16'(882);
			33013: out = 16'(180);
			33014: out = 16'(-396);
			33015: out = 16'(-2423);
			33016: out = 16'(-2326);
			33017: out = 16'(-1299);
			33018: out = 16'(-102);
			33019: out = 16'(669);
			33020: out = 16'(773);
			33021: out = 16'(597);
			33022: out = 16'(10);
			33023: out = 16'(-266);
			33024: out = 16'(-1903);
			33025: out = 16'(-2752);
			33026: out = 16'(-2508);
			33027: out = 16'(-2240);
			33028: out = 16'(-1577);
			33029: out = 16'(-315);
			33030: out = 16'(-23);
			33031: out = 16'(44);
			33032: out = 16'(489);
			33033: out = 16'(554);
			33034: out = 16'(485);
			33035: out = 16'(552);
			33036: out = 16'(86);
			33037: out = 16'(-832);
			33038: out = 16'(-293);
			33039: out = 16'(-52);
			33040: out = 16'(407);
			33041: out = 16'(5);
			33042: out = 16'(396);
			33043: out = 16'(2049);
			33044: out = 16'(1333);
			33045: out = 16'(710);
			33046: out = 16'(-72);
			33047: out = 16'(118);
			33048: out = 16'(531);
			33049: out = 16'(824);
			33050: out = 16'(705);
			33051: out = 16'(322);
			33052: out = 16'(1361);
			33053: out = 16'(920);
			33054: out = 16'(269);
			33055: out = 16'(192);
			33056: out = 16'(-8);
			33057: out = 16'(-495);
			33058: out = 16'(93);
			33059: out = 16'(1);
			33060: out = 16'(-128);
			33061: out = 16'(-1516);
			33062: out = 16'(-2087);
			33063: out = 16'(-2052);
			33064: out = 16'(-635);
			33065: out = 16'(341);
			33066: out = 16'(-286);
			33067: out = 16'(-815);
			33068: out = 16'(-1336);
			33069: out = 16'(209);
			33070: out = 16'(307);
			33071: out = 16'(281);
			33072: out = 16'(336);
			33073: out = 16'(110);
			33074: out = 16'(-100);
			33075: out = 16'(-1115);
			33076: out = 16'(-1068);
			33077: out = 16'(-138);
			33078: out = 16'(1319);
			33079: out = 16'(2136);
			33080: out = 16'(1830);
			33081: out = 16'(719);
			33082: out = 16'(-466);
			33083: out = 16'(82);
			33084: out = 16'(-1055);
			33085: out = 16'(-1275);
			33086: out = 16'(-1063);
			33087: out = 16'(400);
			33088: out = 16'(1563);
			33089: out = 16'(1884);
			33090: out = 16'(1228);
			33091: out = 16'(12);
			33092: out = 16'(-229);
			33093: out = 16'(-350);
			33094: out = 16'(-147);
			33095: out = 16'(130);
			33096: out = 16'(-360);
			33097: out = 16'(-2156);
			33098: out = 16'(-1172);
			33099: out = 16'(-658);
			33100: out = 16'(-93);
			33101: out = 16'(98);
			33102: out = 16'(291);
			33103: out = 16'(-167);
			33104: out = 16'(208);
			33105: out = 16'(409);
			33106: out = 16'(299);
			33107: out = 16'(-55);
			33108: out = 16'(-354);
			33109: out = 16'(-803);
			33110: out = 16'(-454);
			33111: out = 16'(347);
			33112: out = 16'(343);
			33113: out = 16'(300);
			33114: out = 16'(-228);
			33115: out = 16'(-74);
			33116: out = 16'(275);
			33117: out = 16'(2145);
			33118: out = 16'(728);
			33119: out = 16'(448);
			33120: out = 16'(18);
			33121: out = 16'(1878);
			33122: out = 16'(2807);
			33123: out = 16'(2896);
			33124: out = 16'(523);
			33125: out = 16'(-1961);
			33126: out = 16'(-2546);
			33127: out = 16'(-1538);
			33128: out = 16'(659);
			33129: out = 16'(561);
			33130: out = 16'(615);
			33131: out = 16'(-683);
			33132: out = 16'(-163);
			33133: out = 16'(-895);
			33134: out = 16'(-1332);
			33135: out = 16'(-2399);
			33136: out = 16'(-2187);
			33137: out = 16'(-844);
			33138: out = 16'(-428);
			33139: out = 16'(-202);
			33140: out = 16'(-38);
			33141: out = 16'(-104);
			33142: out = 16'(-149);
			33143: out = 16'(-1862);
			33144: out = 16'(-1068);
			33145: out = 16'(61);
			33146: out = 16'(2187);
			33147: out = 16'(1979);
			33148: out = 16'(758);
			33149: out = 16'(-354);
			33150: out = 16'(-1124);
			33151: out = 16'(-1300);
			33152: out = 16'(-563);
			33153: out = 16'(-92);
			33154: out = 16'(-52);
			33155: out = 16'(-504);
			33156: out = 16'(-559);
			33157: out = 16'(480);
			33158: out = 16'(1018);
			33159: out = 16'(1275);
			33160: out = 16'(-730);
			33161: out = 16'(-453);
			33162: out = 16'(-214);
			33163: out = 16'(-228);
			33164: out = 16'(-206);
			33165: out = 16'(-240);
			33166: out = 16'(-595);
			33167: out = 16'(-1089);
			33168: out = 16'(-1773);
			33169: out = 16'(-517);
			33170: out = 16'(101);
			33171: out = 16'(338);
			33172: out = 16'(194);
			33173: out = 16'(12);
			33174: out = 16'(634);
			33175: out = 16'(-601);
			33176: out = 16'(-1239);
			33177: out = 16'(-1217);
			33178: out = 16'(16);
			33179: out = 16'(1367);
			33180: out = 16'(1757);
			33181: out = 16'(2049);
			33182: out = 16'(1710);
			33183: out = 16'(1186);
			33184: out = 16'(159);
			33185: out = 16'(-784);
			33186: out = 16'(-274);
			33187: out = 16'(531);
			33188: out = 16'(1922);
			33189: out = 16'(1424);
			33190: out = 16'(1091);
			33191: out = 16'(234);
			33192: out = 16'(83);
			33193: out = 16'(-457);
			33194: out = 16'(-685);
			33195: out = 16'(-1631);
			33196: out = 16'(-1553);
			33197: out = 16'(-32);
			33198: out = 16'(1381);
			33199: out = 16'(2218);
			33200: out = 16'(1441);
			33201: out = 16'(282);
			33202: out = 16'(-1082);
			33203: out = 16'(-1380);
			33204: out = 16'(-1033);
			33205: out = 16'(-81);
			33206: out = 16'(888);
			33207: out = 16'(1256);
			33208: out = 16'(656);
			33209: out = 16'(46);
			33210: out = 16'(-783);
			33211: out = 16'(-1425);
			33212: out = 16'(-538);
			33213: out = 16'(432);
			33214: out = 16'(671);
			33215: out = 16'(604);
			33216: out = 16'(66);
			33217: out = 16'(-93);
			33218: out = 16'(-201);
			33219: out = 16'(169);
			33220: out = 16'(-1966);
			33221: out = 16'(-1054);
			33222: out = 16'(200);
			33223: out = 16'(434);
			33224: out = 16'(-817);
			33225: out = 16'(-3183);
			33226: out = 16'(-2608);
			33227: out = 16'(-1830);
			33228: out = 16'(-164);
			33229: out = 16'(127);
			33230: out = 16'(351);
			33231: out = 16'(306);
			33232: out = 16'(-22);
			33233: out = 16'(-431);
			33234: out = 16'(-1813);
			33235: out = 16'(-1174);
			33236: out = 16'(-580);
			33237: out = 16'(378);
			33238: out = 16'(-412);
			33239: out = 16'(-1178);
			33240: out = 16'(-878);
			33241: out = 16'(641);
			33242: out = 16'(2527);
			33243: out = 16'(2119);
			33244: out = 16'(892);
			33245: out = 16'(-1356);
			33246: out = 16'(-1694);
			33247: out = 16'(-1271);
			33248: out = 16'(357);
			33249: out = 16'(1705);
			33250: out = 16'(2581);
			33251: out = 16'(2796);
			33252: out = 16'(1086);
			33253: out = 16'(-311);
			33254: out = 16'(377);
			33255: out = 16'(1427);
			33256: out = 16'(2825);
			33257: out = 16'(1241);
			33258: out = 16'(1104);
			33259: out = 16'(550);
			33260: out = 16'(415);
			33261: out = 16'(-297);
			33262: out = 16'(-977);
			33263: out = 16'(-194);
			33264: out = 16'(20);
			33265: out = 16'(-560);
			33266: out = 16'(13);
			33267: out = 16'(-91);
			33268: out = 16'(-370);
			33269: out = 16'(-1457);
			33270: out = 16'(-1812);
			33271: out = 16'(181);
			33272: out = 16'(-199);
			33273: out = 16'(-551);
			33274: out = 16'(-2445);
			33275: out = 16'(-1719);
			33276: out = 16'(-506);
			33277: out = 16'(1465);
			33278: out = 16'(1931);
			33279: out = 16'(1649);
			33280: out = 16'(522);
			33281: out = 16'(-147);
			33282: out = 16'(-353);
			33283: out = 16'(-20);
			33284: out = 16'(130);
			33285: out = 16'(-270);
			33286: out = 16'(-179);
			33287: out = 16'(-167);
			33288: out = 16'(206);
			33289: out = 16'(-202);
			33290: out = 16'(-339);
			33291: out = 16'(-212);
			33292: out = 16'(-189);
			33293: out = 16'(-281);
			33294: out = 16'(-1304);
			33295: out = 16'(-880);
			33296: out = 16'(12);
			33297: out = 16'(-277);
			33298: out = 16'(-39);
			33299: out = 16'(-416);
			33300: out = 16'(1207);
			33301: out = 16'(944);
			33302: out = 16'(238);
			33303: out = 16'(-2203);
			33304: out = 16'(-2765);
			33305: out = 16'(-1209);
			33306: out = 16'(-317);
			33307: out = 16'(436);
			33308: out = 16'(-117);
			33309: out = 16'(221);
			33310: out = 16'(208);
			33311: out = 16'(-759);
			33312: out = 16'(151);
			33313: out = 16'(1007);
			33314: out = 16'(538);
			33315: out = 16'(-473);
			33316: out = 16'(-1859);
			33317: out = 16'(539);
			33318: out = 16'(1633);
			33319: out = 16'(2840);
			33320: out = 16'(908);
			33321: out = 16'(82);
			33322: out = 16'(-264);
			33323: out = 16'(-236);
			33324: out = 16'(5);
			33325: out = 16'(317);
			33326: out = 16'(977);
			33327: out = 16'(1274);
			33328: out = 16'(843);
			33329: out = 16'(-57);
			33330: out = 16'(-998);
			33331: out = 16'(238);
			33332: out = 16'(-181);
			33333: out = 16'(-371);
			33334: out = 16'(-1873);
			33335: out = 16'(-1078);
			33336: out = 16'(381);
			33337: out = 16'(1109);
			33338: out = 16'(1066);
			33339: out = 16'(40);
			33340: out = 16'(-510);
			33341: out = 16'(-774);
			33342: out = 16'(356);
			33343: out = 16'(-618);
			33344: out = 16'(-881);
			33345: out = 16'(-1476);
			33346: out = 16'(-251);
			33347: out = 16'(632);
			33348: out = 16'(1808);
			33349: out = 16'(804);
			33350: out = 16'(-369);
			33351: out = 16'(-710);
			33352: out = 16'(-685);
			33353: out = 16'(-156);
			33354: out = 16'(610);
			33355: out = 16'(1222);
			33356: out = 16'(1769);
			33357: out = 16'(196);
			33358: out = 16'(-185);
			33359: out = 16'(190);
			33360: out = 16'(931);
			33361: out = 16'(1034);
			33362: out = 16'(-377);
			33363: out = 16'(80);
			33364: out = 16'(4);
			33365: out = 16'(-177);
			33366: out = 16'(-650);
			33367: out = 16'(-818);
			33368: out = 16'(229);
			33369: out = 16'(53);
			33370: out = 16'(-431);
			33371: out = 16'(-2173);
			33372: out = 16'(-2594);
			33373: out = 16'(-2293);
			33374: out = 16'(-1207);
			33375: out = 16'(-173);
			33376: out = 16'(372);
			33377: out = 16'(198);
			33378: out = 16'(-863);
			33379: out = 16'(-2946);
			33380: out = 16'(-2205);
			33381: out = 16'(-970);
			33382: out = 16'(1481);
			33383: out = 16'(1276);
			33384: out = 16'(780);
			33385: out = 16'(100);
			33386: out = 16'(-412);
			33387: out = 16'(-842);
			33388: out = 16'(-2276);
			33389: out = 16'(-1383);
			33390: out = 16'(102);
			33391: out = 16'(-83);
			33392: out = 16'(142);
			33393: out = 16'(29);
			33394: out = 16'(1259);
			33395: out = 16'(1560);
			33396: out = 16'(1462);
			33397: out = 16'(431);
			33398: out = 16'(-310);
			33399: out = 16'(-632);
			33400: out = 16'(-1130);
			33401: out = 16'(-959);
			33402: out = 16'(343);
			33403: out = 16'(206);
			33404: out = 16'(-50);
			33405: out = 16'(45);
			33406: out = 16'(-97);
			33407: out = 16'(-71);
			33408: out = 16'(227);
			33409: out = 16'(710);
			33410: out = 16'(956);
			33411: out = 16'(1023);
			33412: out = 16'(563);
			33413: out = 16'(-77);
			33414: out = 16'(-204);
			33415: out = 16'(-62);
			33416: out = 16'(267);
			33417: out = 16'(1396);
			33418: out = 16'(1943);
			33419: out = 16'(1787);
			33420: out = 16'(858);
			33421: out = 16'(-75);
			33422: out = 16'(-243);
			33423: out = 16'(-425);
			33424: out = 16'(-252);
			33425: out = 16'(-228);
			33426: out = 16'(86);
			33427: out = 16'(335);
			33428: out = 16'(-122);
			33429: out = 16'(-210);
			33430: out = 16'(-360);
			33431: out = 16'(-143);
			33432: out = 16'(-93);
			33433: out = 16'(299);
			33434: out = 16'(-677);
			33435: out = 16'(-622);
			33436: out = 16'(-202);
			33437: out = 16'(1514);
			33438: out = 16'(2211);
			33439: out = 16'(1244);
			33440: out = 16'(390);
			33441: out = 16'(-855);
			33442: out = 16'(-2321);
			33443: out = 16'(-2588);
			33444: out = 16'(-2348);
			33445: out = 16'(-1924);
			33446: out = 16'(-1770);
			33447: out = 16'(-1697);
			33448: out = 16'(-897);
			33449: out = 16'(-138);
			33450: out = 16'(608);
			33451: out = 16'(1661);
			33452: out = 16'(1750);
			33453: out = 16'(858);
			33454: out = 16'(575);
			33455: out = 16'(105);
			33456: out = 16'(-3);
			33457: out = 16'(142);
			33458: out = 16'(698);
			33459: out = 16'(1263);
			33460: out = 16'(1462);
			33461: out = 16'(1069);
			33462: out = 16'(30);
			33463: out = 16'(-580);
			33464: out = 16'(-746);
			33465: out = 16'(5);
			33466: out = 16'(384);
			33467: out = 16'(228);
			33468: out = 16'(434);
			33469: out = 16'(-803);
			33470: out = 16'(-2499);
			33471: out = 16'(-2531);
			33472: out = 16'(-1708);
			33473: out = 16'(-29);
			33474: out = 16'(1307);
			33475: out = 16'(1630);
			33476: out = 16'(-331);
			33477: out = 16'(-186);
			33478: out = 16'(-248);
			33479: out = 16'(-36);
			33480: out = 16'(-102);
			33481: out = 16'(-67);
			33482: out = 16'(-74);
			33483: out = 16'(73);
			33484: out = 16'(354);
			33485: out = 16'(-146);
			33486: out = 16'(538);
			33487: out = 16'(1371);
			33488: out = 16'(679);
			33489: out = 16'(-242);
			33490: out = 16'(-1303);
			33491: out = 16'(-1449);
			33492: out = 16'(-869);
			33493: out = 16'(-199);
			33494: out = 16'(1625);
			33495: out = 16'(2208);
			33496: out = 16'(1443);
			33497: out = 16'(-211);
			33498: out = 16'(-1743);
			33499: out = 16'(-2910);
			33500: out = 16'(-2174);
			33501: out = 16'(-1004);
			33502: out = 16'(186);
			33503: out = 16'(-84);
			33504: out = 16'(-776);
			33505: out = 16'(-2112);
			33506: out = 16'(-1552);
			33507: out = 16'(37);
			33508: out = 16'(1219);
			33509: out = 16'(1297);
			33510: out = 16'(532);
			33511: out = 16'(-1421);
			33512: out = 16'(-2405);
			33513: out = 16'(-2253);
			33514: out = 16'(-137);
			33515: out = 16'(1510);
			33516: out = 16'(1980);
			33517: out = 16'(925);
			33518: out = 16'(-250);
			33519: out = 16'(22);
			33520: out = 16'(1130);
			33521: out = 16'(2632);
			33522: out = 16'(2307);
			33523: out = 16'(2027);
			33524: out = 16'(1226);
			33525: out = 16'(120);
			33526: out = 16'(365);
			33527: out = 16'(1948);
			33528: out = 16'(1359);
			33529: out = 16'(781);
			33530: out = 16'(-1032);
			33531: out = 16'(-500);
			33532: out = 16'(-249);
			33533: out = 16'(334);
			33534: out = 16'(183);
			33535: out = 16'(169);
			33536: out = 16'(290);
			33537: out = 16'(247);
			33538: out = 16'(-161);
			33539: out = 16'(-2791);
			33540: out = 16'(-3131);
			33541: out = 16'(-2797);
			33542: out = 16'(-248);
			33543: out = 16'(669);
			33544: out = 16'(893);
			33545: out = 16'(-772);
			33546: out = 16'(-1551);
			33547: out = 16'(-1737);
			33548: out = 16'(-206);
			33549: out = 16'(997);
			33550: out = 16'(1880);
			33551: out = 16'(1037);
			33552: out = 16'(79);
			33553: out = 16'(-626);
			33554: out = 16'(-845);
			33555: out = 16'(-472);
			33556: out = 16'(764);
			33557: out = 16'(1425);
			33558: out = 16'(1825);
			33559: out = 16'(468);
			33560: out = 16'(554);
			33561: out = 16'(900);
			33562: out = 16'(1612);
			33563: out = 16'(1617);
			33564: out = 16'(1199);
			33565: out = 16'(548);
			33566: out = 16'(64);
			33567: out = 16'(-245);
			33568: out = 16'(103);
			33569: out = 16'(268);
			33570: out = 16'(137);
			33571: out = 16'(-837);
			33572: out = 16'(-1432);
			33573: out = 16'(-321);
			33574: out = 16'(-414);
			33575: out = 16'(-329);
			33576: out = 16'(-857);
			33577: out = 16'(-1011);
			33578: out = 16'(-1491);
			33579: out = 16'(-1148);
			33580: out = 16'(-2005);
			33581: out = 16'(-2898);
			33582: out = 16'(-2505);
			33583: out = 16'(-1676);
			33584: out = 16'(-551);
			33585: out = 16'(-93);
			33586: out = 16'(518);
			33587: out = 16'(2149);
			33588: out = 16'(868);
			33589: out = 16'(252);
			33590: out = 16'(-829);
			33591: out = 16'(1704);
			33592: out = 16'(3486);
			33593: out = 16'(3218);
			33594: out = 16'(1586);
			33595: out = 16'(-447);
			33596: out = 16'(296);
			33597: out = 16'(528);
			33598: out = 16'(1416);
			33599: out = 16'(-77);
			33600: out = 16'(-216);
			33601: out = 16'(-411);
			33602: out = 16'(-319);
			33603: out = 16'(-335);
			33604: out = 16'(-141);
			33605: out = 16'(-215);
			33606: out = 16'(-360);
			33607: out = 16'(-1443);
			33608: out = 16'(-955);
			33609: out = 16'(-834);
			33610: out = 16'(-706);
			33611: out = 16'(-1660);
			33612: out = 16'(-2367);
			33613: out = 16'(-1263);
			33614: out = 16'(-1217);
			33615: out = 16'(-1101);
			33616: out = 16'(-759);
			33617: out = 16'(-311);
			33618: out = 16'(116);
			33619: out = 16'(47);
			33620: out = 16'(90);
			33621: out = 16'(44);
			33622: out = 16'(367);
			33623: out = 16'(171);
			33624: out = 16'(-648);
			33625: out = 16'(30);
			33626: out = 16'(770);
			33627: out = 16'(1929);
			33628: out = 16'(1464);
			33629: out = 16'(646);
			33630: out = 16'(-483);
			33631: out = 16'(-848);
			33632: out = 16'(-421);
			33633: out = 16'(609);
			33634: out = 16'(1905);
			33635: out = 16'(2753);
			33636: out = 16'(2888);
			33637: out = 16'(1434);
			33638: out = 16'(-1038);
			33639: out = 16'(-1221);
			33640: out = 16'(-1044);
			33641: out = 16'(337);
			33642: out = 16'(107);
			33643: out = 16'(268);
			33644: out = 16'(120);
			33645: out = 16'(275);
			33646: out = 16'(-16);
			33647: out = 16'(-750);
			33648: out = 16'(-1160);
			33649: out = 16'(-1510);
			33650: out = 16'(-2339);
			33651: out = 16'(-2449);
			33652: out = 16'(-2145);
			33653: out = 16'(42);
			33654: out = 16'(1002);
			33655: out = 16'(1428);
			33656: out = 16'(574);
			33657: out = 16'(178);
			33658: out = 16'(361);
			33659: out = 16'(297);
			33660: out = 16'(758);
			33661: out = 16'(1305);
			33662: out = 16'(2028);
			33663: out = 16'(1987);
			33664: out = 16'(841);
			33665: out = 16'(117);
			33666: out = 16'(-427);
			33667: out = 16'(132);
			33668: out = 16'(177);
			33669: out = 16'(382);
			33670: out = 16'(1133);
			33671: out = 16'(1057);
			33672: out = 16'(623);
			33673: out = 16'(326);
			33674: out = 16'(135);
			33675: out = 16'(235);
			33676: out = 16'(-259);
			33677: out = 16'(-56);
			33678: out = 16'(745);
			33679: out = 16'(-67);
			33680: out = 16'(-278);
			33681: out = 16'(34);
			33682: out = 16'(172);
			33683: out = 16'(-302);
			33684: out = 16'(-3141);
			33685: out = 16'(-3127);
			33686: out = 16'(-2888);
			33687: out = 16'(-373);
			33688: out = 16'(-1313);
			33689: out = 16'(-2479);
			33690: out = 16'(-1399);
			33691: out = 16'(-576);
			33692: out = 16'(637);
			33693: out = 16'(-163);
			33694: out = 16'(-66);
			33695: out = 16'(-58);
			33696: out = 16'(1483);
			33697: out = 16'(1605);
			33698: out = 16'(126);
			33699: out = 16'(336);
			33700: out = 16'(358);
			33701: out = 16'(1524);
			33702: out = 16'(568);
			33703: out = 16'(-28);
			33704: out = 16'(-2017);
			33705: out = 16'(-315);
			33706: out = 16'(1015);
			33707: out = 16'(1397);
			33708: out = 16'(-102);
			33709: out = 16'(-2132);
			33710: out = 16'(-1841);
			33711: out = 16'(-1242);
			33712: out = 16'(123);
			33713: out = 16'(647);
			33714: out = 16'(706);
			33715: out = 16'(-382);
			33716: out = 16'(-553);
			33717: out = 16'(-490);
			33718: out = 16'(1083);
			33719: out = 16'(486);
			33720: out = 16'(217);
			33721: out = 16'(-1419);
			33722: out = 16'(-482);
			33723: out = 16'(-129);
			33724: out = 16'(79);
			33725: out = 16'(-1244);
			33726: out = 16'(-2439);
			33727: out = 16'(-1805);
			33728: out = 16'(-1095);
			33729: out = 16'(140);
			33730: out = 16'(1131);
			33731: out = 16'(2135);
			33732: out = 16'(2813);
			33733: out = 16'(1024);
			33734: out = 16'(242);
			33735: out = 16'(519);
			33736: out = 16'(343);
			33737: out = 16'(55);
			33738: out = 16'(-2038);
			33739: out = 16'(-298);
			33740: out = 16'(683);
			33741: out = 16'(1947);
			33742: out = 16'(343);
			33743: out = 16'(-805);
			33744: out = 16'(284);
			33745: out = 16'(1484);
			33746: out = 16'(2710);
			33747: out = 16'(114);
			33748: out = 16'(-873);
			33749: out = 16'(-2029);
			33750: out = 16'(-519);
			33751: out = 16'(-56);
			33752: out = 16'(470);
			33753: out = 16'(220);
			33754: out = 16'(158);
			33755: out = 16'(-397);
			33756: out = 16'(576);
			33757: out = 16'(931);
			33758: out = 16'(1415);
			33759: out = 16'(27);
			33760: out = 16'(-1274);
			33761: out = 16'(-2945);
			33762: out = 16'(-1921);
			33763: out = 16'(-415);
			33764: out = 16'(49);
			33765: out = 16'(429);
			33766: out = 16'(251);
			33767: out = 16'(1326);
			33768: out = 16'(1342);
			33769: out = 16'(1377);
			33770: out = 16'(434);
			33771: out = 16'(74);
			33772: out = 16'(-187);
			33773: out = 16'(-141);
			33774: out = 16'(-92);
			33775: out = 16'(404);
			33776: out = 16'(-12);
			33777: out = 16'(-483);
			33778: out = 16'(-2507);
			33779: out = 16'(-1453);
			33780: out = 16'(-533);
			33781: out = 16'(883);
			33782: out = 16'(336);
			33783: out = 16'(-457);
			33784: out = 16'(-2725);
			33785: out = 16'(-2071);
			33786: out = 16'(-435);
			33787: out = 16'(1458);
			33788: out = 16'(1738);
			33789: out = 16'(832);
			33790: out = 16'(474);
			33791: out = 16'(513);
			33792: out = 16'(1436);
			33793: out = 16'(1687);
			33794: out = 16'(1382);
			33795: out = 16'(-305);
			33796: out = 16'(-1628);
			33797: out = 16'(-2277);
			33798: out = 16'(274);
			33799: out = 16'(248);
			33800: out = 16'(447);
			33801: out = 16'(-182);
			33802: out = 16'(142);
			33803: out = 16'(174);
			33804: out = 16'(288);
			33805: out = 16'(31);
			33806: out = 16'(-111);
			33807: out = 16'(-1124);
			33808: out = 16'(-1198);
			33809: out = 16'(-730);
			33810: out = 16'(453);
			33811: out = 16'(812);
			33812: out = 16'(-214);
			33813: out = 16'(207);
			33814: out = 16'(471);
			33815: out = 16'(1925);
			33816: out = 16'(837);
			33817: out = 16'(-192);
			33818: out = 16'(-2362);
			33819: out = 16'(-1651);
			33820: out = 16'(-538);
			33821: out = 16'(225);
			33822: out = 16'(488);
			33823: out = 16'(328);
			33824: out = 16'(-517);
			33825: out = 16'(-1179);
			33826: out = 16'(-1830);
			33827: out = 16'(-26);
			33828: out = 16'(558);
			33829: out = 16'(425);
			33830: out = 16'(68);
			33831: out = 16'(303);
			33832: out = 16'(1916);
			33833: out = 16'(1535);
			33834: out = 16'(1152);
			33835: out = 16'(217);
			33836: out = 16'(153);
			33837: out = 16'(172);
			33838: out = 16'(123);
			33839: out = 16'(266);
			33840: out = 16'(325);
			33841: out = 16'(1221);
			33842: out = 16'(656);
			33843: out = 16'(-528);
			33844: out = 16'(-774);
			33845: out = 16'(-461);
			33846: out = 16'(963);
			33847: out = 16'(-572);
			33848: out = 16'(-789);
			33849: out = 16'(-368);
			33850: out = 16'(-202);
			33851: out = 16'(-316);
			33852: out = 16'(-821);
			33853: out = 16'(-917);
			33854: out = 16'(-560);
			33855: out = 16'(742);
			33856: out = 16'(891);
			33857: out = 16'(718);
			33858: out = 16'(314);
			33859: out = 16'(-369);
			33860: out = 16'(-898);
			33861: out = 16'(-886);
			33862: out = 16'(-568);
			33863: out = 16'(-116);
			33864: out = 16'(-164);
			33865: out = 16'(-57);
			33866: out = 16'(269);
			33867: out = 16'(126);
			33868: out = 16'(218);
			33869: out = 16'(-293);
			33870: out = 16'(1178);
			33871: out = 16'(1795);
			33872: out = 16'(1819);
			33873: out = 16'(222);
			33874: out = 16'(-1167);
			33875: out = 16'(-1393);
			33876: out = 16'(-636);
			33877: out = 16'(514);
			33878: out = 16'(666);
			33879: out = 16'(612);
			33880: out = 16'(3);
			33881: out = 16'(178);
			33882: out = 16'(77);
			33883: out = 16'(102);
			33884: out = 16'(-616);
			33885: out = 16'(-1289);
			33886: out = 16'(-1912);
			33887: out = 16'(-2394);
			33888: out = 16'(-1938);
			33889: out = 16'(-113);
			33890: out = 16'(516);
			33891: out = 16'(693);
			33892: out = 16'(-1278);
			33893: out = 16'(-1307);
			33894: out = 16'(-1072);
			33895: out = 16'(773);
			33896: out = 16'(1378);
			33897: out = 16'(1875);
			33898: out = 16'(520);
			33899: out = 16'(364);
			33900: out = 16'(356);
			33901: out = 16'(1164);
			33902: out = 16'(1318);
			33903: out = 16'(1293);
			33904: out = 16'(853);
			33905: out = 16'(869);
			33906: out = 16'(1198);
			33907: out = 16'(967);
			33908: out = 16'(117);
			33909: out = 16'(-1907);
			33910: out = 16'(-2776);
			33911: out = 16'(-2765);
			33912: out = 16'(-365);
			33913: out = 16'(822);
			33914: out = 16'(1786);
			33915: out = 16'(-86);
			33916: out = 16'(-639);
			33917: out = 16'(-1548);
			33918: out = 16'(-350);
			33919: out = 16'(-461);
			33920: out = 16'(-182);
			33921: out = 16'(-1353);
			33922: out = 16'(-731);
			33923: out = 16'(295);
			33924: out = 16'(2192);
			33925: out = 16'(2081);
			33926: out = 16'(-340);
			33927: out = 16'(-1399);
			33928: out = 16'(-1641);
			33929: out = 16'(275);
			33930: out = 16'(1156);
			33931: out = 16'(1728);
			33932: out = 16'(927);
			33933: out = 16'(-511);
			33934: out = 16'(-2247);
			33935: out = 16'(-2894);
			33936: out = 16'(-2004);
			33937: out = 16'(280);
			33938: out = 16'(488);
			33939: out = 16'(1014);
			33940: out = 16'(124);
			33941: out = 16'(1391);
			33942: out = 16'(743);
			33943: out = 16'(-174);
			33944: out = 16'(-2288);
			33945: out = 16'(-2668);
			33946: out = 16'(-735);
			33947: out = 16'(240);
			33948: out = 16'(1033);
			33949: out = 16'(815);
			33950: out = 16'(675);
			33951: out = 16'(306);
			33952: out = 16'(381);
			33953: out = 16'(727);
			33954: out = 16'(1320);
			33955: out = 16'(427);
			33956: out = 16'(-222);
			33957: out = 16'(-1461);
			33958: out = 16'(0);
			33959: out = 16'(130);
			33960: out = 16'(274);
			33961: out = 16'(-1330);
			33962: out = 16'(-1709);
			33963: out = 16'(-1273);
			33964: out = 16'(121);
			33965: out = 16'(1108);
			33966: out = 16'(1262);
			33967: out = 16'(543);
			33968: out = 16'(-249);
			33969: out = 16'(301);
			33970: out = 16'(123);
			33971: out = 16'(222);
			33972: out = 16'(-327);
			33973: out = 16'(-149);
			33974: out = 16'(-129);
			33975: out = 16'(1113);
			33976: out = 16'(816);
			33977: out = 16'(-290);
			33978: out = 16'(184);
			33979: out = 16'(22);
			33980: out = 16'(-123);
			33981: out = 16'(-971);
			33982: out = 16'(-1301);
			33983: out = 16'(-697);
			33984: out = 16'(-833);
			33985: out = 16'(-592);
			33986: out = 16'(-362);
			33987: out = 16'(675);
			33988: out = 16'(1336);
			33989: out = 16'(377);
			33990: out = 16'(324);
			33991: out = 16'(189);
			33992: out = 16'(782);
			33993: out = 16'(764);
			33994: out = 16'(778);
			33995: out = 16'(-35);
			33996: out = 16'(-229);
			33997: out = 16'(-353);
			33998: out = 16'(53);
			33999: out = 16'(124);
			34000: out = 16'(193);
			34001: out = 16'(-880);
			34002: out = 16'(-1316);
			34003: out = 16'(-780);
			34004: out = 16'(-409);
			34005: out = 16'(-187);
			34006: out = 16'(-1291);
			34007: out = 16'(-1013);
			34008: out = 16'(-543);
			34009: out = 16'(697);
			34010: out = 16'(1109);
			34011: out = 16'(1243);
			34012: out = 16'(532);
			34013: out = 16'(-67);
			34014: out = 16'(-806);
			34015: out = 16'(-338);
			34016: out = 16'(76);
			34017: out = 16'(928);
			34018: out = 16'(54);
			34019: out = 16'(-605);
			34020: out = 16'(-1808);
			34021: out = 16'(-725);
			34022: out = 16'(-23);
			34023: out = 16'(444);
			34024: out = 16'(64);
			34025: out = 16'(-216);
			34026: out = 16'(-245);
			34027: out = 16'(352);
			34028: out = 16'(972);
			34029: out = 16'(1291);
			34030: out = 16'(766);
			34031: out = 16'(-236);
			34032: out = 16'(246);
			34033: out = 16'(81);
			34034: out = 16'(-98);
			34035: out = 16'(202);
			34036: out = 16'(378);
			34037: out = 16'(329);
			34038: out = 16'(264);
			34039: out = 16'(190);
			34040: out = 16'(333);
			34041: out = 16'(327);
			34042: out = 16'(168);
			34043: out = 16'(-745);
			34044: out = 16'(-1066);
			34045: out = 16'(-1312);
			34046: out = 16'(-746);
			34047: out = 16'(-976);
			34048: out = 16'(-1177);
			34049: out = 16'(-229);
			34050: out = 16'(151);
			34051: out = 16'(444);
			34052: out = 16'(304);
			34053: out = 16'(133);
			34054: out = 16'(-270);
			34055: out = 16'(266);
			34056: out = 16'(407);
			34057: out = 16'(413);
			34058: out = 16'(-13);
			34059: out = 16'(-226);
			34060: out = 16'(-106);
			34061: out = 16'(659);
			34062: out = 16'(1492);
			34063: out = 16'(1575);
			34064: out = 16'(1758);
			34065: out = 16'(1504);
			34066: out = 16'(1329);
			34067: out = 16'(685);
			34068: out = 16'(199);
			34069: out = 16'(-330);
			34070: out = 16'(-270);
			34071: out = 16'(54);
			34072: out = 16'(119);
			34073: out = 16'(-241);
			34074: out = 16'(-886);
			34075: out = 16'(-1295);
			34076: out = 16'(-1053);
			34077: out = 16'(260);
			34078: out = 16'(560);
			34079: out = 16'(542);
			34080: out = 16'(-811);
			34081: out = 16'(-1120);
			34082: out = 16'(-1311);
			34083: out = 16'(-383);
			34084: out = 16'(-240);
			34085: out = 16'(-134);
			34086: out = 16'(-304);
			34087: out = 16'(-288);
			34088: out = 16'(-324);
			34089: out = 16'(171);
			34090: out = 16'(-501);
			34091: out = 16'(-2477);
			34092: out = 16'(-1078);
			34093: out = 16'(-458);
			34094: out = 16'(527);
			34095: out = 16'(-688);
			34096: out = 16'(-1243);
			34097: out = 16'(-1278);
			34098: out = 16'(-264);
			34099: out = 16'(733);
			34100: out = 16'(2128);
			34101: out = 16'(1563);
			34102: out = 16'(575);
			34103: out = 16'(-1057);
			34104: out = 16'(-775);
			34105: out = 16'(429);
			34106: out = 16'(997);
			34107: out = 16'(1379);
			34108: out = 16'(1125);
			34109: out = 16'(609);
			34110: out = 16'(-142);
			34111: out = 16'(-835);
			34112: out = 16'(-891);
			34113: out = 16'(-638);
			34114: out = 16'(198);
			34115: out = 16'(-478);
			34116: out = 16'(-696);
			34117: out = 16'(321);
			34118: out = 16'(551);
			34119: out = 16'(774);
			34120: out = 16'(172);
			34121: out = 16'(-59);
			34122: out = 16'(-441);
			34123: out = 16'(-696);
			34124: out = 16'(-1091);
			34125: out = 16'(-1203);
			34126: out = 16'(725);
			34127: out = 16'(1585);
			34128: out = 16'(1551);
			34129: out = 16'(724);
			34130: out = 16'(-514);
			34131: out = 16'(-1177);
			34132: out = 16'(-1889);
			34133: out = 16'(-1259);
			34134: out = 16'(135);
			34135: out = 16'(2039);
			34136: out = 16'(2922);
			34137: out = 16'(2195);
			34138: out = 16'(511);
			34139: out = 16'(-1176);
			34140: out = 16'(-1339);
			34141: out = 16'(-928);
			34142: out = 16'(-94);
			34143: out = 16'(181);
			34144: out = 16'(-104);
			34145: out = 16'(-942);
			34146: out = 16'(-1655);
			34147: out = 16'(-1607);
			34148: out = 16'(-721);
			34149: out = 16'(316);
			34150: out = 16'(1203);
			34151: out = 16'(2142);
			34152: out = 16'(874);
			34153: out = 16'(-167);
			34154: out = 16'(-837);
			34155: out = 16'(-307);
			34156: out = 16'(8);
			34157: out = 16'(-1201);
			34158: out = 16'(-2148);
			34159: out = 16'(-2832);
			34160: out = 16'(-1491);
			34161: out = 16'(-285);
			34162: out = 16'(1004);
			34163: out = 16'(497);
			34164: out = 16'(-114);
			34165: out = 16'(-1318);
			34166: out = 16'(-1192);
			34167: out = 16'(-825);
			34168: out = 16'(398);
			34169: out = 16'(262);
			34170: out = 16'(304);
			34171: out = 16'(-66);
			34172: out = 16'(531);
			34173: out = 16'(1086);
			34174: out = 16'(1229);
			34175: out = 16'(1863);
			34176: out = 16'(2131);
			34177: out = 16'(2253);
			34178: out = 16'(718);
			34179: out = 16'(-1082);
			34180: out = 16'(-298);
			34181: out = 16'(-440);
			34182: out = 16'(-305);
			34183: out = 16'(-821);
			34184: out = 16'(-514);
			34185: out = 16'(208);
			34186: out = 16'(-105);
			34187: out = 16'(-183);
			34188: out = 16'(-338);
			34189: out = 16'(5);
			34190: out = 16'(365);
			34191: out = 16'(1306);
			34192: out = 16'(550);
			34193: out = 16'(93);
			34194: out = 16'(90);
			34195: out = 16'(474);
			34196: out = 16'(706);
			34197: out = 16'(318);
			34198: out = 16'(148);
			34199: out = 16'(49);
			34200: out = 16'(-2103);
			34201: out = 16'(-2028);
			34202: out = 16'(-1205);
			34203: out = 16'(398);
			34204: out = 16'(488);
			34205: out = 16'(-891);
			34206: out = 16'(-727);
			34207: out = 16'(-419);
			34208: out = 16'(890);
			34209: out = 16'(1341);
			34210: out = 16'(1739);
			34211: out = 16'(1180);
			34212: out = 16'(525);
			34213: out = 16'(-452);
			34214: out = 16'(-129);
			34215: out = 16'(-774);
			34216: out = 16'(-729);
			34217: out = 16'(-1468);
			34218: out = 16'(-328);
			34219: out = 16'(819);
			34220: out = 16'(905);
			34221: out = 16'(-125);
			34222: out = 16'(-1909);
			34223: out = 16'(-2608);
			34224: out = 16'(-2478);
			34225: out = 16'(-1124);
			34226: out = 16'(-559);
			34227: out = 16'(8);
			34228: out = 16'(340);
			34229: out = 16'(-581);
			34230: out = 16'(-982);
			34231: out = 16'(916);
			34232: out = 16'(1577);
			34233: out = 16'(2258);
			34234: out = 16'(278);
			34235: out = 16'(777);
			34236: out = 16'(1310);
			34237: out = 16'(1324);
			34238: out = 16'(675);
			34239: out = 16'(-424);
			34240: out = 16'(145);
			34241: out = 16'(-16);
			34242: out = 16'(-313);
			34243: out = 16'(-702);
			34244: out = 16'(-595);
			34245: out = 16'(239);
			34246: out = 16'(-41);
			34247: out = 16'(-81);
			34248: out = 16'(337);
			34249: out = 16'(563);
			34250: out = 16'(740);
			34251: out = 16'(-332);
			34252: out = 16'(-161);
			34253: out = 16'(-200);
			34254: out = 16'(842);
			34255: out = 16'(-323);
			34256: out = 16'(-1957);
			34257: out = 16'(-1824);
			34258: out = 16'(-1121);
			34259: out = 16'(391);
			34260: out = 16'(152);
			34261: out = 16'(282);
			34262: out = 16'(195);
			34263: out = 16'(357);
			34264: out = 16'(451);
			34265: out = 16'(812);
			34266: out = 16'(821);
			34267: out = 16'(678);
			34268: out = 16'(263);
			34269: out = 16'(-660);
			34270: out = 16'(-1323);
			34271: out = 16'(-183);
			34272: out = 16'(230);
			34273: out = 16'(899);
			34274: out = 16'(-183);
			34275: out = 16'(437);
			34276: out = 16'(1207);
			34277: out = 16'(188);
			34278: out = 16'(-1089);
			34279: out = 16'(-2954);
			34280: out = 16'(-2090);
			34281: out = 16'(-1215);
			34282: out = 16'(300);
			34283: out = 16'(231);
			34284: out = 16'(236);
			34285: out = 16'(-127);
			34286: out = 16'(216);
			34287: out = 16'(395);
			34288: out = 16'(373);
			34289: out = 16'(574);
			34290: out = 16'(817);
			34291: out = 16'(-172);
			34292: out = 16'(-843);
			34293: out = 16'(-1915);
			34294: out = 16'(108);
			34295: out = 16'(127);
			34296: out = 16'(359);
			34297: out = 16'(-2742);
			34298: out = 16'(-2774);
			34299: out = 16'(-1131);
			34300: out = 16'(1629);
			34301: out = 16'(2488);
			34302: out = 16'(319);
			34303: out = 16'(113);
			34304: out = 16'(-179);
			34305: out = 16'(401);
			34306: out = 16'(1374);
			34307: out = 16'(2366);
			34308: out = 16'(2535);
			34309: out = 16'(1548);
			34310: out = 16'(-78);
			34311: out = 16'(-1013);
			34312: out = 16'(-1321);
			34313: out = 16'(-631);
			34314: out = 16'(-146);
			34315: out = 16'(236);
			34316: out = 16'(-298);
			34317: out = 16'(249);
			34318: out = 16'(-162);
			34319: out = 16'(-748);
			34320: out = 16'(-1216);
			34321: out = 16'(-1022);
			34322: out = 16'(-156);
			34323: out = 16'(487);
			34324: out = 16'(808);
			34325: out = 16'(243);
			34326: out = 16'(-276);
			34327: out = 16'(-793);
			34328: out = 16'(380);
			34329: out = 16'(82);
			34330: out = 16'(-150);
			34331: out = 16'(-1157);
			34332: out = 16'(-750);
			34333: out = 16'(374);
			34334: out = 16'(643);
			34335: out = 16'(1053);
			34336: out = 16'(1229);
			34337: out = 16'(580);
			34338: out = 16'(-377);
			34339: out = 16'(-1805);
			34340: out = 16'(-807);
			34341: out = 16'(518);
			34342: out = 16'(2417);
			34343: out = 16'(2401);
			34344: out = 16'(1815);
			34345: out = 16'(1368);
			34346: out = 16'(335);
			34347: out = 16'(-353);
			34348: out = 16'(-875);
			34349: out = 16'(-721);
			34350: out = 16'(-384);
			34351: out = 16'(-228);
			34352: out = 16'(-316);
			34353: out = 16'(-381);
			34354: out = 16'(-2777);
			34355: out = 16'(-3480);
			34356: out = 16'(-2739);
			34357: out = 16'(-1829);
			34358: out = 16'(-746);
			34359: out = 16'(-97);
			34360: out = 16'(-5);
			34361: out = 16'(-118);
			34362: out = 16'(529);
			34363: out = 16'(353);
			34364: out = 16'(131);
			34365: out = 16'(-2072);
			34366: out = 16'(-1732);
			34367: out = 16'(-906);
			34368: out = 16'(683);
			34369: out = 16'(1072);
			34370: out = 16'(915);
			34371: out = 16'(968);
			34372: out = 16'(1028);
			34373: out = 16'(1417);
			34374: out = 16'(606);
			34375: out = 16'(471);
			34376: out = 16'(894);
			34377: out = 16'(534);
			34378: out = 16'(232);
			34379: out = 16'(-132);
			34380: out = 16'(159);
			34381: out = 16'(286);
			34382: out = 16'(-765);
			34383: out = 16'(-529);
			34384: out = 16'(-94);
			34385: out = 16'(1154);
			34386: out = 16'(1307);
			34387: out = 16'(1169);
			34388: out = 16'(-31);
			34389: out = 16'(-729);
			34390: out = 16'(-1343);
			34391: out = 16'(-125);
			34392: out = 16'(307);
			34393: out = 16'(324);
			34394: out = 16'(7);
			34395: out = 16'(-308);
			34396: out = 16'(-798);
			34397: out = 16'(-754);
			34398: out = 16'(-675);
			34399: out = 16'(317);
			34400: out = 16'(-674);
			34401: out = 16'(-1205);
			34402: out = 16'(-874);
			34403: out = 16'(714);
			34404: out = 16'(2371);
			34405: out = 16'(1746);
			34406: out = 16'(633);
			34407: out = 16'(-1610);
			34408: out = 16'(153);
			34409: out = 16'(-67);
			34410: out = 16'(28);
			34411: out = 16'(-479);
			34412: out = 16'(529);
			34413: out = 16'(2019);
			34414: out = 16'(2820);
			34415: out = 16'(2442);
			34416: out = 16'(1309);
			34417: out = 16'(-830);
			34418: out = 16'(-1948);
			34419: out = 16'(-1017);
			34420: out = 16'(228);
			34421: out = 16'(1158);
			34422: out = 16'(243);
			34423: out = 16'(-1315);
			34424: out = 16'(-3174);
			34425: out = 16'(-2936);
			34426: out = 16'(-1830);
			34427: out = 16'(502);
			34428: out = 16'(-325);
			34429: out = 16'(-284);
			34430: out = 16'(-851);
			34431: out = 16'(-188);
			34432: out = 16'(104);
			34433: out = 16'(938);
			34434: out = 16'(198);
			34435: out = 16'(-371);
			34436: out = 16'(-1765);
			34437: out = 16'(-893);
			34438: out = 16'(-25);
			34439: out = 16'(198);
			34440: out = 16'(112);
			34441: out = 16'(-270);
			34442: out = 16'(460);
			34443: out = 16'(279);
			34444: out = 16'(357);
			34445: out = 16'(121);
			34446: out = 16'(732);
			34447: out = 16'(1253);
			34448: out = 16'(1415);
			34449: out = 16'(729);
			34450: out = 16'(-239);
			34451: out = 16'(-1470);
			34452: out = 16'(-1451);
			34453: out = 16'(-195);
			34454: out = 16'(1333);
			34455: out = 16'(2243);
			34456: out = 16'(2158);
			34457: out = 16'(520);
			34458: out = 16'(-1049);
			34459: out = 16'(161);
			34460: out = 16'(144);
			34461: out = 16'(319);
			34462: out = 16'(180);
			34463: out = 16'(-249);
			34464: out = 16'(-915);
			34465: out = 16'(-2062);
			34466: out = 16'(-1649);
			34467: out = 16'(448);
			34468: out = 16'(-144);
			34469: out = 16'(-19);
			34470: out = 16'(-359);
			34471: out = 16'(566);
			34472: out = 16'(767);
			34473: out = 16'(385);
			34474: out = 16'(-272);
			34475: out = 16'(-770);
			34476: out = 16'(254);
			34477: out = 16'(-21);
			34478: out = 16'(-50);
			34479: out = 16'(-255);
			34480: out = 16'(723);
			34481: out = 16'(1765);
			34482: out = 16'(1686);
			34483: out = 16'(1131);
			34484: out = 16'(12);
			34485: out = 16'(-227);
			34486: out = 16'(-302);
			34487: out = 16'(176);
			34488: out = 16'(487);
			34489: out = 16'(968);
			34490: out = 16'(1545);
			34491: out = 16'(787);
			34492: out = 16'(-221);
			34493: out = 16'(-1241);
			34494: out = 16'(-2057);
			34495: out = 16'(-2369);
			34496: out = 16'(-1886);
			34497: out = 16'(-1571);
			34498: out = 16'(-1140);
			34499: out = 16'(-416);
			34500: out = 16'(-91);
			34501: out = 16'(-88);
			34502: out = 16'(697);
			34503: out = 16'(860);
			34504: out = 16'(821);
			34505: out = 16'(-295);
			34506: out = 16'(-1114);
			34507: out = 16'(-1728);
			34508: out = 16'(-1099);
			34509: out = 16'(-492);
			34510: out = 16'(-277);
			34511: out = 16'(231);
			34512: out = 16'(499);
			34513: out = 16'(872);
			34514: out = 16'(596);
			34515: out = 16'(170);
			34516: out = 16'(303);
			34517: out = 16'(2);
			34518: out = 16'(-343);
			34519: out = 16'(-1449);
			34520: out = 16'(-1972);
			34521: out = 16'(-2142);
			34522: out = 16'(-333);
			34523: out = 16'(1068);
			34524: out = 16'(2236);
			34525: out = 16'(1992);
			34526: out = 16'(1197);
			34527: out = 16'(-766);
			34528: out = 16'(-142);
			34529: out = 16'(405);
			34530: out = 16'(798);
			34531: out = 16'(597);
			34532: out = 16'(286);
			34533: out = 16'(262);
			34534: out = 16'(-70);
			34535: out = 16'(-290);
			34536: out = 16'(-148);
			34537: out = 16'(-141);
			34538: out = 16'(-129);
			34539: out = 16'(-254);
			34540: out = 16'(-225);
			34541: out = 16'(-103);
			34542: out = 16'(-136);
			34543: out = 16'(-132);
			34544: out = 16'(-276);
			34545: out = 16'(-170);
			34546: out = 16'(101);
			34547: out = 16'(1284);
			34548: out = 16'(924);
			34549: out = 16'(627);
			34550: out = 16'(-348);
			34551: out = 16'(-1);
			34552: out = 16'(346);
			34553: out = 16'(1134);
			34554: out = 16'(729);
			34555: out = 16'(-6);
			34556: out = 16'(-172);
			34557: out = 16'(-132);
			34558: out = 16'(234);
			34559: out = 16'(-992);
			34560: out = 16'(-1817);
			34561: out = 16'(-2374);
			34562: out = 16'(-2074);
			34563: out = 16'(-1555);
			34564: out = 16'(-1373);
			34565: out = 16'(-88);
			34566: out = 16'(365);
			34567: out = 16'(-31);
			34568: out = 16'(-144);
			34569: out = 16'(52);
			34570: out = 16'(-276);
			34571: out = 16'(963);
			34572: out = 16'(1741);
			34573: out = 16'(2342);
			34574: out = 16'(445);
			34575: out = 16'(-2047);
			34576: out = 16'(-3193);
			34577: out = 16'(-2358);
			34578: out = 16'(197);
			34579: out = 16'(1557);
			34580: out = 16'(2310);
			34581: out = 16'(1616);
			34582: out = 16'(484);
			34583: out = 16'(-713);
			34584: out = 16'(-1230);
			34585: out = 16'(-357);
			34586: out = 16'(497);
			34587: out = 16'(-238);
			34588: out = 16'(-107);
			34589: out = 16'(-342);
			34590: out = 16'(-54);
			34591: out = 16'(-17);
			34592: out = 16'(306);
			34593: out = 16'(90);
			34594: out = 16'(678);
			34595: out = 16'(1277);
			34596: out = 16'(452);
			34597: out = 16'(-632);
			34598: out = 16'(-2490);
			34599: out = 16'(-639);
			34600: out = 16'(150);
			34601: out = 16'(893);
			34602: out = 16'(-518);
			34603: out = 16'(-1760);
			34604: out = 16'(-3387);
			34605: out = 16'(-1832);
			34606: out = 16'(-238);
			34607: out = 16'(350);
			34608: out = 16'(505);
			34609: out = 16'(297);
			34610: out = 16'(315);
			34611: out = 16'(940);
			34612: out = 16'(1993);
			34613: out = 16'(2054);
			34614: out = 16'(1993);
			34615: out = 16'(1078);
			34616: out = 16'(1058);
			34617: out = 16'(392);
			34618: out = 16'(298);
			34619: out = 16'(-1449);
			34620: out = 16'(-1382);
			34621: out = 16'(290);
			34622: out = 16'(1207);
			34623: out = 16'(1449);
			34624: out = 16'(-333);
			34625: out = 16'(-639);
			34626: out = 16'(-802);
			34627: out = 16'(-225);
			34628: out = 16'(6);
			34629: out = 16'(111);
			34630: out = 16'(-207);
			34631: out = 16'(-968);
			34632: out = 16'(-1893);
			34633: out = 16'(-1810);
			34634: out = 16'(-1148);
			34635: out = 16'(432);
			34636: out = 16'(131);
			34637: out = 16'(349);
			34638: out = 16'(156);
			34639: out = 16'(1635);
			34640: out = 16'(2254);
			34641: out = 16'(2108);
			34642: out = 16'(999);
			34643: out = 16'(-275);
			34644: out = 16'(-636);
			34645: out = 16'(-1297);
			34646: out = 16'(-1190);
			34647: out = 16'(-1512);
			34648: out = 16'(4);
			34649: out = 16'(1454);
			34650: out = 16'(2406);
			34651: out = 16'(2066);
			34652: out = 16'(1058);
			34653: out = 16'(70);
			34654: out = 16'(-366);
			34655: out = 16'(-383);
			34656: out = 16'(-232);
			34657: out = 16'(-234);
			34658: out = 16'(251);
			34659: out = 16'(-1967);
			34660: out = 16'(-2962);
			34661: out = 16'(-2375);
			34662: out = 16'(-528);
			34663: out = 16'(1080);
			34664: out = 16'(279);
			34665: out = 16'(162);
			34666: out = 16'(-368);
			34667: out = 16'(-53);
			34668: out = 16'(-6);
			34669: out = 16'(287);
			34670: out = 16'(187);
			34671: out = 16'(53);
			34672: out = 16'(-324);
			34673: out = 16'(-1027);
			34674: out = 16'(-1071);
			34675: out = 16'(-133);
			34676: out = 16'(24);
			34677: out = 16'(297);
			34678: out = 16'(-171);
			34679: out = 16'(295);
			34680: out = 16'(414);
			34681: out = 16'(914);
			34682: out = 16'(262);
			34683: out = 16'(-89);
			34684: out = 16'(283);
			34685: out = 16'(975);
			34686: out = 16'(1751);
			34687: out = 16'(845);
			34688: out = 16'(534);
			34689: out = 16'(109);
			34690: out = 16'(1355);
			34691: out = 16'(2012);
			34692: out = 16'(2888);
			34693: out = 16'(413);
			34694: out = 16'(-1262);
			34695: out = 16'(-3068);
			34696: out = 16'(-1674);
			34697: out = 16'(-536);
			34698: out = 16'(21);
			34699: out = 16'(5);
			34700: out = 16'(-505);
			34701: out = 16'(-1705);
			34702: out = 16'(-2160);
			34703: out = 16'(-2151);
			34704: out = 16'(-312);
			34705: out = 16'(71);
			34706: out = 16'(255);
			34707: out = 16'(-680);
			34708: out = 16'(-153);
			34709: out = 16'(980);
			34710: out = 16'(1826);
			34711: out = 16'(2008);
			34712: out = 16'(1085);
			34713: out = 16'(287);
			34714: out = 16'(-919);
			34715: out = 16'(-1685);
			34716: out = 16'(-1969);
			34717: out = 16'(-1551);
			34718: out = 16'(-1427);
			34719: out = 16'(-457);
			34720: out = 16'(95);
			34721: out = 16'(1780);
			34722: out = 16'(970);
			34723: out = 16'(208);
			34724: out = 16'(-375);
			34725: out = 16'(942);
			34726: out = 16'(2663);
			34727: out = 16'(2602);
			34728: out = 16'(1400);
			34729: out = 16'(-1087);
			34730: out = 16'(-1578);
			34731: out = 16'(-1746);
			34732: out = 16'(-769);
			34733: out = 16'(-261);
			34734: out = 16'(300);
			34735: out = 16'(227);
			34736: out = 16'(-24);
			34737: out = 16'(-596);
			34738: out = 16'(-1704);
			34739: out = 16'(-1010);
			34740: out = 16'(-213);
			34741: out = 16'(-1180);
			34742: out = 16'(-1578);
			34743: out = 16'(-2162);
			34744: out = 16'(-407);
			34745: out = 16'(16);
			34746: out = 16'(375);
			34747: out = 16'(302);
			34748: out = 16'(968);
			34749: out = 16'(2165);
			34750: out = 16'(1461);
			34751: out = 16'(896);
			34752: out = 16'(-208);
			34753: out = 16'(767);
			34754: out = 16'(1112);
			34755: out = 16'(243);
			34756: out = 16'(-8);
			34757: out = 16'(-379);
			34758: out = 16'(224);
			34759: out = 16'(-380);
			34760: out = 16'(-779);
			34761: out = 16'(-411);
			34762: out = 16'(345);
			34763: out = 16'(1241);
			34764: out = 16'(357);
			34765: out = 16'(240);
			34766: out = 16'(90);
			34767: out = 16'(141);
			34768: out = 16'(-36);
			34769: out = 16'(-345);
			34770: out = 16'(-664);
			34771: out = 16'(-840);
			34772: out = 16'(-756);
			34773: out = 16'(-818);
			34774: out = 16'(-644);
			34775: out = 16'(-166);
			34776: out = 16'(346);
			34777: out = 16'(816);
			34778: out = 16'(124);
			34779: out = 16'(489);
			34780: out = 16'(758);
			34781: out = 16'(1137);
			34782: out = 16'(765);
			34783: out = 16'(-23);
			34784: out = 16'(-567);
			34785: out = 16'(-1340);
			34786: out = 16'(-2276);
			34787: out = 16'(-518);
			34788: out = 16'(691);
			34789: out = 16'(1583);
			34790: out = 16'(1344);
			34791: out = 16'(840);
			34792: out = 16'(-200);
			34793: out = 16'(-200);
			34794: out = 16'(-250);
			34795: out = 16'(-287);
			34796: out = 16'(-638);
			34797: out = 16'(-776);
			34798: out = 16'(-863);
			34799: out = 16'(-336);
			34800: out = 16'(243);
			34801: out = 16'(1438);
			34802: out = 16'(1122);
			34803: out = 16'(129);
			34804: out = 16'(-896);
			34805: out = 16'(-1291);
			34806: out = 16'(-690);
			34807: out = 16'(-84);
			34808: out = 16'(419);
			34809: out = 16'(197);
			34810: out = 16'(59);
			34811: out = 16'(-229);
			34812: out = 16'(267);
			34813: out = 16'(-464);
			34814: out = 16'(-770);
			34815: out = 16'(-843);
			34816: out = 16'(-202);
			34817: out = 16'(334);
			34818: out = 16'(-124);
			34819: out = 16'(-23);
			34820: out = 16'(205);
			34821: out = 16'(-163);
			34822: out = 16'(31);
			34823: out = 16'(285);
			34824: out = 16'(697);
			34825: out = 16'(340);
			34826: out = 16'(-799);
			34827: out = 16'(-1119);
			34828: out = 16'(-960);
			34829: out = 16'(352);
			34830: out = 16'(301);
			34831: out = 16'(267);
			34832: out = 16'(-257);
			34833: out = 16'(-517);
			34834: out = 16'(-693);
			34835: out = 16'(294);
			34836: out = 16'(322);
			34837: out = 16'(320);
			34838: out = 16'(-206);
			34839: out = 16'(-112);
			34840: out = 16'(200);
			34841: out = 16'(193);
			34842: out = 16'(-100);
			34843: out = 16'(-814);
			34844: out = 16'(-384);
			34845: out = 16'(-36);
			34846: out = 16'(864);
			34847: out = 16'(657);
			34848: out = 16'(982);
			34849: out = 16'(1458);
			34850: out = 16'(2115);
			34851: out = 16'(2084);
			34852: out = 16'(826);
			34853: out = 16'(-425);
			34854: out = 16'(-1673);
			34855: out = 16'(-3112);
			34856: out = 16'(-3212);
			34857: out = 16'(-2483);
			34858: out = 16'(115);
			34859: out = 16'(1436);
			34860: out = 16'(1986);
			34861: out = 16'(374);
			34862: out = 16'(-203);
			34863: out = 16'(416);
			34864: out = 16'(182);
			34865: out = 16'(271);
			34866: out = 16'(-292);
			34867: out = 16'(166);
			34868: out = 16'(-383);
			34869: out = 16'(-2595);
			34870: out = 16'(-2830);
			34871: out = 16'(-2337);
			34872: out = 16'(-464);
			34873: out = 16'(434);
			34874: out = 16'(903);
			34875: out = 16'(1292);
			34876: out = 16'(904);
			34877: out = 16'(265);
			34878: out = 16'(-1231);
			34879: out = 16'(-1917);
			34880: out = 16'(-2079);
			34881: out = 16'(-695);
			34882: out = 16'(27);
			34883: out = 16'(-225);
			34884: out = 16'(594);
			34885: out = 16'(1113);
			34886: out = 16'(1711);
			34887: out = 16'(1481);
			34888: out = 16'(1110);
			34889: out = 16'(883);
			34890: out = 16'(226);
			34891: out = 16'(-379);
			34892: out = 16'(-683);
			34893: out = 16'(-360);
			34894: out = 16'(262);
			34895: out = 16'(-652);
			34896: out = 16'(-698);
			34897: out = 16'(-688);
			34898: out = 16'(-174);
			34899: out = 16'(-58);
			34900: out = 16'(-66);
			34901: out = 16'(-74);
			34902: out = 16'(-51);
			34903: out = 16'(-86);
			34904: out = 16'(240);
			34905: out = 16'(402);
			34906: out = 16'(382);
			34907: out = 16'(68);
			34908: out = 16'(-244);
			34909: out = 16'(229);
			34910: out = 16'(292);
			34911: out = 16'(246);
			34912: out = 16'(-1437);
			34913: out = 16'(-2084);
			34914: out = 16'(-2629);
			34915: out = 16'(-536);
			34916: out = 16'(130);
			34917: out = 16'(542);
			34918: out = 16'(30);
			34919: out = 16'(342);
			34920: out = 16'(864);
			34921: out = 16'(1575);
			34922: out = 16'(1511);
			34923: out = 16'(962);
			34924: out = 16'(-450);
			34925: out = 16'(-1124);
			34926: out = 16'(-739);
			34927: out = 16'(648);
			34928: out = 16'(1899);
			34929: out = 16'(2038);
			34930: out = 16'(1117);
			34931: out = 16'(-323);
			34932: out = 16'(273);
			34933: out = 16'(176);
			34934: out = 16'(348);
			34935: out = 16'(-62);
			34936: out = 16'(-320);
			34937: out = 16'(-768);
			34938: out = 16'(-1411);
			34939: out = 16'(-1702);
			34940: out = 16'(-1610);
			34941: out = 16'(-599);
			34942: out = 16'(247);
			34943: out = 16'(819);
			34944: out = 16'(378);
			34945: out = 16'(-42);
			34946: out = 16'(844);
			34947: out = 16'(990);
			34948: out = 16'(1206);
			34949: out = 16'(-581);
			34950: out = 16'(-511);
			34951: out = 16'(-191);
			34952: out = 16'(290);
			34953: out = 16'(224);
			34954: out = 16'(-135);
			34955: out = 16'(201);
			34956: out = 16'(-139);
			34957: out = 16'(-1269);
			34958: out = 16'(-62);
			34959: out = 16'(765);
			34960: out = 16'(2107);
			34961: out = 16'(673);
			34962: out = 16'(-233);
			34963: out = 16'(370);
			34964: out = 16'(254);
			34965: out = 16'(149);
			34966: out = 16'(-1580);
			34967: out = 16'(-1734);
			34968: out = 16'(-1507);
			34969: out = 16'(62);
			34970: out = 16'(810);
			34971: out = 16'(1226);
			34972: out = 16'(891);
			34973: out = 16'(590);
			34974: out = 16'(157);
			34975: out = 16'(169);
			34976: out = 16'(160);
			34977: out = 16'(173);
			34978: out = 16'(-404);
			34979: out = 16'(-942);
			34980: out = 16'(-1139);
			34981: out = 16'(-1510);
			34982: out = 16'(-1575);
			34983: out = 16'(-1212);
			34984: out = 16'(-559);
			34985: out = 16'(191);
			34986: out = 16'(1086);
			34987: out = 16'(1709);
			34988: out = 16'(2006);
			34989: out = 16'(579);
			34990: out = 16'(-519);
			34991: out = 16'(-1767);
			34992: out = 16'(-863);
			34993: out = 16'(-465);
			34994: out = 16'(351);
			34995: out = 16'(-818);
			34996: out = 16'(-1040);
			34997: out = 16'(-701);
			34998: out = 16'(605);
			34999: out = 16'(1439);
			35000: out = 16'(1675);
			35001: out = 16'(680);
			35002: out = 16'(-550);
			35003: out = 16'(-1579);
			35004: out = 16'(-923);
			35005: out = 16'(448);
			35006: out = 16'(-208);
			35007: out = 16'(136);
			35008: out = 16'(157);
			35009: out = 16'(277);
			35010: out = 16'(54);
			35011: out = 16'(-60);
			35012: out = 16'(162);
			35013: out = 16'(342);
			35014: out = 16'(-259);
			35015: out = 16'(870);
			35016: out = 16'(955);
			35017: out = 16'(-92);
			35018: out = 16'(-1083);
			35019: out = 16'(-1653);
			35020: out = 16'(-271);
			35021: out = 16'(23);
			35022: out = 16'(386);
			35023: out = 16'(-705);
			35024: out = 16'(-458);
			35025: out = 16'(-265);
			35026: out = 16'(-174);
			35027: out = 16'(-599);
			35028: out = 16'(-1165);
			35029: out = 16'(-476);
			35030: out = 16'(324);
			35031: out = 16'(1305);
			35032: out = 16'(1297);
			35033: out = 16'(929);
			35034: out = 16'(-139);
			35035: out = 16'(103);
			35036: out = 16'(175);
			35037: out = 16'(-163);
			35038: out = 16'(410);
			35039: out = 16'(761);
			35040: out = 16'(313);
			35041: out = 16'(96);
			35042: out = 16'(-138);
			35043: out = 16'(655);
			35044: out = 16'(897);
			35045: out = 16'(1167);
			35046: out = 16'(291);
			35047: out = 16'(-84);
			35048: out = 16'(-390);
			35049: out = 16'(-193);
			35050: out = 16'(-259);
			35051: out = 16'(-307);
			35052: out = 16'(-709);
			35053: out = 16'(-653);
			35054: out = 16'(-180);
			35055: out = 16'(633);
			35056: out = 16'(1218);
			35057: out = 16'(649);
			35058: out = 16'(496);
			35059: out = 16'(356);
			35060: out = 16'(2669);
			35061: out = 16'(2097);
			35062: out = 16'(1126);
			35063: out = 16'(-2342);
			35064: out = 16'(-2873);
			35065: out = 16'(-2167);
			35066: out = 16'(-460);
			35067: out = 16'(217);
			35068: out = 16'(-334);
			35069: out = 16'(571);
			35070: out = 16'(536);
			35071: out = 16'(101);
			35072: out = 16'(-817);
			35073: out = 16'(-1379);
			35074: out = 16'(-658);
			35075: out = 16'(-1729);
			35076: out = 16'(-2310);
			35077: out = 16'(-2745);
			35078: out = 16'(-1642);
			35079: out = 16'(-383);
			35080: out = 16'(134);
			35081: out = 16'(257);
			35082: out = 16'(-11);
			35083: out = 16'(727);
			35084: out = 16'(1489);
			35085: out = 16'(2596);
			35086: out = 16'(1489);
			35087: out = 16'(642);
			35088: out = 16'(-896);
			35089: out = 16'(-304);
			35090: out = 16'(-452);
			35091: out = 16'(-653);
			35092: out = 16'(-1417);
			35093: out = 16'(-1443);
			35094: out = 16'(-250);
			35095: out = 16'(-66);
			35096: out = 16'(-56);
			35097: out = 16'(359);
			35098: out = 16'(-677);
			35099: out = 16'(-1705);
			35100: out = 16'(-1157);
			35101: out = 16'(-546);
			35102: out = 16'(442);
			35103: out = 16'(-93);
			35104: out = 16'(-518);
			35105: out = 16'(-1650);
			35106: out = 16'(119);
			35107: out = 16'(873);
			35108: out = 16'(1892);
			35109: out = 16'(714);
			35110: out = 16'(346);
			35111: out = 16'(400);
			35112: out = 16'(1000);
			35113: out = 16'(1181);
			35114: out = 16'(337);
			35115: out = 16'(-273);
			35116: out = 16'(-638);
			35117: out = 16'(-149);
			35118: out = 16'(570);
			35119: out = 16'(1376);
			35120: out = 16'(1600);
			35121: out = 16'(1185);
			35122: out = 16'(197);
			35123: out = 16'(243);
			35124: out = 16'(412);
			35125: out = 16'(1304);
			35126: out = 16'(1633);
			35127: out = 16'(2015);
			35128: out = 16'(1274);
			35129: out = 16'(1944);
			35130: out = 16'(1291);
			35131: out = 16'(-97);
			35132: out = 16'(-2226);
			35133: out = 16'(-3443);
			35134: out = 16'(-2395);
			35135: out = 16'(-1111);
			35136: out = 16'(258);
			35137: out = 16'(-1244);
			35138: out = 16'(-1356);
			35139: out = 16'(-1732);
			35140: out = 16'(-19);
			35141: out = 16'(141);
			35142: out = 16'(-120);
			35143: out = 16'(-509);
			35144: out = 16'(-1094);
			35145: out = 16'(-2225);
			35146: out = 16'(-730);
			35147: out = 16'(-13);
			35148: out = 16'(-41);
			35149: out = 16'(205);
			35150: out = 16'(304);
			35151: out = 16'(-79);
			35152: out = 16'(933);
			35153: out = 16'(1788);
			35154: out = 16'(1239);
			35155: out = 16'(697);
			35156: out = 16'(-288);
			35157: out = 16'(445);
			35158: out = 16'(22);
			35159: out = 16'(-47);
			35160: out = 16'(-1499);
			35161: out = 16'(-1325);
			35162: out = 16'(-685);
			35163: out = 16'(156);
			35164: out = 16'(567);
			35165: out = 16'(1401);
			35166: out = 16'(-121);
			35167: out = 16'(-930);
			35168: out = 16'(-2324);
			35169: out = 16'(227);
			35170: out = 16'(1951);
			35171: out = 16'(2562);
			35172: out = 16'(137);
			35173: out = 16'(-2585);
			35174: out = 16'(-2536);
			35175: out = 16'(-1543);
			35176: out = 16'(621);
			35177: out = 16'(-279);
			35178: out = 16'(-186);
			35179: out = 16'(-731);
			35180: out = 16'(321);
			35181: out = 16'(334);
			35182: out = 16'(-27);
			35183: out = 16'(628);
			35184: out = 16'(810);
			35185: out = 16'(421);
			35186: out = 16'(-520);
			35187: out = 16'(-1142);
			35188: out = 16'(-107);
			35189: out = 16'(74);
			35190: out = 16'(552);
			35191: out = 16'(150);
			35192: out = 16'(635);
			35193: out = 16'(908);
			35194: out = 16'(2349);
			35195: out = 16'(1960);
			35196: out = 16'(1103);
			35197: out = 16'(1506);
			35198: out = 16'(1654);
			35199: out = 16'(1890);
			35200: out = 16'(353);
			35201: out = 16'(-966);
			35202: out = 16'(-2302);
			35203: out = 16'(-2407);
			35204: out = 16'(-1928);
			35205: out = 16'(-826);
			35206: out = 16'(-325);
			35207: out = 16'(-123);
			35208: out = 16'(-209);
			35209: out = 16'(-791);
			35210: out = 16'(-1095);
			35211: out = 16'(238);
			35212: out = 16'(604);
			35213: out = 16'(687);
			35214: out = 16'(-848);
			35215: out = 16'(-1664);
			35216: out = 16'(-2086);
			35217: out = 16'(-1434);
			35218: out = 16'(-626);
			35219: out = 16'(-42);
			35220: out = 16'(1646);
			35221: out = 16'(1865);
			35222: out = 16'(310);
			35223: out = 16'(368);
			35224: out = 16'(295);
			35225: out = 16'(845);
			35226: out = 16'(773);
			35227: out = 16'(697);
			35228: out = 16'(-92);
			35229: out = 16'(51);
			35230: out = 16'(177);
			35231: out = 16'(-268);
			35232: out = 16'(-261);
			35233: out = 16'(-259);
			35234: out = 16'(160);
			35235: out = 16'(15);
			35236: out = 16'(-235);
			35237: out = 16'(-221);
			35238: out = 16'(498);
			35239: out = 16'(2092);
			35240: out = 16'(1169);
			35241: out = 16'(212);
			35242: out = 16'(-1220);
			35243: out = 16'(-1585);
			35244: out = 16'(-1766);
			35245: out = 16'(-2241);
			35246: out = 16'(-1356);
			35247: out = 16'(-396);
			35248: out = 16'(755);
			35249: out = 16'(486);
			35250: out = 16'(-179);
			35251: out = 16'(-510);
			35252: out = 16'(-712);
			35253: out = 16'(-614);
			35254: out = 16'(-644);
			35255: out = 16'(-620);
			35256: out = 16'(-610);
			35257: out = 16'(-947);
			35258: out = 16'(-1160);
			35259: out = 16'(-1557);
			35260: out = 16'(-545);
			35261: out = 16'(138);
			35262: out = 16'(559);
			35263: out = 16'(485);
			35264: out = 16'(675);
			35265: out = 16'(777);
			35266: out = 16'(2062);
			35267: out = 16'(3027);
			35268: out = 16'(2999);
			35269: out = 16'(1528);
			35270: out = 16'(-560);
			35271: out = 16'(-563);
			35272: out = 16'(-539);
			35273: out = 16'(291);
			35274: out = 16'(-1331);
			35275: out = 16'(-2008);
			35276: out = 16'(-2686);
			35277: out = 16'(-1616);
			35278: out = 16'(-613);
			35279: out = 16'(413);
			35280: out = 16'(1572);
			35281: out = 16'(2040);
			35282: out = 16'(342);
			35283: out = 16'(441);
			35284: out = 16'(129);
			35285: out = 16'(561);
			35286: out = 16'(-460);
			35287: out = 16'(-1117);
			35288: out = 16'(-445);
			35289: out = 16'(969);
			35290: out = 16'(2588);
			35291: out = 16'(1434);
			35292: out = 16'(718);
			35293: out = 16'(-206);
			35294: out = 16'(108);
			35295: out = 16'(169);
			35296: out = 16'(107);
			35297: out = 16'(241);
			35298: out = 16'(-457);
			35299: out = 16'(-2702);
			35300: out = 16'(-2773);
			35301: out = 16'(-2174);
			35302: out = 16'(270);
			35303: out = 16'(1129);
			35304: out = 16'(1670);
			35305: out = 16'(14);
			35306: out = 16'(-79);
			35307: out = 16'(-7);
			35308: out = 16'(1450);
			35309: out = 16'(1675);
			35310: out = 16'(1550);
			35311: out = 16'(146);
			35312: out = 16'(-836);
			35313: out = 16'(-1758);
			35314: out = 16'(-662);
			35315: out = 16'(-170);
			35316: out = 16'(-301);
			35317: out = 16'(-510);
			35318: out = 16'(-708);
			35319: out = 16'(-170);
			35320: out = 16'(-39);
			35321: out = 16'(325);
			35322: out = 16'(-192);
			35323: out = 16'(467);
			35324: out = 16'(728);
			35325: out = 16'(520);
			35326: out = 16'(-565);
			35327: out = 16'(-1747);
			35328: out = 16'(-1710);
			35329: out = 16'(-781);
			35330: out = 16'(1016);
			35331: out = 16'(81);
			35332: out = 16'(-74);
			35333: out = 16'(-191);
			35334: out = 16'(111);
			35335: out = 16'(329);
			35336: out = 16'(184);
			35337: out = 16'(932);
			35338: out = 16'(1456);
			35339: out = 16'(2502);
			35340: out = 16'(1204);
			35341: out = 16'(-233);
			35342: out = 16'(-1558);
			35343: out = 16'(-1174);
			35344: out = 16'(-34);
			35345: out = 16'(-30);
			35346: out = 16'(531);
			35347: out = 16'(768);
			35348: out = 16'(1848);
			35349: out = 16'(1498);
			35350: out = 16'(63);
			35351: out = 16'(-39);
			35352: out = 16'(-682);
			35353: out = 16'(-637);
			35354: out = 16'(-2608);
			35355: out = 16'(-3140);
			35356: out = 16'(-2246);
			35357: out = 16'(-622);
			35358: out = 16'(751);
			35359: out = 16'(1622);
			35360: out = 16'(829);
			35361: out = 16'(-353);
			35362: out = 16'(-1026);
			35363: out = 16'(-860);
			35364: out = 16'(26);
			35365: out = 16'(1314);
			35366: out = 16'(1677);
			35367: out = 16'(1032);
			35368: out = 16'(-93);
			35369: out = 16'(-1505);
			35370: out = 16'(-2563);
			35371: out = 16'(-2379);
			35372: out = 16'(-1504);
			35373: out = 16'(-142);
			35374: out = 16'(38);
			35375: out = 16'(90);
			35376: out = 16'(562);
			35377: out = 16'(176);
			35378: out = 16'(71);
			35379: out = 16'(-85);
			35380: out = 16'(935);
			35381: out = 16'(1720);
			35382: out = 16'(555);
			35383: out = 16'(-881);
			35384: out = 16'(-2740);
			35385: out = 16'(-823);
			35386: out = 16'(-366);
			35387: out = 16'(154);
			35388: out = 16'(-481);
			35389: out = 16'(-212);
			35390: out = 16'(510);
			35391: out = 16'(815);
			35392: out = 16'(794);
			35393: out = 16'(8);
			35394: out = 16'(39);
			35395: out = 16'(-118);
			35396: out = 16'(-1044);
			35397: out = 16'(-364);
			35398: out = 16'(609);
			35399: out = 16'(1184);
			35400: out = 16'(1255);
			35401: out = 16'(765);
			35402: out = 16'(1372);
			35403: out = 16'(844);
			35404: out = 16'(420);
			35405: out = 16'(245);
			35406: out = 16'(937);
			35407: out = 16'(2008);
			35408: out = 16'(1535);
			35409: out = 16'(464);
			35410: out = 16'(-1158);
			35411: out = 16'(-2588);
			35412: out = 16'(-3201);
			35413: out = 16'(-2688);
			35414: out = 16'(-1169);
			35415: out = 16'(354);
			35416: out = 16'(712);
			35417: out = 16'(989);
			35418: out = 16'(821);
			35419: out = 16'(870);
			35420: out = 16'(1006);
			35421: out = 16'(1231);
			35422: out = 16'(144);
			35423: out = 16'(-86);
			35424: out = 16'(306);
			35425: out = 16'(-1273);
			35426: out = 16'(-1670);
			35427: out = 16'(-1657);
			35428: out = 16'(100);
			35429: out = 16'(1074);
			35430: out = 16'(1265);
			35431: out = 16'(680);
			35432: out = 16'(135);
			35433: out = 16'(-108);
			35434: out = 16'(611);
			35435: out = 16'(1259);
			35436: out = 16'(809);
			35437: out = 16'(305);
			35438: out = 16'(-421);
			35439: out = 16'(-1456);
			35440: out = 16'(-1721);
			35441: out = 16'(-1582);
			35442: out = 16'(621);
			35443: out = 16'(1737);
			35444: out = 16'(2475);
			35445: out = 16'(521);
			35446: out = 16'(-751);
			35447: out = 16'(-1723);
			35448: out = 16'(-107);
			35449: out = 16'(1010);
			35450: out = 16'(1179);
			35451: out = 16'(-98);
			35452: out = 16'(-1632);
			35453: out = 16'(-2032);
			35454: out = 16'(-2324);
			35455: out = 16'(-1907);
			35456: out = 16'(97);
			35457: out = 16'(313);
			35458: out = 16'(-128);
			35459: out = 16'(-122);
			35460: out = 16'(120);
			35461: out = 16'(945);
			35462: out = 16'(779);
			35463: out = 16'(712);
			35464: out = 16'(168);
			35465: out = 16'(48);
			35466: out = 16'(-160);
			35467: out = 16'(-85);
			35468: out = 16'(66);
			35469: out = 16'(255);
			35470: out = 16'(151);
			35471: out = 16'(328);
			35472: out = 16'(260);
			35473: out = 16'(-195);
			35474: out = 16'(-328);
			35475: out = 16'(-126);
			35476: out = 16'(952);
			35477: out = 16'(1452);
			35478: out = 16'(1465);
			35479: out = 16'(201);
			35480: out = 16'(-1126);
			35481: out = 16'(-2232);
			35482: out = 16'(-2687);
			35483: out = 16'(-2201);
			35484: out = 16'(-642);
			35485: out = 16'(304);
			35486: out = 16'(1041);
			35487: out = 16'(727);
			35488: out = 16'(1175);
			35489: out = 16'(1229);
			35490: out = 16'(1693);
			35491: out = 16'(879);
			35492: out = 16'(-177);
			35493: out = 16'(-2428);
			35494: out = 16'(-2429);
			35495: out = 16'(-1428);
			35496: out = 16'(-980);
			35497: out = 16'(-306);
			35498: out = 16'(-269);
			35499: out = 16'(811);
			35500: out = 16'(542);
			35501: out = 16'(17);
			35502: out = 16'(-928);
			35503: out = 16'(-747);
			35504: out = 16'(375);
			35505: out = 16'(1579);
			35506: out = 16'(1916);
			35507: out = 16'(390);
			35508: out = 16'(-468);
			35509: out = 16'(-1330);
			35510: out = 16'(-1121);
			35511: out = 16'(-670);
			35512: out = 16'(83);
			35513: out = 16'(-222);
			35514: out = 16'(-310);
			35515: out = 16'(-667);
			35516: out = 16'(663);
			35517: out = 16'(907);
			35518: out = 16'(821);
			35519: out = 16'(103);
			35520: out = 16'(-454);
			35521: out = 16'(-594);
			35522: out = 16'(-1072);
			35523: out = 16'(-815);
			35524: out = 16'(247);
			35525: out = 16'(652);
			35526: out = 16'(784);
			35527: out = 16'(410);
			35528: out = 16'(570);
			35529: out = 16'(785);
			35530: out = 16'(-108);
			35531: out = 16'(162);
			35532: out = 16'(203);
			35533: out = 16'(1543);
			35534: out = 16'(838);
			35535: out = 16'(-197);
			35536: out = 16'(-2162);
			35537: out = 16'(-1922);
			35538: out = 16'(-34);
			35539: out = 16'(491);
			35540: out = 16'(746);
			35541: out = 16'(199);
			35542: out = 16'(-94);
			35543: out = 16'(-102);
			35544: out = 16'(286);
			35545: out = 16'(1522);
			35546: out = 16'(2437);
			35547: out = 16'(2259);
			35548: out = 16'(1208);
			35549: out = 16'(-318);
			35550: out = 16'(-1876);
			35551: out = 16'(-1726);
			35552: out = 16'(-496);
			35553: out = 16'(-856);
			35554: out = 16'(-725);
			35555: out = 16'(-1224);
			35556: out = 16'(127);
			35557: out = 16'(650);
			35558: out = 16'(1688);
			35559: out = 16'(256);
			35560: out = 16'(-118);
			35561: out = 16'(-198);
			35562: out = 16'(752);
			35563: out = 16'(924);
			35564: out = 16'(-206);
			35565: out = 16'(-822);
			35566: out = 16'(-1123);
			35567: out = 16'(-780);
			35568: out = 16'(-215);
			35569: out = 16'(201);
			35570: out = 16'(297);
			35571: out = 16'(-574);
			35572: out = 16'(-1600);
			35573: out = 16'(-1258);
			35574: out = 16'(-161);
			35575: out = 16'(1687);
			35576: out = 16'(1033);
			35577: out = 16'(-2);
			35578: out = 16'(-2085);
			35579: out = 16'(-2349);
			35580: out = 16'(-2058);
			35581: out = 16'(-91);
			35582: out = 16'(209);
			35583: out = 16'(478);
			35584: out = 16'(-29);
			35585: out = 16'(45);
			35586: out = 16'(67);
			35587: out = 16'(792);
			35588: out = 16'(860);
			35589: out = 16'(782);
			35590: out = 16'(504);
			35591: out = 16'(-7);
			35592: out = 16'(-654);
			35593: out = 16'(-1002);
			35594: out = 16'(-710);
			35595: out = 16'(417);
			35596: out = 16'(282);
			35597: out = 16'(762);
			35598: out = 16'(1560);
			35599: out = 16'(1871);
			35600: out = 16'(1748);
			35601: out = 16'(712);
			35602: out = 16'(275);
			35603: out = 16'(-364);
			35604: out = 16'(-535);
			35605: out = 16'(-1488);
			35606: out = 16'(-2068);
			35607: out = 16'(-2124);
			35608: out = 16'(-1142);
			35609: out = 16'(89);
			35610: out = 16'(-28);
			35611: out = 16'(-311);
			35612: out = 16'(-1096);
			35613: out = 16'(-662);
			35614: out = 16'(-374);
			35615: out = 16'(49);
			35616: out = 16'(866);
			35617: out = 16'(1215);
			35618: out = 16'(337);
			35619: out = 16'(425);
			35620: out = 16'(195);
			35621: out = 16'(486);
			35622: out = 16'(19);
			35623: out = 16'(-135);
			35624: out = 16'(-296);
			35625: out = 16'(681);
			35626: out = 16'(1646);
			35627: out = 16'(858);
			35628: out = 16'(381);
			35629: out = 16'(-315);
			35630: out = 16'(-65);
			35631: out = 16'(-152);
			35632: out = 16'(-229);
			35633: out = 16'(-266);
			35634: out = 16'(10);
			35635: out = 16'(798);
			35636: out = 16'(155);
			35637: out = 16'(-142);
			35638: out = 16'(-151);
			35639: out = 16'(593);
			35640: out = 16'(1142);
			35641: out = 16'(105);
			35642: out = 16'(259);
			35643: out = 16'(270);
			35644: out = 16'(1090);
			35645: out = 16'(299);
			35646: out = 16'(-922);
			35647: out = 16'(-672);
			35648: out = 16'(-691);
			35649: out = 16'(-213);
			35650: out = 16'(-1783);
			35651: out = 16'(-1746);
			35652: out = 16'(-577);
			35653: out = 16'(-299);
			35654: out = 16'(83);
			35655: out = 16'(172);
			35656: out = 16'(611);
			35657: out = 16'(666);
			35658: out = 16'(-110);
			35659: out = 16'(97);
			35660: out = 16'(205);
			35661: out = 16'(358);
			35662: out = 16'(45);
			35663: out = 16'(-256);
			35664: out = 16'(-165);
			35665: out = 16'(384);
			35666: out = 16'(1235);
			35667: out = 16'(1390);
			35668: out = 16'(1307);
			35669: out = 16'(507);
			35670: out = 16'(393);
			35671: out = 16'(-308);
			35672: out = 16'(-664);
			35673: out = 16'(-1802);
			35674: out = 16'(-1946);
			35675: out = 16'(-1232);
			35676: out = 16'(-304);
			35677: out = 16'(246);
			35678: out = 16'(249);
			35679: out = 16'(-729);
			35680: out = 16'(-1738);
			35681: out = 16'(-1964);
			35682: out = 16'(-1078);
			35683: out = 16'(625);
			35684: out = 16'(877);
			35685: out = 16'(1728);
			35686: out = 16'(1809);
			35687: out = 16'(1834);
			35688: out = 16'(696);
			35689: out = 16'(-693);
			35690: out = 16'(-2119);
			35691: out = 16'(-2493);
			35692: out = 16'(-2029);
			35693: out = 16'(-214);
			35694: out = 16'(1226);
			35695: out = 16'(1442);
			35696: out = 16'(1688);
			35697: out = 16'(1314);
			35698: out = 16'(483);
			35699: out = 16'(-258);
			35700: out = 16'(-698);
			35701: out = 16'(106);
			35702: out = 16'(71);
			35703: out = 16'(-125);
			35704: out = 16'(123);
			35705: out = 16'(374);
			35706: out = 16'(759);
			35707: out = 16'(1270);
			35708: out = 16'(1645);
			35709: out = 16'(1807);
			35710: out = 16'(1551);
			35711: out = 16'(1164);
			35712: out = 16'(562);
			35713: out = 16'(265);
			35714: out = 16'(-311);
			35715: out = 16'(-1212);
			35716: out = 16'(-1859);
			35717: out = 16'(-2236);
			35718: out = 16'(-2192);
			35719: out = 16'(-1722);
			35720: out = 16'(-987);
			35721: out = 16'(-69);
			35722: out = 16'(501);
			35723: out = 16'(682);
			35724: out = 16'(73);
			35725: out = 16'(-503);
			35726: out = 16'(-1168);
			35727: out = 16'(-811);
			35728: out = 16'(-499);
			35729: out = 16'(-55);
			35730: out = 16'(-174);
			35731: out = 16'(-512);
			35732: out = 16'(-2110);
			35733: out = 16'(-911);
			35734: out = 16'(126);
			35735: out = 16'(1189);
			35736: out = 16'(528);
			35737: out = 16'(-323);
			35738: out = 16'(-575);
			35739: out = 16'(-51);
			35740: out = 16'(924);
			35741: out = 16'(-26);
			35742: out = 16'(102);
			35743: out = 16'(224);
			35744: out = 16'(384);
			35745: out = 16'(78);
			35746: out = 16'(-704);
			35747: out = 16'(16);
			35748: out = 16'(281);
			35749: out = 16'(404);
			35750: out = 16'(-299);
			35751: out = 16'(-600);
			35752: out = 16'(-66);
			35753: out = 16'(601);
			35754: out = 16'(1280);
			35755: out = 16'(668);
			35756: out = 16'(822);
			35757: out = 16'(587);
			35758: out = 16'(376);
			35759: out = 16'(-663);
			35760: out = 16'(-1657);
			35761: out = 16'(-867);
			35762: out = 16'(-329);
			35763: out = 16'(227);
			35764: out = 16'(632);
			35765: out = 16'(751);
			35766: out = 16'(738);
			35767: out = 16'(391);
			35768: out = 16'(587);
			35769: out = 16'(1888);
			35770: out = 16'(1410);
			35771: out = 16'(467);
			35772: out = 16'(-2503);
			35773: out = 16'(-2440);
			35774: out = 16'(-1806);
			35775: out = 16'(-99);
			35776: out = 16'(729);
			35777: out = 16'(1197);
			35778: out = 16'(1452);
			35779: out = 16'(1359);
			35780: out = 16'(1013);
			35781: out = 16'(1075);
			35782: out = 16'(992);
			35783: out = 16'(1005);
			35784: out = 16'(396);
			35785: out = 16'(-131);
			35786: out = 16'(-879);
			35787: out = 16'(-1088);
			35788: out = 16'(-1592);
			35789: out = 16'(-2572);
			35790: out = 16'(-2708);
			35791: out = 16'(-2151);
			35792: out = 16'(-7);
			35793: out = 16'(960);
			35794: out = 16'(1606);
			35795: out = 16'(1164);
			35796: out = 16'(630);
			35797: out = 16'(-332);
			35798: out = 16'(307);
			35799: out = 16'(-741);
			35800: out = 16'(-2152);
			35801: out = 16'(-1387);
			35802: out = 16'(-757);
			35803: out = 16'(-64);
			35804: out = 16'(220);
			35805: out = 16'(603);
			35806: out = 16'(1635);
			35807: out = 16'(466);
			35808: out = 16'(-293);
			35809: out = 16'(-674);
			35810: out = 16'(-216);
			35811: out = 16'(184);
			35812: out = 16'(-186);
			35813: out = 16'(-873);
			35814: out = 16'(-1697);
			35815: out = 16'(-1526);
			35816: out = 16'(-903);
			35817: out = 16'(499);
			35818: out = 16'(-153);
			35819: out = 16'(490);
			35820: out = 16'(1194);
			35821: out = 16'(1855);
			35822: out = 16'(1641);
			35823: out = 16'(692);
			35824: out = 16'(445);
			35825: out = 16'(249);
			35826: out = 16'(198);
			35827: out = 16'(-322);
			35828: out = 16'(-818);
			35829: out = 16'(-570);
			35830: out = 16'(-1212);
			35831: out = 16'(-1570);
			35832: out = 16'(-2043);
			35833: out = 16'(-1146);
			35834: out = 16'(66);
			35835: out = 16'(665);
			35836: out = 16'(871);
			35837: out = 16'(808);
			35838: out = 16'(122);
			35839: out = 16'(179);
			35840: out = 16'(831);
			35841: out = 16'(1344);
			35842: out = 16'(1336);
			35843: out = 16'(135);
			35844: out = 16'(-326);
			35845: out = 16'(-665);
			35846: out = 16'(268);
			35847: out = 16'(-117);
			35848: out = 16'(-266);
			35849: out = 16'(-666);
			35850: out = 16'(-632);
			35851: out = 16'(-619);
			35852: out = 16'(144);
			35853: out = 16'(451);
			35854: out = 16'(786);
			35855: out = 16'(-821);
			35856: out = 16'(-1104);
			35857: out = 16'(-1071);
			35858: out = 16'(363);
			35859: out = 16'(785);
			35860: out = 16'(328);
			35861: out = 16'(312);
			35862: out = 16'(248);
			35863: out = 16'(348);
			35864: out = 16'(812);
			35865: out = 16'(1261);
			35866: out = 16'(1479);
			35867: out = 16'(1116);
			35868: out = 16'(511);
			35869: out = 16'(236);
			35870: out = 16'(-78);
			35871: out = 16'(-150);
			35872: out = 16'(41);
			35873: out = 16'(136);
			35874: out = 16'(48);
			35875: out = 16'(-210);
			35876: out = 16'(-380);
			35877: out = 16'(-279);
			35878: out = 16'(44);
			35879: out = 16'(311);
			35880: out = 16'(23);
			35881: out = 16'(198);
			35882: out = 16'(-22);
			35883: out = 16'(262);
			35884: out = 16'(-1240);
			35885: out = 16'(-2071);
			35886: out = 16'(-809);
			35887: out = 16'(-196);
			35888: out = 16'(270);
			35889: out = 16'(-939);
			35890: out = 16'(-1546);
			35891: out = 16'(-1970);
			35892: out = 16'(-460);
			35893: out = 16'(612);
			35894: out = 16'(1611);
			35895: out = 16'(1607);
			35896: out = 16'(1164);
			35897: out = 16'(141);
			35898: out = 16'(-701);
			35899: out = 16'(-1189);
			35900: out = 16'(-577);
			35901: out = 16'(-1022);
			35902: out = 16'(-907);
			35903: out = 16'(-149);
			35904: out = 16'(379);
			35905: out = 16'(840);
			35906: out = 16'(305);
			35907: out = 16'(741);
			35908: out = 16'(1105);
			35909: out = 16'(422);
			35910: out = 16'(19);
			35911: out = 16'(-321);
			35912: out = 16'(-1053);
			35913: out = 16'(-835);
			35914: out = 16'(257);
			35915: out = 16'(205);
			35916: out = 16'(327);
			35917: out = 16'(99);
			35918: out = 16'(275);
			35919: out = 16'(358);
			35920: out = 16'(1144);
			35921: out = 16'(334);
			35922: out = 16'(-335);
			35923: out = 16'(-711);
			35924: out = 16'(-590);
			35925: out = 16'(-216);
			35926: out = 16'(60);
			35927: out = 16'(60);
			35928: out = 16'(-192);
			35929: out = 16'(569);
			35930: out = 16'(672);
			35931: out = 16'(662);
			35932: out = 16'(316);
			35933: out = 16'(104);
			35934: out = 16'(-259);
			35935: out = 16'(690);
			35936: out = 16'(1090);
			35937: out = 16'(1008);
			35938: out = 16'(444);
			35939: out = 16'(-157);
			35940: out = 16'(-338);
			35941: out = 16'(-379);
			35942: out = 16'(-155);
			35943: out = 16'(59);
			35944: out = 16'(411);
			35945: out = 16'(525);
			35946: out = 16'(157);
			35947: out = 16'(-532);
			35948: out = 16'(-1403);
			35949: out = 16'(-1248);
			35950: out = 16'(-1181);
			35951: out = 16'(-707);
			35952: out = 16'(-1519);
			35953: out = 16'(-1426);
			35954: out = 16'(-695);
			35955: out = 16'(-35);
			35956: out = 16'(220);
			35957: out = 16'(-747);
			35958: out = 16'(-657);
			35959: out = 16'(-608);
			35960: out = 16'(234);
			35961: out = 16'(-79);
			35962: out = 16'(-239);
			35963: out = 16'(-684);
			35964: out = 16'(-229);
			35965: out = 16'(229);
			35966: out = 16'(12);
			35967: out = 16'(-312);
			35968: out = 16'(-650);
			35969: out = 16'(-1073);
			35970: out = 16'(-671);
			35971: out = 16'(325);
			35972: out = 16'(658);
			35973: out = 16'(732);
			35974: out = 16'(352);
			35975: out = 16'(95);
			35976: out = 16'(-101);
			35977: out = 16'(-87);
			35978: out = 16'(381);
			35979: out = 16'(882);
			35980: out = 16'(1117);
			35981: out = 16'(772);
			35982: out = 16'(182);
			35983: out = 16'(243);
			35984: out = 16'(-88);
			35985: out = 16'(-274);
			35986: out = 16'(71);
			35987: out = 16'(228);
			35988: out = 16'(270);
			35989: out = 16'(-64);
			35990: out = 16'(-186);
			35991: out = 16'(-142);
			35992: out = 16'(-170);
			35993: out = 16'(-156);
			35994: out = 16'(-278);
			35995: out = 16'(-307);
			35996: out = 16'(-202);
			35997: out = 16'(163);
			35998: out = 16'(6);
			35999: out = 16'(-8);
			36000: out = 16'(1425);
			36001: out = 16'(1466);
			36002: out = 16'(1413);
			36003: out = 16'(306);
			36004: out = 16'(525);
			36005: out = 16'(1032);
			36006: out = 16'(704);
			36007: out = 16'(221);
			36008: out = 16'(-445);
			36009: out = 16'(-1367);
			36010: out = 16'(-2005);
			36011: out = 16'(-2635);
			36012: out = 16'(-1096);
			36013: out = 16'(257);
			36014: out = 16'(1466);
			36015: out = 16'(824);
			36016: out = 16'(81);
			36017: out = 16'(-78);
			36018: out = 16'(-220);
			36019: out = 16'(-112);
			36020: out = 16'(107);
			36021: out = 16'(-42);
			36022: out = 16'(-411);
			36023: out = 16'(-1396);
			36024: out = 16'(-1550);
			36025: out = 16'(-1016);
			36026: out = 16'(-383);
			36027: out = 16'(171);
			36028: out = 16'(275);
			36029: out = 16'(415);
			36030: out = 16'(148);
			36031: out = 16'(-162);
			36032: out = 16'(-856);
			36033: out = 16'(-939);
			36034: out = 16'(227);
			36035: out = 16'(308);
			36036: out = 16'(322);
			36037: out = 16'(-207);
			36038: out = 16'(-184);
			36039: out = 16'(-224);
			36040: out = 16'(-49);
			36041: out = 16'(-106);
			36042: out = 16'(-9);
			36043: out = 16'(111);
			36044: out = 16'(484);
			36045: out = 16'(726);
			36046: out = 16'(1437);
			36047: out = 16'(1078);
			36048: out = 16'(-174);
			36049: out = 16'(-812);
			36050: out = 16'(-1159);
			36051: out = 16'(-660);
			36052: out = 16'(-198);
			36053: out = 16'(263);
			36054: out = 16'(-315);
			36055: out = 16'(121);
			36056: out = 16'(399);
			36057: out = 16'(1099);
			36058: out = 16'(941);
			36059: out = 16'(639);
			36060: out = 16'(345);
			36061: out = 16'(56);
			36062: out = 16'(-344);
			36063: out = 16'(75);
			36064: out = 16'(30);
			36065: out = 16'(-153);
			36066: out = 16'(-272);
			36067: out = 16'(-151);
			36068: out = 16'(236);
			36069: out = 16'(813);
			36070: out = 16'(928);
			36071: out = 16'(-229);
			36072: out = 16'(12);
			36073: out = 16'(143);
			36074: out = 16'(675);
			36075: out = 16'(161);
			36076: out = 16'(-529);
			36077: out = 16'(-1496);
			36078: out = 16'(-1396);
			36079: out = 16'(-556);
			36080: out = 16'(-505);
			36081: out = 16'(80);
			36082: out = 16'(181);
			36083: out = 16'(1083);
			36084: out = 16'(538);
			36085: out = 16'(-702);
			36086: out = 16'(-1776);
			36087: out = 16'(-1663);
			36088: out = 16'(184);
			36089: out = 16'(810);
			36090: out = 16'(1068);
			36091: out = 16'(315);
			36092: out = 16'(-230);
			36093: out = 16'(-862);
			36094: out = 16'(-1560);
			36095: out = 16'(-862);
			36096: out = 16'(387);
			36097: out = 16'(86);
			36098: out = 16'(98);
			36099: out = 16'(-358);
			36100: out = 16'(-41);
			36101: out = 16'(-53);
			36102: out = 16'(436);
			36103: out = 16'(-105);
			36104: out = 16'(144);
			36105: out = 16'(662);
			36106: out = 16'(1083);
			36107: out = 16'(751);
			36108: out = 16'(-642);
			36109: out = 16'(-1554);
			36110: out = 16'(-2020);
			36111: out = 16'(-677);
			36112: out = 16'(-404);
			36113: out = 16'(155);
			36114: out = 16'(971);
			36115: out = 16'(1449);
			36116: out = 16'(1434);
			36117: out = 16'(1293);
			36118: out = 16'(557);
			36119: out = 16'(-223);
			36120: out = 16'(-1299);
			36121: out = 16'(-1836);
			36122: out = 16'(-2071);
			36123: out = 16'(-694);
			36124: out = 16'(351);
			36125: out = 16'(1123);
			36126: out = 16'(695);
			36127: out = 16'(152);
			36128: out = 16'(-40);
			36129: out = 16'(-173);
			36130: out = 16'(-86);
			36131: out = 16'(-134);
			36132: out = 16'(-128);
			36133: out = 16'(-307);
			36134: out = 16'(-609);
			36135: out = 16'(-568);
			36136: out = 16'(-99);
			36137: out = 16'(-215);
			36138: out = 16'(412);
			36139: out = 16'(1169);
			36140: out = 16'(1760);
			36141: out = 16'(1801);
			36142: out = 16'(1475);
			36143: out = 16'(617);
			36144: out = 16'(32);
			36145: out = 16'(-204);
			36146: out = 16'(-14);
			36147: out = 16'(-78);
			36148: out = 16'(-1214);
			36149: out = 16'(-1259);
			36150: out = 16'(-1070);
			36151: out = 16'(-285);
			36152: out = 16'(265);
			36153: out = 16'(700);
			36154: out = 16'(329);
			36155: out = 16'(220);
			36156: out = 16'(274);
			36157: out = 16'(-231);
			36158: out = 16'(-296);
			36159: out = 16'(-379);
			36160: out = 16'(-188);
			36161: out = 16'(-889);
			36162: out = 16'(-2558);
			36163: out = 16'(-2637);
			36164: out = 16'(-1887);
			36165: out = 16'(711);
			36166: out = 16'(1521);
			36167: out = 16'(1885);
			36168: out = 16'(371);
			36169: out = 16'(299);
			36170: out = 16'(32);
			36171: out = 16'(-1386);
			36172: out = 16'(-1472);
			36173: out = 16'(-938);
			36174: out = 16'(62);
			36175: out = 16'(628);
			36176: out = 16'(742);
			36177: out = 16'(802);
			36178: out = 16'(904);
			36179: out = 16'(1639);
			36180: out = 16'(582);
			36181: out = 16'(232);
			36182: out = 16'(91);
			36183: out = 16'(1000);
			36184: out = 16'(1360);
			36185: out = 16'(91);
			36186: out = 16'(-337);
			36187: out = 16'(-880);
			36188: out = 16'(-220);
			36189: out = 16'(-1011);
			36190: out = 16'(-1672);
			36191: out = 16'(-1261);
			36192: out = 16'(-632);
			36193: out = 16'(308);
			36194: out = 16'(127);
			36195: out = 16'(106);
			36196: out = 16'(-306);
			36197: out = 16'(543);
			36198: out = 16'(832);
			36199: out = 16'(1161);
			36200: out = 16'(234);
			36201: out = 16'(-167);
			36202: out = 16'(161);
			36203: out = 16'(115);
			36204: out = 16'(111);
			36205: out = 16'(156);
			36206: out = 16'(-323);
			36207: out = 16'(-812);
			36208: out = 16'(-744);
			36209: out = 16'(-309);
			36210: out = 16'(393);
			36211: out = 16'(-164);
			36212: out = 16'(14);
			36213: out = 16'(142);
			36214: out = 16'(605);
			36215: out = 16'(801);
			36216: out = 16'(1114);
			36217: out = 16'(128);
			36218: out = 16'(-179);
			36219: out = 16'(281);
			36220: out = 16'(175);
			36221: out = 16'(374);
			36222: out = 16'(986);
			36223: out = 16'(1470);
			36224: out = 16'(1677);
			36225: out = 16'(157);
			36226: out = 16'(151);
			36227: out = 16'(-152);
			36228: out = 16'(-44);
			36229: out = 16'(-1582);
			36230: out = 16'(-3318);
			36231: out = 16'(-2805);
			36232: out = 16'(-1699);
			36233: out = 16'(335);
			36234: out = 16'(-123);
			36235: out = 16'(-108);
			36236: out = 16'(-292);
			36237: out = 16'(21);
			36238: out = 16'(338);
			36239: out = 16'(678);
			36240: out = 16'(982);
			36241: out = 16'(919);
			36242: out = 16'(-127);
			36243: out = 16'(-482);
			36244: out = 16'(-754);
			36245: out = 16'(-341);
			36246: out = 16'(-96);
			36247: out = 16'(146);
			36248: out = 16'(-253);
			36249: out = 16'(-316);
			36250: out = 16'(-261);
			36251: out = 16'(25);
			36252: out = 16'(387);
			36253: out = 16'(679);
			36254: out = 16'(1016);
			36255: out = 16'(956);
			36256: out = 16'(656);
			36257: out = 16'(25);
			36258: out = 16'(-726);
			36259: out = 16'(-2161);
			36260: out = 16'(-1115);
			36261: out = 16'(-90);
			36262: out = 16'(-243);
			36263: out = 16'(133);
			36264: out = 16'(277);
			36265: out = 16'(287);
			36266: out = 16'(232);
			36267: out = 16'(82);
			36268: out = 16'(-53);
			36269: out = 16'(-407);
			36270: out = 16'(-763);
			36271: out = 16'(-1813);
			36272: out = 16'(-1996);
			36273: out = 16'(-1442);
			36274: out = 16'(-647);
			36275: out = 16'(106);
			36276: out = 16'(187);
			36277: out = 16'(725);
			36278: out = 16'(885);
			36279: out = 16'(1677);
			36280: out = 16'(629);
			36281: out = 16'(-150);
			36282: out = 16'(239);
			36283: out = 16'(255);
			36284: out = 16'(363);
			36285: out = 16'(678);
			36286: out = 16'(591);
			36287: out = 16'(238);
			36288: out = 16'(-127);
			36289: out = 16'(-321);
			36290: out = 16'(-208);
			36291: out = 16'(418);
			36292: out = 16'(916);
			36293: out = 16'(1040);
			36294: out = 16'(1361);
			36295: out = 16'(1546);
			36296: out = 16'(2239);
			36297: out = 16'(982);
			36298: out = 16'(-205);
			36299: out = 16'(-1149);
			36300: out = 16'(-1377);
			36301: out = 16'(-1250);
			36302: out = 16'(-1694);
			36303: out = 16'(-1464);
			36304: out = 16'(-1088);
			36305: out = 16'(-318);
			36306: out = 16'(34);
			36307: out = 16'(140);
			36308: out = 16'(-126);
			36309: out = 16'(-447);
			36310: out = 16'(-674);
			36311: out = 16'(-1058);
			36312: out = 16'(-798);
			36313: out = 16'(353);
			36314: out = 16'(788);
			36315: out = 16'(862);
			36316: out = 16'(-1136);
			36317: out = 16'(-731);
			36318: out = 16'(-632);
			36319: out = 16'(325);
			36320: out = 16'(-897);
			36321: out = 16'(-1795);
			36322: out = 16'(-112);
			36323: out = 16'(1166);
			36324: out = 16'(2191);
			36325: out = 16'(1706);
			36326: out = 16'(291);
			36327: out = 16'(-2082);
			36328: out = 16'(-2251);
			36329: out = 16'(-1772);
			36330: out = 16'(396);
			36331: out = 16'(238);
			36332: out = 16'(475);
			36333: out = 16'(285);
			36334: out = 16'(633);
			36335: out = 16'(816);
			36336: out = 16'(1433);
			36337: out = 16'(1619);
			36338: out = 16'(1675);
			36339: out = 16'(251);
			36340: out = 16'(-227);
			36341: out = 16'(-822);
			36342: out = 16'(-80);
			36343: out = 16'(-716);
			36344: out = 16'(-1526);
			36345: out = 16'(-1946);
			36346: out = 16'(-1237);
			36347: out = 16'(426);
			36348: out = 16'(1116);
			36349: out = 16'(1229);
			36350: out = 16'(-212);
			36351: out = 16'(-46);
			36352: out = 16'(59);
			36353: out = 16'(1487);
			36354: out = 16'(920);
			36355: out = 16'(463);
			36356: out = 16'(-1066);
			36357: out = 16'(-738);
			36358: out = 16'(-217);
			36359: out = 16'(207);
			36360: out = 16'(16);
			36361: out = 16'(-286);
			36362: out = 16'(4);
			36363: out = 16'(237);
			36364: out = 16'(186);
			36365: out = 16'(1150);
			36366: out = 16'(1159);
			36367: out = 16'(588);
			36368: out = 16'(-879);
			36369: out = 16'(-1946);
			36370: out = 16'(-2434);
			36371: out = 16'(-1483);
			36372: out = 16'(-204);
			36373: out = 16'(896);
			36374: out = 16'(1160);
			36375: out = 16'(896);
			36376: out = 16'(244);
			36377: out = 16'(40);
			36378: out = 16'(143);
			36379: out = 16'(-159);
			36380: out = 16'(-188);
			36381: out = 16'(-352);
			36382: out = 16'(-590);
			36383: out = 16'(-763);
			36384: out = 16'(-628);
			36385: out = 16'(-1049);
			36386: out = 16'(-885);
			36387: out = 16'(-220);
			36388: out = 16'(-452);
			36389: out = 16'(-893);
			36390: out = 16'(-1873);
			36391: out = 16'(-1458);
			36392: out = 16'(-640);
			36393: out = 16'(195);
			36394: out = 16'(1276);
			36395: out = 16'(1811);
			36396: out = 16'(564);
			36397: out = 16'(-280);
			36398: out = 16'(-1052);
			36399: out = 16'(-209);
			36400: out = 16'(387);
			36401: out = 16'(1192);
			36402: out = 16'(403);
			36403: out = 16'(144);
			36404: out = 16'(231);
			36405: out = 16'(263);
			36406: out = 16'(261);
			36407: out = 16'(-165);
			36408: out = 16'(210);
			36409: out = 16'(377);
			36410: out = 16'(1153);
			36411: out = 16'(75);
			36412: out = 16'(-885);
			36413: out = 16'(-1910);
			36414: out = 16'(-969);
			36415: out = 16'(389);
			36416: out = 16'(-142);
			36417: out = 16'(114);
			36418: out = 16'(215);
			36419: out = 16'(288);
			36420: out = 16'(581);
			36421: out = 16'(1115);
			36422: out = 16'(1083);
			36423: out = 16'(734);
			36424: out = 16'(-194);
			36425: out = 16'(-470);
			36426: out = 16'(-698);
			36427: out = 16'(-203);
			36428: out = 16'(-545);
			36429: out = 16'(-767);
			36430: out = 16'(-1521);
			36431: out = 16'(-838);
			36432: out = 16'(35);
			36433: out = 16'(549);
			36434: out = 16'(1000);
			36435: out = 16'(1010);
			36436: out = 16'(832);
			36437: out = 16'(280);
			36438: out = 16'(-144);
			36439: out = 16'(-1248);
			36440: out = 16'(-1542);
			36441: out = 16'(-1466);
			36442: out = 16'(114);
			36443: out = 16'(1062);
			36444: out = 16'(1438);
			36445: out = 16'(1002);
			36446: out = 16'(441);
			36447: out = 16'(-198);
			36448: out = 16'(-298);
			36449: out = 16'(-81);
			36450: out = 16'(1023);
			36451: out = 16'(822);
			36452: out = 16'(510);
			36453: out = 16'(-984);
			36454: out = 16'(-791);
			36455: out = 16'(-190);
			36456: out = 16'(204);
			36457: out = 16'(83);
			36458: out = 16'(-278);
			36459: out = 16'(-1582);
			36460: out = 16'(-1762);
			36461: out = 16'(-947);
			36462: out = 16'(164);
			36463: out = 16'(1055);
			36464: out = 16'(1438);
			36465: out = 16'(517);
			36466: out = 16'(-612);
			36467: out = 16'(-1322);
			36468: out = 16'(-1356);
			36469: out = 16'(-729);
			36470: out = 16'(30);
			36471: out = 16'(611);
			36472: out = 16'(673);
			36473: out = 16'(402);
			36474: out = 16'(-330);
			36475: out = 16'(-1003);
			36476: out = 16'(-261);
			36477: out = 16'(284);
			36478: out = 16'(748);
			36479: out = 16'(441);
			36480: out = 16'(-156);
			36481: out = 16'(-1006);
			36482: out = 16'(-1051);
			36483: out = 16'(-863);
			36484: out = 16'(-603);
			36485: out = 16'(62);
			36486: out = 16'(503);
			36487: out = 16'(777);
			36488: out = 16'(531);
			36489: out = 16'(167);
			36490: out = 16'(-533);
			36491: out = 16'(-161);
			36492: out = 16'(479);
			36493: out = 16'(1017);
			36494: out = 16'(896);
			36495: out = 16'(245);
			36496: out = 16'(288);
			36497: out = 16'(51);
			36498: out = 16'(-225);
			36499: out = 16'(-99);
			36500: out = 16'(-98);
			36501: out = 16'(-59);
			36502: out = 16'(58);
			36503: out = 16'(369);
			36504: out = 16'(590);
			36505: out = 16'(1206);
			36506: out = 16'(1243);
			36507: out = 16'(336);
			36508: out = 16'(-759);
			36509: out = 16'(-1547);
			36510: out = 16'(-1180);
			36511: out = 16'(-609);
			36512: out = 16'(-25);
			36513: out = 16'(1247);
			36514: out = 16'(1303);
			36515: out = 16'(1062);
			36516: out = 16'(-957);
			36517: out = 16'(-1181);
			36518: out = 16'(219);
			36519: out = 16'(1505);
			36520: out = 16'(1904);
			36521: out = 16'(172);
			36522: out = 16'(-509);
			36523: out = 16'(-1305);
			36524: out = 16'(-1036);
			36525: out = 16'(-965);
			36526: out = 16'(-524);
			36527: out = 16'(-328);
			36528: out = 16'(-14);
			36529: out = 16'(192);
			36530: out = 16'(-213);
			36531: out = 16'(-150);
			36532: out = 16'(-74);
			36533: out = 16'(1757);
			36534: out = 16'(1793);
			36535: out = 16'(492);
			36536: out = 16'(-228);
			36537: out = 16'(-889);
			36538: out = 16'(-577);
			36539: out = 16'(-1070);
			36540: out = 16'(-855);
			36541: out = 16'(98);
			36542: out = 16'(686);
			36543: out = 16'(1042);
			36544: out = 16'(211);
			36545: out = 16'(276);
			36546: out = 16'(-62);
			36547: out = 16'(-74);
			36548: out = 16'(-1482);
			36549: out = 16'(-3001);
			36550: out = 16'(-2930);
			36551: out = 16'(-1905);
			36552: out = 16'(54);
			36553: out = 16'(200);
			36554: out = 16'(578);
			36555: out = 16'(774);
			36556: out = 16'(252);
			36557: out = 16'(-109);
			36558: out = 16'(-140);
			36559: out = 16'(392);
			36560: out = 16'(944);
			36561: out = 16'(1450);
			36562: out = 16'(908);
			36563: out = 16'(155);
			36564: out = 16'(300);
			36565: out = 16'(-279);
			36566: out = 16'(-667);
			36567: out = 16'(-644);
			36568: out = 16'(-430);
			36569: out = 16'(4);
			36570: out = 16'(-192);
			36571: out = 16'(247);
			36572: out = 16'(690);
			36573: out = 16'(1846);
			36574: out = 16'(1996);
			36575: out = 16'(1359);
			36576: out = 16'(297);
			36577: out = 16'(-559);
			36578: out = 16'(-667);
			36579: out = 16'(-317);
			36580: out = 16'(229);
			36581: out = 16'(134);
			36582: out = 16'(295);
			36583: out = 16'(94);
			36584: out = 16'(-162);
			36585: out = 16'(-746);
			36586: out = 16'(-1129);
			36587: out = 16'(-429);
			36588: out = 16'(-347);
			36589: out = 16'(-764);
			36590: out = 16'(-267);
			36591: out = 16'(-221);
			36592: out = 16'(271);
			36593: out = 16'(-1122);
			36594: out = 16'(-1333);
			36595: out = 16'(-652);
			36596: out = 16'(35);
			36597: out = 16'(348);
			36598: out = 16'(382);
			36599: out = 16'(-30);
			36600: out = 16'(-124);
			36601: out = 16'(-246);
			36602: out = 16'(1092);
			36603: out = 16'(2192);
			36604: out = 16'(1574);
			36605: out = 16'(486);
			36606: out = 16'(-865);
			36607: out = 16'(-2581);
			36608: out = 16'(-2269);
			36609: out = 16'(-435);
			36610: out = 16'(888);
			36611: out = 16'(1341);
			36612: out = 16'(8);
			36613: out = 16'(-283);
			36614: out = 16'(-704);
			36615: out = 16'(38);
			36616: out = 16'(-50);
			36617: out = 16'(312);
			36618: out = 16'(32);
			36619: out = 16'(568);
			36620: out = 16'(557);
			36621: out = 16'(333);
			36622: out = 16'(-667);
			36623: out = 16'(-1618);
			36624: out = 16'(-1859);
			36625: out = 16'(-1907);
			36626: out = 16'(-1830);
			36627: out = 16'(-469);
			36628: out = 16'(70);
			36629: out = 16'(298);
			36630: out = 16'(-43);
			36631: out = 16'(115);
			36632: out = 16'(788);
			36633: out = 16'(1097);
			36634: out = 16'(705);
			36635: out = 16'(-1356);
			36636: out = 16'(-1958);
			36637: out = 16'(-1979);
			36638: out = 16'(721);
			36639: out = 16'(1011);
			36640: out = 16'(1206);
			36641: out = 16'(311);
			36642: out = 16'(504);
			36643: out = 16'(863);
			36644: out = 16'(2278);
			36645: out = 16'(2505);
			36646: out = 16'(1983);
			36647: out = 16'(506);
			36648: out = 16'(-791);
			36649: out = 16'(-1431);
			36650: out = 16'(-1733);
			36651: out = 16'(-904);
			36652: out = 16'(574);
			36653: out = 16'(1698);
			36654: out = 16'(1933);
			36655: out = 16'(711);
			36656: out = 16'(-125);
			36657: out = 16'(-816);
			36658: out = 16'(-720);
			36659: out = 16'(-344);
			36660: out = 16'(175);
			36661: out = 16'(-117);
			36662: out = 16'(-215);
			36663: out = 16'(-288);
			36664: out = 16'(-991);
			36665: out = 16'(-974);
			36666: out = 16'(-647);
			36667: out = 16'(-307);
			36668: out = 16'(-213);
			36669: out = 16'(0);
			36670: out = 16'(-826);
			36671: out = 16'(-837);
			36672: out = 16'(-320);
			36673: out = 16'(1538);
			36674: out = 16'(2470);
			36675: out = 16'(1143);
			36676: out = 16'(-460);
			36677: out = 16'(-2149);
			36678: out = 16'(-224);
			36679: out = 16'(-279);
			36680: out = 16'(37);
			36681: out = 16'(-283);
			36682: out = 16'(794);
			36683: out = 16'(2213);
			36684: out = 16'(681);
			36685: out = 16'(-452);
			36686: out = 16'(-2094);
			36687: out = 16'(-428);
			36688: out = 16'(221);
			36689: out = 16'(-151);
			36690: out = 16'(-183);
			36691: out = 16'(-129);
			36692: out = 16'(704);
			36693: out = 16'(245);
			36694: out = 16'(-278);
			36695: out = 16'(-544);
			36696: out = 16'(-936);
			36697: out = 16'(-1068);
			36698: out = 16'(-1935);
			36699: out = 16'(-1098);
			36700: out = 16'(85);
			36701: out = 16'(346);
			36702: out = 16'(-297);
			36703: out = 16'(-2026);
			36704: out = 16'(-1103);
			36705: out = 16'(-581);
			36706: out = 16'(559);
			36707: out = 16'(77);
			36708: out = 16'(-80);
			36709: out = 16'(-1011);
			36710: out = 16'(-105);
			36711: out = 16'(445);
			36712: out = 16'(853);
			36713: out = 16'(561);
			36714: out = 16'(516);
			36715: out = 16'(1036);
			36716: out = 16'(1718);
			36717: out = 16'(2186);
			36718: out = 16'(1614);
			36719: out = 16'(880);
			36720: out = 16'(79);
			36721: out = 16'(-581);
			36722: out = 16'(-260);
			36723: out = 16'(716);
			36724: out = 16'(692);
			36725: out = 16'(137);
			36726: out = 16'(-1565);
			36727: out = 16'(-1801);
			36728: out = 16'(-1586);
			36729: out = 16'(389);
			36730: out = 16'(290);
			36731: out = 16'(233);
			36732: out = 16'(-1018);
			36733: out = 16'(-770);
			36734: out = 16'(-546);
			36735: out = 16'(-149);
			36736: out = 16'(-341);
			36737: out = 16'(-574);
			36738: out = 16'(-926);
			36739: out = 16'(-675);
			36740: out = 16'(-33);
			36741: out = 16'(299);
			36742: out = 16'(354);
			36743: out = 16'(-46);
			36744: out = 16'(-3);
			36745: out = 16'(-250);
			36746: out = 16'(-493);
			36747: out = 16'(-286);
			36748: out = 16'(-32);
			36749: out = 16'(-176);
			36750: out = 16'(36);
			36751: out = 16'(199);
			36752: out = 16'(2191);
			36753: out = 16'(2056);
			36754: out = 16'(1697);
			36755: out = 16'(-719);
			36756: out = 16'(-922);
			36757: out = 16'(-535);
			36758: out = 16'(1127);
			36759: out = 16'(1280);
			36760: out = 16'(647);
			36761: out = 16'(-599);
			36762: out = 16'(-992);
			36763: out = 16'(-146);
			36764: out = 16'(131);
			36765: out = 16'(192);
			36766: out = 16'(-603);
			36767: out = 16'(-1375);
			36768: out = 16'(-1833);
			36769: out = 16'(-565);
			36770: out = 16'(-306);
			36771: out = 16'(81);
			36772: out = 16'(-169);
			36773: out = 16'(65);
			36774: out = 16'(272);
			36775: out = 16'(-77);
			36776: out = 16'(-4);
			36777: out = 16'(318);
			36778: out = 16'(340);
			36779: out = 16'(491);
			36780: out = 16'(777);
			36781: out = 16'(445);
			36782: out = 16'(432);
			36783: out = 16'(706);
			36784: out = 16'(732);
			36785: out = 16'(546);
			36786: out = 16'(-47);
			36787: out = 16'(-193);
			36788: out = 16'(-406);
			36789: out = 16'(-2306);
			36790: out = 16'(-1936);
			36791: out = 16'(-1127);
			36792: out = 16'(1833);
			36793: out = 16'(2169);
			36794: out = 16'(1720);
			36795: out = 16'(-178);
			36796: out = 16'(-487);
			36797: out = 16'(257);
			36798: out = 16'(1099);
			36799: out = 16'(1225);
			36800: out = 16'(171);
			36801: out = 16'(-31);
			36802: out = 16'(-366);
			36803: out = 16'(-237);
			36804: out = 16'(16);
			36805: out = 16'(408);
			36806: out = 16'(973);
			36807: out = 16'(377);
			36808: out = 16'(-548);
			36809: out = 16'(-1011);
			36810: out = 16'(-1059);
			36811: out = 16'(-571);
			36812: out = 16'(-811);
			36813: out = 16'(-381);
			36814: out = 16'(-107);
			36815: out = 16'(1105);
			36816: out = 16'(1457);
			36817: out = 16'(1355);
			36818: out = 16'(577);
			36819: out = 16'(-12);
			36820: out = 16'(-175);
			36821: out = 16'(-247);
			36822: out = 16'(-125);
			36823: out = 16'(49);
			36824: out = 16'(-136);
			36825: out = 16'(-398);
			36826: out = 16'(-128);
			36827: out = 16'(-323);
			36828: out = 16'(-331);
			36829: out = 16'(-1552);
			36830: out = 16'(-935);
			36831: out = 16'(-102);
			36832: out = 16'(-108);
			36833: out = 16'(-481);
			36834: out = 16'(-1134);
			36835: out = 16'(-2100);
			36836: out = 16'(-2194);
			36837: out = 16'(-1370);
			36838: out = 16'(54);
			36839: out = 16'(1091);
			36840: out = 16'(1039);
			36841: out = 16'(740);
			36842: out = 16'(-101);
			36843: out = 16'(-392);
			36844: out = 16'(-1408);
			36845: out = 16'(-1817);
			36846: out = 16'(-1498);
			36847: out = 16'(-580);
			36848: out = 16'(538);
			36849: out = 16'(1025);
			36850: out = 16'(1554);
			36851: out = 16'(1855);
			36852: out = 16'(680);
			36853: out = 16'(216);
			36854: out = 16'(280);
			36855: out = 16'(-58);
			36856: out = 16'(-57);
			36857: out = 16'(-251);
			36858: out = 16'(131);
			36859: out = 16'(26);
			36860: out = 16'(-560);
			36861: out = 16'(-1147);
			36862: out = 16'(-1299);
			36863: out = 16'(-74);
			36864: out = 16'(183);
			36865: out = 16'(353);
			36866: out = 16'(-513);
			36867: out = 16'(-320);
			36868: out = 16'(33);
			36869: out = 16'(-164);
			36870: out = 16'(-113);
			36871: out = 16'(-129);
			36872: out = 16'(936);
			36873: out = 16'(973);
			36874: out = 16'(294);
			36875: out = 16'(87);
			36876: out = 16'(31);
			36877: out = 16'(827);
			36878: out = 16'(150);
			36879: out = 16'(-76);
			36880: out = 16'(-108);
			36881: out = 16'(177);
			36882: out = 16'(263);
			36883: out = 16'(-12);
			36884: out = 16'(-554);
			36885: out = 16'(-1138);
			36886: out = 16'(-1399);
			36887: out = 16'(-977);
			36888: out = 16'(60);
			36889: out = 16'(139);
			36890: out = 16'(1043);
			36891: out = 16'(1849);
			36892: out = 16'(1964);
			36893: out = 16'(1224);
			36894: out = 16'(-155);
			36895: out = 16'(-1068);
			36896: out = 16'(-1458);
			36897: out = 16'(-554);
			36898: out = 16'(-694);
			36899: out = 16'(-538);
			36900: out = 16'(-677);
			36901: out = 16'(-88);
			36902: out = 16'(102);
			36903: out = 16'(-1286);
			36904: out = 16'(-1856);
			36905: out = 16'(-2183);
			36906: out = 16'(20);
			36907: out = 16'(608);
			36908: out = 16'(882);
			36909: out = 16'(81);
			36910: out = 16'(-89);
			36911: out = 16'(-67);
			36912: out = 16'(609);
			36913: out = 16'(1024);
			36914: out = 16'(1605);
			36915: out = 16'(1247);
			36916: out = 16'(1119);
			36917: out = 16'(617);
			36918: out = 16'(1491);
			36919: out = 16'(1558);
			36920: out = 16'(370);
			36921: out = 16'(-1240);
			36922: out = 16'(-2355);
			36923: out = 16'(-302);
			36924: out = 16'(790);
			36925: out = 16'(1907);
			36926: out = 16'(1140);
			36927: out = 16'(734);
			36928: out = 16'(43);
			36929: out = 16'(-491);
			36930: out = 16'(-603);
			36931: out = 16'(-60);
			36932: out = 16'(633);
			36933: out = 16'(1006);
			36934: out = 16'(89);
			36935: out = 16'(597);
			36936: out = 16'(433);
			36937: out = 16'(235);
			36938: out = 16'(-930);
			36939: out = 16'(-1519);
			36940: out = 16'(-359);
			36941: out = 16'(-80);
			36942: out = 16'(69);
			36943: out = 16'(-969);
			36944: out = 16'(-1150);
			36945: out = 16'(-1029);
			36946: out = 16'(-1122);
			36947: out = 16'(-738);
			36948: out = 16'(-145);
			36949: out = 16'(805);
			36950: out = 16'(1095);
			36951: out = 16'(624);
			36952: out = 16'(506);
			36953: out = 16'(108);
			36954: out = 16'(-30);
			36955: out = 16'(-500);
			36956: out = 16'(-572);
			36957: out = 16'(-291);
			36958: out = 16'(297);
			36959: out = 16'(709);
			36960: out = 16'(312);
			36961: out = 16'(241);
			36962: out = 16'(138);
			36963: out = 16'(143);
			36964: out = 16'(204);
			36965: out = 16'(265);
			36966: out = 16'(-119);
			36967: out = 16'(-559);
			36968: out = 16'(-1114);
			36969: out = 16'(-787);
			36970: out = 16'(-416);
			36971: out = 16'(180);
			36972: out = 16'(204);
			36973: out = 16'(-30);
			36974: out = 16'(-1056);
			36975: out = 16'(-824);
			36976: out = 16'(-372);
			36977: out = 16'(1024);
			36978: out = 16'(1121);
			36979: out = 16'(982);
			36980: out = 16'(0);
			36981: out = 16'(-168);
			36982: out = 16'(-268);
			36983: out = 16'(-222);
			36984: out = 16'(-397);
			36985: out = 16'(-646);
			36986: out = 16'(-680);
			36987: out = 16'(-329);
			36988: out = 16'(342);
			36989: out = 16'(863);
			36990: out = 16'(990);
			36991: out = 16'(237);
			36992: out = 16'(239);
			36993: out = 16'(89);
			36994: out = 16'(158);
			36995: out = 16'(173);
			36996: out = 16'(244);
			36997: out = 16'(-285);
			36998: out = 16'(-92);
			36999: out = 16'(215);
			37000: out = 16'(1225);
			37001: out = 16'(1414);
			37002: out = 16'(1283);
			37003: out = 16'(439);
			37004: out = 16'(-79);
			37005: out = 16'(-348);
			37006: out = 16'(-384);
			37007: out = 16'(-344);
			37008: out = 16'(-371);
			37009: out = 16'(-347);
			37010: out = 16'(-322);
			37011: out = 16'(-174);
			37012: out = 16'(-224);
			37013: out = 16'(-246);
			37014: out = 16'(-718);
			37015: out = 16'(-918);
			37016: out = 16'(-1110);
			37017: out = 16'(96);
			37018: out = 16'(-248);
			37019: out = 16'(-689);
			37020: out = 16'(-715);
			37021: out = 16'(-292);
			37022: out = 16'(341);
			37023: out = 16'(1214);
			37024: out = 16'(1017);
			37025: out = 16'(-261);
			37026: out = 16'(-121);
			37027: out = 16'(107);
			37028: out = 16'(1503);
			37029: out = 16'(567);
			37030: out = 16'(108);
			37031: out = 16'(-230);
			37032: out = 16'(255);
			37033: out = 16'(591);
			37034: out = 16'(83);
			37035: out = 16'(-60);
			37036: out = 16'(-197);
			37037: out = 16'(523);
			37038: out = 16'(413);
			37039: out = 16'(127);
			37040: out = 16'(102);
			37041: out = 16'(-113);
			37042: out = 16'(-388);
			37043: out = 16'(-345);
			37044: out = 16'(-381);
			37045: out = 16'(-314);
			37046: out = 16'(-675);
			37047: out = 16'(-580);
			37048: out = 16'(62);
			37049: out = 16'(429);
			37050: out = 16'(498);
			37051: out = 16'(-312);
			37052: out = 16'(-755);
			37053: out = 16'(-1152);
			37054: out = 16'(83);
			37055: out = 16'(-282);
			37056: out = 16'(-745);
			37057: out = 16'(-724);
			37058: out = 16'(-479);
			37059: out = 16'(-68);
			37060: out = 16'(65);
			37061: out = 16'(222);
			37062: out = 16'(250);
			37063: out = 16'(558);
			37064: out = 16'(647);
			37065: out = 16'(619);
			37066: out = 16'(321);
			37067: out = 16'(-182);
			37068: out = 16'(-1115);
			37069: out = 16'(-935);
			37070: out = 16'(-534);
			37071: out = 16'(-250);
			37072: out = 16'(485);
			37073: out = 16'(1102);
			37074: out = 16'(1010);
			37075: out = 16'(533);
			37076: out = 16'(-328);
			37077: out = 16'(160);
			37078: out = 16'(-172);
			37079: out = 16'(-276);
			37080: out = 16'(-1083);
			37081: out = 16'(-795);
			37082: out = 16'(126);
			37083: out = 16'(510);
			37084: out = 16'(499);
			37085: out = 16'(138);
			37086: out = 16'(-714);
			37087: out = 16'(-1027);
			37088: out = 16'(99);
			37089: out = 16'(403);
			37090: out = 16'(618);
			37091: out = 16'(134);
			37092: out = 16'(83);
			37093: out = 16'(98);
			37094: out = 16'(62);
			37095: out = 16'(169);
			37096: out = 16'(211);
			37097: out = 16'(1192);
			37098: out = 16'(1092);
			37099: out = 16'(521);
			37100: out = 16'(184);
			37101: out = 16'(-193);
			37102: out = 16'(-835);
			37103: out = 16'(-157);
			37104: out = 16'(-21);
			37105: out = 16'(142);
			37106: out = 16'(-1221);
			37107: out = 16'(-1954);
			37108: out = 16'(-1559);
			37109: out = 16'(-182);
			37110: out = 16'(1199);
			37111: out = 16'(1509);
			37112: out = 16'(1064);
			37113: out = 16'(-102);
			37114: out = 16'(-779);
			37115: out = 16'(-1393);
			37116: out = 16'(-1381);
			37117: out = 16'(-638);
			37118: out = 16'(122);
			37119: out = 16'(572);
			37120: out = 16'(314);
			37121: out = 16'(-70);
			37122: out = 16'(-246);
			37123: out = 16'(-79);
			37124: out = 16'(121);
			37125: out = 16'(-360);
			37126: out = 16'(7);
			37127: out = 16'(57);
			37128: out = 16'(194);
			37129: out = 16'(-548);
			37130: out = 16'(-1013);
			37131: out = 16'(-426);
			37132: out = 16'(593);
			37133: out = 16'(1749);
			37134: out = 16'(1017);
			37135: out = 16'(645);
			37136: out = 16'(-15);
			37137: out = 16'(209);
			37138: out = 16'(105);
			37139: out = 16'(87);
			37140: out = 16'(-525);
			37141: out = 16'(-608);
			37142: out = 16'(115);
			37143: out = 16'(4);
			37144: out = 16'(96);
			37145: out = 16'(-284);
			37146: out = 16'(468);
			37147: out = 16'(848);
			37148: out = 16'(131);
			37149: out = 16'(-365);
			37150: out = 16'(-662);
			37151: out = 16'(331);
			37152: out = 16'(867);
			37153: out = 16'(1180);
			37154: out = 16'(1266);
			37155: out = 16'(756);
			37156: out = 16'(97);
			37157: out = 16'(-655);
			37158: out = 16'(-409);
			37159: out = 16'(835);
			37160: out = 16'(1279);
			37161: out = 16'(1241);
			37162: out = 16'(-2);
			37163: out = 16'(-21);
			37164: out = 16'(-200);
			37165: out = 16'(-877);
			37166: out = 16'(-450);
			37167: out = 16'(-8);
			37168: out = 16'(419);
			37169: out = 16'(21);
			37170: out = 16'(-542);
			37171: out = 16'(-1855);
			37172: out = 16'(-1415);
			37173: out = 16'(-113);
			37174: out = 16'(0);
			37175: out = 16'(141);
			37176: out = 16'(1);
			37177: out = 16'(-830);
			37178: out = 16'(-1025);
			37179: out = 16'(-312);
			37180: out = 16'(220);
			37181: out = 16'(406);
			37182: out = 16'(-724);
			37183: out = 16'(-1128);
			37184: out = 16'(-1423);
			37185: out = 16'(61);
			37186: out = 16'(69);
			37187: out = 16'(108);
			37188: out = 16'(-175);
			37189: out = 16'(-32);
			37190: out = 16'(76);
			37191: out = 16'(-231);
			37192: out = 16'(-310);
			37193: out = 16'(-263);
			37194: out = 16'(-317);
			37195: out = 16'(-118);
			37196: out = 16'(226);
			37197: out = 16'(469);
			37198: out = 16'(320);
			37199: out = 16'(-1149);
			37200: out = 16'(-322);
			37201: out = 16'(366);
			37202: out = 16'(1609);
			37203: out = 16'(873);
			37204: out = 16'(-177);
			37205: out = 16'(-2040);
			37206: out = 16'(-2407);
			37207: out = 16'(-2074);
			37208: out = 16'(-125);
			37209: out = 16'(546);
			37210: out = 16'(608);
			37211: out = 16'(289);
			37212: out = 16'(258);
			37213: out = 16'(670);
			37214: out = 16'(91);
			37215: out = 16'(-540);
			37216: out = 16'(-1867);
			37217: out = 16'(-1539);
			37218: out = 16'(-1083);
			37219: out = 16'(213);
			37220: out = 16'(266);
			37221: out = 16'(428);
			37222: out = 16'(593);
			37223: out = 16'(1058);
			37224: out = 16'(1292);
			37225: out = 16'(304);
			37226: out = 16'(-66);
			37227: out = 16'(-206);
			37228: out = 16'(445);
			37229: out = 16'(679);
			37230: out = 16'(537);
			37231: out = 16'(918);
			37232: out = 16'(873);
			37233: out = 16'(972);
			37234: out = 16'(37);
			37235: out = 16'(56);
			37236: out = 16'(1200);
			37237: out = 16'(1473);
			37238: out = 16'(1110);
			37239: out = 16'(-1061);
			37240: out = 16'(-1642);
			37241: out = 16'(-1888);
			37242: out = 16'(-833);
			37243: out = 16'(-276);
			37244: out = 16'(254);
			37245: out = 16'(146);
			37246: out = 16'(70);
			37247: out = 16'(-239);
			37248: out = 16'(-571);
			37249: out = 16'(-633);
			37250: out = 16'(-218);
			37251: out = 16'(-231);
			37252: out = 16'(-128);
			37253: out = 16'(-324);
			37254: out = 16'(0);
			37255: out = 16'(49);
			37256: out = 16'(-152);
			37257: out = 16'(-219);
			37258: out = 16'(-84);
			37259: out = 16'(136);
			37260: out = 16'(432);
			37261: out = 16'(500);
			37262: out = 16'(181);
			37263: out = 16'(-465);
			37264: out = 16'(-1169);
			37265: out = 16'(-1075);
			37266: out = 16'(-706);
			37267: out = 16'(256);
			37268: out = 16'(387);
			37269: out = 16'(817);
			37270: out = 16'(839);
			37271: out = 16'(1258);
			37272: out = 16'(1078);
			37273: out = 16'(987);
			37274: out = 16'(-220);
			37275: out = 16'(-824);
			37276: out = 16'(-792);
			37277: out = 16'(176);
			37278: out = 16'(918);
			37279: out = 16'(148);
			37280: out = 16'(-249);
			37281: out = 16'(-879);
			37282: out = 16'(-1028);
			37283: out = 16'(-1177);
			37284: out = 16'(-1038);
			37285: out = 16'(-347);
			37286: out = 16'(-112);
			37287: out = 16'(-186);
			37288: out = 16'(-816);
			37289: out = 16'(-937);
			37290: out = 16'(-145);
			37291: out = 16'(-234);
			37292: out = 16'(102);
			37293: out = 16'(523);
			37294: out = 16'(1108);
			37295: out = 16'(1111);
			37296: out = 16'(-95);
			37297: out = 16'(-448);
			37298: out = 16'(-654);
			37299: out = 16'(76);
			37300: out = 16'(-20);
			37301: out = 16'(-180);
			37302: out = 16'(-599);
			37303: out = 16'(-662);
			37304: out = 16'(-629);
			37305: out = 16'(-14);
			37306: out = 16'(103);
			37307: out = 16'(-143);
			37308: out = 16'(87);
			37309: out = 16'(111);
			37310: out = 16'(-162);
			37311: out = 16'(588);
			37312: out = 16'(1155);
			37313: out = 16'(1616);
			37314: out = 16'(1030);
			37315: out = 16'(309);
			37316: out = 16'(-212);
			37317: out = 16'(-415);
			37318: out = 16'(-234);
			37319: out = 16'(71);
			37320: out = 16'(87);
			37321: out = 16'(-333);
			37322: out = 16'(-153);
			37323: out = 16'(-851);
			37324: out = 16'(-1470);
			37325: out = 16'(-2215);
			37326: out = 16'(-1695);
			37327: out = 16'(-164);
			37328: out = 16'(158);
			37329: out = 16'(80);
			37330: out = 16'(-1020);
			37331: out = 16'(-734);
			37332: out = 16'(-385);
			37333: out = 16'(276);
			37334: out = 16'(560);
			37335: out = 16'(703);
			37336: out = 16'(1069);
			37337: out = 16'(409);
			37338: out = 16'(-320);
			37339: out = 16'(-597);
			37340: out = 16'(9);
			37341: out = 16'(1109);
			37342: out = 16'(25);
			37343: out = 16'(-393);
			37344: out = 16'(-1089);
			37345: out = 16'(-292);
			37346: out = 16'(127);
			37347: out = 16'(667);
			37348: out = 16'(384);
			37349: out = 16'(236);
			37350: out = 16'(154);
			37351: out = 16'(107);
			37352: out = 16'(273);
			37353: out = 16'(953);
			37354: out = 16'(793);
			37355: out = 16'(451);
			37356: out = 16'(-138);
			37357: out = 16'(-497);
			37358: out = 16'(-638);
			37359: out = 16'(-685);
			37360: out = 16'(-449);
			37361: out = 16'(-232);
			37362: out = 16'(213);
			37363: out = 16'(144);
			37364: out = 16'(-135);
			37365: out = 16'(-1318);
			37366: out = 16'(-2016);
			37367: out = 16'(-2144);
			37368: out = 16'(-1200);
			37369: out = 16'(42);
			37370: out = 16'(1307);
			37371: out = 16'(1733);
			37372: out = 16'(1513);
			37373: out = 16'(361);
			37374: out = 16'(-629);
			37375: out = 16'(-1365);
			37376: out = 16'(217);
			37377: out = 16'(439);
			37378: out = 16'(718);
			37379: out = 16'(-476);
			37380: out = 16'(-133);
			37381: out = 16'(718);
			37382: out = 16'(969);
			37383: out = 16'(672);
			37384: out = 16'(-261);
			37385: out = 16'(-784);
			37386: out = 16'(-788);
			37387: out = 16'(332);
			37388: out = 16'(680);
			37389: out = 16'(999);
			37390: out = 16'(192);
			37391: out = 16'(319);
			37392: out = 16'(158);
			37393: out = 16'(232);
			37394: out = 16'(-148);
			37395: out = 16'(-182);
			37396: out = 16'(-257);
			37397: out = 16'(371);
			37398: out = 16'(965);
			37399: out = 16'(1294);
			37400: out = 16'(742);
			37401: out = 16'(-359);
			37402: out = 16'(-1473);
			37403: out = 16'(-1809);
			37404: out = 16'(-965);
			37405: out = 16'(-337);
			37406: out = 16'(292);
			37407: out = 16'(-251);
			37408: out = 16'(410);
			37409: out = 16'(653);
			37410: out = 16'(1010);
			37411: out = 16'(355);
			37412: out = 16'(-235);
			37413: out = 16'(-211);
			37414: out = 16'(-451);
			37415: out = 16'(-654);
			37416: out = 16'(29);
			37417: out = 16'(8);
			37418: out = 16'(-311);
			37419: out = 16'(-815);
			37420: out = 16'(-1096);
			37421: out = 16'(-940);
			37422: out = 16'(-776);
			37423: out = 16'(-358);
			37424: out = 16'(-140);
			37425: out = 16'(480);
			37426: out = 16'(570);
			37427: out = 16'(-52);
			37428: out = 16'(45);
			37429: out = 16'(262);
			37430: out = 16'(74);
			37431: out = 16'(669);
			37432: out = 16'(933);
			37433: out = 16'(451);
			37434: out = 16'(-459);
			37435: out = 16'(-1491);
			37436: out = 16'(-1752);
			37437: out = 16'(-1398);
			37438: out = 16'(-469);
			37439: out = 16'(-164);
			37440: out = 16'(-9);
			37441: out = 16'(-1);
			37442: out = 16'(-908);
			37443: out = 16'(-1324);
			37444: out = 16'(-894);
			37445: out = 16'(-151);
			37446: out = 16'(534);
			37447: out = 16'(338);
			37448: out = 16'(226);
			37449: out = 16'(27);
			37450: out = 16'(1069);
			37451: out = 16'(931);
			37452: out = 16'(653);
			37453: out = 16'(48);
			37454: out = 16'(153);
			37455: out = 16'(795);
			37456: out = 16'(-29);
			37457: out = 16'(95);
			37458: out = 16'(236);
			37459: out = 16'(1411);
			37460: out = 16'(1389);
			37461: out = 16'(247);
			37462: out = 16'(-571);
			37463: out = 16'(-1170);
			37464: out = 16'(-1413);
			37465: out = 16'(-553);
			37466: out = 16'(481);
			37467: out = 16'(1219);
			37468: out = 16'(1570);
			37469: out = 16'(1536);
			37470: out = 16'(-85);
			37471: out = 16'(-236);
			37472: out = 16'(-136);
			37473: out = 16'(1139);
			37474: out = 16'(523);
			37475: out = 16'(-1258);
			37476: out = 16'(-1617);
			37477: out = 16'(-1838);
			37478: out = 16'(-1344);
			37479: out = 16'(-633);
			37480: out = 16'(-12);
			37481: out = 16'(-151);
			37482: out = 16'(175);
			37483: out = 16'(126);
			37484: out = 16'(-180);
			37485: out = 16'(86);
			37486: out = 16'(329);
			37487: out = 16'(229);
			37488: out = 16'(-342);
			37489: out = 16'(-1041);
			37490: out = 16'(-239);
			37491: out = 16'(-133);
			37492: out = 16'(-16);
			37493: out = 16'(-83);
			37494: out = 16'(-23);
			37495: out = 16'(-74);
			37496: out = 16'(186);
			37497: out = 16'(186);
			37498: out = 16'(236);
			37499: out = 16'(-82);
			37500: out = 16'(-182);
			37501: out = 16'(-199);
			37502: out = 16'(-65);
			37503: out = 16'(-54);
			37504: out = 16'(282);
			37505: out = 16'(-437);
			37506: out = 16'(-930);
			37507: out = 16'(-279);
			37508: out = 16'(404);
			37509: out = 16'(1136);
			37510: out = 16'(1044);
			37511: out = 16'(643);
			37512: out = 16'(-315);
			37513: out = 16'(142);
			37514: out = 16'(175);
			37515: out = 16'(318);
			37516: out = 16'(-21);
			37517: out = 16'(-55);
			37518: out = 16'(165);
			37519: out = 16'(144);
			37520: out = 16'(153);
			37521: out = 16'(134);
			37522: out = 16'(147);
			37523: out = 16'(119);
			37524: out = 16'(146);
			37525: out = 16'(100);
			37526: out = 16'(156);
			37527: out = 16'(171);
			37528: out = 16'(668);
			37529: out = 16'(1303);
			37530: out = 16'(410);
			37531: out = 16'(-359);
			37532: out = 16'(-1586);
			37533: out = 16'(-514);
			37534: out = 16'(-344);
			37535: out = 16'(-654);
			37536: out = 16'(-661);
			37537: out = 16'(-383);
			37538: out = 16'(648);
			37539: out = 16'(607);
			37540: out = 16'(538);
			37541: out = 16'(-168);
			37542: out = 16'(91);
			37543: out = 16'(181);
			37544: out = 16'(-149);
			37545: out = 16'(-823);
			37546: out = 16'(-1449);
			37547: out = 16'(-391);
			37548: out = 16'(-39);
			37549: out = 16'(167);
			37550: out = 16'(-12);
			37551: out = 16'(-171);
			37552: out = 16'(-178);
			37553: out = 16'(-816);
			37554: out = 16'(-805);
			37555: out = 16'(-23);
			37556: out = 16'(144);
			37557: out = 16'(305);
			37558: out = 16'(-243);
			37559: out = 16'(154);
			37560: out = 16'(279);
			37561: out = 16'(241);
			37562: out = 16'(-243);
			37563: out = 16'(-486);
			37564: out = 16'(862);
			37565: out = 16'(1185);
			37566: out = 16'(1270);
			37567: out = 16'(133);
			37568: out = 16'(-266);
			37569: out = 16'(-201);
			37570: out = 16'(-631);
			37571: out = 16'(-447);
			37572: out = 16'(-156);
			37573: out = 16'(473);
			37574: out = 16'(233);
			37575: out = 16'(-1444);
			37576: out = 16'(-1419);
			37577: out = 16'(-1130);
			37578: out = 16'(305);
			37579: out = 16'(108);
			37580: out = 16'(-63);
			37581: out = 16'(224);
			37582: out = 16'(63);
			37583: out = 16'(-86);
			37584: out = 16'(-517);
			37585: out = 16'(-421);
			37586: out = 16'(-129);
			37587: out = 16'(546);
			37588: out = 16'(505);
			37589: out = 16'(-152);
			37590: out = 16'(-357);
			37591: out = 16'(-827);
			37592: out = 16'(-1326);
			37593: out = 16'(-869);
			37594: out = 16'(-112);
			37595: out = 16'(1033);
			37596: out = 16'(1313);
			37597: out = 16'(1330);
			37598: out = 16'(673);
			37599: out = 16'(513);
			37600: out = 16'(75);
			37601: out = 16'(-755);
			37602: out = 16'(-1817);
			37603: out = 16'(-2600);
			37604: out = 16'(-900);
			37605: out = 16'(298);
			37606: out = 16'(1517);
			37607: out = 16'(871);
			37608: out = 16'(354);
			37609: out = 16'(-629);
			37610: out = 16'(-525);
			37611: out = 16'(-428);
			37612: out = 16'(312);
			37613: out = 16'(-60);
			37614: out = 16'(-362);
			37615: out = 16'(-1822);
			37616: out = 16'(-784);
			37617: out = 16'(137);
			37618: out = 16'(1415);
			37619: out = 16'(945);
			37620: out = 16'(288);
			37621: out = 16'(-74);
			37622: out = 16'(66);
			37623: out = 16'(446);
			37624: out = 16'(1834);
			37625: out = 16'(1573);
			37626: out = 16'(127);
			37627: out = 16'(-9);
			37628: out = 16'(-95);
			37629: out = 16'(778);
			37630: out = 16'(288);
			37631: out = 16'(381);
			37632: out = 16'(554);
			37633: out = 16'(446);
			37634: out = 16'(125);
			37635: out = 16'(233);
			37636: out = 16'(-191);
			37637: out = 16'(-238);
			37638: out = 16'(-731);
			37639: out = 16'(-2);
			37640: out = 16'(619);
			37641: out = 16'(669);
			37642: out = 16'(-35);
			37643: out = 16'(-1193);
			37644: out = 16'(-1972);
			37645: out = 16'(-2322);
			37646: out = 16'(-2134);
			37647: out = 16'(-1051);
			37648: out = 16'(-136);
			37649: out = 16'(338);
			37650: out = 16'(414);
			37651: out = 16'(417);
			37652: out = 16'(729);
			37653: out = 16'(709);
			37654: out = 16'(652);
			37655: out = 16'(252);
			37656: out = 16'(-1);
			37657: out = 16'(-200);
			37658: out = 16'(-190);
			37659: out = 16'(-4);
			37660: out = 16'(199);
			37661: out = 16'(-105);
			37662: out = 16'(-206);
			37663: out = 16'(-138);
			37664: out = 16'(166);
			37665: out = 16'(410);
			37666: out = 16'(219);
			37667: out = 16'(1113);
			37668: out = 16'(1392);
			37669: out = 16'(1776);
			37670: out = 16'(-47);
			37671: out = 16'(-1346);
			37672: out = 16'(-1811);
			37673: out = 16'(-752);
			37674: out = 16'(579);
			37675: out = 16'(815);
			37676: out = 16'(944);
			37677: out = 16'(480);
			37678: out = 16'(724);
			37679: out = 16'(179);
			37680: out = 16'(-296);
			37681: out = 16'(-944);
			37682: out = 16'(-744);
			37683: out = 16'(216);
			37684: out = 16'(-1035);
			37685: out = 16'(-1649);
			37686: out = 16'(-2258);
			37687: out = 16'(-603);
			37688: out = 16'(429);
			37689: out = 16'(107);
			37690: out = 16'(310);
			37691: out = 16'(257);
			37692: out = 16'(1113);
			37693: out = 16'(941);
			37694: out = 16'(1028);
			37695: out = 16'(-144);
			37696: out = 16'(581);
			37697: out = 16'(1308);
			37698: out = 16'(1128);
			37699: out = 16'(47);
			37700: out = 16'(-1547);
			37701: out = 16'(-1480);
			37702: out = 16'(-1037);
			37703: out = 16'(-69);
			37704: out = 16'(669);
			37705: out = 16'(826);
			37706: out = 16'(-206);
			37707: out = 16'(-405);
			37708: out = 16'(-581);
			37709: out = 16'(295);
			37710: out = 16'(202);
			37711: out = 16'(227);
			37712: out = 16'(-244);
			37713: out = 16'(-256);
			37714: out = 16'(-249);
			37715: out = 16'(97);
			37716: out = 16'(135);
			37717: out = 16'(85);
			37718: out = 16'(-148);
			37719: out = 16'(-550);
			37720: out = 16'(-1064);
			37721: out = 16'(-717);
			37722: out = 16'(-568);
			37723: out = 16'(-631);
			37724: out = 16'(-317);
			37725: out = 16'(55);
			37726: out = 16'(1103);
			37727: out = 16'(478);
			37728: out = 16'(-51);
			37729: out = 16'(-1411);
			37730: out = 16'(-536);
			37731: out = 16'(342);
			37732: out = 16'(617);
			37733: out = 16'(490);
			37734: out = 16'(349);
			37735: out = 16'(811);
			37736: out = 16'(1591);
			37737: out = 16'(2306);
			37738: out = 16'(2364);
			37739: out = 16'(1431);
			37740: out = 16'(-367);
			37741: out = 16'(-1130);
			37742: out = 16'(-1951);
			37743: out = 16'(-2832);
			37744: out = 16'(-1192);
			37745: out = 16'(279);
			37746: out = 16'(1581);
			37747: out = 16'(880);
			37748: out = 16'(-48);
			37749: out = 16'(-583);
			37750: out = 16'(-366);
			37751: out = 16'(176);
			37752: out = 16'(-192);
			37753: out = 16'(-191);
			37754: out = 16'(-348);
			37755: out = 16'(-1277);
			37756: out = 16'(-1231);
			37757: out = 16'(-521);
			37758: out = 16'(-79);
			37759: out = 16'(254);
			37760: out = 16'(95);
			37761: out = 16'(199);
			37762: out = 16'(104);
			37763: out = 16'(189);
			37764: out = 16'(-42);
			37765: out = 16'(-111);
			37766: out = 16'(-128);
			37767: out = 16'(-140);
			37768: out = 16'(-357);
			37769: out = 16'(-952);
			37770: out = 16'(-861);
			37771: out = 16'(-424);
			37772: out = 16'(-26);
			37773: out = 16'(773);
			37774: out = 16'(1377);
			37775: out = 16'(1397);
			37776: out = 16'(941);
			37777: out = 16'(169);
			37778: out = 16'(192);
			37779: out = 16'(-213);
			37780: out = 16'(-1162);
			37781: out = 16'(-188);
			37782: out = 16'(101);
			37783: out = 16'(-106);
			37784: out = 16'(-709);
			37785: out = 16'(-1006);
			37786: out = 16'(-668);
			37787: out = 16'(252);
			37788: out = 16'(1072);
			37789: out = 16'(262);
			37790: out = 16'(236);
			37791: out = 16'(83);
			37792: out = 16'(-72);
			37793: out = 16'(-55);
			37794: out = 16'(153);
			37795: out = 16'(115);
			37796: out = 16'(18);
			37797: out = 16'(-282);
			37798: out = 16'(28);
			37799: out = 16'(101);
			37800: out = 16'(-165);
			37801: out = 16'(-103);
			37802: out = 16'(-133);
			37803: out = 16'(227);
			37804: out = 16'(-611);
			37805: out = 16'(-832);
			37806: out = 16'(542);
			37807: out = 16'(1013);
			37808: out = 16'(1309);
			37809: out = 16'(1046);
			37810: out = 16'(265);
			37811: out = 16'(-768);
			37812: out = 16'(-190);
			37813: out = 16'(-70);
			37814: out = 16'(276);
			37815: out = 16'(-207);
			37816: out = 16'(-230);
			37817: out = 16'(-153);
			37818: out = 16'(-168);
			37819: out = 16'(-242);
			37820: out = 16'(-666);
			37821: out = 16'(-393);
			37822: out = 16'(-245);
			37823: out = 16'(-242);
			37824: out = 16'(-444);
			37825: out = 16'(-612);
			37826: out = 16'(-247);
			37827: out = 16'(-217);
			37828: out = 16'(-219);
			37829: out = 16'(-208);
			37830: out = 16'(-83);
			37831: out = 16'(236);
			37832: out = 16'(222);
			37833: out = 16'(341);
			37834: out = 16'(217);
			37835: out = 16'(873);
			37836: out = 16'(848);
			37837: out = 16'(660);
			37838: out = 16'(-1292);
			37839: out = 16'(-2519);
			37840: out = 16'(-2096);
			37841: out = 16'(-2073);
			37842: out = 16'(-1326);
			37843: out = 16'(66);
			37844: out = 16'(800);
			37845: out = 16'(1109);
			37846: out = 16'(1122);
			37847: out = 16'(749);
			37848: out = 16'(274);
			37849: out = 16'(648);
			37850: out = 16'(654);
			37851: out = 16'(644);
			37852: out = 16'(-32);
			37853: out = 16'(-227);
			37854: out = 16'(-82);
			37855: out = 16'(156);
			37856: out = 16'(218);
			37857: out = 16'(-271);
			37858: out = 16'(-103);
			37859: out = 16'(-88);
			37860: out = 16'(223);
			37861: out = 16'(-309);
			37862: out = 16'(-608);
			37863: out = 16'(-233);
			37864: out = 16'(-132);
			37865: out = 16'(-60);
			37866: out = 16'(173);
			37867: out = 16'(5);
			37868: out = 16'(-210);
			37869: out = 16'(92);
			37870: out = 16'(277);
			37871: out = 16'(266);
			37872: out = 16'(1084);
			37873: out = 16'(1364);
			37874: out = 16'(1287);
			37875: out = 16'(804);
			37876: out = 16'(553);
			37877: out = 16'(935);
			37878: out = 16'(476);
			37879: out = 16'(-204);
			37880: out = 16'(-1818);
			37881: out = 16'(-1978);
			37882: out = 16'(-1771);
			37883: out = 16'(-1546);
			37884: out = 16'(-760);
			37885: out = 16'(30);
			37886: out = 16'(868);
			37887: out = 16'(799);
			37888: out = 16'(178);
			37889: out = 16'(292);
			37890: out = 16'(194);
			37891: out = 16'(264);
			37892: out = 16'(-124);
			37893: out = 16'(-452);
			37894: out = 16'(-1051);
			37895: out = 16'(-716);
			37896: out = 16'(-582);
			37897: out = 16'(-581);
			37898: out = 16'(-583);
			37899: out = 16'(-474);
			37900: out = 16'(-107);
			37901: out = 16'(128);
			37902: out = 16'(308);
			37903: out = 16'(-46);
			37904: out = 16'(-77);
			37905: out = 16'(-65);
			37906: out = 16'(-54);
			37907: out = 16'(-81);
			37908: out = 16'(-46);
			37909: out = 16'(151);
			37910: out = 16'(113);
			37911: out = 16'(-234);
			37912: out = 16'(671);
			37913: out = 16'(1109);
			37914: out = 16'(1282);
			37915: out = 16'(463);
			37916: out = 16'(-376);
			37917: out = 16'(-453);
			37918: out = 16'(-1327);
			37919: out = 16'(-1709);
			37920: out = 16'(-1040);
			37921: out = 16'(-331);
			37922: out = 16'(441);
			37923: out = 16'(164);
			37924: out = 16'(237);
			37925: out = 16'(153);
			37926: out = 16'(356);
			37927: out = 16'(120);
			37928: out = 16'(-180);
			37929: out = 16'(-225);
			37930: out = 16'(-15);
			37931: out = 16'(279);
			37932: out = 16'(754);
			37933: out = 16'(1067);
			37934: out = 16'(1308);
			37935: out = 16'(464);
			37936: out = 16'(-392);
			37937: out = 16'(-862);
			37938: out = 16'(-1270);
			37939: out = 16'(-1248);
			37940: out = 16'(-351);
			37941: out = 16'(215);
			37942: out = 16'(704);
			37943: out = 16'(582);
			37944: out = 16'(785);
			37945: out = 16'(964);
			37946: out = 16'(1971);
			37947: out = 16'(2157);
			37948: out = 16'(1767);
			37949: out = 16'(671);
			37950: out = 16'(-793);
			37951: out = 16'(-2677);
			37952: out = 16'(-2523);
			37953: out = 16'(-1806);
			37954: out = 16'(-215);
			37955: out = 16'(61);
			37956: out = 16'(46);
			37957: out = 16'(-947);
			37958: out = 16'(-461);
			37959: out = 16'(266);
			37960: out = 16'(-132);
			37961: out = 16'(-65);
			37962: out = 16'(-272);
			37963: out = 16'(-26);
			37964: out = 16'(-172);
			37965: out = 16'(-153);
			37966: out = 16'(-865);
			37967: out = 16'(-672);
			37968: out = 16'(-66);
			37969: out = 16'(680);
			37970: out = 16'(1096);
			37971: out = 16'(1323);
			37972: out = 16'(861);
			37973: out = 16'(461);
			37974: out = 16'(-153);
			37975: out = 16'(40);
			37976: out = 16'(22);
			37977: out = 16'(241);
			37978: out = 16'(-844);
			37979: out = 16'(-1867);
			37980: out = 16'(-2239);
			37981: out = 16'(-940);
			37982: out = 16'(1247);
			37983: out = 16'(2199);
			37984: out = 16'(2230);
			37985: out = 16'(727);
			37986: out = 16'(457);
			37987: out = 16'(-71);
			37988: out = 16'(323);
			37989: out = 16'(-128);
			37990: out = 16'(-458);
			37991: out = 16'(-2317);
			37992: out = 16'(-1894);
			37993: out = 16'(-1708);
			37994: out = 16'(-458);
			37995: out = 16'(-1588);
			37996: out = 16'(-2594);
			37997: out = 16'(-2535);
			37998: out = 16'(-1445);
			37999: out = 16'(218);
			38000: out = 16'(279);
			38001: out = 16'(538);
			38002: out = 16'(255);
			38003: out = 16'(477);
			38004: out = 16'(638);
			38005: out = 16'(1569);
			38006: out = 16'(568);
			38007: out = 16'(47);
			38008: out = 16'(-972);
			38009: out = 16'(419);
			38010: out = 16'(1169);
			38011: out = 16'(1073);
			38012: out = 16'(454);
			38013: out = 16'(-92);
			38014: out = 16'(336);
			38015: out = 16'(310);
			38016: out = 16'(352);
			38017: out = 16'(1269);
			38018: out = 16'(917);
			38019: out = 16'(154);
			38020: out = 16'(-1043);
			38021: out = 16'(-1088);
			38022: out = 16'(-32);
			38023: out = 16'(64);
			38024: out = 16'(584);
			38025: out = 16'(914);
			38026: out = 16'(1260);
			38027: out = 16'(1005);
			38028: out = 16'(-134);
			38029: out = 16'(22);
			38030: out = 16'(135);
			38031: out = 16'(238);
			38032: out = 16'(-20);
			38033: out = 16'(-396);
			38034: out = 16'(-1283);
			38035: out = 16'(-1269);
			38036: out = 16'(-895);
			38037: out = 16'(-346);
			38038: out = 16'(-71);
			38039: out = 16'(-87);
			38040: out = 16'(218);
			38041: out = 16'(408);
			38042: out = 16'(650);
			38043: out = 16'(1078);
			38044: out = 16'(1411);
			38045: out = 16'(1544);
			38046: out = 16'(985);
			38047: out = 16'(180);
			38048: out = 16'(-546);
			38049: out = 16'(-1224);
			38050: out = 16'(-1271);
			38051: out = 16'(-401);
			38052: out = 16'(220);
			38053: out = 16'(605);
			38054: out = 16'(926);
			38055: out = 16'(437);
			38056: out = 16'(-235);
			38057: out = 16'(-265);
			38058: out = 16'(-167);
			38059: out = 16'(83);
			38060: out = 16'(-194);
			38061: out = 16'(-366);
			38062: out = 16'(-218);
			38063: out = 16'(-1104);
			38064: out = 16'(-1580);
			38065: out = 16'(-2258);
			38066: out = 16'(-1369);
			38067: out = 16'(-835);
			38068: out = 16'(-433);
			38069: out = 16'(-1181);
			38070: out = 16'(-1541);
			38071: out = 16'(-1038);
			38072: out = 16'(489);
			38073: out = 16'(1819);
			38074: out = 16'(963);
			38075: out = 16'(-378);
			38076: out = 16'(-2166);
			38077: out = 16'(-2078);
			38078: out = 16'(-1006);
			38079: out = 16'(1347);
			38080: out = 16'(1547);
			38081: out = 16'(1560);
			38082: out = 16'(164);
			38083: out = 16'(405);
			38084: out = 16'(612);
			38085: out = 16'(2077);
			38086: out = 16'(1776);
			38087: out = 16'(1435);
			38088: out = 16'(-32);
			38089: out = 16'(-323);
			38090: out = 16'(-615);
			38091: out = 16'(149);
			38092: out = 16'(-45);
			38093: out = 16'(-132);
			38094: out = 16'(377);
			38095: out = 16'(1367);
			38096: out = 16'(2531);
			38097: out = 16'(1549);
			38098: out = 16'(494);
			38099: out = 16'(-1145);
			38100: out = 16'(-1064);
			38101: out = 16'(-825);
			38102: out = 16'(280);
			38103: out = 16'(-94);
			38104: out = 16'(-375);
			38105: out = 16'(-1817);
			38106: out = 16'(-1527);
			38107: out = 16'(-1215);
			38108: out = 16'(259);
			38109: out = 16'(-154);
			38110: out = 16'(-520);
			38111: out = 16'(-695);
			38112: out = 16'(399);
			38113: out = 16'(1724);
			38114: out = 16'(1717);
			38115: out = 16'(659);
			38116: out = 16'(-1545);
			38117: out = 16'(-1942);
			38118: out = 16'(-1695);
			38119: out = 16'(366);
			38120: out = 16'(53);
			38121: out = 16'(319);
			38122: out = 16'(63);
			38123: out = 16'(757);
			38124: out = 16'(925);
			38125: out = 16'(681);
			38126: out = 16'(175);
			38127: out = 16'(-422);
			38128: out = 16'(-1577);
			38129: out = 16'(-1798);
			38130: out = 16'(-1550);
			38131: out = 16'(273);
			38132: out = 16'(1166);
			38133: out = 16'(1648);
			38134: out = 16'(273);
			38135: out = 16'(-616);
			38136: out = 16'(-1313);
			38137: out = 16'(-555);
			38138: out = 16'(51);
			38139: out = 16'(140);
			38140: out = 16'(346);
			38141: out = 16'(361);
			38142: out = 16'(1082);
			38143: out = 16'(302);
			38144: out = 16'(-355);
			38145: out = 16'(-1287);
			38146: out = 16'(-800);
			38147: out = 16'(-28);
			38148: out = 16'(240);
			38149: out = 16'(210);
			38150: out = 16'(-103);
			38151: out = 16'(-41);
			38152: out = 16'(124);
			38153: out = 16'(715);
			38154: out = 16'(311);
			38155: out = 16'(292);
			38156: out = 16'(218);
			38157: out = 16'(775);
			38158: out = 16'(827);
			38159: out = 16'(99);
			38160: out = 16'(-88);
			38161: out = 16'(-292);
			38162: out = 16'(178);
			38163: out = 16'(-155);
			38164: out = 16'(-181);
			38165: out = 16'(-247);
			38166: out = 16'(543);
			38167: out = 16'(1321);
			38168: out = 16'(1242);
			38169: out = 16'(822);
			38170: out = 16'(71);
			38171: out = 16'(-107);
			38172: out = 16'(-166);
			38173: out = 16'(68);
			38174: out = 16'(21);
			38175: out = 16'(44);
			38176: out = 16'(36);
			38177: out = 16'(-198);
			38178: out = 16'(-528);
			38179: out = 16'(-1496);
			38180: out = 16'(-586);
			38181: out = 16'(343);
			38182: out = 16'(1143);
			38183: out = 16'(761);
			38184: out = 16'(-76);
			38185: out = 16'(-837);
			38186: out = 16'(-1343);
			38187: out = 16'(-1369);
			38188: out = 16'(-1177);
			38189: out = 16'(-549);
			38190: out = 16'(183);
			38191: out = 16'(219);
			38192: out = 16'(242);
			38193: out = 16'(118);
			38194: out = 16'(216);
			38195: out = 16'(285);
			38196: out = 16'(630);
			38197: out = 16'(-173);
			38198: out = 16'(-744);
			38199: out = 16'(-580);
			38200: out = 16'(-668);
			38201: out = 16'(-551);
			38202: out = 16'(-648);
			38203: out = 16'(-310);
			38204: out = 16'(-50);
			38205: out = 16'(154);
			38206: out = 16'(64);
			38207: out = 16'(-61);
			38208: out = 16'(491);
			38209: out = 16'(570);
			38210: out = 16'(165);
			38211: out = 16'(331);
			38212: out = 16'(130);
			38213: out = 16'(232);
			38214: out = 16'(-1245);
			38215: out = 16'(-1818);
			38216: out = 16'(-1827);
			38217: out = 16'(-39);
			38218: out = 16'(1142);
			38219: out = 16'(231);
			38220: out = 16'(139);
			38221: out = 16'(-251);
			38222: out = 16'(355);
			38223: out = 16'(36);
			38224: out = 16'(-169);
			38225: out = 16'(83);
			38226: out = 16'(386);
			38227: out = 16'(629);
			38228: out = 16'(-9);
			38229: out = 16'(-578);
			38230: out = 16'(-1407);
			38231: out = 16'(-215);
			38232: out = 16'(452);
			38233: out = 16'(1027);
			38234: out = 16'(265);
			38235: out = 16'(-169);
			38236: out = 16'(-190);
			38237: out = 16'(85);
			38238: out = 16'(256);
			38239: out = 16'(-69);
			38240: out = 16'(-335);
			38241: out = 16'(-597);
			38242: out = 16'(-587);
			38243: out = 16'(-389);
			38244: out = 16'(-164);
			38245: out = 16'(-35);
			38246: out = 16'(-109);
			38247: out = 16'(14);
			38248: out = 16'(-528);
			38249: out = 16'(-141);
			38250: out = 16'(673);
			38251: out = 16'(1640);
			38252: out = 16'(1845);
			38253: out = 16'(1333);
			38254: out = 16'(-368);
			38255: out = 16'(-1641);
			38256: out = 16'(-1705);
			38257: out = 16'(-968);
			38258: out = 16'(46);
			38259: out = 16'(-167);
			38260: out = 16'(33);
			38261: out = 16'(-118);
			38262: out = 16'(-4);
			38263: out = 16'(26);
			38264: out = 16'(260);
			38265: out = 16'(-59);
			38266: out = 16'(89);
			38267: out = 16'(305);
			38268: out = 16'(-24);
			38269: out = 16'(-398);
			38270: out = 16'(-949);
			38271: out = 16'(-320);
			38272: out = 16'(104);
			38273: out = 16'(304);
			38274: out = 16'(69);
			38275: out = 16'(-175);
			38276: out = 16'(270);
			38277: out = 16'(-33);
			38278: out = 16'(-128);
			38279: out = 16'(-82);
			38280: out = 16'(279);
			38281: out = 16'(693);
			38282: out = 16'(268);
			38283: out = 16'(46);
			38284: out = 16'(-217);
			38285: out = 16'(130);
			38286: out = 16'(186);
			38287: out = 16'(168);
			38288: out = 16'(170);
			38289: out = 16'(215);
			38290: out = 16'(261);
			38291: out = 16'(715);
			38292: out = 16'(973);
			38293: out = 16'(521);
			38294: out = 16'(832);
			38295: out = 16'(839);
			38296: out = 16'(621);
			38297: out = 16'(112);
			38298: out = 16'(-447);
			38299: out = 16'(-1664);
			38300: out = 16'(-1712);
			38301: out = 16'(-1266);
			38302: out = 16'(-793);
			38303: out = 16'(-250);
			38304: out = 16'(198);
			38305: out = 16'(154);
			38306: out = 16'(189);
			38307: out = 16'(144);
			38308: out = 16'(528);
			38309: out = 16'(553);
			38310: out = 16'(286);
			38311: out = 16'(-265);
			38312: out = 16'(-661);
			38313: out = 16'(-555);
			38314: out = 16'(-578);
			38315: out = 16'(-542);
			38316: out = 16'(-212);
			38317: out = 16'(-39);
			38318: out = 16'(281);
			38319: out = 16'(-157);
			38320: out = 16'(521);
			38321: out = 16'(1338);
			38322: out = 16'(1636);
			38323: out = 16'(902);
			38324: out = 16'(-711);
			38325: out = 16'(-1480);
			38326: out = 16'(-1446);
			38327: out = 16'(290);
			38328: out = 16'(50);
			38329: out = 16'(215);
			38330: out = 16'(-212);
			38331: out = 16'(593);
			38332: out = 16'(861);
			38333: out = 16'(-85);
			38334: out = 16'(-143);
			38335: out = 16'(-89);
			38336: out = 16'(197);
			38337: out = 16'(206);
			38338: out = 16'(64);
			38339: out = 16'(-520);
			38340: out = 16'(-548);
			38341: out = 16'(-179);
			38342: out = 16'(-220);
			38343: out = 16'(20);
			38344: out = 16'(217);
			38345: out = 16'(218);
			38346: out = 16'(-63);
			38347: out = 16'(-603);
			38348: out = 16'(-202);
			38349: out = 16'(322);
			38350: out = 16'(501);
			38351: out = 16'(864);
			38352: out = 16'(779);
			38353: out = 16'(279);
			38354: out = 16'(-887);
			38355: out = 16'(-1885);
			38356: out = 16'(-1433);
			38357: out = 16'(-908);
			38358: out = 16'(-120);
			38359: out = 16'(-526);
			38360: out = 16'(-658);
			38361: out = 16'(-930);
			38362: out = 16'(-280);
			38363: out = 16'(356);
			38364: out = 16'(1394);
			38365: out = 16'(1111);
			38366: out = 16'(882);
			38367: out = 16'(635);
			38368: out = 16'(172);
			38369: out = 16'(-187);
			38370: out = 16'(-100);
			38371: out = 16'(38);
			38372: out = 16'(259);
			38373: out = 16'(-227);
			38374: out = 16'(-225);
			38375: out = 16'(-207);
			38376: out = 16'(828);
			38377: out = 16'(677);
			38378: out = 16'(-21);
			38379: out = 16'(-1331);
			38380: out = 16'(-1850);
			38381: out = 16'(-1170);
			38382: out = 16'(-1522);
			38383: out = 16'(-822);
			38384: out = 16'(-174);
			38385: out = 16'(1428);
			38386: out = 16'(1824);
			38387: out = 16'(711);
			38388: out = 16'(103);
			38389: out = 16'(-51);
			38390: out = 16'(833);
			38391: out = 16'(1351);
			38392: out = 16'(1497);
			38393: out = 16'(1448);
			38394: out = 16'(17);
			38395: out = 16'(-1606);
			38396: out = 16'(-2839);
			38397: out = 16'(-2134);
			38398: out = 16'(9);
			38399: out = 16'(889);
			38400: out = 16'(1097);
			38401: out = 16'(-275);
			38402: out = 16'(220);
			38403: out = 16'(472);
			38404: out = 16'(1654);
			38405: out = 16'(1323);
			38406: out = 16'(1067);
			38407: out = 16'(180);
			38408: out = 16'(97);
			38409: out = 16'(42);
			38410: out = 16'(135);
			38411: out = 16'(144);
			38412: out = 16'(108);
			38413: out = 16'(112);
			38414: out = 16'(-446);
			38415: out = 16'(-1159);
			38416: out = 16'(-1389);
			38417: out = 16'(-1219);
			38418: out = 16'(-583);
			38419: out = 16'(-664);
			38420: out = 16'(-525);
			38421: out = 16'(-212);
			38422: out = 16'(-731);
			38423: out = 16'(-1290);
			38424: out = 16'(-2616);
			38425: out = 16'(-1386);
			38426: out = 16'(-54);
			38427: out = 16'(1566);
			38428: out = 16'(1586);
			38429: out = 16'(1190);
			38430: out = 16'(399);
			38431: out = 16'(238);
			38432: out = 16'(245);
			38433: out = 16'(221);
			38434: out = 16'(-164);
			38435: out = 16'(-649);
			38436: out = 16'(-1830);
			38437: out = 16'(-2192);
			38438: out = 16'(-2092);
			38439: out = 16'(-449);
			38440: out = 16'(477);
			38441: out = 16'(306);
			38442: out = 16'(399);
			38443: out = 16'(512);
			38444: out = 16'(1372);
			38445: out = 16'(1524);
			38446: out = 16'(1666);
			38447: out = 16'(1290);
			38448: out = 16'(1142);
			38449: out = 16'(766);
			38450: out = 16'(-62);
			38451: out = 16'(-805);
			38452: out = 16'(-1419);
			38453: out = 16'(-8);
			38454: out = 16'(270);
			38455: out = 16'(208);
			38456: out = 16'(-693);
			38457: out = 16'(-993);
			38458: out = 16'(-520);
			38459: out = 16'(-317);
			38460: out = 16'(208);
			38461: out = 16'(920);
			38462: out = 16'(598);
			38463: out = 16'(-81);
			38464: out = 16'(-1250);
			38465: out = 16'(-1464);
			38466: out = 16'(-1138);
			38467: out = 16'(-364);
			38468: out = 16'(467);
			38469: out = 16'(1007);
			38470: out = 16'(396);
			38471: out = 16'(113);
			38472: out = 16'(-61);
			38473: out = 16'(458);
			38474: out = 16'(596);
			38475: out = 16'(150);
			38476: out = 16'(372);
			38477: out = 16'(12);
			38478: out = 16'(-109);
			38479: out = 16'(-1368);
			38480: out = 16'(-1541);
			38481: out = 16'(-660);
			38482: out = 16'(792);
			38483: out = 16'(1781);
			38484: out = 16'(1629);
			38485: out = 16'(756);
			38486: out = 16'(-343);
			38487: out = 16'(-503);
			38488: out = 16'(-689);
			38489: out = 16'(-580);
			38490: out = 16'(-160);
			38491: out = 16'(-404);
			38492: out = 16'(-1036);
			38493: out = 16'(-2248);
			38494: out = 16'(-1984);
			38495: out = 16'(69);
			38496: out = 16'(-518);
			38497: out = 16'(-480);
			38498: out = 16'(-942);
			38499: out = 16'(185);
			38500: out = 16'(1073);
			38501: out = 16'(1969);
			38502: out = 16'(2079);
			38503: out = 16'(1823);
			38504: out = 16'(1096);
			38505: out = 16'(348);
			38506: out = 16'(-349);
			38507: out = 16'(-186);
			38508: out = 16'(-572);
			38509: out = 16'(-1014);
			38510: out = 16'(-372);
			38511: out = 16'(172);
			38512: out = 16'(1068);
			38513: out = 16'(47);
			38514: out = 16'(-16);
			38515: out = 16'(77);
			38516: out = 16'(1169);
			38517: out = 16'(1673);
			38518: out = 16'(1920);
			38519: out = 16'(540);
			38520: out = 16'(-673);
			38521: out = 16'(-1412);
			38522: out = 16'(-850);
			38523: out = 16'(6);
			38524: out = 16'(420);
			38525: out = 16'(448);
			38526: out = 16'(108);
			38527: out = 16'(128);
			38528: out = 16'(41);
			38529: out = 16'(75);
			38530: out = 16'(189);
			38531: out = 16'(31);
			38532: out = 16'(-339);
			38533: out = 16'(-1406);
			38534: out = 16'(-1832);
			38535: out = 16'(-1301);
			38536: out = 16'(-1191);
			38537: out = 16'(-677);
			38538: out = 16'(121);
			38539: out = 16'(290);
			38540: out = 16'(287);
			38541: out = 16'(276);
			38542: out = 16'(594);
			38543: out = 16'(1085);
			38544: out = 16'(1159);
			38545: out = 16'(1331);
			38546: out = 16'(1064);
			38547: out = 16'(193);
			38548: out = 16'(-1016);
			38549: out = 16'(-2268);
			38550: out = 16'(-1967);
			38551: out = 16'(-1200);
			38552: out = 16'(216);
			38553: out = 16'(164);
			38554: out = 16'(23);
			38555: out = 16'(-582);
			38556: out = 16'(-352);
			38557: out = 16'(-1);
			38558: out = 16'(571);
			38559: out = 16'(1029);
			38560: out = 16'(1232);
			38561: out = 16'(306);
			38562: out = 16'(162);
			38563: out = 16'(109);
			38564: out = 16'(111);
			38565: out = 16'(115);
			38566: out = 16'(112);
			38567: out = 16'(474);
			38568: out = 16'(679);
			38569: out = 16'(909);
			38570: out = 16'(353);
			38571: out = 16'(133);
			38572: out = 16'(141);
			38573: out = 16'(141);
			38574: out = 16'(-197);
			38575: out = 16'(-1017);
			38576: out = 16'(-1316);
			38577: out = 16'(-1364);
			38578: out = 16'(-1056);
			38579: out = 16'(-613);
			38580: out = 16'(-87);
			38581: out = 16'(524);
			38582: out = 16'(626);
			38583: out = 16'(571);
			38584: out = 16'(191);
			38585: out = 16'(38);
			38586: out = 16'(-193);
			38587: out = 16'(237);
			38588: out = 16'(-256);
			38589: out = 16'(-1432);
			38590: out = 16'(-1940);
			38591: out = 16'(-1962);
			38592: out = 16'(-863);
			38593: out = 16'(-732);
			38594: out = 16'(-180);
			38595: out = 16'(987);
			38596: out = 16'(873);
			38597: out = 16'(457);
			38598: out = 16'(-1189);
			38599: out = 16'(-648);
			38600: out = 16'(436);
			38601: out = 16'(508);
			38602: out = 16'(779);
			38603: out = 16'(527);
			38604: out = 16'(214);
			38605: out = 16'(-690);
			38606: out = 16'(-1700);
			38607: out = 16'(-1187);
			38608: out = 16'(-313);
			38609: out = 16'(1053);
			38610: out = 16'(1041);
			38611: out = 16'(934);
			38612: out = 16'(662);
			38613: out = 16'(409);
			38614: out = 16'(178);
			38615: out = 16'(-92);
			38616: out = 16'(-101);
			38617: out = 16'(-123);
			38618: out = 16'(-163);
			38619: out = 16'(-573);
			38620: out = 16'(-976);
			38621: out = 16'(-199);
			38622: out = 16'(80);
			38623: out = 16'(301);
			38624: out = 16'(208);
			38625: out = 16'(83);
			38626: out = 16'(-86);
			38627: out = 16'(97);
			38628: out = 16'(114);
			38629: out = 16'(-261);
			38630: out = 16'(159);
			38631: out = 16'(189);
			38632: out = 16'(-38);
			38633: out = 16'(-605);
			38634: out = 16'(-1023);
			38635: out = 16'(-955);
			38636: out = 16'(-519);
			38637: out = 16'(139);
			38638: out = 16'(841);
			38639: out = 16'(1081);
			38640: out = 16'(908);
			38641: out = 16'(373);
			38642: out = 16'(-169);
			38643: out = 16'(-600);
			38644: out = 16'(-30);
			38645: out = 16'(252);
			38646: out = 16'(245);
			38647: out = 16'(222);
			38648: out = 16'(-29);
			38649: out = 16'(-606);
			38650: out = 16'(-587);
			38651: out = 16'(-482);
			38652: out = 16'(165);
			38653: out = 16'(211);
			38654: out = 16'(329);
			38655: out = 16'(219);
			38656: out = 16'(479);
			38657: out = 16'(543);
			38658: out = 16'(398);
			38659: out = 16'(-317);
			38660: out = 16'(-1026);
			38661: out = 16'(-1346);
			38662: out = 16'(-972);
			38663: out = 16'(-145);
			38664: out = 16'(107);
			38665: out = 16'(166);
			38666: out = 16'(232);
			38667: out = 16'(-634);
			38668: out = 16'(-743);
			38669: out = 16'(157);
			38670: out = 16'(912);
			38671: out = 16'(1407);
			38672: out = 16'(1695);
			38673: out = 16'(477);
			38674: out = 16'(-866);
			38675: out = 16'(-1281);
			38676: out = 16'(-598);
			38677: out = 16'(922);
			38678: out = 16'(1002);
			38679: out = 16'(1660);
			38680: out = 16'(1725);
			38681: out = 16'(1837);
			38682: out = 16'(1411);
			38683: out = 16'(1069);
			38684: out = 16'(256);
			38685: out = 16'(-95);
			38686: out = 16'(-29);
			38687: out = 16'(-184);
			38688: out = 16'(-379);
			38689: out = 16'(-683);
			38690: out = 16'(-948);
			38691: out = 16'(-948);
			38692: out = 16'(-44);
			38693: out = 16'(-129);
			38694: out = 16'(-376);
			38695: out = 16'(-304);
			38696: out = 16'(-212);
			38697: out = 16'(46);
			38698: out = 16'(-1192);
			38699: out = 16'(-1354);
			38700: out = 16'(-1359);
			38701: out = 16'(-157);
			38702: out = 16'(-147);
			38703: out = 16'(-969);
			38704: out = 16'(-1446);
			38705: out = 16'(-1379);
			38706: out = 16'(-131);
			38707: out = 16'(31);
			38708: out = 16'(174);
			38709: out = 16'(-181);
			38710: out = 16'(-157);
			38711: out = 16'(20);
			38712: out = 16'(1123);
			38713: out = 16'(1553);
			38714: out = 16'(1707);
			38715: out = 16'(173);
			38716: out = 16'(-634);
			38717: out = 16'(-1324);
			38718: out = 16'(-989);
			38719: out = 16'(-545);
			38720: out = 16'(241);
			38721: out = 16'(183);
			38722: out = 16'(462);
			38723: out = 16'(908);
			38724: out = 16'(465);
			38725: out = 16'(213);
			38726: out = 16'(610);
			38727: out = 16'(261);
			38728: out = 16'(-102);
			38729: out = 16'(-1672);
			38730: out = 16'(-834);
			38731: out = 16'(44);
			38732: out = 16'(187);
			38733: out = 16'(-176);
			38734: out = 16'(-1010);
			38735: out = 16'(-191);
			38736: out = 16'(-232);
			38737: out = 16'(-106);
			38738: out = 16'(-246);
			38739: out = 16'(108);
			38740: out = 16'(587);
			38741: out = 16'(419);
			38742: out = 16'(70);
			38743: out = 16'(-104);
			38744: out = 16'(-901);
			38745: out = 16'(-1359);
			38746: out = 16'(-2013);
			38747: out = 16'(-683);
			38748: out = 16'(709);
			38749: out = 16'(1717);
			38750: out = 16'(1657);
			38751: out = 16'(1139);
			38752: out = 16'(1547);
			38753: out = 16'(1436);
			38754: out = 16'(1410);
			38755: out = 16'(114);
			38756: out = 16'(-389);
			38757: out = 16'(-612);
			38758: out = 16'(-665);
			38759: out = 16'(-463);
			38760: out = 16'(-154);
			38761: out = 16'(307);
			38762: out = 16'(556);
			38763: out = 16'(492);
			38764: out = 16'(129);
			38765: out = 16'(-249);
			38766: out = 16'(-133);
			38767: out = 16'(-217);
			38768: out = 16'(-125);
			38769: out = 16'(-295);
			38770: out = 16'(-73);
			38771: out = 16'(-13);
			38772: out = 16'(-764);
			38773: out = 16'(-1399);
			38774: out = 16'(-2063);
			38775: out = 16'(-1403);
			38776: out = 16'(-1092);
			38777: out = 16'(-826);
			38778: out = 16'(-270);
			38779: out = 16'(341);
			38780: out = 16'(1286);
			38781: out = 16'(647);
			38782: out = 16'(188);
			38783: out = 16'(235);
			38784: out = 16'(129);
			38785: out = 16'(118);
			38786: out = 16'(-535);
			38787: out = 16'(-277);
			38788: out = 16'(128);
			38789: out = 16'(1878);
			38790: out = 16'(2160);
			38791: out = 16'(1955);
			38792: out = 16'(788);
			38793: out = 16'(245);
			38794: out = 16'(56);
			38795: out = 16'(78);
			38796: out = 16'(197);
			38797: out = 16'(445);
			38798: out = 16'(-518);
			38799: out = 16'(-1530);
			38800: out = 16'(-2844);
			38801: out = 16'(-2210);
			38802: out = 16'(-1262);
			38803: out = 16'(-214);
			38804: out = 16'(138);
			38805: out = 16'(122);
			38806: out = 16'(209);
			38807: out = 16'(101);
			38808: out = 16'(195);
			38809: out = 16'(-233);
			38810: out = 16'(49);
			38811: out = 16'(216);
			38812: out = 16'(602);
			38813: out = 16'(-6);
			38814: out = 16'(-1345);
			38815: out = 16'(-2067);
			38816: out = 16'(-2269);
			38817: out = 16'(-1461);
			38818: out = 16'(-668);
			38819: out = 16'(231);
			38820: out = 16'(213);
			38821: out = 16'(1231);
			38822: out = 16'(1553);
			38823: out = 16'(1035);
			38824: out = 16'(567);
			38825: out = 16'(128);
			38826: out = 16'(-29);
			38827: out = 16'(206);
			38828: out = 16'(661);
			38829: out = 16'(260);
			38830: out = 16'(385);
			38831: out = 16'(577);
			38832: out = 16'(328);
			38833: out = 16'(80);
			38834: out = 16'(-210);
			38835: out = 16'(-140);
			38836: out = 16'(-22);
			38837: out = 16'(123);
			38838: out = 16'(133);
			38839: out = 16'(77);
			38840: out = 16'(-74);
			38841: out = 16'(-354);
			38842: out = 16'(-630);
			38843: out = 16'(-881);
			38844: out = 16'(-756);
			38845: out = 16'(-402);
			38846: out = 16'(17);
			38847: out = 16'(649);
			38848: out = 16'(1247);
			38849: out = 16'(704);
			38850: out = 16'(296);
			38851: out = 16'(-261);
			38852: out = 16'(-112);
			38853: out = 16'(-47);
			38854: out = 16'(277);
			38855: out = 16'(-331);
			38856: out = 16'(-719);
			38857: out = 16'(-1289);
			38858: out = 16'(-809);
			38859: out = 16'(-424);
			38860: out = 16'(-172);
			38861: out = 16'(-112);
			38862: out = 16'(69);
			38863: out = 16'(480);
			38864: out = 16'(1103);
			38865: out = 16'(1532);
			38866: out = 16'(1569);
			38867: out = 16'(814);
			38868: out = 16'(-380);
			38869: out = 16'(-785);
			38870: out = 16'(-813);
			38871: out = 16'(-152);
			38872: out = 16'(-283);
			38873: out = 16'(-243);
			38874: out = 16'(-622);
			38875: out = 16'(-507);
			38876: out = 16'(-589);
			38877: out = 16'(-488);
			38878: out = 16'(-583);
			38879: out = 16'(-294);
			38880: out = 16'(814);
			38881: out = 16'(983);
			38882: out = 16'(761);
			38883: out = 16'(313);
			38884: out = 16'(-408);
			38885: out = 16'(-951);
			38886: out = 16'(-1277);
			38887: out = 16'(-605);
			38888: out = 16'(762);
			38889: out = 16'(1007);
			38890: out = 16'(1143);
			38891: out = 16'(415);
			38892: out = 16'(455);
			38893: out = 16'(-32);
			38894: out = 16'(31);
			38895: out = 16'(-1199);
			38896: out = 16'(-1648);
			38897: out = 16'(-1736);
			38898: out = 16'(-173);
			38899: out = 16'(1184);
			38900: out = 16'(1469);
			38901: out = 16'(963);
			38902: out = 16'(122);
			38903: out = 16'(569);
			38904: out = 16'(626);
			38905: out = 16'(890);
			38906: out = 16'(808);
			38907: out = 16'(732);
			38908: out = 16'(445);
			38909: out = 16'(167);
			38910: out = 16'(-20);
			38911: out = 16'(54);
			38912: out = 16'(-118);
			38913: out = 16'(-304);
			38914: out = 16'(-626);
			38915: out = 16'(-1072);
			38916: out = 16'(-1388);
			38917: out = 16'(-1302);
			38918: out = 16'(-976);
			38919: out = 16'(-347);
			38920: out = 16'(400);
			38921: out = 16'(793);
			38922: out = 16'(787);
			38923: out = 16'(358);
			38924: out = 16'(-14);
			38925: out = 16'(-253);
			38926: out = 16'(-827);
			38927: out = 16'(-840);
			38928: out = 16'(-545);
			38929: out = 16'(-4);
			38930: out = 16'(438);
			38931: out = 16'(875);
			38932: out = 16'(440);
			38933: out = 16'(-270);
			38934: out = 16'(-1598);
			38935: out = 16'(-1674);
			38936: out = 16'(-1522);
			38937: out = 16'(-908);
			38938: out = 16'(-651);
			38939: out = 16'(-399);
			38940: out = 16'(-188);
			38941: out = 16'(2);
			38942: out = 16'(-17);
			38943: out = 16'(615);
			38944: out = 16'(415);
			38945: out = 16'(-22);
			38946: out = 16'(-384);
			38947: out = 16'(-329);
			38948: out = 16'(-15);
			38949: out = 16'(478);
			38950: out = 16'(508);
			38951: out = 16'(-104);
			38952: out = 16'(-1000);
			38953: out = 16'(-1582);
			38954: out = 16'(-747);
			38955: out = 16'(-656);
			38956: out = 16'(-245);
			38957: out = 16'(275);
			38958: out = 16'(437);
			38959: out = 16'(354);
			38960: out = 16'(672);
			38961: out = 16'(880);
			38962: out = 16'(1343);
			38963: out = 16'(375);
			38964: out = 16'(0);
			38965: out = 16'(-577);
			38966: out = 16'(877);
			38967: out = 16'(1134);
			38968: out = 16'(571);
			38969: out = 16'(-116);
			38970: out = 16'(-647);
			38971: out = 16'(-490);
			38972: out = 16'(-356);
			38973: out = 16'(-86);
			38974: out = 16'(-183);
			38975: out = 16'(-118);
			38976: out = 16'(-160);
			38977: out = 16'(-126);
			38978: out = 16'(-5);
			38979: out = 16'(252);
			38980: out = 16'(168);
			38981: out = 16'(159);
			38982: out = 16'(-53);
			38983: out = 16'(737);
			38984: out = 16'(1129);
			38985: out = 16'(1552);
			38986: out = 16'(829);
			38987: out = 16'(390);
			38988: out = 16'(123);
			38989: out = 16'(-46);
			38990: out = 16'(-121);
			38991: out = 16'(225);
			38992: out = 16'(-54);
			38993: out = 16'(-364);
			38994: out = 16'(-1280);
			38995: out = 16'(-788);
			38996: out = 16'(-70);
			38997: out = 16'(144);
			38998: out = 16'(277);
			38999: out = 16'(194);
			39000: out = 16'(-52);
			39001: out = 16'(79);
			39002: out = 16'(604);
			39003: out = 16'(537);
			39004: out = 16'(294);
			39005: out = 16'(-674);
			39006: out = 16'(-56);
			39007: out = 16'(173);
			39008: out = 16'(593);
			39009: out = 16'(-158);
			39010: out = 16'(-686);
			39011: out = 16'(-928);
			39012: out = 16'(-547);
			39013: out = 16'(-259);
			39014: out = 16'(-1162);
			39015: out = 16'(-1425);
			39016: out = 16'(-1492);
			39017: out = 16'(-298);
			39018: out = 16'(514);
			39019: out = 16'(1310);
			39020: out = 16'(490);
			39021: out = 16'(120);
			39022: out = 16'(-175);
			39023: out = 16'(-163);
			39024: out = 16'(-163);
			39025: out = 16'(-174);
			39026: out = 16'(58);
			39027: out = 16'(206);
			39028: out = 16'(150);
			39029: out = 16'(244);
			39030: out = 16'(394);
			39031: out = 16'(1470);
			39032: out = 16'(1072);
			39033: out = 16'(331);
			39034: out = 16'(-684);
			39035: out = 16'(-1071);
			39036: out = 16'(-761);
			39037: out = 16'(-494);
			39038: out = 16'(530);
			39039: out = 16'(1487);
			39040: out = 16'(2020);
			39041: out = 16'(1424);
			39042: out = 16'(-343);
			39043: out = 16'(-997);
			39044: out = 16'(-1133);
			39045: out = 16'(264);
			39046: out = 16'(-47);
			39047: out = 16'(-389);
			39048: out = 16'(-2010);
			39049: out = 16'(-2013);
			39050: out = 16'(-1883);
			39051: out = 16'(-569);
			39052: out = 16'(-625);
			39053: out = 16'(-829);
			39054: out = 16'(-1150);
			39055: out = 16'(-625);
			39056: out = 16'(421);
			39057: out = 16'(765);
			39058: out = 16'(1289);
			39059: out = 16'(1517);
			39060: out = 16'(1186);
			39061: out = 16'(645);
			39062: out = 16'(325);
			39063: out = 16'(-335);
			39064: out = 16'(-657);
			39065: out = 16'(-1328);
			39066: out = 16'(-330);
			39067: out = 16'(387);
			39068: out = 16'(601);
			39069: out = 16'(65);
			39070: out = 16'(-675);
			39071: out = 16'(-1150);
			39072: out = 16'(-970);
			39073: out = 16'(-373);
			39074: out = 16'(122);
			39075: out = 16'(684);
			39076: out = 16'(1296);
			39077: out = 16'(189);
			39078: out = 16'(-19);
			39079: out = 16'(151);
			39080: out = 16'(946);
			39081: out = 16'(981);
			39082: out = 16'(-127);
			39083: out = 16'(-577);
			39084: out = 16'(-873);
			39085: out = 16'(-57);
			39086: out = 16'(-115);
			39087: out = 16'(-32);
			39088: out = 16'(144);
			39089: out = 16'(-9);
			39090: out = 16'(-308);
			39091: out = 16'(-1417);
			39092: out = 16'(-1664);
			39093: out = 16'(-1497);
			39094: out = 16'(-704);
			39095: out = 16'(-150);
			39096: out = 16'(296);
			39097: out = 16'(521);
			39098: out = 16'(922);
			39099: out = 16'(1226);
			39100: out = 16'(1926);
			39101: out = 16'(2130);
			39102: out = 16'(2129);
			39103: out = 16'(901);
			39104: out = 16'(-338);
			39105: out = 16'(-1624);
			39106: out = 16'(-1025);
			39107: out = 16'(-21);
			39108: out = 16'(74);
			39109: out = 16'(269);
			39110: out = 16'(0);
			39111: out = 16'(-135);
			39112: out = 16'(-264);
			39113: out = 16'(-52);
			39114: out = 16'(-205);
			39115: out = 16'(23);
			39116: out = 16'(172);
			39117: out = 16'(265);
			39118: out = 16'(70);
			39119: out = 16'(-195);
			39120: out = 16'(-947);
			39121: out = 16'(-1284);
			39122: out = 16'(-890);
			39123: out = 16'(-699);
			39124: out = 16'(-432);
			39125: out = 16'(-213);
			39126: out = 16'(33);
			39127: out = 16'(162);
			39128: out = 16'(-452);
			39129: out = 16'(-635);
			39130: out = 16'(-858);
			39131: out = 16'(-88);
			39132: out = 16'(25);
			39133: out = 16'(286);
			39134: out = 16'(-1280);
			39135: out = 16'(-1085);
			39136: out = 16'(322);
			39137: out = 16'(771);
			39138: out = 16'(848);
			39139: out = 16'(-48);
			39140: out = 16'(-81);
			39141: out = 16'(0);
			39142: out = 16'(606);
			39143: out = 16'(1161);
			39144: out = 16'(1554);
			39145: out = 16'(953);
			39146: out = 16'(431);
			39147: out = 16'(-214);
			39148: out = 16'(-63);
			39149: out = 16'(-140);
			39150: out = 16'(-74);
			39151: out = 16'(147);
			39152: out = 16'(254);
			39153: out = 16'(208);
			39154: out = 16'(151);
			39155: out = 16'(140);
			39156: out = 16'(227);
			39157: out = 16'(432);
			39158: out = 16'(481);
			39159: out = 16'(104);
			39160: out = 16'(-283);
			39161: out = 16'(-756);
			39162: out = 16'(-1187);
			39163: out = 16'(-1499);
			39164: out = 16'(-1568);
			39165: out = 16'(-1255);
			39166: out = 16'(-675);
			39167: out = 16'(124);
			39168: out = 16'(-496);
			39169: out = 16'(-104);
			39170: out = 16'(224);
			39171: out = 16'(939);
			39172: out = 16'(518);
			39173: out = 16'(-475);
			39174: out = 16'(-1034);
			39175: out = 16'(-823);
			39176: out = 16'(366);
			39177: out = 16'(948);
			39178: out = 16'(1256);
			39179: out = 16'(619);
			39180: out = 16'(237);
			39181: out = 16'(-288);
			39182: out = 16'(-442);
			39183: out = 16'(-376);
			39184: out = 16'(-80);
			39185: out = 16'(-51);
			39186: out = 16'(-50);
			39187: out = 16'(-146);
			39188: out = 16'(-46);
			39189: out = 16'(188);
			39190: out = 16'(674);
			39191: out = 16'(278);
			39192: out = 16'(129);
			39193: out = 16'(-59);
			39194: out = 16'(-45);
			39195: out = 16'(-70);
			39196: out = 16'(-153);
			39197: out = 16'(-168);
			39198: out = 16'(-46);
			39199: out = 16'(632);
			39200: out = 16'(247);
			39201: out = 16'(-224);
			39202: out = 16'(-1109);
			39203: out = 16'(-939);
			39204: out = 16'(-346);
			39205: out = 16'(-144);
			39206: out = 16'(168);
			39207: out = 16'(316);
			39208: out = 16'(851);
			39209: out = 16'(954);
			39210: out = 16'(920);
			39211: out = 16'(196);
			39212: out = 16'(-188);
			39213: out = 16'(-140);
			39214: out = 16'(-169);
			39215: out = 16'(140);
			39216: out = 16'(854);
			39217: out = 16'(1091);
			39218: out = 16'(1101);
			39219: out = 16'(551);
			39220: out = 16'(315);
			39221: out = 16'(-25);
			39222: out = 16'(-517);
			39223: out = 16'(-660);
			39224: out = 16'(-533);
			39225: out = 16'(-253);
			39226: out = 16'(153);
			39227: out = 16'(529);
			39228: out = 16'(46);
			39229: out = 16'(-494);
			39230: out = 16'(-1308);
			39231: out = 16'(-1040);
			39232: out = 16'(-671);
			39233: out = 16'(174);
			39234: out = 16'(-58);
			39235: out = 16'(-299);
			39236: out = 16'(-868);
			39237: out = 16'(-691);
			39238: out = 16'(-404);
			39239: out = 16'(-82);
			39240: out = 16'(97);
			39241: out = 16'(130);
			39242: out = 16'(-1027);
			39243: out = 16'(-1244);
			39244: out = 16'(-1142);
			39245: out = 16'(-622);
			39246: out = 16'(-174);
			39247: out = 16'(294);
			39248: out = 16'(534);
			39249: out = 16'(812);
			39250: out = 16'(934);
			39251: out = 16'(1211);
			39252: out = 16'(1160);
			39253: out = 16'(974);
			39254: out = 16'(42);
			39255: out = 16'(-608);
			39256: out = 16'(-193);
			39257: out = 16'(180);
			39258: out = 16'(629);
			39259: out = 16'(-106);
			39260: out = 16'(-51);
			39261: out = 16'(-124);
			39262: out = 16'(537);
			39263: out = 16'(301);
			39264: out = 16'(-110);
			39265: out = 16'(131);
			39266: out = 16'(346);
			39267: out = 16'(522);
			39268: out = 16'(115);
			39269: out = 16'(-267);
			39270: out = 16'(-112);
			39271: out = 16'(-1223);
			39272: out = 16'(-1727);
			39273: out = 16'(-2070);
			39274: out = 16'(-726);
			39275: out = 16'(497);
			39276: out = 16'(1177);
			39277: out = 16'(794);
			39278: out = 16'(52);
			39279: out = 16'(-24);
			39280: out = 16'(405);
			39281: out = 16'(1324);
			39282: out = 16'(320);
			39283: out = 16'(117);
			39284: out = 16'(-294);
			39285: out = 16'(99);
			39286: out = 16'(84);
			39287: out = 16'(162);
			39288: out = 16'(-182);
			39289: out = 16'(-133);
			39290: out = 16'(76);
			39291: out = 16'(421);
			39292: out = 16'(574);
			39293: out = 16'(891);
			39294: out = 16'(241);
			39295: out = 16'(-340);
			39296: out = 16'(-237);
			39297: out = 16'(-70);
			39298: out = 16'(148);
			39299: out = 16'(-1102);
			39300: out = 16'(-1764);
			39301: out = 16'(-2404);
			39302: out = 16'(-236);
			39303: out = 16'(766);
			39304: out = 16'(1582);
			39305: out = 16'(309);
			39306: out = 16'(-123);
			39307: out = 16'(207);
			39308: out = 16'(369);
			39309: out = 16'(609);
			39310: out = 16'(496);
			39311: out = 16'(231);
			39312: out = 16'(-378);
			39313: out = 16'(-770);
			39314: out = 16'(-1421);
			39315: out = 16'(-1464);
			39316: out = 16'(-435);
			39317: out = 16'(565);
			39318: out = 16'(1232);
			39319: out = 16'(1553);
			39320: out = 16'(977);
			39321: out = 16'(142);
			39322: out = 16'(-1002);
			39323: out = 16'(-942);
			39324: out = 16'(323);
			39325: out = 16'(625);
			39326: out = 16'(787);
			39327: out = 16'(23);
			39328: out = 16'(-78);
			39329: out = 16'(-453);
			39330: out = 16'(-911);
			39331: out = 16'(-786);
			39332: out = 16'(-452);
			39333: out = 16'(45);
			39334: out = 16'(8);
			39335: out = 16'(-255);
			39336: out = 16'(-59);
			39337: out = 16'(-51);
			39338: out = 16'(166);
			39339: out = 16'(-1070);
			39340: out = 16'(-1266);
			39341: out = 16'(-1222);
			39342: out = 16'(-149);
			39343: out = 16'(305);
			39344: out = 16'(281);
			39345: out = 16'(311);
			39346: out = 16'(223);
			39347: out = 16'(-73);
			39348: out = 16'(354);
			39349: out = 16'(545);
			39350: out = 16'(-57);
			39351: out = 16'(-278);
			39352: out = 16'(-531);
			39353: out = 16'(164);
			39354: out = 16'(-5);
			39355: out = 16'(-191);
			39356: out = 16'(-498);
			39357: out = 16'(-262);
			39358: out = 16'(246);
			39359: out = 16'(-56);
			39360: out = 16'(144);
			39361: out = 16'(643);
			39362: out = 16'(583);
			39363: out = 16'(447);
			39364: out = 16'(-264);
			39365: out = 16'(146);
			39366: out = 16'(320);
			39367: out = 16'(959);
			39368: out = 16'(20);
			39369: out = 16'(-690);
			39370: out = 16'(-907);
			39371: out = 16'(-501);
			39372: out = 16'(-53);
			39373: out = 16'(-463);
			39374: out = 16'(-832);
			39375: out = 16'(-1199);
			39376: out = 16'(-44);
			39377: out = 16'(428);
			39378: out = 16'(621);
			39379: out = 16'(1374);
			39380: out = 16'(1460);
			39381: out = 16'(1166);
			39382: out = 16'(202);
			39383: out = 16'(-285);
			39384: out = 16'(168);
			39385: out = 16'(116);
			39386: out = 16'(188);
			39387: out = 16'(-290);
			39388: out = 16'(207);
			39389: out = 16'(542);
			39390: out = 16'(172);
			39391: out = 16'(161);
			39392: out = 16'(77);
			39393: out = 16'(797);
			39394: out = 16'(413);
			39395: out = 16'(-286);
			39396: out = 16'(-793);
			39397: out = 16'(-1067);
			39398: out = 16'(-930);
			39399: out = 16'(-1241);
			39400: out = 16'(-1198);
			39401: out = 16'(-872);
			39402: out = 16'(-478);
			39403: out = 16'(32);
			39404: out = 16'(186);
			39405: out = 16'(743);
			39406: out = 16'(808);
			39407: out = 16'(697);
			39408: out = 16'(-609);
			39409: out = 16'(-1831);
			39410: out = 16'(-1931);
			39411: out = 16'(-1521);
			39412: out = 16'(-629);
			39413: out = 16'(-3);
			39414: out = 16'(340);
			39415: out = 16'(154);
			39416: out = 16'(107);
			39417: out = 16'(-6);
			39418: out = 16'(321);
			39419: out = 16'(-51);
			39420: out = 16'(474);
			39421: out = 16'(1883);
			39422: out = 16'(1668);
			39423: out = 16'(1329);
			39424: out = 16'(576);
			39425: out = 16'(726);
			39426: out = 16'(845);
			39427: out = 16'(475);
			39428: out = 16'(849);
			39429: out = 16'(1059);
			39430: out = 16'(250);
			39431: out = 16'(-194);
			39432: out = 16'(-740);
			39433: out = 16'(-874);
			39434: out = 16'(-1165);
			39435: out = 16'(-1280);
			39436: out = 16'(-1072);
			39437: out = 16'(-631);
			39438: out = 16'(-98);
			39439: out = 16'(109);
			39440: out = 16'(-58);
			39441: out = 16'(-916);
			39442: out = 16'(-876);
			39443: out = 16'(-822);
			39444: out = 16'(-501);
			39445: out = 16'(-265);
			39446: out = 16'(50);
			39447: out = 16'(-97);
			39448: out = 16'(147);
			39449: out = 16'(184);
			39450: out = 16'(643);
			39451: out = 16'(442);
			39452: out = 16'(285);
			39453: out = 16'(-995);
			39454: out = 16'(-1029);
			39455: out = 16'(-429);
			39456: out = 16'(569);
			39457: out = 16'(1041);
			39458: out = 16'(914);
			39459: out = 16'(473);
			39460: out = 16'(342);
			39461: out = 16'(875);
			39462: out = 16'(1582);
			39463: out = 16'(1962);
			39464: out = 16'(499);
			39465: out = 16'(187);
			39466: out = 16'(-320);
			39467: out = 16'(-74);
			39468: out = 16'(-724);
			39469: out = 16'(-1358);
			39470: out = 16'(-1799);
			39471: out = 16'(-1814);
			39472: out = 16'(-1422);
			39473: out = 16'(-763);
			39474: out = 16'(-160);
			39475: out = 16'(116);
			39476: out = 16'(541);
			39477: out = 16'(383);
			39478: out = 16'(-81);
			39479: out = 16'(-1041);
			39480: out = 16'(-1263);
			39481: out = 16'(182);
			39482: out = 16'(402);
			39483: out = 16'(609);
			39484: out = 16'(283);
			39485: out = 16'(133);
			39486: out = 16'(-73);
			39487: out = 16'(190);
			39488: out = 16'(78);
			39489: out = 16'(-53);
			39490: out = 16'(211);
			39491: out = 16'(166);
			39492: out = 16'(-76);
			39493: out = 16'(130);
			39494: out = 16'(102);
			39495: out = 16'(-66);
			39496: out = 16'(328);
			39497: out = 16'(603);
			39498: out = 16'(487);
			39499: out = 16'(722);
			39500: out = 16'(838);
			39501: out = 16'(1061);
			39502: out = 16'(890);
			39503: out = 16'(732);
			39504: out = 16'(728);
			39505: out = 16'(718);
			39506: out = 16'(585);
			39507: out = 16'(-382);
			39508: out = 16'(-1201);
			39509: out = 16'(-2056);
			39510: out = 16'(-1685);
			39511: out = 16'(-1286);
			39512: out = 16'(-476);
			39513: out = 16'(-1055);
			39514: out = 16'(-1098);
			39515: out = 16'(-828);
			39516: out = 16'(-325);
			39517: out = 16'(11);
			39518: out = 16'(-180);
			39519: out = 16'(46);
			39520: out = 16'(158);
			39521: out = 16'(-36);
			39522: out = 16'(-85);
			39523: out = 16'(-130);
			39524: out = 16'(134);
			39525: out = 16'(209);
			39526: out = 16'(282);
			39527: out = 16'(168);
			39528: out = 16'(100);
			39529: out = 16'(-96);
			39530: out = 16'(889);
			39531: out = 16'(990);
			39532: out = 16'(472);
			39533: out = 16'(54);
			39534: out = 16'(-313);
			39535: out = 16'(-147);
			39536: out = 16'(-30);
			39537: out = 16'(438);
			39538: out = 16'(962);
			39539: out = 16'(1283);
			39540: out = 16'(1236);
			39541: out = 16'(1107);
			39542: out = 16'(530);
			39543: out = 16'(31);
			39544: out = 16'(-193);
			39545: out = 16'(-237);
			39546: out = 16'(-379);
			39547: out = 16'(-476);
			39548: out = 16'(-1230);
			39549: out = 16'(-2359);
			39550: out = 16'(-2338);
			39551: out = 16'(-1673);
			39552: out = 16'(239);
			39553: out = 16'(-39);
			39554: out = 16'(-97);
			39555: out = 16'(-513);
			39556: out = 16'(-93);
			39557: out = 16'(308);
			39558: out = 16'(804);
			39559: out = 16'(998);
			39560: out = 16'(1054);
			39561: out = 16'(265);
			39562: out = 16'(151);
			39563: out = 16'(74);
			39564: out = 16'(206);
			39565: out = 16'(47);
			39566: out = 16'(-145);
			39567: out = 16'(-209);
			39568: out = 16'(-149);
			39569: out = 16'(114);
			39570: out = 16'(141);
			39571: out = 16'(247);
			39572: out = 16'(489);
			39573: out = 16'(264);
			39574: out = 16'(190);
			39575: out = 16'(431);
			39576: out = 16'(768);
			39577: out = 16'(969);
			39578: out = 16'(50);
			39579: out = 16'(-410);
			39580: out = 16'(-1044);
			39581: out = 16'(68);
			39582: out = 16'(-451);
			39583: out = 16'(-945);
			39584: out = 16'(-2170);
			39585: out = 16'(-1504);
			39586: out = 16'(275);
			39587: out = 16'(589);
			39588: out = 16'(743);
			39589: out = 16'(0);
			39590: out = 16'(-247);
			39591: out = 16'(-739);
			39592: out = 16'(-742);
			39593: out = 16'(-1141);
			39594: out = 16'(-946);
			39595: out = 16'(-264);
			39596: out = 16'(448);
			39597: out = 16'(958);
			39598: out = 16'(1387);
			39599: out = 16'(1130);
			39600: out = 16'(738);
			39601: out = 16'(808);
			39602: out = 16'(641);
			39603: out = 16'(387);
			39604: out = 16'(-58);
			39605: out = 16'(-644);
			39606: out = 16'(-1248);
			39607: out = 16'(-1499);
			39608: out = 16'(-1351);
			39609: out = 16'(-817);
			39610: out = 16'(-183);
			39611: out = 16'(256);
			39612: out = 16'(97);
			39613: out = 16'(571);
			39614: out = 16'(1038);
			39615: out = 16'(1852);
			39616: out = 16'(1807);
			39617: out = 16'(1351);
			39618: out = 16'(78);
			39619: out = 16'(-741);
			39620: out = 16'(-1319);
			39621: out = 16'(-1833);
			39622: out = 16'(-1897);
			39623: out = 16'(-1862);
			39624: out = 16'(-516);
			39625: out = 16'(42);
			39626: out = 16'(299);
			39627: out = 16'(-281);
			39628: out = 16'(-398);
			39629: out = 16'(-165);
			39630: out = 16'(552);
			39631: out = 16'(790);
			39632: out = 16'(313);
			39633: out = 16'(-513);
			39634: out = 16'(-1230);
			39635: out = 16'(-1102);
			39636: out = 16'(-619);
			39637: out = 16'(199);
			39638: out = 16'(953);
			39639: out = 16'(1361);
			39640: out = 16'(1353);
			39641: out = 16'(431);
			39642: out = 16'(-251);
			39643: out = 16'(-846);
			39644: out = 16'(190);
			39645: out = 16'(689);
			39646: out = 16'(797);
			39647: out = 16'(-13);
			39648: out = 16'(-902);
			39649: out = 16'(-1817);
			39650: out = 16'(-1497);
			39651: out = 16'(-803);
			39652: out = 16'(188);
			39653: out = 16'(486);
			39654: out = 16'(624);
			39655: out = 16'(816);
			39656: out = 16'(1125);
			39657: out = 16'(1416);
			39658: out = 16'(1125);
			39659: out = 16'(753);
			39660: out = 16'(70);
			39661: out = 16'(238);
			39662: out = 16'(0);
			39663: out = 16'(-122);
			39664: out = 16'(-721);
			39665: out = 16'(-776);
			39666: out = 16'(-205);
			39667: out = 16'(-149);
			39668: out = 16'(-117);
			39669: out = 16'(-214);
			39670: out = 16'(-155);
			39671: out = 16'(33);
			39672: out = 16'(1006);
			39673: out = 16'(1093);
			39674: out = 16'(945);
			39675: out = 16'(204);
			39676: out = 16'(-391);
			39677: out = 16'(-943);
			39678: out = 16'(-82);
			39679: out = 16'(122);
			39680: out = 16'(161);
			39681: out = 16'(-160);
			39682: out = 16'(-278);
			39683: out = 16'(-238);
			39684: out = 16'(-44);
			39685: out = 16'(117);
			39686: out = 16'(142);
			39687: out = 16'(177);
			39688: out = 16'(124);
			39689: out = 16'(79);
			39690: out = 16'(-56);
			39691: out = 16'(-204);
			39692: out = 16'(-225);
			39693: out = 16'(-576);
			39694: out = 16'(-938);
			39695: out = 16'(-582);
			39696: out = 16'(-472);
			39697: out = 16'(-155);
			39698: out = 16'(-301);
			39699: out = 16'(-9);
			39700: out = 16'(159);
			39701: out = 16'(930);
			39702: out = 16'(827);
			39703: out = 16'(86);
			39704: out = 16'(-1035);
			39705: out = 16'(-1398);
			39706: out = 16'(166);
			39707: out = 16'(-61);
			39708: out = 16'(-125);
			39709: out = 16'(-550);
			39710: out = 16'(-345);
			39711: out = 16'(-203);
			39712: out = 16'(-466);
			39713: out = 16'(-659);
			39714: out = 16'(-793);
			39715: out = 16'(14);
			39716: out = 16'(184);
			39717: out = 16'(132);
			39718: out = 16'(-337);
			39719: out = 16'(-444);
			39720: out = 16'(-90);
			39721: out = 16'(-403);
			39722: out = 16'(-525);
			39723: out = 16'(-823);
			39724: out = 16'(-269);
			39725: out = 16'(32);
			39726: out = 16'(-35);
			39727: out = 16'(93);
			39728: out = 16'(360);
			39729: out = 16'(1355);
			39730: out = 16'(1586);
			39731: out = 16'(1634);
			39732: out = 16'(1166);
			39733: out = 16'(816);
			39734: out = 16'(386);
			39735: out = 16'(-26);
			39736: out = 16'(-227);
			39737: out = 16'(-117);
			39738: out = 16'(-282);
			39739: out = 16'(-283);
			39740: out = 16'(-640);
			39741: out = 16'(193);
			39742: out = 16'(536);
			39743: out = 16'(793);
			39744: out = 16'(144);
			39745: out = 16'(-469);
			39746: out = 16'(-1221);
			39747: out = 16'(-710);
			39748: out = 16'(-193);
			39749: out = 16'(-523);
			39750: out = 16'(-964);
			39751: out = 16'(-1544);
			39752: out = 16'(-626);
			39753: out = 16'(-93);
			39754: out = 16'(647);
			39755: out = 16'(257);
			39756: out = 16'(245);
			39757: out = 16'(107);
			39758: out = 16'(163);
			39759: out = 16'(-46);
			39760: out = 16'(-506);
			39761: out = 16'(-116);
			39762: out = 16'(343);
			39763: out = 16'(765);
			39764: out = 16'(867);
			39765: out = 16'(700);
			39766: out = 16'(563);
			39767: out = 16'(229);
			39768: out = 16'(70);
			39769: out = 16'(-303);
			39770: out = 16'(330);
			39771: out = 16'(1088);
			39772: out = 16'(805);
			39773: out = 16'(377);
			39774: out = 16'(-350);
			39775: out = 16'(-210);
			39776: out = 16'(-32);
			39777: out = 16'(444);
			39778: out = 16'(-11);
			39779: out = 16'(-348);
			39780: out = 16'(-550);
			39781: out = 16'(-1286);
			39782: out = 16'(-1494);
			39783: out = 16'(-584);
			39784: out = 16'(-144);
			39785: out = 16'(265);
			39786: out = 16'(65);
			39787: out = 16'(31);
			39788: out = 16'(-140);
			39789: out = 16'(475);
			39790: out = 16'(97);
			39791: out = 16'(-640);
			39792: out = 16'(-506);
			39793: out = 16'(-416);
			39794: out = 16'(204);
			39795: out = 16'(-729);
			39796: out = 16'(-567);
			39797: out = 16'(63);
			39798: out = 16'(1011);
			39799: out = 16'(1365);
			39800: out = 16'(1066);
			39801: out = 16'(464);
			39802: out = 16'(-67);
			39803: out = 16'(-263);
			39804: out = 16'(-109);
			39805: out = 16'(41);
			39806: out = 16'(93);
			39807: out = 16'(-276);
			39808: out = 16'(-548);
			39809: out = 16'(-438);
			39810: out = 16'(422);
			39811: out = 16'(1335);
			39812: out = 16'(1404);
			39813: out = 16'(479);
			39814: out = 16'(-1351);
			39815: out = 16'(-1808);
			39816: out = 16'(-1534);
			39817: out = 16'(116);
			39818: out = 16'(148);
			39819: out = 16'(124);
			39820: out = 16'(178);
			39821: out = 16'(-905);
			39822: out = 16'(-1652);
			39823: out = 16'(-1934);
			39824: out = 16'(-663);
			39825: out = 16'(751);
			39826: out = 16'(817);
			39827: out = 16'(-47);
			39828: out = 16'(-1729);
			39829: out = 16'(-1362);
			39830: out = 16'(-1225);
			39831: out = 16'(-264);
			39832: out = 16'(-554);
			39833: out = 16'(-178);
			39834: out = 16'(-46);
			39835: out = 16'(475);
			39836: out = 16'(685);
			39837: out = 16'(926);
			39838: out = 16'(854);
			39839: out = 16'(858);
			39840: out = 16'(521);
			39841: out = 16'(736);
			39842: out = 16'(798);
			39843: out = 16'(872);
			39844: out = 16'(331);
			39845: out = 16'(-189);
			39846: out = 16'(-121);
			39847: out = 16'(-23);
			39848: out = 16'(219);
			39849: out = 16'(91);
			39850: out = 16'(84);
			39851: out = 16'(77);
			39852: out = 16'(91);
			39853: out = 16'(-56);
			39854: out = 16'(-621);
			39855: out = 16'(-83);
			39856: out = 16'(29);
			39857: out = 16'(-182);
			39858: out = 16'(-819);
			39859: out = 16'(-1082);
			39860: out = 16'(80);
			39861: out = 16'(334);
			39862: out = 16'(496);
			39863: out = 16'(-151);
			39864: out = 16'(-221);
			39865: out = 16'(-172);
			39866: out = 16'(152);
			39867: out = 16'(217);
			39868: out = 16'(163);
			39869: out = 16'(243);
			39870: out = 16'(47);
			39871: out = 16'(-177);
			39872: out = 16'(-935);
			39873: out = 16'(-1126);
			39874: out = 16'(-811);
			39875: out = 16'(-206);
			39876: out = 16'(228);
			39877: out = 16'(-92);
			39878: out = 16'(-30);
			39879: out = 16'(-36);
			39880: out = 16'(256);
			39881: out = 16'(246);
			39882: out = 16'(285);
			39883: out = 16'(487);
			39884: out = 16'(562);
			39885: out = 16'(493);
			39886: out = 16'(222);
			39887: out = 16'(-127);
			39888: out = 16'(-535);
			39889: out = 16'(-182);
			39890: out = 16'(-75);
			39891: out = 16'(-88);
			39892: out = 16'(53);
			39893: out = 16'(126);
			39894: out = 16'(-122);
			39895: out = 16'(115);
			39896: out = 16'(206);
			39897: out = 16'(241);
			39898: out = 16'(134);
			39899: out = 16'(72);
			39900: out = 16'(-878);
			39901: out = 16'(-73);
			39902: out = 16'(932);
			39903: out = 16'(1022);
			39904: out = 16'(679);
			39905: out = 16'(-265);
			39906: out = 16'(131);
			39907: out = 16'(-180);
			39908: out = 16'(-535);
			39909: out = 16'(-136);
			39910: out = 16'(189);
			39911: out = 16'(100);
			39912: out = 16'(247);
			39913: out = 16'(19);
			39914: out = 16'(-118);
			39915: out = 16'(-1055);
			39916: out = 16'(-1524);
			39917: out = 16'(-903);
			39918: out = 16'(-504);
			39919: out = 16'(-129);
			39920: out = 16'(-177);
			39921: out = 16'(-121);
			39922: out = 16'(-19);
			39923: out = 16'(-131);
			39924: out = 16'(282);
			39925: out = 16'(850);
			39926: out = 16'(872);
			39927: out = 16'(442);
			39928: out = 16'(-555);
			39929: out = 16'(-1402);
			39930: out = 16'(-1972);
			39931: out = 16'(-1729);
			39932: out = 16'(-1464);
			39933: out = 16'(-764);
			39934: out = 16'(-97);
			39935: out = 16'(437);
			39936: out = 16'(699);
			39937: out = 16'(1184);
			39938: out = 16'(1058);
			39939: out = 16'(798);
			39940: out = 16'(-238);
			39941: out = 16'(-751);
			39942: out = 16'(-1117);
			39943: out = 16'(-217);
			39944: out = 16'(207);
			39945: out = 16'(616);
			39946: out = 16'(-135);
			39947: out = 16'(-709);
			39948: out = 16'(-1460);
			39949: out = 16'(-557);
			39950: out = 16'(234);
			39951: out = 16'(1210);
			39952: out = 16'(712);
			39953: out = 16'(87);
			39954: out = 16'(-1048);
			39955: out = 16'(-490);
			39956: out = 16'(396);
			39957: out = 16'(794);
			39958: out = 16'(563);
			39959: out = 16'(-145);
			39960: out = 16'(291);
			39961: out = 16'(400);
			39962: out = 16'(961);
			39963: out = 16'(286);
			39964: out = 16'(377);
			39965: out = 16'(467);
			39966: out = 16'(1200);
			39967: out = 16'(1046);
			39968: out = 16'(-147);
			39969: out = 16'(-390);
			39970: out = 16'(-501);
			39971: out = 16'(96);
			39972: out = 16'(-96);
			39973: out = 16'(-262);
			39974: out = 16'(-197);
			39975: out = 16'(-397);
			39976: out = 16'(-501);
			39977: out = 16'(-282);
			39978: out = 16'(223);
			39979: out = 16'(863);
			39980: out = 16'(527);
			39981: out = 16'(278);
			39982: out = 16'(-292);
			39983: out = 16'(-198);
			39984: out = 16'(-166);
			39985: out = 16'(238);
			39986: out = 16'(-115);
			39987: out = 16'(-510);
			39988: out = 16'(-1977);
			39989: out = 16'(-999);
			39990: out = 16'(-416);
			39991: out = 16'(-120);
			39992: out = 16'(-861);
			39993: out = 16'(-1492);
			39994: out = 16'(-834);
			39995: out = 16'(-126);
			39996: out = 16'(726);
			39997: out = 16'(558);
			39998: out = 16'(521);
			39999: out = 16'(109);
			40000: out = 16'(56);
			40001: out = 16'(80);
			40002: out = 16'(677);
			40003: out = 16'(0);
			40004: out = 16'(-286);
			40005: out = 16'(-868);
			40006: out = 16'(161);
			40007: out = 16'(649);
			40008: out = 16'(549);
			40009: out = 16'(212);
			40010: out = 16'(-75);
			40011: out = 16'(270);
			40012: out = 16'(219);
			40013: out = 16'(221);
			40014: out = 16'(-62);
			40015: out = 16'(40);
			40016: out = 16'(252);
			40017: out = 16'(-74);
			40018: out = 16'(7);
			40019: out = 16'(128);
			40020: out = 16'(144);
			40021: out = 16'(3);
			40022: out = 16'(-179);
			40023: out = 16'(-678);
			40024: out = 16'(-697);
			40025: out = 16'(-48);
			40026: out = 16'(-66);
			40027: out = 16'(-209);
			40028: out = 16'(-1119);
			40029: out = 16'(-1335);
			40030: out = 16'(-1295);
			40031: out = 16'(121);
			40032: out = 16'(543);
			40033: out = 16'(966);
			40034: out = 16'(212);
			40035: out = 16'(293);
			40036: out = 16'(258);
			40037: out = 16'(1334);
			40038: out = 16'(922);
			40039: out = 16'(-133);
			40040: out = 16'(75);
			40041: out = 16'(419);
			40042: out = 16'(1104);
			40043: out = 16'(1118);
			40044: out = 16'(841);
			40045: out = 16'(131);
			40046: out = 16'(-942);
			40047: out = 16'(-1692);
			40048: out = 16'(-1494);
			40049: out = 16'(-1041);
			40050: out = 16'(-317);
			40051: out = 16'(-277);
			40052: out = 16'(-78);
			40053: out = 16'(-184);
			40054: out = 16'(288);
			40055: out = 16'(115);
			40056: out = 16'(-9);
			40057: out = 16'(89);
			40058: out = 16'(266);
			40059: out = 16'(217);
			40060: out = 16'(543);
			40061: out = 16'(363);
			40062: out = 16'(-145);
			40063: out = 16'(-814);
			40064: out = 16'(-1179);
			40065: out = 16'(-1119);
			40066: out = 16'(-362);
			40067: out = 16'(306);
			40068: out = 16'(-71);
			40069: out = 16'(50);
			40070: out = 16'(-29);
			40071: out = 16'(234);
			40072: out = 16'(152);
			40073: out = 16'(241);
			40074: out = 16'(-37);
			40075: out = 16'(210);
			40076: out = 16'(588);
			40077: out = 16'(367);
			40078: out = 16'(136);
			40079: out = 16'(-43);
			40080: out = 16'(-78);
			40081: out = 16'(47);
			40082: out = 16'(216);
			40083: out = 16'(468);
			40084: out = 16'(443);
			40085: out = 16'(-23);
			40086: out = 16'(-312);
			40087: out = 16'(-496);
			40088: out = 16'(-512);
			40089: out = 16'(-178);
			40090: out = 16'(177);
			40091: out = 16'(-127);
			40092: out = 16'(-44);
			40093: out = 16'(228);
			40094: out = 16'(161);
			40095: out = 16'(500);
			40096: out = 16'(798);
			40097: out = 16'(1110);
			40098: out = 16'(743);
			40099: out = 16'(-85);
			40100: out = 16'(-668);
			40101: out = 16'(-716);
			40102: out = 16'(-153);
			40103: out = 16'(470);
			40104: out = 16'(702);
			40105: out = 16'(-93);
			40106: out = 16'(-1087);
			40107: out = 16'(-1915);
			40108: out = 16'(-1234);
			40109: out = 16'(-502);
			40110: out = 16'(410);
			40111: out = 16'(769);
			40112: out = 16'(568);
			40113: out = 16'(-249);
			40114: out = 16'(191);
			40115: out = 16'(630);
			40116: out = 16'(1769);
			40117: out = 16'(822);
			40118: out = 16'(165);
			40119: out = 16'(-913);
			40120: out = 16'(-259);
			40121: out = 16'(246);
			40122: out = 16'(454);
			40123: out = 16'(334);
			40124: out = 16'(-115);
			40125: out = 16'(-737);
			40126: out = 16'(-1109);
			40127: out = 16'(-1043);
			40128: out = 16'(-427);
			40129: out = 16'(351);
			40130: out = 16'(807);
			40131: out = 16'(900);
			40132: out = 16'(406);
			40133: out = 16'(-211);
			40134: out = 16'(-995);
			40135: out = 16'(-1021);
			40136: out = 16'(-515);
			40137: out = 16'(616);
			40138: out = 16'(1193);
			40139: out = 16'(1092);
			40140: out = 16'(132);
			40141: out = 16'(-792);
			40142: out = 16'(-1131);
			40143: out = 16'(-891);
			40144: out = 16'(-417);
			40145: out = 16'(-154);
			40146: out = 16'(-58);
			40147: out = 16'(-126);
			40148: out = 16'(-1004);
			40149: out = 16'(-1045);
			40150: out = 16'(-724);
			40151: out = 16'(565);
			40152: out = 16'(778);
			40153: out = 16'(200);
			40154: out = 16'(-224);
			40155: out = 16'(-430);
			40156: out = 16'(-6);
			40157: out = 16'(302);
			40158: out = 16'(649);
			40159: out = 16'(506);
			40160: out = 16'(405);
			40161: out = 16'(120);
			40162: out = 16'(-20);
			40163: out = 16'(-152);
			40164: out = 16'(-260);
			40165: out = 16'(-1026);
			40166: out = 16'(-1455);
			40167: out = 16'(-1800);
			40168: out = 16'(-957);
			40169: out = 16'(-242);
			40170: out = 16'(743);
			40171: out = 16'(992);
			40172: out = 16'(1236);
			40173: out = 16'(742);
			40174: out = 16'(1205);
			40175: out = 16'(682);
			40176: out = 16'(-374);
			40177: out = 16'(-1658);
			40178: out = 16'(-2086);
			40179: out = 16'(-1177);
			40180: out = 16'(26);
			40181: out = 16'(1016);
			40182: out = 16'(217);
			40183: out = 16'(-338);
			40184: out = 16'(-1210);
			40185: out = 16'(-382);
			40186: out = 16'(-474);
			40187: out = 16'(-314);
			40188: out = 16'(-746);
			40189: out = 16'(-446);
			40190: out = 16'(-48);
			40191: out = 16'(527);
			40192: out = 16'(716);
			40193: out = 16'(996);
			40194: out = 16'(279);
			40195: out = 16'(-13);
			40196: out = 16'(-35);
			40197: out = 16'(708);
			40198: out = 16'(1341);
			40199: out = 16'(1680);
			40200: out = 16'(1293);
			40201: out = 16'(633);
			40202: out = 16'(-72);
			40203: out = 16'(-137);
			40204: out = 16'(209);
			40205: out = 16'(653);
			40206: out = 16'(747);
			40207: out = 16'(377);
			40208: out = 16'(-7);
			40209: out = 16'(-438);
			40210: out = 16'(-493);
			40211: out = 16'(-414);
			40212: out = 16'(-86);
			40213: out = 16'(-233);
			40214: out = 16'(1069);
			40215: out = 16'(1645);
			40216: out = 16'(1315);
			40217: out = 16'(622);
			40218: out = 16'(-287);
			40219: out = 16'(-1111);
			40220: out = 16'(-1501);
			40221: out = 16'(-1528);
			40222: out = 16'(-986);
			40223: out = 16'(-697);
			40224: out = 16'(-538);
			40225: out = 16'(-1038);
			40226: out = 16'(-1291);
			40227: out = 16'(-1457);
			40228: out = 16'(-243);
			40229: out = 16'(619);
			40230: out = 16'(1483);
			40231: out = 16'(649);
			40232: out = 16'(82);
			40233: out = 16'(-132);
			40234: out = 16'(-3);
			40235: out = 16'(153);
			40236: out = 16'(-90);
			40237: out = 16'(105);
			40238: out = 16'(224);
			40239: out = 16'(-63);
			40240: out = 16'(-118);
			40241: out = 16'(-162);
			40242: out = 16'(472);
			40243: out = 16'(618);
			40244: out = 16'(832);
			40245: out = 16'(-588);
			40246: out = 16'(-713);
			40247: out = 16'(-147);
			40248: out = 16'(128);
			40249: out = 16'(131);
			40250: out = 16'(-212);
			40251: out = 16'(-599);
			40252: out = 16'(-986);
			40253: out = 16'(-1486);
			40254: out = 16'(-902);
			40255: out = 16'(-171);
			40256: out = 16'(1117);
			40257: out = 16'(597);
			40258: out = 16'(-214);
			40259: out = 16'(-613);
			40260: out = 16'(-480);
			40261: out = 16'(79);
			40262: out = 16'(-117);
			40263: out = 16'(122);
			40264: out = 16'(127);
			40265: out = 16'(-19);
			40266: out = 16'(-263);
			40267: out = 16'(-359);
			40268: out = 16'(-196);
			40269: out = 16'(346);
			40270: out = 16'(1307);
			40271: out = 16'(1329);
			40272: out = 16'(1210);
			40273: out = 16'(1028);
			40274: out = 16'(674);
			40275: out = 16'(342);
			40276: out = 16'(117);
			40277: out = 16'(-250);
			40278: out = 16'(-549);
			40279: out = 16'(26);
			40280: out = 16'(-18);
			40281: out = 16'(-126);
			40282: out = 16'(-236);
			40283: out = 16'(-115);
			40284: out = 16'(69);
			40285: out = 16'(378);
			40286: out = 16'(335);
			40287: out = 16'(54);
			40288: out = 16'(-171);
			40289: out = 16'(-207);
			40290: out = 16'(-159);
			40291: out = 16'(78);
			40292: out = 16'(-51);
			40293: out = 16'(-1021);
			40294: out = 16'(-1656);
			40295: out = 16'(-2003);
			40296: out = 16'(-1137);
			40297: out = 16'(-626);
			40298: out = 16'(-46);
			40299: out = 16'(-404);
			40300: out = 16'(-265);
			40301: out = 16'(-76);
			40302: out = 16'(-28);
			40303: out = 16'(82);
			40304: out = 16'(198);
			40305: out = 16'(264);
			40306: out = 16'(318);
			40307: out = 16'(576);
			40308: out = 16'(271);
			40309: out = 16'(548);
			40310: out = 16'(1768);
			40311: out = 16'(1799);
			40312: out = 16'(1581);
			40313: out = 16'(1044);
			40314: out = 16'(327);
			40315: out = 16'(-231);
			40316: out = 16'(10);
			40317: out = 16'(0);
			40318: out = 16'(2);
			40319: out = 16'(367);
			40320: out = 16'(258);
			40321: out = 16'(83);
			40322: out = 16'(-900);
			40323: out = 16'(-1126);
			40324: out = 16'(-823);
			40325: out = 16'(-200);
			40326: out = 16'(-58);
			40327: out = 16'(-862);
			40328: out = 16'(-591);
			40329: out = 16'(-378);
			40330: out = 16'(70);
			40331: out = 16'(19);
			40332: out = 16'(-105);
			40333: out = 16'(529);
			40334: out = 16'(-159);
			40335: out = 16'(-913);
			40336: out = 16'(-1917);
			40337: out = 16'(-1554);
			40338: out = 16'(-548);
			40339: out = 16'(501);
			40340: out = 16'(749);
			40341: out = 16'(144);
			40342: out = 16'(66);
			40343: out = 16'(-295);
			40344: out = 16'(-358);
			40345: out = 16'(-118);
			40346: out = 16'(442);
			40347: out = 16'(971);
			40348: out = 16'(968);
			40349: out = 16'(500);
			40350: out = 16'(-314);
			40351: out = 16'(-875);
			40352: out = 16'(-921);
			40353: out = 16'(-224);
			40354: out = 16'(388);
			40355: out = 16'(742);
			40356: out = 16'(620);
			40357: out = 16'(-131);
			40358: out = 16'(-1113);
			40359: out = 16'(-1585);
			40360: out = 16'(-1193);
			40361: out = 16'(312);
			40362: out = 16'(-24);
			40363: out = 16'(69);
			40364: out = 16'(182);
			40365: out = 16'(171);
			40366: out = 16'(161);
			40367: out = 16'(177);
			40368: out = 16'(79);
			40369: out = 16'(-16);
			40370: out = 16'(543);
			40371: out = 16'(215);
			40372: out = 16'(-60);
			40373: out = 16'(-424);
			40374: out = 16'(-126);
			40375: out = 16'(281);
			40376: out = 16'(1157);
			40377: out = 16'(1124);
			40378: out = 16'(728);
			40379: out = 16'(55);
			40380: out = 16'(96);
			40381: out = 16'(722);
			40382: out = 16'(1269);
			40383: out = 16'(1206);
			40384: out = 16'(134);
			40385: out = 16'(-644);
			40386: out = 16'(-1172);
			40387: out = 16'(-541);
			40388: out = 16'(-176);
			40389: out = 16'(225);
			40390: out = 16'(407);
			40391: out = 16'(-100);
			40392: out = 16'(-946);
			40393: out = 16'(-784);
			40394: out = 16'(-476);
			40395: out = 16'(278);
			40396: out = 16'(-137);
			40397: out = 16'(-64);
			40398: out = 16'(-263);
			40399: out = 16'(68);
			40400: out = 16'(0);
			40401: out = 16'(-166);
			40402: out = 16'(-412);
			40403: out = 16'(-488);
			40404: out = 16'(-505);
			40405: out = 16'(-83);
			40406: out = 16'(226);
			40407: out = 16'(188);
			40408: out = 16'(-114);
			40409: out = 16'(-518);
			40410: out = 16'(85);
			40411: out = 16'(107);
			40412: out = 16'(172);
			40413: out = 16'(-1450);
			40414: out = 16'(-1644);
			40415: out = 16'(-1275);
			40416: out = 16'(254);
			40417: out = 16'(1109);
			40418: out = 16'(1245);
			40419: out = 16'(1364);
			40420: out = 16'(941);
			40421: out = 16'(-119);
			40422: out = 16'(-158);
			40423: out = 16'(-218);
			40424: out = 16'(-83);
			40425: out = 16'(-148);
			40426: out = 16'(-135);
			40427: out = 16'(-824);
			40428: out = 16'(-335);
			40429: out = 16'(139);
			40430: out = 16'(233);
			40431: out = 16'(-205);
			40432: out = 16'(-854);
			40433: out = 16'(-1270);
			40434: out = 16'(-1128);
			40435: out = 16'(-321);
			40436: out = 16'(23);
			40437: out = 16'(416);
			40438: out = 16'(474);
			40439: out = 16'(568);
			40440: out = 16'(462);
			40441: out = 16'(533);
			40442: out = 16'(311);
			40443: out = 16'(106);
			40444: out = 16'(-449);
			40445: out = 16'(-471);
			40446: out = 16'(-421);
			40447: out = 16'(-91);
			40448: out = 16'(23);
			40449: out = 16'(162);
			40450: out = 16'(83);
			40451: out = 16'(393);
			40452: out = 16'(759);
			40453: out = 16'(94);
			40454: out = 16'(-413);
			40455: out = 16'(-1107);
			40456: out = 16'(-431);
			40457: out = 16'(12);
			40458: out = 16'(185);
			40459: out = 16'(218);
			40460: out = 16'(-130);
			40461: out = 16'(-990);
			40462: out = 16'(-1268);
			40463: out = 16'(-1195);
			40464: out = 16'(-195);
			40465: out = 16'(125);
			40466: out = 16'(271);
			40467: out = 16'(-57);
			40468: out = 16'(-222);
			40469: out = 16'(-397);
			40470: out = 16'(106);
			40471: out = 16'(162);
			40472: out = 16'(-34);
			40473: out = 16'(25);
			40474: out = 16'(-55);
			40475: out = 16'(-57);
			40476: out = 16'(-100);
			40477: out = 16'(272);
			40478: out = 16'(1057);
			40479: out = 16'(1255);
			40480: out = 16'(1289);
			40481: out = 16'(1314);
			40482: out = 16'(667);
			40483: out = 16'(-22);
			40484: out = 16'(-699);
			40485: out = 16'(-703);
			40486: out = 16'(-398);
			40487: out = 16'(77);
			40488: out = 16'(214);
			40489: out = 16'(46);
			40490: out = 16'(-102);
			40491: out = 16'(-203);
			40492: out = 16'(-45);
			40493: out = 16'(-205);
			40494: out = 16'(-79);
			40495: out = 16'(76);
			40496: out = 16'(209);
			40497: out = 16'(145);
			40498: out = 16'(149);
			40499: out = 16'(-277);
			40500: out = 16'(-555);
			40501: out = 16'(-781);
			40502: out = 16'(-585);
			40503: out = 16'(-486);
			40504: out = 16'(-669);
			40505: out = 16'(-1020);
			40506: out = 16'(-1265);
			40507: out = 16'(-309);
			40508: out = 16'(431);
			40509: out = 16'(1140);
			40510: out = 16'(1103);
			40511: out = 16'(750);
			40512: out = 16'(-100);
			40513: out = 16'(130);
			40514: out = 16'(212);
			40515: out = 16'(536);
			40516: out = 16'(481);
			40517: out = 16'(447);
			40518: out = 16'(116);
			40519: out = 16'(111);
			40520: out = 16'(129);
			40521: out = 16'(465);
			40522: out = 16'(332);
			40523: out = 16'(136);
			40524: out = 16'(207);
			40525: out = 16'(100);
			40526: out = 16'(48);
			40527: out = 16'(-920);
			40528: out = 16'(-1113);
			40529: out = 16'(-1067);
			40530: out = 16'(-384);
			40531: out = 16'(-98);
			40532: out = 16'(-154);
			40533: out = 16'(-98);
			40534: out = 16'(123);
			40535: out = 16'(786);
			40536: out = 16'(445);
			40537: out = 16'(159);
			40538: out = 16'(541);
			40539: out = 16'(115);
			40540: out = 16'(-116);
			40541: out = 16'(-515);
			40542: out = 16'(-113);
			40543: out = 16'(180);
			40544: out = 16'(280);
			40545: out = 16'(-461);
			40546: out = 16'(-1422);
			40547: out = 16'(-1445);
			40548: out = 16'(-637);
			40549: out = 16'(898);
			40550: out = 16'(1511);
			40551: out = 16'(1740);
			40552: out = 16'(1210);
			40553: out = 16'(378);
			40554: out = 16'(-226);
			40555: out = 16'(127);
			40556: out = 16'(365);
			40557: out = 16'(761);
			40558: out = 16'(345);
			40559: out = 16'(189);
			40560: out = 16'(-338);
			40561: out = 16'(-363);
			40562: out = 16'(-1032);
			40563: out = 16'(-1410);
			40564: out = 16'(-1541);
			40565: out = 16'(-814);
			40566: out = 16'(177);
			40567: out = 16'(207);
			40568: out = 16'(87);
			40569: out = 16'(-160);
			40570: out = 16'(-1224);
			40571: out = 16'(-1865);
			40572: out = 16'(-1944);
			40573: out = 16'(-1219);
			40574: out = 16'(-412);
			40575: out = 16'(-161);
			40576: out = 16'(87);
			40577: out = 16'(129);
			40578: out = 16'(1391);
			40579: out = 16'(975);
			40580: out = 16'(434);
			40581: out = 16'(-517);
			40582: out = 16'(-726);
			40583: out = 16'(-648);
			40584: out = 16'(-198);
			40585: out = 16'(-2);
			40586: out = 16'(23);
			40587: out = 16'(238);
			40588: out = 16'(254);
			40589: out = 16'(-37);
			40590: out = 16'(751);
			40591: out = 16'(1228);
			40592: out = 16'(1575);
			40593: out = 16'(780);
			40594: out = 16'(59);
			40595: out = 16'(191);
			40596: out = 16'(223);
			40597: out = 16'(535);
			40598: out = 16'(48);
			40599: out = 16'(152);
			40600: out = 16'(10);
			40601: out = 16'(544);
			40602: out = 16'(-285);
			40603: out = 16'(-1500);
			40604: out = 16'(-1674);
			40605: out = 16'(-1280);
			40606: out = 16'(-20);
			40607: out = 16'(-126);
			40608: out = 16'(10);
			40609: out = 16'(-175);
			40610: out = 16'(103);
			40611: out = 16'(180);
			40612: out = 16'(260);
			40613: out = 16'(189);
			40614: out = 16'(101);
			40615: out = 16'(-433);
			40616: out = 16'(-235);
			40617: out = 16'(97);
			40618: out = 16'(1391);
			40619: out = 16'(1580);
			40620: out = 16'(1436);
			40621: out = 16'(149);
			40622: out = 16'(-140);
			40623: out = 16'(135);
			40624: out = 16'(88);
			40625: out = 16'(324);
			40626: out = 16'(687);
			40627: out = 16'(321);
			40628: out = 16'(-1);
			40629: out = 16'(-213);
			40630: out = 16'(-275);
			40631: out = 16'(-354);
			40632: out = 16'(-1138);
			40633: out = 16'(-664);
			40634: out = 16'(48);
			40635: out = 16'(1317);
			40636: out = 16'(1547);
			40637: out = 16'(1247);
			40638: out = 16'(-206);
			40639: out = 16'(-1165);
			40640: out = 16'(-1806);
			40641: out = 16'(-1558);
			40642: out = 16'(-1114);
			40643: out = 16'(-437);
			40644: out = 16'(-68);
			40645: out = 16'(114);
			40646: out = 16'(-233);
			40647: out = 16'(122);
			40648: out = 16'(325);
			40649: out = 16'(1030);
			40650: out = 16'(652);
			40651: out = 16'(369);
			40652: out = 16'(-130);
			40653: out = 16'(-104);
			40654: out = 16'(-179);
			40655: out = 16'(166);
			40656: out = 16'(-504);
			40657: out = 16'(-1123);
			40658: out = 16'(-1184);
			40659: out = 16'(-286);
			40660: out = 16'(1121);
			40661: out = 16'(1001);
			40662: out = 16'(664);
			40663: out = 16'(-279);
			40664: out = 16'(-812);
			40665: out = 16'(-1130);
			40666: out = 16'(-713);
			40667: out = 16'(-638);
			40668: out = 16'(-281);
			40669: out = 16'(78);
			40670: out = 16'(174);
			40671: out = 16'(77);
			40672: out = 16'(-134);
			40673: out = 16'(14);
			40674: out = 16'(290);
			40675: out = 16'(417);
			40676: out = 16'(412);
			40677: out = 16'(116);
			40678: out = 16'(199);
			40679: out = 16'(-236);
			40680: out = 16'(-819);
			40681: out = 16'(-786);
			40682: out = 16'(-534);
			40683: out = 16'(179);
			40684: out = 16'(-93);
			40685: out = 16'(-141);
			40686: out = 16'(-174);
			40687: out = 16'(266);
			40688: out = 16'(543);
			40689: out = 16'(483);
			40690: out = 16'(195);
			40691: out = 16'(-156);
			40692: out = 16'(-30);
			40693: out = 16'(-155);
			40694: out = 16'(-137);
			40695: out = 16'(-146);
			40696: out = 16'(265);
			40697: out = 16'(771);
			40698: out = 16'(252);
			40699: out = 16'(-200);
			40700: out = 16'(-835);
			40701: out = 16'(-327);
			40702: out = 16'(-104);
			40703: out = 16'(-95);
			40704: out = 16'(-74);
			40705: out = 16'(-2);
			40706: out = 16'(510);
			40707: out = 16'(302);
			40708: out = 16'(157);
			40709: out = 16'(-127);
			40710: out = 16'(339);
			40711: out = 16'(743);
			40712: out = 16'(134);
			40713: out = 16'(-158);
			40714: out = 16'(-505);
			40715: out = 16'(555);
			40716: out = 16'(658);
			40717: out = 16'(363);
			40718: out = 16'(194);
			40719: out = 16'(-31);
			40720: out = 16'(105);
			40721: out = 16'(-627);
			40722: out = 16'(-777);
			40723: out = 16'(-537);
			40724: out = 16'(-114);
			40725: out = 16'(-29);
			40726: out = 16'(-776);
			40727: out = 16'(-827);
			40728: out = 16'(-662);
			40729: out = 16'(-174);
			40730: out = 16'(475);
			40731: out = 16'(1058);
			40732: out = 16'(768);
			40733: out = 16'(491);
			40734: out = 16'(13);
			40735: out = 16'(102);
			40736: out = 16'(-47);
			40737: out = 16'(-238);
			40738: out = 16'(-402);
			40739: out = 16'(-708);
			40740: out = 16'(-1052);
			40741: out = 16'(-1356);
			40742: out = 16'(-1173);
			40743: out = 16'(-465);
			40744: out = 16'(322);
			40745: out = 16'(939);
			40746: out = 16'(982);
			40747: out = 16'(927);
			40748: out = 16'(721);
			40749: out = 16'(993);
			40750: out = 16'(945);
			40751: out = 16'(908);
			40752: out = 16'(246);
			40753: out = 16'(-141);
			40754: out = 16'(-589);
			40755: out = 16'(-85);
			40756: out = 16'(157);
			40757: out = 16'(429);
			40758: out = 16'(113);
			40759: out = 16'(35);
			40760: out = 16'(99);
			40761: out = 16'(118);
			40762: out = 16'(-17);
			40763: out = 16'(-558);
			40764: out = 16'(-574);
			40765: out = 16'(-522);
			40766: out = 16'(-270);
			40767: out = 16'(-363);
			40768: out = 16'(-537);
			40769: out = 16'(-196);
			40770: out = 16'(-361);
			40771: out = 16'(-486);
			40772: out = 16'(-789);
			40773: out = 16'(-511);
			40774: out = 16'(-29);
			40775: out = 16'(755);
			40776: out = 16'(942);
			40777: out = 16'(368);
			40778: out = 16'(282);
			40779: out = 16'(-132);
			40780: out = 16'(-444);
			40781: out = 16'(-570);
			40782: out = 16'(-328);
			40783: out = 16'(112);
			40784: out = 16'(498);
			40785: out = 16'(790);
			40786: out = 16'(1190);
			40787: out = 16'(1200);
			40788: out = 16'(1098);
			40789: out = 16'(-49);
			40790: out = 16'(-144);
			40791: out = 16'(23);
			40792: out = 16'(302);
			40793: out = 16'(265);
			40794: out = 16'(-46);
			40795: out = 16'(-853);
			40796: out = 16'(-1284);
			40797: out = 16'(-1100);
			40798: out = 16'(-1204);
			40799: out = 16'(-969);
			40800: out = 16'(-528);
			40801: out = 16'(-303);
			40802: out = 16'(-202);
			40803: out = 16'(-467);
			40804: out = 16'(-444);
			40805: out = 16'(-482);
			40806: out = 16'(-404);
			40807: out = 16'(-712);
			40808: out = 16'(-1047);
			40809: out = 16'(-776);
			40810: out = 16'(-375);
			40811: out = 16'(245);
			40812: out = 16'(-281);
			40813: out = 16'(-489);
			40814: out = 16'(-679);
			40815: out = 16'(10);
			40816: out = 16'(438);
			40817: out = 16'(509);
			40818: out = 16'(768);
			40819: out = 16'(864);
			40820: out = 16'(1358);
			40821: out = 16'(833);
			40822: out = 16'(347);
			40823: out = 16'(-399);
			40824: out = 16'(-231);
			40825: out = 16'(165);
			40826: out = 16'(87);
			40827: out = 16'(122);
			40828: out = 16'(92);
			40829: out = 16'(-45);
			40830: out = 16'(-124);
			40831: out = 16'(-170);
			40832: out = 16'(106);
			40833: out = 16'(259);
			40834: out = 16'(485);
			40835: out = 16'(-165);
			40836: out = 16'(-652);
			40837: out = 16'(-1077);
			40838: out = 16'(-707);
			40839: out = 16'(-443);
			40840: out = 16'(-732);
			40841: out = 16'(-731);
			40842: out = 16'(-623);
			40843: out = 16'(-214);
			40844: out = 16'(430);
			40845: out = 16'(1204);
			40846: out = 16'(1671);
			40847: out = 16'(1759);
			40848: out = 16'(1374);
			40849: out = 16'(303);
			40850: out = 16'(-425);
			40851: out = 16'(-392);
			40852: out = 16'(-888);
			40853: out = 16'(-553);
			40854: out = 16'(-209);
			40855: out = 16'(973);
			40856: out = 16'(1441);
			40857: out = 16'(980);
			40858: out = 16'(400);
			40859: out = 16'(35);
			40860: out = 16'(588);
			40861: out = 16'(1021);
			40862: out = 16'(1337);
			40863: out = 16'(115);
			40864: out = 16'(-453);
			40865: out = 16'(-986);
			40866: out = 16'(-667);
			40867: out = 16'(-603);
			40868: out = 16'(-584);
			40869: out = 16'(355);
			40870: out = 16'(698);
			40871: out = 16'(578);
			40872: out = 16'(14);
			40873: out = 16'(-377);
			40874: out = 16'(38);
			40875: out = 16'(-249);
			40876: out = 16'(-418);
			40877: out = 16'(-1239);
			40878: out = 16'(-827);
			40879: out = 16'(-665);
			40880: out = 16'(-1681);
			40881: out = 16'(-2078);
			40882: out = 16'(-2273);
			40883: out = 16'(-448);
			40884: out = 16'(82);
			40885: out = 16'(254);
			40886: out = 16'(-61);
			40887: out = 16'(-123);
			40888: out = 16'(-38);
			40889: out = 16'(-42);
			40890: out = 16'(13);
			40891: out = 16'(257);
			40892: out = 16'(215);
			40893: out = 16'(144);
			40894: out = 16'(-504);
			40895: out = 16'(157);
			40896: out = 16'(670);
			40897: out = 16'(1540);
			40898: out = 16'(805);
			40899: out = 16'(-117);
			40900: out = 16'(-675);
			40901: out = 16'(-722);
			40902: out = 16'(-402);
			40903: out = 16'(-17);
			40904: out = 16'(151);
			40905: out = 16'(57);
			40906: out = 16'(-559);
			40907: out = 16'(-847);
			40908: out = 16'(-712);
			40909: out = 16'(-358);
			40910: out = 16'(-63);
			40911: out = 16'(-196);
			40912: out = 16'(97);
			40913: out = 16'(150);
			40914: out = 16'(257);
			40915: out = 16'(210);
			40916: out = 16'(229);
			40917: out = 16'(-100);
			40918: out = 16'(235);
			40919: out = 16'(515);
			40920: out = 16'(499);
			40921: out = 16'(321);
			40922: out = 16'(58);
			40923: out = 16'(-625);
			40924: out = 16'(-829);
			40925: out = 16'(-728);
			40926: out = 16'(-96);
			40927: out = 16'(302);
			40928: out = 16'(497);
			40929: out = 16'(654);
			40930: out = 16'(900);
			40931: out = 16'(1210);
			40932: out = 16'(1298);
			40933: out = 16'(934);
			40934: out = 16'(-132);
			40935: out = 16'(-964);
			40936: out = 16'(-1497);
			40937: out = 16'(-1156);
			40938: out = 16'(-710);
			40939: out = 16'(-84);
			40940: out = 16'(21);
			40941: out = 16'(75);
			40942: out = 16'(-136);
			40943: out = 16'(187);
			40944: out = 16'(150);
			40945: out = 16'(108);
			40946: out = 16'(-359);
			40947: out = 16'(-427);
			40948: out = 16'(-167);
			40949: out = 16'(-188);
			40950: out = 16'(-204);
			40951: out = 16'(-492);
			40952: out = 16'(-272);
			40953: out = 16'(-110);
			40954: out = 16'(-37);
			40955: out = 16'(59);
			40956: out = 16'(289);
			40957: out = 16'(170);
			40958: out = 16'(410);
			40959: out = 16'(479);
			40960: out = 16'(1238);
			40961: out = 16'(836);
			40962: out = 16'(122);
			40963: out = 16'(-612);
			40964: out = 16'(-593);
			40965: out = 16'(156);
			40966: out = 16'(164);
			40967: out = 16'(-24);
			40968: out = 16'(-818);
			40969: out = 16'(-593);
			40970: out = 16'(-322);
			40971: out = 16'(162);
			40972: out = 16'(382);
			40973: out = 16'(399);
			40974: out = 16'(-34);
			40975: out = 16'(-297);
			40976: out = 16'(-524);
			40977: out = 16'(-1336);
			40978: out = 16'(-1003);
			40979: out = 16'(-338);
			40980: out = 16'(365);
			40981: out = 16'(459);
			40982: out = 16'(104);
			40983: out = 16'(-532);
			40984: out = 16'(-563);
			40985: out = 16'(222);
			40986: out = 16'(377);
			40987: out = 16'(562);
			40988: out = 16'(490);
			40989: out = 16'(-31);
			40990: out = 16'(-676);
			40991: out = 16'(-1270);
			40992: out = 16'(-1084);
			40993: out = 16'(-433);
			40994: out = 16'(596);
			40995: out = 16'(1043);
			40996: out = 16'(992);
			40997: out = 16'(1127);
			40998: out = 16'(559);
			40999: out = 16'(-130);
			41000: out = 16'(-142);
			41001: out = 16'(-181);
			41002: out = 16'(-189);
			41003: out = 16'(-178);
			41004: out = 16'(-155);
			41005: out = 16'(-48);
			41006: out = 16'(30);
			41007: out = 16'(163);
			41008: out = 16'(41);
			41009: out = 16'(547);
			41010: out = 16'(666);
			41011: out = 16'(181);
			41012: out = 16'(-533);
			41013: out = 16'(-1115);
			41014: out = 16'(-524);
			41015: out = 16'(-279);
			41016: out = 16'(-36);
			41017: out = 16'(398);
			41018: out = 16'(494);
			41019: out = 16'(482);
			41020: out = 16'(0);
			41021: out = 16'(-18);
			41022: out = 16'(169);
			41023: out = 16'(784);
			41024: out = 16'(775);
			41025: out = 16'(-139);
			41026: out = 16'(-351);
			41027: out = 16'(-437);
			41028: out = 16'(150);
			41029: out = 16'(307);
			41030: out = 16'(416);
			41031: out = 16'(111);
			41032: out = 16'(-213);
			41033: out = 16'(-533);
			41034: out = 16'(-278);
			41035: out = 16'(158);
			41036: out = 16'(746);
			41037: out = 16'(250);
			41038: out = 16'(-250);
			41039: out = 16'(-1210);
			41040: out = 16'(-431);
			41041: out = 16'(-172);
			41042: out = 16'(-116);
			41043: out = 16'(-342);
			41044: out = 16'(-648);
			41045: out = 16'(-1075);
			41046: out = 16'(-895);
			41047: out = 16'(-682);
			41048: out = 16'(-992);
			41049: out = 16'(-757);
			41050: out = 16'(-607);
			41051: out = 16'(160);
			41052: out = 16'(-84);
			41053: out = 16'(-346);
			41054: out = 16'(-405);
			41055: out = 16'(94);
			41056: out = 16'(810);
			41057: out = 16'(1154);
			41058: out = 16'(946);
			41059: out = 16'(167);
			41060: out = 16'(-192);
			41061: out = 16'(-417);
			41062: out = 16'(-94);
			41063: out = 16'(68);
			41064: out = 16'(295);
			41065: out = 16'(431);
			41066: out = 16'(319);
			41067: out = 16'(203);
			41068: out = 16'(409);
			41069: out = 16'(779);
			41070: out = 16'(1198);
			41071: out = 16'(1107);
			41072: out = 16'(752);
			41073: out = 16'(-38);
			41074: out = 16'(-55);
			41075: out = 16'(-705);
			41076: out = 16'(-1313);
			41077: out = 16'(-1176);
			41078: out = 16'(-571);
			41079: out = 16'(420);
			41080: out = 16'(612);
			41081: out = 16'(532);
			41082: out = 16'(88);
			41083: out = 16'(-588);
			41084: out = 16'(-1119);
			41085: out = 16'(-927);
			41086: out = 16'(-1041);
			41087: out = 16'(-891);
			41088: out = 16'(-757);
			41089: out = 16'(-253);
			41090: out = 16'(260);
			41091: out = 16'(821);
			41092: out = 16'(1184);
			41093: out = 16'(1377);
			41094: out = 16'(638);
			41095: out = 16'(109);
			41096: out = 16'(-481);
			41097: out = 16'(169);
			41098: out = 16'(616);
			41099: out = 16'(1137);
			41100: out = 16'(278);
			41101: out = 16'(-551);
			41102: out = 16'(-1239);
			41103: out = 16'(-1377);
			41104: out = 16'(-1159);
			41105: out = 16'(-792);
			41106: out = 16'(-355);
			41107: out = 16'(-97);
			41108: out = 16'(117);
			41109: out = 16'(57);
			41110: out = 16'(-46);
			41111: out = 16'(-61);
			41112: out = 16'(-27);
			41113: out = 16'(-63);
			41114: out = 16'(381);
			41115: out = 16'(391);
			41116: out = 16'(188);
			41117: out = 16'(-415);
			41118: out = 16'(-758);
			41119: out = 16'(-635);
			41120: out = 16'(-510);
			41121: out = 16'(-471);
			41122: out = 16'(-1229);
			41123: out = 16'(-886);
			41124: out = 16'(-441);
			41125: out = 16'(438);
			41126: out = 16'(664);
			41127: out = 16'(799);
			41128: out = 16'(733);
			41129: out = 16'(757);
			41130: out = 16'(688);
			41131: out = 16'(754);
			41132: out = 16'(498);
			41133: out = 16'(185);
			41134: out = 16'(-102);
			41135: out = 16'(-79);
			41136: out = 16'(186);
			41137: out = 16'(350);
			41138: out = 16'(366);
			41139: out = 16'(86);
			41140: out = 16'(71);
			41141: out = 16'(62);
			41142: out = 16'(-120);
			41143: out = 16'(14);
			41144: out = 16'(61);
			41145: out = 16'(95);
			41146: out = 16'(-174);
			41147: out = 16'(-493);
			41148: out = 16'(-718);
			41149: out = 16'(-491);
			41150: out = 16'(-10);
			41151: out = 16'(508);
			41152: out = 16'(523);
			41153: out = 16'(-194);
			41154: out = 16'(-24);
			41155: out = 16'(-178);
			41156: out = 16'(-26);
			41157: out = 16'(-532);
			41158: out = 16'(-838);
			41159: out = 16'(-1595);
			41160: out = 16'(-1171);
			41161: out = 16'(-905);
			41162: out = 16'(-576);
			41163: out = 16'(-1074);
			41164: out = 16'(-1412);
			41165: out = 16'(-992);
			41166: out = 16'(-97);
			41167: out = 16'(973);
			41168: out = 16'(1171);
			41169: out = 16'(1329);
			41170: out = 16'(1211);
			41171: out = 16'(510);
			41172: out = 16'(11);
			41173: out = 16'(-370);
			41174: out = 16'(49);
			41175: out = 16'(325);
			41176: out = 16'(499);
			41177: out = 16'(-69);
			41178: out = 16'(-390);
			41179: out = 16'(-26);
			41180: out = 16'(361);
			41181: out = 16'(729);
			41182: out = 16'(-56);
			41183: out = 16'(-39);
			41184: out = 16'(-180);
			41185: out = 16'(142);
			41186: out = 16'(26);
			41187: out = 16'(-19);
			41188: out = 16'(-109);
			41189: out = 16'(138);
			41190: out = 16'(429);
			41191: out = 16'(492);
			41192: out = 16'(256);
			41193: out = 16'(-119);
			41194: out = 16'(-765);
			41195: out = 16'(-792);
			41196: out = 16'(213);
			41197: out = 16'(356);
			41198: out = 16'(321);
			41199: out = 16'(-647);
			41200: out = 16'(-824);
			41201: out = 16'(-953);
			41202: out = 16'(-676);
			41203: out = 16'(-528);
			41204: out = 16'(-292);
			41205: out = 16'(145);
			41206: out = 16'(386);
			41207: out = 16'(482);
			41208: out = 16'(96);
			41209: out = 16'(-58);
			41210: out = 16'(-7);
			41211: out = 16'(104);
			41212: out = 16'(118);
			41213: out = 16'(-168);
			41214: out = 16'(82);
			41215: out = 16'(122);
			41216: out = 16'(-5);
			41217: out = 16'(-63);
			41218: out = 16'(-137);
			41219: out = 16'(-368);
			41220: out = 16'(-116);
			41221: out = 16'(226);
			41222: out = 16'(128);
			41223: out = 16'(233);
			41224: out = 16'(222);
			41225: out = 16'(466);
			41226: out = 16'(307);
			41227: out = 16'(-65);
			41228: out = 16'(340);
			41229: out = 16'(490);
			41230: out = 16'(437);
			41231: out = 16'(83);
			41232: out = 16'(-259);
			41233: out = 16'(-49);
			41234: out = 16'(-876);
			41235: out = 16'(-1303);
			41236: out = 16'(-1547);
			41237: out = 16'(-698);
			41238: out = 16'(199);
			41239: out = 16'(662);
			41240: out = 16'(597);
			41241: out = 16'(119);
			41242: out = 16'(-440);
			41243: out = 16'(-911);
			41244: out = 16'(-1145);
			41245: out = 16'(-116);
			41246: out = 16'(546);
			41247: out = 16'(1017);
			41248: out = 16'(677);
			41249: out = 16'(344);
			41250: out = 16'(-30);
			41251: out = 16'(-15);
			41252: out = 16'(-53);
			41253: out = 16'(-58);
			41254: out = 16'(-299);
			41255: out = 16'(-288);
			41256: out = 16'(-87);
			41257: out = 16'(409);
			41258: out = 16'(753);
			41259: out = 16'(779);
			41260: out = 16'(342);
			41261: out = 16'(-213);
			41262: out = 16'(-1073);
			41263: out = 16'(-992);
			41264: out = 16'(-258);
			41265: out = 16'(427);
			41266: out = 16'(854);
			41267: out = 16'(645);
			41268: out = 16'(404);
			41269: out = 16'(-101);
			41270: out = 16'(-325);
			41271: out = 16'(-630);
			41272: out = 16'(-630);
			41273: out = 16'(-709);
			41274: out = 16'(-192);
			41275: out = 16'(211);
			41276: out = 16'(-33);
			41277: out = 16'(117);
			41278: out = 16'(241);
			41279: out = 16'(189);
			41280: out = 16'(-46);
			41281: out = 16'(-415);
			41282: out = 16'(74);
			41283: out = 16'(201);
			41284: out = 16'(235);
			41285: out = 16'(200);
			41286: out = 16'(256);
			41287: out = 16'(184);
			41288: out = 16'(719);
			41289: out = 16'(960);
			41290: out = 16'(920);
			41291: out = 16'(615);
			41292: out = 16'(422);
			41293: out = 16'(874);
			41294: out = 16'(737);
			41295: out = 16'(541);
			41296: out = 16'(176);
			41297: out = 16'(-79);
			41298: out = 16'(-267);
			41299: out = 16'(-514);
			41300: out = 16'(-198);
			41301: out = 16'(394);
			41302: out = 16'(107);
			41303: out = 16'(-463);
			41304: out = 16'(-1766);
			41305: out = 16'(-768);
			41306: out = 16'(-393);
			41307: out = 16'(-175);
			41308: out = 16'(-914);
			41309: out = 16'(-1215);
			41310: out = 16'(-109);
			41311: out = 16'(-211);
			41312: out = 16'(-204);
			41313: out = 16'(-1300);
			41314: out = 16'(-544);
			41315: out = 16'(296);
			41316: out = 16'(1103);
			41317: out = 16'(717);
			41318: out = 16'(-215);
			41319: out = 16'(-714);
			41320: out = 16'(-1065);
			41321: out = 16'(-884);
			41322: out = 16'(-998);
			41323: out = 16'(-654);
			41324: out = 16'(-76);
			41325: out = 16'(151);
			41326: out = 16'(321);
			41327: out = 16'(224);
			41328: out = 16'(426);
			41329: out = 16'(552);
			41330: out = 16'(1019);
			41331: out = 16'(530);
			41332: out = 16'(155);
			41333: out = 16'(-79);
			41334: out = 16'(398);
			41335: out = 16'(980);
			41336: out = 16'(921);
			41337: out = 16'(536);
			41338: out = 16'(-224);
			41339: out = 16'(-109);
			41340: out = 16'(-335);
			41341: out = 16'(-447);
			41342: out = 16'(-450);
			41343: out = 16'(-645);
			41344: out = 16'(-1308);
			41345: out = 16'(-878);
			41346: out = 16'(-471);
			41347: out = 16'(206);
			41348: out = 16'(234);
			41349: out = 16'(187);
			41350: out = 16'(-92);
			41351: out = 16'(-265);
			41352: out = 16'(-431);
			41353: out = 16'(-357);
			41354: out = 16'(-394);
			41355: out = 16'(-341);
			41356: out = 16'(-410);
			41357: out = 16'(-139);
			41358: out = 16'(216);
			41359: out = 16'(821);
			41360: out = 16'(959);
			41361: out = 16'(689);
			41362: out = 16'(350);
			41363: out = 16'(-2);
			41364: out = 16'(0);
			41365: out = 16'(-326);
			41366: out = 16'(-350);
			41367: out = 16'(-194);
			41368: out = 16'(484);
			41369: out = 16'(1051);
			41370: out = 16'(1096);
			41371: out = 16'(981);
			41372: out = 16'(483);
			41373: out = 16'(-24);
			41374: out = 16'(-642);
			41375: out = 16'(-989);
			41376: out = 16'(-404);
			41377: out = 16'(180);
			41378: out = 16'(636);
			41379: out = 16'(108);
			41380: out = 16'(-743);
			41381: out = 16'(-1888);
			41382: out = 16'(-1939);
			41383: out = 16'(-1442);
			41384: out = 16'(-120);
			41385: out = 16'(451);
			41386: out = 16'(892);
			41387: out = 16'(1431);
			41388: out = 16'(944);
			41389: out = 16'(246);
			41390: out = 16'(-566);
			41391: out = 16'(-765);
			41392: out = 16'(-620);
			41393: out = 16'(-218);
			41394: out = 16'(-96);
			41395: out = 16'(-118);
			41396: out = 16'(149);
			41397: out = 16'(537);
			41398: out = 16'(1225);
			41399: out = 16'(647);
			41400: out = 16'(189);
			41401: out = 16'(-433);
			41402: out = 16'(-277);
			41403: out = 16'(74);
			41404: out = 16'(902);
			41405: out = 16'(1073);
			41406: out = 16'(1044);
			41407: out = 16'(418);
			41408: out = 16'(79);
			41409: out = 16'(-255);
			41410: out = 16'(142);
			41411: out = 16'(64);
			41412: out = 16'(13);
			41413: out = 16'(-664);
			41414: out = 16'(-689);
			41415: out = 16'(-438);
			41416: out = 16'(-269);
			41417: out = 16'(-167);
			41418: out = 16'(-208);
			41419: out = 16'(-172);
			41420: out = 16'(-132);
			41421: out = 16'(103);
			41422: out = 16'(-278);
			41423: out = 16'(-383);
			41424: out = 16'(100);
			41425: out = 16'(102);
			41426: out = 16'(237);
			41427: out = 16'(357);
			41428: out = 16'(675);
			41429: out = 16'(856);
			41430: out = 16'(454);
			41431: out = 16'(120);
			41432: out = 16'(-277);
			41433: out = 16'(-198);
			41434: out = 16'(-209);
			41435: out = 16'(-115);
			41436: out = 16'(-2);
			41437: out = 16'(-51);
			41438: out = 16'(-540);
			41439: out = 16'(-80);
			41440: out = 16'(92);
			41441: out = 16'(141);
			41442: out = 16'(-77);
			41443: out = 16'(-250);
			41444: out = 16'(-490);
			41445: out = 16'(-154);
			41446: out = 16'(271);
			41447: out = 16'(789);
			41448: out = 16'(692);
			41449: out = 16'(224);
			41450: out = 16'(-535);
			41451: out = 16'(-1082);
			41452: out = 16'(-1262);
			41453: out = 16'(-1152);
			41454: out = 16'(-601);
			41455: out = 16'(120);
			41456: out = 16'(185);
			41457: out = 16'(87);
			41458: out = 16'(-143);
			41459: out = 16'(-512);
			41460: out = 16'(-737);
			41461: out = 16'(-660);
			41462: out = 16'(-549);
			41463: out = 16'(-287);
			41464: out = 16'(-67);
			41465: out = 16'(87);
			41466: out = 16'(108);
			41467: out = 16'(-329);
			41468: out = 16'(-287);
			41469: out = 16'(-67);
			41470: out = 16'(-379);
			41471: out = 16'(-254);
			41472: out = 16'(-75);
			41473: out = 16'(365);
			41474: out = 16'(519);
			41475: out = 16'(487);
			41476: out = 16'(264);
			41477: out = 16'(120);
			41478: out = 16'(224);
			41479: out = 16'(55);
			41480: out = 16'(-122);
			41481: out = 16'(-384);
			41482: out = 16'(-411);
			41483: out = 16'(-348);
			41484: out = 16'(-187);
			41485: out = 16'(180);
			41486: out = 16'(515);
			41487: out = 16'(453);
			41488: out = 16'(279);
			41489: out = 16'(-130);
			41490: out = 16'(125);
			41491: out = 16'(-32);
			41492: out = 16'(-124);
			41493: out = 16'(-217);
			41494: out = 16'(166);
			41495: out = 16'(911);
			41496: out = 16'(1089);
			41497: out = 16'(1001);
			41498: out = 16'(397);
			41499: out = 16'(70);
			41500: out = 16'(-69);
			41501: out = 16'(844);
			41502: out = 16'(720);
			41503: out = 16'(517);
			41504: out = 16'(-111);
			41505: out = 16'(-115);
			41506: out = 16'(27);
			41507: out = 16'(-20);
			41508: out = 16'(-48);
			41509: out = 16'(-202);
			41510: out = 16'(251);
			41511: out = 16'(340);
			41512: out = 16'(318);
			41513: out = 16'(-100);
			41514: out = 16'(-415);
			41515: out = 16'(-829);
			41516: out = 16'(-469);
			41517: out = 16'(-33);
			41518: out = 16'(821);
			41519: out = 16'(431);
			41520: out = 16'(-185);
			41521: out = 16'(-1519);
			41522: out = 16'(-1701);
			41523: out = 16'(-1482);
			41524: out = 16'(-398);
			41525: out = 16'(15);
			41526: out = 16'(176);
			41527: out = 16'(-351);
			41528: out = 16'(-451);
			41529: out = 16'(-427);
			41530: out = 16'(36);
			41531: out = 16'(269);
			41532: out = 16'(450);
			41533: out = 16'(189);
			41534: out = 16'(63);
			41535: out = 16'(-150);
			41536: out = 16'(548);
			41537: out = 16'(867);
			41538: out = 16'(439);
			41539: out = 16'(-221);
			41540: out = 16'(-869);
			41541: out = 16'(-966);
			41542: out = 16'(-785);
			41543: out = 16'(-344);
			41544: out = 16'(-10);
			41545: out = 16'(146);
			41546: out = 16'(58);
			41547: out = 16'(-734);
			41548: out = 16'(-1062);
			41549: out = 16'(-891);
			41550: out = 16'(-572);
			41551: out = 16'(-406);
			41552: out = 16'(-1005);
			41553: out = 16'(-322);
			41554: out = 16'(52);
			41555: out = 16'(543);
			41556: out = 16'(308);
			41557: out = 16'(118);
			41558: out = 16'(-374);
			41559: out = 16'(-70);
			41560: out = 16'(166);
			41561: out = 16'(34);
			41562: out = 16'(-68);
			41563: out = 16'(-44);
			41564: out = 16'(41);
			41565: out = 16'(607);
			41566: out = 16'(1227);
			41567: out = 16'(1408);
			41568: out = 16'(1100);
			41569: out = 16'(422);
			41570: out = 16'(147);
			41571: out = 16'(160);
			41572: out = 16'(344);
			41573: out = 16'(1036);
			41574: out = 16'(1134);
			41575: out = 16'(190);
			41576: out = 16'(-872);
			41577: out = 16'(-1720);
			41578: out = 16'(-1060);
			41579: out = 16'(-525);
			41580: out = 16'(194);
			41581: out = 16'(27);
			41582: out = 16'(66);
			41583: out = 16'(-144);
			41584: out = 16'(139);
			41585: out = 16'(235);
			41586: out = 16'(422);
			41587: out = 16'(401);
			41588: out = 16'(250);
			41589: out = 16'(-229);
			41590: out = 16'(-553);
			41591: out = 16'(-712);
			41592: out = 16'(-141);
			41593: out = 16'(-189);
			41594: out = 16'(103);
			41595: out = 16'(793);
			41596: out = 16'(1181);
			41597: out = 16'(1185);
			41598: out = 16'(-64);
			41599: out = 16'(-641);
			41600: out = 16'(-1058);
			41601: out = 16'(-244);
			41602: out = 16'(-63);
			41603: out = 16'(93);
			41604: out = 16'(-226);
			41605: out = 16'(134);
			41606: out = 16'(922);
			41607: out = 16'(991);
			41608: out = 16'(1002);
			41609: out = 16'(531);
			41610: out = 16'(621);
			41611: out = 16'(368);
			41612: out = 16'(-250);
			41613: out = 16'(-632);
			41614: out = 16'(-796);
			41615: out = 16'(-183);
			41616: out = 16'(-359);
			41617: out = 16'(-643);
			41618: out = 16'(-1516);
			41619: out = 16'(-1659);
			41620: out = 16'(-1551);
			41621: out = 16'(-1120);
			41622: out = 16'(-738);
			41623: out = 16'(-376);
			41624: out = 16'(-417);
			41625: out = 16'(-216);
			41626: out = 16'(163);
			41627: out = 16'(562);
			41628: out = 16'(761);
			41629: out = 16'(681);
			41630: out = 16'(386);
			41631: out = 16'(-64);
			41632: out = 16'(-358);
			41633: out = 16'(-350);
			41634: out = 16'(-46);
			41635: out = 16'(-179);
			41636: out = 16'(459);
			41637: out = 16'(890);
			41638: out = 16'(327);
			41639: out = 16'(-333);
			41640: out = 16'(-995);
			41641: out = 16'(-288);
			41642: out = 16'(379);
			41643: out = 16'(1174);
			41644: out = 16'(1336);
			41645: out = 16'(1212);
			41646: out = 16'(858);
			41647: out = 16'(111);
			41648: out = 16'(-321);
			41649: out = 16'(-248);
			41650: out = 16'(249);
			41651: out = 16'(596);
			41652: out = 16'(77);
			41653: out = 16'(-74);
			41654: out = 16'(-249);
			41655: out = 16'(565);
			41656: out = 16'(356);
			41657: out = 16'(-21);
			41658: out = 16'(-421);
			41659: out = 16'(-525);
			41660: out = 16'(-216);
			41661: out = 16'(-1430);
			41662: out = 16'(-1580);
			41663: out = 16'(-1329);
			41664: out = 16'(108);
			41665: out = 16'(897);
			41666: out = 16'(1096);
			41667: out = 16'(346);
			41668: out = 16'(-217);
			41669: out = 16'(121);
			41670: out = 16'(0);
			41671: out = 16'(19);
			41672: out = 16'(-494);
			41673: out = 16'(-346);
			41674: out = 16'(-156);
			41675: out = 16'(98);
			41676: out = 16'(161);
			41677: out = 16'(82);
			41678: out = 16'(-44);
			41679: out = 16'(-367);
			41680: out = 16'(-737);
			41681: out = 16'(-978);
			41682: out = 16'(-709);
			41683: out = 16'(124);
			41684: out = 16'(170);
			41685: out = 16'(106);
			41686: out = 16'(-140);
			41687: out = 16'(-663);
			41688: out = 16'(-1039);
			41689: out = 16'(-912);
			41690: out = 16'(-964);
			41691: out = 16'(-817);
			41692: out = 16'(-186);
			41693: out = 16'(-11);
			41694: out = 16'(24);
			41695: out = 16'(150);
			41696: out = 16'(248);
			41697: out = 16'(217);
			41698: out = 16'(701);
			41699: out = 16'(480);
			41700: out = 16'(-138);
			41701: out = 16'(-708);
			41702: out = 16'(-863);
			41703: out = 16'(-311);
			41704: out = 16'(-159);
			41705: out = 16'(134);
			41706: out = 16'(464);
			41707: out = 16'(510);
			41708: out = 16'(516);
			41709: out = 16'(697);
			41710: out = 16'(939);
			41711: out = 16'(1165);
			41712: out = 16'(714);
			41713: out = 16'(430);
			41714: out = 16'(-22);
			41715: out = 16'(-331);
			41716: out = 16'(-627);
			41717: out = 16'(-674);
			41718: out = 16'(-373);
			41719: out = 16'(146);
			41720: out = 16'(657);
			41721: out = 16'(858);
			41722: out = 16'(710);
			41723: out = 16'(151);
			41724: out = 16'(-76);
			41725: out = 16'(-218);
			41726: out = 16'(61);
			41727: out = 16'(39);
			41728: out = 16'(28);
			41729: out = 16'(-217);
			41730: out = 16'(-95);
			41731: out = 16'(102);
			41732: out = 16'(300);
			41733: out = 16'(675);
			41734: out = 16'(1093);
			41735: out = 16'(483);
			41736: out = 16'(140);
			41737: out = 16'(-218);
			41738: out = 16'(-153);
			41739: out = 16'(-285);
			41740: out = 16'(-509);
			41741: out = 16'(-724);
			41742: out = 16'(-697);
			41743: out = 16'(-218);
			41744: out = 16'(-241);
			41745: out = 16'(-159);
			41746: out = 16'(121);
			41747: out = 16'(96);
			41748: out = 16'(-55);
			41749: out = 16'(-945);
			41750: out = 16'(-853);
			41751: out = 16'(-375);
			41752: out = 16'(-70);
			41753: out = 16'(87);
			41754: out = 16'(-183);
			41755: out = 16'(932);
			41756: out = 16'(1043);
			41757: out = 16'(875);
			41758: out = 16'(-513);
			41759: out = 16'(-1142);
			41760: out = 16'(-705);
			41761: out = 16'(-485);
			41762: out = 16'(-184);
			41763: out = 16'(-831);
			41764: out = 16'(-57);
			41765: out = 16'(563);
			41766: out = 16'(1064);
			41767: out = 16'(916);
			41768: out = 16'(503);
			41769: out = 16'(242);
			41770: out = 16'(-309);
			41771: out = 16'(-830);
			41772: out = 16'(-806);
			41773: out = 16'(-469);
			41774: out = 16'(192);
			41775: out = 16'(-97);
			41776: out = 16'(-258);
			41777: out = 16'(-798);
			41778: out = 16'(-362);
			41779: out = 16'(-57);
			41780: out = 16'(455);
			41781: out = 16'(43);
			41782: out = 16'(-93);
			41783: out = 16'(51);
			41784: out = 16'(90);
			41785: out = 16'(12);
			41786: out = 16'(136);
			41787: out = 16'(-361);
			41788: out = 16'(-744);
			41789: out = 16'(-541);
			41790: out = 16'(-81);
			41791: out = 16'(449);
			41792: out = 16'(657);
			41793: out = 16'(309);
			41794: out = 16'(-506);
			41795: out = 16'(-889);
			41796: out = 16'(-809);
			41797: out = 16'(-59);
			41798: out = 16'(273);
			41799: out = 16'(222);
			41800: out = 16'(-999);
			41801: out = 16'(-1138);
			41802: out = 16'(-1093);
			41803: out = 16'(171);
			41804: out = 16'(563);
			41805: out = 16'(1059);
			41806: out = 16'(853);
			41807: out = 16'(1090);
			41808: out = 16'(1080);
			41809: out = 16'(1199);
			41810: out = 16'(838);
			41811: out = 16'(608);
			41812: out = 16'(-748);
			41813: out = 16'(-1047);
			41814: out = 16'(-780);
			41815: out = 16'(379);
			41816: out = 16'(862);
			41817: out = 16'(302);
			41818: out = 16'(-281);
			41819: out = 16'(-1041);
			41820: out = 16'(-1240);
			41821: out = 16'(-1419);
			41822: out = 16'(-1070);
			41823: out = 16'(-259);
			41824: out = 16'(480);
			41825: out = 16'(889);
			41826: out = 16'(16);
			41827: out = 16'(-129);
			41828: out = 16'(-90);
			41829: out = 16'(-371);
			41830: out = 16'(-708);
			41831: out = 16'(-1330);
			41832: out = 16'(-101);
			41833: out = 16'(380);
			41834: out = 16'(731);
			41835: out = 16'(-64);
			41836: out = 16'(-459);
			41837: out = 16'(-358);
			41838: out = 16'(-40);
			41839: out = 16'(227);
			41840: out = 16'(160);
			41841: out = 16'(55);
			41842: out = 16'(-53);
			41843: out = 16'(384);
			41844: out = 16'(489);
			41845: out = 16'(637);
			41846: out = 16'(361);
			41847: out = 16'(460);
			41848: out = 16'(578);
			41849: out = 16'(394);
			41850: out = 16'(253);
			41851: out = 16'(-8);
			41852: out = 16'(67);
			41853: out = 16'(-149);
			41854: out = 16'(-703);
			41855: out = 16'(-986);
			41856: out = 16'(-1288);
			41857: out = 16'(-1350);
			41858: out = 16'(-1441);
			41859: out = 16'(-1159);
			41860: out = 16'(-172);
			41861: out = 16'(24);
			41862: out = 16'(-25);
			41863: out = 16'(-8);
			41864: out = 16'(-129);
			41865: out = 16'(-9);
			41866: out = 16'(-64);
			41867: out = 16'(170);
			41868: out = 16'(181);
			41869: out = 16'(1006);
			41870: out = 16'(759);
			41871: out = 16'(-16);
			41872: out = 16'(-994);
			41873: out = 16'(-1202);
			41874: out = 16'(-297);
			41875: out = 16'(671);
			41876: out = 16'(1476);
			41877: out = 16'(1212);
			41878: out = 16'(1000);
			41879: out = 16'(459);
			41880: out = 16'(489);
			41881: out = 16'(79);
			41882: out = 16'(-83);
			41883: out = 16'(-134);
			41884: out = 16'(24);
			41885: out = 16'(96);
			41886: out = 16'(-66);
			41887: out = 16'(-304);
			41888: out = 16'(-368);
			41889: out = 16'(-302);
			41890: out = 16'(61);
			41891: out = 16'(328);
			41892: out = 16'(843);
			41893: out = 16'(926);
			41894: out = 16'(604);
			41895: out = 16'(-176);
			41896: out = 16'(-952);
			41897: out = 16'(-1898);
			41898: out = 16'(-1718);
			41899: out = 16'(-1262);
			41900: out = 16'(-698);
			41901: out = 16'(-465);
			41902: out = 16'(-252);
			41903: out = 16'(20);
			41904: out = 16'(578);
			41905: out = 16'(1119);
			41906: out = 16'(1457);
			41907: out = 16'(1008);
			41908: out = 16'(-136);
			41909: out = 16'(-810);
			41910: out = 16'(-1071);
			41911: out = 16'(-295);
			41912: out = 16'(-269);
			41913: out = 16'(-1);
			41914: out = 16'(69);
			41915: out = 16'(206);
			41916: out = 16'(204);
			41917: out = 16'(636);
			41918: out = 16'(605);
			41919: out = 16'(603);
			41920: out = 16'(172);
			41921: out = 16'(168);
			41922: out = 16'(87);
			41923: out = 16'(191);
			41924: out = 16'(-154);
			41925: out = 16'(-680);
			41926: out = 16'(-1046);
			41927: out = 16'(-1169);
			41928: out = 16'(-1114);
			41929: out = 16'(-598);
			41930: out = 16'(-262);
			41931: out = 16'(-370);
			41932: out = 16'(-154);
			41933: out = 16'(-63);
			41934: out = 16'(16);
			41935: out = 16'(-56);
			41936: out = 16'(-67);
			41937: out = 16'(-7);
			41938: out = 16'(-25);
			41939: out = 16'(-6);
			41940: out = 16'(-91);
			41941: out = 16'(126);
			41942: out = 16'(488);
			41943: out = 16'(217);
			41944: out = 16'(222);
			41945: out = 16'(123);
			41946: out = 16'(661);
			41947: out = 16'(948);
			41948: out = 16'(1040);
			41949: out = 16'(761);
			41950: out = 16'(523);
			41951: out = 16'(625);
			41952: out = 16'(273);
			41953: out = 16'(71);
			41954: out = 16'(-146);
			41955: out = 16'(-14);
			41956: out = 16'(77);
			41957: out = 16'(-85);
			41958: out = 16'(-282);
			41959: out = 16'(-454);
			41960: out = 16'(-910);
			41961: out = 16'(-589);
			41962: out = 16'(150);
			41963: out = 16'(433);
			41964: out = 16'(683);
			41965: out = 16'(758);
			41966: out = 16'(311);
			41967: out = 16'(-265);
			41968: out = 16'(-926);
			41969: out = 16'(-954);
			41970: out = 16'(-904);
			41971: out = 16'(-909);
			41972: out = 16'(-749);
			41973: out = 16'(-529);
			41974: out = 16'(23);
			41975: out = 16'(405);
			41976: out = 16'(665);
			41977: out = 16'(636);
			41978: out = 16'(397);
			41979: out = 16'(34);
			41980: out = 16'(103);
			41981: out = 16'(53);
			41982: out = 16'(69);
			41983: out = 16'(-300);
			41984: out = 16'(-431);
			41985: out = 16'(-373);
			41986: out = 16'(-225);
			41987: out = 16'(109);
			41988: out = 16'(585);
			41989: out = 16'(623);
			41990: out = 16'(555);
			41991: out = 16'(618);
			41992: out = 16'(192);
			41993: out = 16'(-218);
			41994: out = 16'(-636);
			41995: out = 16'(-692);
			41996: out = 16'(-687);
			41997: out = 16'(-857);
			41998: out = 16'(-1012);
			41999: out = 16'(-1097);
			42000: out = 16'(-770);
			42001: out = 16'(-319);
			42002: out = 16'(152);
			42003: out = 16'(692);
			42004: out = 16'(977);
			42005: out = 16'(1316);
			42006: out = 16'(514);
			42007: out = 16'(50);
			42008: out = 16'(-108);
			42009: out = 16'(326);
			42010: out = 16'(545);
			42011: out = 16'(-54);
			42012: out = 16'(-519);
			42013: out = 16'(-921);
			42014: out = 16'(-451);
			42015: out = 16'(-145);
			42016: out = 16'(218);
			42017: out = 16'(534);
			42018: out = 16'(544);
			42019: out = 16'(327);
			42020: out = 16'(-585);
			42021: out = 16'(-1137);
			42022: out = 16'(-1407);
			42023: out = 16'(-392);
			42024: out = 16'(403);
			42025: out = 16'(807);
			42026: out = 16'(604);
			42027: out = 16'(216);
			42028: out = 16'(-352);
			42029: out = 16'(-161);
			42030: out = 16'(155);
			42031: out = 16'(121);
			42032: out = 16'(168);
			42033: out = 16'(22);
			42034: out = 16'(119);
			42035: out = 16'(-55);
			42036: out = 16'(-166);
			42037: out = 16'(-368);
			42038: out = 16'(-340);
			42039: out = 16'(-135);
			42040: out = 16'(-691);
			42041: out = 16'(-876);
			42042: out = 16'(-561);
			42043: out = 16'(-505);
			42044: out = 16'(-168);
			42045: out = 16'(55);
			42046: out = 16'(884);
			42047: out = 16'(1290);
			42048: out = 16'(1083);
			42049: out = 16'(557);
			42050: out = 16'(-25);
			42051: out = 16'(174);
			42052: out = 16'(190);
			42053: out = 16'(346);
			42054: out = 16'(-768);
			42055: out = 16'(-870);
			42056: out = 16'(-589);
			42057: out = 16'(-237);
			42058: out = 16'(111);
			42059: out = 16'(369);
			42060: out = 16'(591);
			42061: out = 16'(423);
			42062: out = 16'(-194);
			42063: out = 16'(-168);
			42064: out = 16'(-86);
			42065: out = 16'(368);
			42066: out = 16'(214);
			42067: out = 16'(-84);
			42068: out = 16'(-861);
			42069: out = 16'(-822);
			42070: out = 16'(-555);
			42071: out = 16'(-165);
			42072: out = 16'(71);
			42073: out = 16'(178);
			42074: out = 16'(548);
			42075: out = 16'(676);
			42076: out = 16'(836);
			42077: out = 16'(260);
			42078: out = 16'(-38);
			42079: out = 16'(-467);
			42080: out = 16'(-225);
			42081: out = 16'(-174);
			42082: out = 16'(147);
			42083: out = 16'(-638);
			42084: out = 16'(-757);
			42085: out = 16'(-16);
			42086: out = 16'(768);
			42087: out = 16'(1156);
			42088: out = 16'(234);
			42089: out = 16'(-494);
			42090: out = 16'(-1261);
			42091: out = 16'(-936);
			42092: out = 16'(-625);
			42093: out = 16'(-55);
			42094: out = 16'(273);
			42095: out = 16'(430);
			42096: out = 16'(354);
			42097: out = 16'(-333);
			42098: out = 16'(-838);
			42099: out = 16'(-1127);
			42100: out = 16'(-447);
			42101: out = 16'(228);
			42102: out = 16'(820);
			42103: out = 16'(626);
			42104: out = 16'(289);
			42105: out = 16'(220);
			42106: out = 16'(-5);
			42107: out = 16'(-243);
			42108: out = 16'(-566);
			42109: out = 16'(-776);
			42110: out = 16'(-852);
			42111: out = 16'(-903);
			42112: out = 16'(-560);
			42113: out = 16'(-25);
			42114: out = 16'(490);
			42115: out = 16'(818);
			42116: out = 16'(1083);
			42117: out = 16'(256);
			42118: out = 16'(-105);
			42119: out = 16'(142);
			42120: out = 16'(97);
			42121: out = 16'(266);
			42122: out = 16'(595);
			42123: out = 16'(357);
			42124: out = 16'(26);
			42125: out = 16'(-579);
			42126: out = 16'(-677);
			42127: out = 16'(-504);
			42128: out = 16'(660);
			42129: out = 16'(874);
			42130: out = 16'(736);
			42131: out = 16'(-346);
			42132: out = 16'(-910);
			42133: out = 16'(-1126);
			42134: out = 16'(-413);
			42135: out = 16'(37);
			42136: out = 16'(158);
			42137: out = 16'(55);
			42138: out = 16'(-206);
			42139: out = 16'(-577);
			42140: out = 16'(-643);
			42141: out = 16'(-494);
			42142: out = 16'(-142);
			42143: out = 16'(-28);
			42144: out = 16'(-23);
			42145: out = 16'(-17);
			42146: out = 16'(61);
			42147: out = 16'(263);
			42148: out = 16'(163);
			42149: out = 16'(302);
			42150: out = 16'(413);
			42151: out = 16'(452);
			42152: out = 16'(211);
			42153: out = 16'(-135);
			42154: out = 16'(-506);
			42155: out = 16'(-479);
			42156: out = 16'(152);
			42157: out = 16'(151);
			42158: out = 16'(187);
			42159: out = 16'(111);
			42160: out = 16'(139);
			42161: out = 16'(228);
			42162: out = 16'(356);
			42163: out = 16'(419);
			42164: out = 16'(374);
			42165: out = 16'(825);
			42166: out = 16'(392);
			42167: out = 16'(-189);
			42168: out = 16'(-992);
			42169: out = 16'(-1046);
			42170: out = 16'(-553);
			42171: out = 16'(-263);
			42172: out = 16'(181);
			42173: out = 16'(629);
			42174: out = 16'(469);
			42175: out = 16'(238);
			42176: out = 16'(-452);
			42177: out = 16'(-190);
			42178: out = 16'(-175);
			42179: out = 16'(192);
			42180: out = 16'(-925);
			42181: out = 16'(-1741);
			42182: out = 16'(-1678);
			42183: out = 16'(-770);
			42184: out = 16'(468);
			42185: out = 16'(1101);
			42186: out = 16'(1322);
			42187: out = 16'(986);
			42188: out = 16'(570);
			42189: out = 16'(386);
			42190: out = 16'(656);
			42191: out = 16'(249);
			42192: out = 16'(-66);
			42193: out = 16'(-676);
			42194: out = 16'(-652);
			42195: out = 16'(-551);
			42196: out = 16'(-59);
			42197: out = 16'(30);
			42198: out = 16'(62);
			42199: out = 16'(-374);
			42200: out = 16'(-253);
			42201: out = 16'(-104);
			42202: out = 16'(66);
			42203: out = 16'(71);
			42204: out = 16'(-77);
			42205: out = 16'(165);
			42206: out = 16'(58);
			42207: out = 16'(-77);
			42208: out = 16'(-702);
			42209: out = 16'(-927);
			42210: out = 16'(-837);
			42211: out = 16'(-350);
			42212: out = 16'(-30);
			42213: out = 16'(-158);
			42214: out = 16'(-41);
			42215: out = 16'(-232);
			42216: out = 16'(-502);
			42217: out = 16'(-900);
			42218: out = 16'(-1005);
			42219: out = 16'(-121);
			42220: out = 16'(10);
			42221: out = 16'(32);
			42222: out = 16'(-45);
			42223: out = 16'(23);
			42224: out = 16'(244);
			42225: out = 16'(387);
			42226: out = 16'(592);
			42227: out = 16'(668);
			42228: out = 16'(1032);
			42229: out = 16'(1013);
			42230: out = 16'(859);
			42231: out = 16'(326);
			42232: out = 16'(15);
			42233: out = 16'(-88);
			42234: out = 16'(340);
			42235: out = 16'(579);
			42236: out = 16'(129);
			42237: out = 16'(107);
			42238: out = 16'(40);
			42239: out = 16'(51);
			42240: out = 16'(64);
			42241: out = 16'(55);
			42242: out = 16'(323);
			42243: out = 16'(325);
			42244: out = 16'(349);
			42245: out = 16'(-81);
			42246: out = 16'(24);
			42247: out = 16'(312);
			42248: out = 16'(373);
			42249: out = 16'(35);
			42250: out = 16'(-678);
			42251: out = 16'(-1091);
			42252: out = 16'(-1012);
			42253: out = 16'(-236);
			42254: out = 16'(411);
			42255: out = 16'(851);
			42256: out = 16'(805);
			42257: out = 16'(187);
			42258: out = 16'(-598);
			42259: out = 16'(-631);
			42260: out = 16'(-436);
			42261: out = 16'(134);
			42262: out = 16'(-231);
			42263: out = 16'(-53);
			42264: out = 16'(38);
			42265: out = 16'(137);
			42266: out = 16'(82);
			42267: out = 16'(57);
			42268: out = 16'(-311);
			42269: out = 16'(-415);
			42270: out = 16'(-149);
			42271: out = 16'(-200);
			42272: out = 16'(-195);
			42273: out = 16'(-451);
			42274: out = 16'(-116);
			42275: out = 16'(119);
			42276: out = 16'(383);
			42277: out = 16'(142);
			42278: out = 16'(-159);
			42279: out = 16'(-360);
			42280: out = 16'(-427);
			42281: out = 16'(-351);
			42282: out = 16'(418);
			42283: out = 16'(710);
			42284: out = 16'(778);
			42285: out = 16'(82);
			42286: out = 16'(-329);
			42287: out = 16'(-406);
			42288: out = 16'(-292);
			42289: out = 16'(-226);
			42290: out = 16'(-725);
			42291: out = 16'(-454);
			42292: out = 16'(-425);
			42293: out = 16'(-352);
			42294: out = 16'(-570);
			42295: out = 16'(-504);
			42296: out = 16'(67);
			42297: out = 16'(536);
			42298: out = 16'(826);
			42299: out = 16'(704);
			42300: out = 16'(275);
			42301: out = 16'(-182);
			42302: out = 16'(-223);
			42303: out = 16'(174);
			42304: out = 16'(828);
			42305: out = 16'(661);
			42306: out = 16'(355);
			42307: out = 16'(-177);
			42308: out = 16'(-565);
			42309: out = 16'(-534);
			42310: out = 16'(22);
			42311: out = 16'(630);
			42312: out = 16'(1057);
			42313: out = 16'(986);
			42314: out = 16'(544);
			42315: out = 16'(-49);
			42316: out = 16'(-82);
			42317: out = 16'(-207);
			42318: out = 16'(-135);
			42319: out = 16'(-10);
			42320: out = 16'(-145);
			42321: out = 16'(-496);
			42322: out = 16'(-274);
			42323: out = 16'(-179);
			42324: out = 16'(-143);
			42325: out = 16'(23);
			42326: out = 16'(-245);
			42327: out = 16'(-1207);
			42328: out = 16'(-1197);
			42329: out = 16'(-1002);
			42330: out = 16'(-182);
			42331: out = 16'(-134);
			42332: out = 16'(-141);
			42333: out = 16'(-123);
			42334: out = 16'(-261);
			42335: out = 16'(-388);
			42336: out = 16'(-599);
			42337: out = 16'(-432);
			42338: out = 16'(-58);
			42339: out = 16'(137);
			42340: out = 16'(351);
			42341: out = 16'(672);
			42342: out = 16'(271);
			42343: out = 16'(117);
			42344: out = 16'(-98);
			42345: out = 16'(282);
			42346: out = 16'(339);
			42347: out = 16'(204);
			42348: out = 16'(-344);
			42349: out = 16'(-637);
			42350: out = 16'(-417);
			42351: out = 16'(162);
			42352: out = 16'(722);
			42353: out = 16'(776);
			42354: out = 16'(645);
			42355: out = 16'(276);
			42356: out = 16'(-259);
			42357: out = 16'(-642);
			42358: out = 16'(-906);
			42359: out = 16'(-116);
			42360: out = 16'(82);
			42361: out = 16'(-101);
			42362: out = 16'(-453);
			42363: out = 16'(-684);
			42364: out = 16'(-601);
			42365: out = 16'(-188);
			42366: out = 16'(193);
			42367: out = 16'(-102);
			42368: out = 16'(134);
			42369: out = 16'(100);
			42370: out = 16'(-287);
			42371: out = 16'(-624);
			42372: out = 16'(-768);
			42373: out = 16'(505);
			42374: out = 16'(689);
			42375: out = 16'(604);
			42376: out = 16'(9);
			42377: out = 16'(-107);
			42378: out = 16'(151);
			42379: out = 16'(-120);
			42380: out = 16'(-165);
			42381: out = 16'(-411);
			42382: out = 16'(332);
			42383: out = 16'(811);
			42384: out = 16'(1239);
			42385: out = 16'(978);
			42386: out = 16'(728);
			42387: out = 16'(808);
			42388: out = 16'(512);
			42389: out = 16'(225);
			42390: out = 16'(-127);
			42391: out = 16'(-72);
			42392: out = 16'(93);
			42393: out = 16'(-184);
			42394: out = 16'(-142);
			42395: out = 16'(-217);
			42396: out = 16'(-93);
			42397: out = 16'(-533);
			42398: out = 16'(-1240);
			42399: out = 16'(-1437);
			42400: out = 16'(-1161);
			42401: out = 16'(-109);
			42402: out = 16'(-134);
			42403: out = 16'(-11);
			42404: out = 16'(78);
			42405: out = 16'(83);
			42406: out = 16'(72);
			42407: out = 16'(-96);
			42408: out = 16'(264);
			42409: out = 16'(613);
			42410: out = 16'(-79);
			42411: out = 16'(-79);
			42412: out = 16'(-105);
			42413: out = 16'(322);
			42414: out = 16'(197);
			42415: out = 16'(-149);
			42416: out = 16'(-301);
			42417: out = 16'(-474);
			42418: out = 16'(-364);
			42419: out = 16'(-629);
			42420: out = 16'(-512);
			42421: out = 16'(-157);
			42422: out = 16'(226);
			42423: out = 16'(394);
			42424: out = 16'(147);
			42425: out = 16'(138);
			42426: out = 16'(43);
			42427: out = 16'(-110);
			42428: out = 16'(-404);
			42429: out = 16'(-654);
			42430: out = 16'(-86);
			42431: out = 16'(-4);
			42432: out = 16'(112);
			42433: out = 16'(-761);
			42434: out = 16'(-623);
			42435: out = 16'(-97);
			42436: out = 16'(97);
			42437: out = 16'(-186);
			42438: out = 16'(-1155);
			42439: out = 16'(-1238);
			42440: out = 16'(-1370);
			42441: out = 16'(-1301);
			42442: out = 16'(-732);
			42443: out = 16'(101);
			42444: out = 16'(1260);
			42445: out = 16'(1442);
			42446: out = 16'(1181);
			42447: out = 16'(394);
			42448: out = 16'(-184);
			42449: out = 16'(-571);
			42450: out = 16'(-96);
			42451: out = 16'(240);
			42452: out = 16'(734);
			42453: out = 16'(57);
			42454: out = 16'(48);
			42455: out = 16'(188);
			42456: out = 16'(736);
			42457: out = 16'(657);
			42458: out = 16'(-76);
			42459: out = 16'(-244);
			42460: out = 16'(-310);
			42461: out = 16'(182);
			42462: out = 16'(423);
			42463: out = 16'(650);
			42464: out = 16'(387);
			42465: out = 16'(174);
			42466: out = 16'(-169);
			42467: out = 16'(-94);
			42468: out = 16'(-205);
			42469: out = 16'(-107);
			42470: out = 16'(-144);
			42471: out = 16'(65);
			42472: out = 16'(91);
			42473: out = 16'(187);
			42474: out = 16'(-245);
			42475: out = 16'(-877);
			42476: out = 16'(-1118);
			42477: out = 16'(-880);
			42478: out = 16'(-62);
			42479: out = 16'(538);
			42480: out = 16'(815);
			42481: out = 16'(182);
			42482: out = 16'(27);
			42483: out = 16'(-180);
			42484: out = 16'(-132);
			42485: out = 16'(10);
			42486: out = 16'(183);
			42487: out = 16'(-23);
			42488: out = 16'(-277);
			42489: out = 16'(-655);
			42490: out = 16'(-192);
			42491: out = 16'(-91);
			42492: out = 16'(-33);
			42493: out = 16'(-257);
			42494: out = 16'(-498);
			42495: out = 16'(-845);
			42496: out = 16'(-670);
			42497: out = 16'(-527);
			42498: out = 16'(-605);
			42499: out = 16'(71);
			42500: out = 16'(648);
			42501: out = 16'(1063);
			42502: out = 16'(821);
			42503: out = 16'(291);
			42504: out = 16'(88);
			42505: out = 16'(-245);
			42506: out = 16'(-346);
			42507: out = 16'(-1051);
			42508: out = 16'(-801);
			42509: out = 16'(-273);
			42510: out = 16'(39);
			42511: out = 16'(136);
			42512: out = 16'(-96);
			42513: out = 16'(-7);
			42514: out = 16'(140);
			42515: out = 16'(714);
			42516: out = 16'(514);
			42517: out = 16'(308);
			42518: out = 16'(-322);
			42519: out = 16'(-359);
			42520: out = 16'(-212);
			42521: out = 16'(597);
			42522: out = 16'(867);
			42523: out = 16'(1049);
			42524: out = 16'(11);
			42525: out = 16'(13);
			42526: out = 16'(81);
			42527: out = 16'(219);
			42528: out = 16'(-210);
			42529: out = 16'(-910);
			42530: out = 16'(-901);
			42531: out = 16'(-524);
			42532: out = 16'(488);
			42533: out = 16'(250);
			42534: out = 16'(93);
			42535: out = 16'(-379);
			42536: out = 16'(-194);
			42537: out = 16'(-134);
			42538: out = 16'(-360);
			42539: out = 16'(-168);
			42540: out = 16'(65);
			42541: out = 16'(588);
			42542: out = 16'(576);
			42543: out = 16'(367);
			42544: out = 16'(227);
			42545: out = 16'(44);
			42546: out = 16'(-58);
			42547: out = 16'(60);
			42548: out = 16'(131);
			42549: out = 16'(151);
			42550: out = 16'(4);
			42551: out = 16'(-270);
			42552: out = 16'(-898);
			42553: out = 16'(-558);
			42554: out = 16'(-219);
			42555: out = 16'(174);
			42556: out = 16'(156);
			42557: out = 16'(117);
			42558: out = 16'(105);
			42559: out = 16'(251);
			42560: out = 16'(412);
			42561: out = 16'(182);
			42562: out = 16'(146);
			42563: out = 16'(61);
			42564: out = 16'(-34);
			42565: out = 16'(-127);
			42566: out = 16'(-61);
			42567: out = 16'(-509);
			42568: out = 16'(-791);
			42569: out = 16'(-1152);
			42570: out = 16'(-569);
			42571: out = 16'(-212);
			42572: out = 16'(-3);
			42573: out = 16'(93);
			42574: out = 16'(183);
			42575: out = 16'(108);
			42576: out = 16'(251);
			42577: out = 16'(151);
			42578: out = 16'(260);
			42579: out = 16'(-621);
			42580: out = 16'(-1390);
			42581: out = 16'(-1140);
			42582: out = 16'(-505);
			42583: out = 16'(377);
			42584: out = 16'(783);
			42585: out = 16'(825);
			42586: out = 16'(402);
			42587: out = 16'(136);
			42588: out = 16'(-65);
			42589: out = 16'(14);
			42590: out = 16'(412);
			42591: out = 16'(743);
			42592: out = 16'(598);
			42593: out = 16'(282);
			42594: out = 16'(-207);
			42595: out = 16'(-251);
			42596: out = 16'(-683);
			42597: out = 16'(-840);
			42598: out = 16'(-1150);
			42599: out = 16'(-516);
			42600: out = 16'(285);
			42601: out = 16'(396);
			42602: out = 16'(336);
			42603: out = 16'(-84);
			42604: out = 16'(253);
			42605: out = 16'(90);
			42606: out = 16'(-60);
			42607: out = 16'(-654);
			42608: out = 16'(-634);
			42609: out = 16'(205);
			42610: out = 16'(202);
			42611: out = 16'(136);
			42612: out = 16'(-569);
			42613: out = 16'(-285);
			42614: out = 16'(58);
			42615: out = 16'(629);
			42616: out = 16'(808);
			42617: out = 16'(865);
			42618: out = 16'(668);
			42619: out = 16'(545);
			42620: out = 16'(364);
			42621: out = 16'(180);
			42622: out = 16'(-107);
			42623: out = 16'(-393);
			42624: out = 16'(-220);
			42625: out = 16'(-50);
			42626: out = 16'(81);
			42627: out = 16'(259);
			42628: out = 16'(394);
			42629: out = 16'(532);
			42630: out = 16'(283);
			42631: out = 16'(35);
			42632: out = 16'(-54);
			42633: out = 16'(-357);
			42634: out = 16'(-655);
			42635: out = 16'(-767);
			42636: out = 16'(-722);
			42637: out = 16'(-513);
			42638: out = 16'(-990);
			42639: out = 16'(-633);
			42640: out = 16'(-14);
			42641: out = 16'(294);
			42642: out = 16'(325);
			42643: out = 16'(-89);
			42644: out = 16'(-161);
			42645: out = 16'(-322);
			42646: out = 16'(-5);
			42647: out = 16'(-558);
			42648: out = 16'(-691);
			42649: out = 16'(-527);
			42650: out = 16'(-56);
			42651: out = 16'(296);
			42652: out = 16'(396);
			42653: out = 16'(295);
			42654: out = 16'(115);
			42655: out = 16'(-61);
			42656: out = 16'(4);
			42657: out = 16'(153);
			42658: out = 16'(511);
			42659: out = 16'(659);
			42660: out = 16'(757);
			42661: out = 16'(123);
			42662: out = 16'(-66);
			42663: out = 16'(103);
			42664: out = 16'(388);
			42665: out = 16'(579);
			42666: out = 16'(508);
			42667: out = 16'(259);
			42668: out = 16'(-53);
			42669: out = 16'(-136);
			42670: out = 16'(-208);
			42671: out = 16'(-144);
			42672: out = 16'(-187);
			42673: out = 16'(-113);
			42674: out = 16'(-94);
			42675: out = 16'(73);
			42676: out = 16'(-215);
			42677: out = 16'(-619);
			42678: out = 16'(-35);
			42679: out = 16'(105);
			42680: out = 16'(126);
			42681: out = 16'(-38);
			42682: out = 16'(-94);
			42683: out = 16'(-168);
			42684: out = 16'(1);
			42685: out = 16'(123);
			42686: out = 16'(333);
			42687: out = 16'(200);
			42688: out = 16'(52);
			42689: out = 16'(-368);
			42690: out = 16'(-367);
			42691: out = 16'(-367);
			42692: out = 16'(-132);
			42693: out = 16'(-261);
			42694: out = 16'(-359);
			42695: out = 16'(-782);
			42696: out = 16'(-447);
			42697: out = 16'(154);
			42698: out = 16'(614);
			42699: out = 16'(770);
			42700: out = 16'(735);
			42701: out = 16'(269);
			42702: out = 16'(189);
			42703: out = 16'(503);
			42704: out = 16'(794);
			42705: out = 16'(561);
			42706: out = 16'(-1087);
			42707: out = 16'(-1214);
			42708: out = 16'(-1210);
			42709: out = 16'(-397);
			42710: out = 16'(-166);
			42711: out = 16'(144);
			42712: out = 16'(29);
			42713: out = 16'(314);
			42714: out = 16'(531);
			42715: out = 16'(381);
			42716: out = 16'(217);
			42717: out = 16'(28);
			42718: out = 16'(-101);
			42719: out = 16'(-242);
			42720: out = 16'(-385);
			42721: out = 16'(-239);
			42722: out = 16'(7);
			42723: out = 16'(557);
			42724: out = 16'(359);
			42725: out = 16'(317);
			42726: out = 16'(266);
			42727: out = 16'(545);
			42728: out = 16'(591);
			42729: out = 16'(-64);
			42730: out = 16'(-386);
			42731: out = 16'(-641);
			42732: out = 16'(-238);
			42733: out = 16'(-113);
			42734: out = 16'(24);
			42735: out = 16'(-687);
			42736: out = 16'(-879);
			42737: out = 16'(-777);
			42738: out = 16'(-209);
			42739: out = 16'(352);
			42740: out = 16'(668);
			42741: out = 16'(913);
			42742: out = 16'(653);
			42743: out = 16'(-69);
			42744: out = 16'(-712);
			42745: out = 16'(-1098);
			42746: out = 16'(-825);
			42747: out = 16'(-474);
			42748: out = 16'(-54);
			42749: out = 16'(-196);
			42750: out = 16'(-60);
			42751: out = 16'(-68);
			42752: out = 16'(110);
			42753: out = 16'(-97);
			42754: out = 16'(-338);
			42755: out = 16'(48);
			42756: out = 16'(307);
			42757: out = 16'(556);
			42758: out = 16'(413);
			42759: out = 16'(263);
			42760: out = 16'(146);
			42761: out = 16'(-22);
			42762: out = 16'(-109);
			42763: out = 16'(-133);
			42764: out = 16'(-38);
			42765: out = 16'(41);
			42766: out = 16'(-364);
			42767: out = 16'(-254);
			42768: out = 16'(-62);
			42769: out = 16'(637);
			42770: out = 16'(738);
			42771: out = 16'(673);
			42772: out = 16'(9);
			42773: out = 16'(-94);
			42774: out = 16'(62);
			42775: out = 16'(-147);
			42776: out = 16'(-303);
			42777: out = 16'(-625);
			42778: out = 16'(-301);
			42779: out = 16'(-78);
			42780: out = 16'(112);
			42781: out = 16'(237);
			42782: out = 16'(385);
			42783: out = 16'(687);
			42784: out = 16'(582);
			42785: out = 16'(391);
			42786: out = 16'(-74);
			42787: out = 16'(-173);
			42788: out = 16'(-99);
			42789: out = 16'(23);
			42790: out = 16'(90);
			42791: out = 16'(47);
			42792: out = 16'(55);
			42793: out = 16'(-75);
			42794: out = 16'(-195);
			42795: out = 16'(-70);
			42796: out = 16'(20);
			42797: out = 16'(-185);
			42798: out = 16'(14);
			42799: out = 16'(-93);
			42800: out = 16'(-117);
			42801: out = 16'(-885);
			42802: out = 16'(-1392);
			42803: out = 16'(-1544);
			42804: out = 16'(-931);
			42805: out = 16'(-215);
			42806: out = 16'(-168);
			42807: out = 16'(-243);
			42808: out = 16'(-574);
			42809: out = 16'(-67);
			42810: out = 16'(-46);
			42811: out = 16'(-1);
			42812: out = 16'(117);
			42813: out = 16'(365);
			42814: out = 16'(794);
			42815: out = 16'(265);
			42816: out = 16'(17);
			42817: out = 16'(-127);
			42818: out = 16'(72);
			42819: out = 16'(109);
			42820: out = 16'(-102);
			42821: out = 16'(-276);
			42822: out = 16'(-218);
			42823: out = 16'(461);
			42824: out = 16'(852);
			42825: out = 16'(1100);
			42826: out = 16'(924);
			42827: out = 16'(627);
			42828: out = 16'(240);
			42829: out = 16'(72);
			42830: out = 16'(-46);
			42831: out = 16'(-172);
			42832: out = 16'(24);
			42833: out = 16'(-286);
			42834: out = 16'(-1107);
			42835: out = 16'(-952);
			42836: out = 16'(-560);
			42837: out = 16'(293);
			42838: out = 16'(571);
			42839: out = 16'(586);
			42840: out = 16'(-114);
			42841: out = 16'(-533);
			42842: out = 16'(-899);
			42843: out = 16'(-1039);
			42844: out = 16'(-950);
			42845: out = 16'(-739);
			42846: out = 16'(-210);
			42847: out = 16'(-161);
			42848: out = 16'(-341);
			42849: out = 16'(-179);
			42850: out = 16'(135);
			42851: out = 16'(607);
			42852: out = 16'(827);
			42853: out = 16'(910);
			42854: out = 16'(714);
			42855: out = 16'(351);
			42856: out = 16'(-48);
			42857: out = 16'(-329);
			42858: out = 16'(-415);
			42859: out = 16'(-304);
			42860: out = 16'(13);
			42861: out = 16'(115);
			42862: out = 16'(134);
			42863: out = 16'(288);
			42864: out = 16'(335);
			42865: out = 16'(287);
			42866: out = 16'(328);
			42867: out = 16'(147);
			42868: out = 16'(-159);
			42869: out = 16'(-491);
			42870: out = 16'(-650);
			42871: out = 16'(-581);
			42872: out = 16'(-307);
			42873: out = 16'(-62);
			42874: out = 16'(25);
			42875: out = 16'(-23);
			42876: out = 16'(-298);
			42877: out = 16'(-737);
			42878: out = 16'(-847);
			42879: out = 16'(-654);
			42880: out = 16'(-154);
			42881: out = 16'(383);
			42882: out = 16'(776);
			42883: out = 16'(590);
			42884: out = 16'(371);
			42885: out = 16'(96);
			42886: out = 16'(-42);
			42887: out = 16'(-106);
			42888: out = 16'(-149);
			42889: out = 16'(27);
			42890: out = 16'(44);
			42891: out = 16'(69);
			42892: out = 16'(-101);
			42893: out = 16'(-115);
			42894: out = 16'(-112);
			42895: out = 16'(614);
			42896: out = 16'(1210);
			42897: out = 16'(1366);
			42898: out = 16'(1056);
			42899: out = 16'(490);
			42900: out = 16'(165);
			42901: out = 16'(-147);
			42902: out = 16'(-286);
			42903: out = 16'(-1425);
			42904: out = 16'(-1483);
			42905: out = 16'(-991);
			42906: out = 16'(-770);
			42907: out = 16'(-379);
			42908: out = 16'(-189);
			42909: out = 16'(249);
			42910: out = 16'(267);
			42911: out = 16'(103);
			42912: out = 16'(-793);
			42913: out = 16'(-1337);
			42914: out = 16'(-964);
			42915: out = 16'(-1028);
			42916: out = 16'(-939);
			42917: out = 16'(-977);
			42918: out = 16'(-615);
			42919: out = 16'(-145);
			42920: out = 16'(-100);
			42921: out = 16'(665);
			42922: out = 16'(1455);
			42923: out = 16'(1356);
			42924: out = 16'(1135);
			42925: out = 16'(717);
			42926: out = 16'(257);
			42927: out = 16'(37);
			42928: out = 16'(166);
			42929: out = 16'(-39);
			42930: out = 16'(-65);
			42931: out = 16'(101);
			42932: out = 16'(-236);
			42933: out = 16'(-339);
			42934: out = 16'(-429);
			42935: out = 16'(361);
			42936: out = 16'(1025);
			42937: out = 16'(1059);
			42938: out = 16'(572);
			42939: out = 16'(-272);
			42940: out = 16'(166);
			42941: out = 16'(-79);
			42942: out = 16'(-85);
			42943: out = 16'(-770);
			42944: out = 16'(-614);
			42945: out = 16'(-168);
			42946: out = 16'(21);
			42947: out = 16'(-168);
			42948: out = 16'(-818);
			42949: out = 16'(-984);
			42950: out = 16'(-855);
			42951: out = 16'(-57);
			42952: out = 16'(188);
			42953: out = 16'(351);
			42954: out = 16'(-121);
			42955: out = 16'(-311);
			42956: out = 16'(-588);
			42957: out = 16'(-99);
			42958: out = 16'(-70);
			42959: out = 16'(144);
			42960: out = 16'(-717);
			42961: out = 16'(-415);
			42962: out = 16'(160);
			42963: out = 16'(933);
			42964: out = 16'(1177);
			42965: out = 16'(1110);
			42966: out = 16'(413);
			42967: out = 16'(40);
			42968: out = 16'(45);
			42969: out = 16'(343);
			42970: out = 16'(503);
			42971: out = 16'(315);
			42972: out = 16'(-324);
			42973: out = 16'(-979);
			42974: out = 16'(-988);
			42975: out = 16'(-900);
			42976: out = 16'(-433);
			42977: out = 16'(-200);
			42978: out = 16'(182);
			42979: out = 16'(318);
			42980: out = 16'(398);
			42981: out = 16'(166);
			42982: out = 16'(-69);
			42983: out = 16'(-296);
			42984: out = 16'(-306);
			42985: out = 16'(-146);
			42986: out = 16'(26);
			42987: out = 16'(-34);
			42988: out = 16'(-583);
			42989: out = 16'(-450);
			42990: out = 16'(-205);
			42991: out = 16'(333);
			42992: out = 16'(477);
			42993: out = 16'(517);
			42994: out = 16'(173);
			42995: out = 16'(103);
			42996: out = 16'(43);
			42997: out = 16'(-124);
			42998: out = 16'(-119);
			42999: out = 16'(-73);
			43000: out = 16'(-72);
			43001: out = 16'(-167);
			43002: out = 16'(-360);
			43003: out = 16'(-54);
			43004: out = 16'(272);
			43005: out = 16'(730);
			43006: out = 16'(606);
			43007: out = 16'(371);
			43008: out = 16'(-90);
			43009: out = 16'(-108);
			43010: out = 16'(-78);
			43011: out = 16'(26);
			43012: out = 16'(-61);
			43013: out = 16'(-202);
			43014: out = 16'(-60);
			43015: out = 16'(-234);
			43016: out = 16'(-408);
			43017: out = 16'(-962);
			43018: out = 16'(-815);
			43019: out = 16'(-274);
			43020: out = 16'(-56);
			43021: out = 16'(176);
			43022: out = 16'(106);
			43023: out = 16'(466);
			43024: out = 16'(463);
			43025: out = 16'(103);
			43026: out = 16'(-4);
			43027: out = 16'(-241);
			43028: out = 16'(-299);
			43029: out = 16'(-621);
			43030: out = 16'(-755);
			43031: out = 16'(-599);
			43032: out = 16'(-177);
			43033: out = 16'(282);
			43034: out = 16'(664);
			43035: out = 16'(879);
			43036: out = 16'(897);
			43037: out = 16'(776);
			43038: out = 16'(503);
			43039: out = 16'(45);
			43040: out = 16'(-14);
			43041: out = 16'(-275);
			43042: out = 16'(-574);
			43043: out = 16'(-792);
			43044: out = 16'(-645);
			43045: out = 16'(-103);
			43046: out = 16'(423);
			43047: out = 16'(754);
			43048: out = 16'(520);
			43049: out = 16'(311);
			43050: out = 16'(-3);
			43051: out = 16'(-518);
			43052: out = 16'(-633);
			43053: out = 16'(-540);
			43054: out = 16'(-157);
			43055: out = 16'(-56);
			43056: out = 16'(-84);
			43057: out = 16'(56);
			43058: out = 16'(82);
			43059: out = 16'(62);
			43060: out = 16'(252);
			43061: out = 16'(382);
			43062: out = 16'(524);
			43063: out = 16'(377);
			43064: out = 16'(256);
			43065: out = 16'(74);
			43066: out = 16'(115);
			43067: out = 16'(44);
			43068: out = 16'(78);
			43069: out = 16'(-535);
			43070: out = 16'(-1141);
			43071: out = 16'(-1047);
			43072: out = 16'(-779);
			43073: out = 16'(-247);
			43074: out = 16'(-53);
			43075: out = 16'(186);
			43076: out = 16'(104);
			43077: out = 16'(487);
			43078: out = 16'(527);
			43079: out = 16'(542);
			43080: out = 16'(87);
			43081: out = 16'(-176);
			43082: out = 16'(-368);
			43083: out = 16'(-503);
			43084: out = 16'(-595);
			43085: out = 16'(-286);
			43086: out = 16'(-740);
			43087: out = 16'(-1022);
			43088: out = 16'(-1019);
			43089: out = 16'(-529);
			43090: out = 16'(86);
			43091: out = 16'(327);
			43092: out = 16'(277);
			43093: out = 16'(-131);
			43094: out = 16'(119);
			43095: out = 16'(171);
			43096: out = 16'(435);
			43097: out = 16'(19);
			43098: out = 16'(-155);
			43099: out = 16'(-334);
			43100: out = 16'(146);
			43101: out = 16'(445);
			43102: out = 16'(325);
			43103: out = 16'(394);
			43104: out = 16'(345);
			43105: out = 16'(599);
			43106: out = 16'(268);
			43107: out = 16'(41);
			43108: out = 16'(-84);
			43109: out = 16'(187);
			43110: out = 16'(496);
			43111: out = 16'(-178);
			43112: out = 16'(-761);
			43113: out = 16'(-1294);
			43114: out = 16'(-1131);
			43115: out = 16'(-714);
			43116: out = 16'(-93);
			43117: out = 16'(393);
			43118: out = 16'(638);
			43119: out = 16'(754);
			43120: out = 16'(369);
			43121: out = 16'(124);
			43122: out = 16'(336);
			43123: out = 16'(433);
			43124: out = 16'(484);
			43125: out = 16'(108);
			43126: out = 16'(-390);
			43127: out = 16'(-867);
			43128: out = 16'(-403);
			43129: out = 16'(-178);
			43130: out = 16'(218);
			43131: out = 16'(384);
			43132: out = 16'(708);
			43133: out = 16'(863);
			43134: out = 16'(920);
			43135: out = 16'(633);
			43136: out = 16'(37);
			43137: out = 16'(-102);
			43138: out = 16'(-296);
			43139: out = 16'(-419);
			43140: out = 16'(-332);
			43141: out = 16'(-114);
			43142: out = 16'(25);
			43143: out = 16'(307);
			43144: out = 16'(427);
			43145: out = 16'(-91);
			43146: out = 16'(-192);
			43147: out = 16'(-199);
			43148: out = 16'(-26);
			43149: out = 16'(-34);
			43150: out = 16'(-155);
			43151: out = 16'(-6);
			43152: out = 16'(-71);
			43153: out = 16'(-212);
			43154: out = 16'(-511);
			43155: out = 16'(-763);
			43156: out = 16'(-1075);
			43157: out = 16'(-783);
			43158: out = 16'(-357);
			43159: out = 16'(539);
			43160: out = 16'(300);
			43161: out = 16'(64);
			43162: out = 16'(-140);
			43163: out = 16'(-27);
			43164: out = 16'(140);
			43165: out = 16'(-90);
			43166: out = 16'(-100);
			43167: out = 16'(-86);
			43168: out = 16'(-94);
			43169: out = 16'(-36);
			43170: out = 16'(60);
			43171: out = 16'(-44);
			43172: out = 16'(-107);
			43173: out = 16'(-76);
			43174: out = 16'(-156);
			43175: out = 16'(-75);
			43176: out = 16'(96);
			43177: out = 16'(509);
			43178: out = 16'(680);
			43179: out = 16'(297);
			43180: out = 16'(-44);
			43181: out = 16'(-535);
			43182: out = 16'(-733);
			43183: out = 16'(-900);
			43184: out = 16'(-728);
			43185: out = 16'(-689);
			43186: out = 16'(-284);
			43187: out = 16'(-68);
			43188: out = 16'(361);
			43189: out = 16'(107);
			43190: out = 16'(-312);
			43191: out = 16'(-731);
			43192: out = 16'(-463);
			43193: out = 16'(377);
			43194: out = 16'(802);
			43195: out = 16'(820);
			43196: out = 16'(381);
			43197: out = 16'(-338);
			43198: out = 16'(-846);
			43199: out = 16'(-575);
			43200: out = 16'(2);
			43201: out = 16'(681);
			43202: out = 16'(499);
			43203: out = 16'(327);
			43204: out = 16'(-166);
			43205: out = 16'(177);
			43206: out = 16'(0);
			43207: out = 16'(-53);
			43208: out = 16'(-349);
			43209: out = 16'(-205);
			43210: out = 16'(160);
			43211: out = 16'(-31);
			43212: out = 16'(-57);
			43213: out = 16'(98);
			43214: out = 16'(51);
			43215: out = 16'(88);
			43216: out = 16'(52);
			43217: out = 16'(16);
			43218: out = 16'(-71);
			43219: out = 16'(358);
			43220: out = 16'(74);
			43221: out = 16'(-210);
			43222: out = 16'(-755);
			43223: out = 16'(-528);
			43224: out = 16'(-89);
			43225: out = 16'(-297);
			43226: out = 16'(-551);
			43227: out = 16'(-1032);
			43228: out = 16'(-630);
			43229: out = 16'(-355);
			43230: out = 16'(18);
			43231: out = 16'(273);
			43232: out = 16'(398);
			43233: out = 16'(158);
			43234: out = 16'(213);
			43235: out = 16'(153);
			43236: out = 16'(199);
			43237: out = 16'(135);
			43238: out = 16'(60);
			43239: out = 16'(-529);
			43240: out = 16'(-337);
			43241: out = 16'(-14);
			43242: out = 16'(658);
			43243: out = 16'(720);
			43244: out = 16'(515);
			43245: out = 16'(59);
			43246: out = 16'(-121);
			43247: out = 16'(-110);
			43248: out = 16'(8);
			43249: out = 16'(81);
			43250: out = 16'(-95);
			43251: out = 16'(-70);
			43252: out = 16'(-276);
			43253: out = 16'(-759);
			43254: out = 16'(-553);
			43255: out = 16'(-124);
			43256: out = 16'(459);
			43257: out = 16'(897);
			43258: out = 16'(1122);
			43259: out = 16'(1123);
			43260: out = 16'(823);
			43261: out = 16'(419);
			43262: out = 16'(-21);
			43263: out = 16'(-108);
			43264: out = 16'(109);
			43265: out = 16'(-475);
			43266: out = 16'(-846);
			43267: out = 16'(-1318);
			43268: out = 16'(-508);
			43269: out = 16'(66);
			43270: out = 16'(283);
			43271: out = 16'(368);
			43272: out = 16'(233);
			43273: out = 16'(122);
			43274: out = 16'(-464);
			43275: out = 16'(-799);
			43276: out = 16'(-382);
			43277: out = 16'(-131);
			43278: out = 16'(188);
			43279: out = 16'(60);
			43280: out = 16'(87);
			43281: out = 16'(50);
			43282: out = 16'(319);
			43283: out = 16'(199);
			43284: out = 16'(-126);
			43285: out = 16'(-87);
			43286: out = 16'(-304);
			43287: out = 16'(-583);
			43288: out = 16'(-448);
			43289: out = 16'(-210);
			43290: out = 16'(119);
			43291: out = 16'(299);
			43292: out = 16'(269);
			43293: out = 16'(-42);
			43294: out = 16'(-223);
			43295: out = 16'(-366);
			43296: out = 16'(-574);
			43297: out = 16'(-339);
			43298: out = 16'(-2);
			43299: out = 16'(290);
			43300: out = 16'(297);
			43301: out = 16'(123);
			43302: out = 16'(93);
			43303: out = 16'(3);
			43304: out = 16'(-156);
			43305: out = 16'(90);
			43306: out = 16'(73);
			43307: out = 16'(-45);
			43308: out = 16'(-696);
			43309: out = 16'(-1088);
			43310: out = 16'(-978);
			43311: out = 16'(-640);
			43312: out = 16'(-183);
			43313: out = 16'(-60);
			43314: out = 16'(9);
			43315: out = 16'(-16);
			43316: out = 16'(143);
			43317: out = 16'(61);
			43318: out = 16'(-7);
			43319: out = 16'(334);
			43320: out = 16'(271);
			43321: out = 16'(-56);
			43322: out = 16'(-60);
			43323: out = 16'(-176);
			43324: out = 16'(-302);
			43325: out = 16'(-126);
			43326: out = 16'(197);
			43327: out = 16'(978);
			43328: out = 16'(714);
			43329: out = 16'(428);
			43330: out = 16'(-342);
			43331: out = 16'(-120);
			43332: out = 16'(162);
			43333: out = 16'(717);
			43334: out = 16'(366);
			43335: out = 16'(-198);
			43336: out = 16'(-887);
			43337: out = 16'(-994);
			43338: out = 16'(-705);
			43339: out = 16'(-206);
			43340: out = 16'(85);
			43341: out = 16'(161);
			43342: out = 16'(-21);
			43343: out = 16'(-56);
			43344: out = 16'(202);
			43345: out = 16'(134);
			43346: out = 16'(-86);
			43347: out = 16'(-1011);
			43348: out = 16'(-851);
			43349: out = 16'(-593);
			43350: out = 16'(166);
			43351: out = 16'(206);
			43352: out = 16'(195);
			43353: out = 16'(153);
			43354: out = 16'(71);
			43355: out = 16'(-26);
			43356: out = 16'(-15);
			43357: out = 16'(-34);
			43358: out = 16'(-3);
			43359: out = 16'(130);
			43360: out = 16'(310);
			43361: out = 16'(590);
			43362: out = 16'(439);
			43363: out = 16'(244);
			43364: out = 16'(-57);
			43365: out = 16'(181);
			43366: out = 16'(493);
			43367: out = 16'(859);
			43368: out = 16'(950);
			43369: out = 16'(746);
			43370: out = 16'(-18);
			43371: out = 16'(-301);
			43372: out = 16'(-356);
			43373: out = 16'(-188);
			43374: out = 16'(96);
			43375: out = 16'(275);
			43376: out = 16'(142);
			43377: out = 16'(-302);
			43378: out = 16'(-842);
			43379: out = 16'(-1035);
			43380: out = 16'(-918);
			43381: out = 16'(-581);
			43382: out = 16'(-82);
			43383: out = 16'(67);
			43384: out = 16'(-101);
			43385: out = 16'(-528);
			43386: out = 16'(-772);
			43387: out = 16'(-563);
			43388: out = 16'(-172);
			43389: out = 16'(232);
			43390: out = 16'(737);
			43391: out = 16'(597);
			43392: out = 16'(297);
			43393: out = 16'(-640);
			43394: out = 16'(-472);
			43395: out = 16'(181);
			43396: out = 16'(468);
			43397: out = 16'(455);
			43398: out = 16'(58);
			43399: out = 16'(-395);
			43400: out = 16'(-443);
			43401: out = 16'(122);
			43402: out = 16'(269);
			43403: out = 16'(307);
			43404: out = 16'(-61);
			43405: out = 16'(-322);
			43406: out = 16'(-583);
			43407: out = 16'(-333);
			43408: out = 16'(-90);
			43409: out = 16'(237);
			43410: out = 16'(131);
			43411: out = 16'(175);
			43412: out = 16'(39);
			43413: out = 16'(-201);
			43414: out = 16'(-417);
			43415: out = 16'(-464);
			43416: out = 16'(-339);
			43417: out = 16'(-250);
			43418: out = 16'(-293);
			43419: out = 16'(-242);
			43420: out = 16'(-231);
			43421: out = 16'(-39);
			43422: out = 16'(-197);
			43423: out = 16'(-263);
			43424: out = 16'(-484);
			43425: out = 16'(25);
			43426: out = 16'(440);
			43427: out = 16'(333);
			43428: out = 16'(289);
			43429: out = 16'(80);
			43430: out = 16'(349);
			43431: out = 16'(315);
			43432: out = 16'(345);
			43433: out = 16'(-202);
			43434: out = 16'(-164);
			43435: out = 16'(120);
			43436: out = 16'(499);
			43437: out = 16'(801);
			43438: out = 16'(952);
			43439: out = 16'(777);
			43440: out = 16'(453);
			43441: out = 16'(111);
			43442: out = 16'(-62);
			43443: out = 16'(-52);
			43444: out = 16'(238);
			43445: out = 16'(166);
			43446: out = 16'(-4);
			43447: out = 16'(-478);
			43448: out = 16'(-587);
			43449: out = 16'(-519);
			43450: out = 16'(-726);
			43451: out = 16'(-757);
			43452: out = 16'(-917);
			43453: out = 16'(-189);
			43454: out = 16'(19);
			43455: out = 16'(110);
			43456: out = 16'(-496);
			43457: out = 16'(-524);
			43458: out = 16'(135);
			43459: out = 16'(124);
			43460: out = 16'(159);
			43461: out = 16'(89);
			43462: out = 16'(91);
			43463: out = 16'(124);
			43464: out = 16'(287);
			43465: out = 16'(496);
			43466: out = 16'(600);
			43467: out = 16'(216);
			43468: out = 16'(-344);
			43469: out = 16'(-952);
			43470: out = 16'(-563);
			43471: out = 16'(-274);
			43472: out = 16'(190);
			43473: out = 16'(93);
			43474: out = 16'(180);
			43475: out = 16'(101);
			43476: out = 16'(630);
			43477: out = 16'(848);
			43478: out = 16'(782);
			43479: out = 16'(593);
			43480: out = 16'(315);
			43481: out = 16'(-61);
			43482: out = 16'(-261);
			43483: out = 16'(-379);
			43484: out = 16'(-520);
			43485: out = 16'(-532);
			43486: out = 16'(-521);
			43487: out = 16'(-502);
			43488: out = 16'(-513);
			43489: out = 16'(-482);
			43490: out = 16'(-628);
			43491: out = 16'(-737);
			43492: out = 16'(-847);
			43493: out = 16'(-407);
			43494: out = 16'(-154);
			43495: out = 16'(-47);
			43496: out = 16'(-46);
			43497: out = 16'(-17);
			43498: out = 16'(140);
			43499: out = 16'(270);
			43500: out = 16'(400);
			43501: out = 16'(316);
			43502: out = 16'(369);
			43503: out = 16'(320);
			43504: out = 16'(529);
			43505: out = 16'(323);
			43506: out = 16'(112);
			43507: out = 16'(-39);
			43508: out = 16'(77);
			43509: out = 16'(318);
			43510: out = 16'(0);
			43511: out = 16'(-426);
			43512: out = 16'(-1123);
			43513: out = 16'(-665);
			43514: out = 16'(-234);
			43515: out = 16'(332);
			43516: out = 16'(347);
			43517: out = 16'(300);
			43518: out = 16'(107);
			43519: out = 16'(69);
			43520: out = 16'(145);
			43521: out = 16'(458);
			43522: out = 16'(500);
			43523: out = 16'(372);
			43524: out = 16'(-332);
			43525: out = 16'(-810);
			43526: out = 16'(-1060);
			43527: out = 16'(-307);
			43528: out = 16'(121);
			43529: out = 16'(289);
			43530: out = 16'(379);
			43531: out = 16'(171);
			43532: out = 16'(-67);
			43533: out = 16'(-679);
			43534: out = 16'(-707);
			43535: out = 16'(90);
			43536: out = 16'(536);
			43537: out = 16'(922);
			43538: out = 16'(955);
			43539: out = 16'(737);
			43540: out = 16'(345);
			43541: out = 16'(115);
			43542: out = 16'(-174);
			43543: out = 16'(-325);
			43544: out = 16'(-10);
			43545: out = 16'(0);
			43546: out = 16'(-106);
			43547: out = 16'(21);
			43548: out = 16'(8);
			43549: out = 16'(-118);
			43550: out = 16'(72);
			43551: out = 16'(23);
			43552: out = 16'(-136);
			43553: out = 16'(-509);
			43554: out = 16'(-829);
			43555: out = 16'(-1086);
			43556: out = 16'(-1106);
			43557: out = 16'(-1008);
			43558: out = 16'(-459);
			43559: out = 16'(-466);
			43560: out = 16'(-402);
			43561: out = 16'(-877);
			43562: out = 16'(-288);
			43563: out = 16'(467);
			43564: out = 16'(835);
			43565: out = 16'(582);
			43566: out = 16'(-128);
			43567: out = 16'(-342);
			43568: out = 16'(-344);
			43569: out = 16'(193);
			43570: out = 16'(238);
			43571: out = 16'(467);
			43572: out = 16'(659);
			43573: out = 16'(598);
			43574: out = 16'(463);
			43575: out = 16'(491);
			43576: out = 16'(646);
			43577: out = 16'(763);
			43578: out = 16'(100);
			43579: out = 16'(21);
			43580: out = 16'(-155);
			43581: out = 16'(-65);
			43582: out = 16'(-580);
			43583: out = 16'(-1164);
			43584: out = 16'(-642);
			43585: out = 16'(-156);
			43586: out = 16'(543);
			43587: out = 16'(152);
			43588: out = 16'(-18);
			43589: out = 16'(-353);
			43590: out = 16'(16);
			43591: out = 16'(128);
			43592: out = 16'(126);
			43593: out = 16'(0);
			43594: out = 16'(-95);
			43595: out = 16'(-307);
			43596: out = 16'(-118);
			43597: out = 16'(155);
			43598: out = 16'(776);
			43599: out = 16'(508);
			43600: out = 16'(-10);
			43601: out = 16'(-738);
			43602: out = 16'(-852);
			43603: out = 16'(-402);
			43604: out = 16'(-217);
			43605: out = 16'(189);
			43606: out = 16'(455);
			43607: out = 16'(647);
			43608: out = 16'(484);
			43609: out = 16'(105);
			43610: out = 16'(-53);
			43611: out = 16'(-187);
			43612: out = 16'(-335);
			43613: out = 16'(-181);
			43614: out = 16'(-26);
			43615: out = 16'(267);
			43616: out = 16'(109);
			43617: out = 16'(-99);
			43618: out = 16'(51);
			43619: out = 16'(31);
			43620: out = 16'(16);
			43621: out = 16'(-257);
			43622: out = 16'(-368);
			43623: out = 16'(-318);
			43624: out = 16'(-771);
			43625: out = 16'(-1027);
			43626: out = 16'(-1337);
			43627: out = 16'(-829);
			43628: out = 16'(-562);
			43629: out = 16'(-432);
			43630: out = 16'(-437);
			43631: out = 16'(-318);
			43632: out = 16'(-11);
			43633: out = 16'(439);
			43634: out = 16'(777);
			43635: out = 16'(713);
			43636: out = 16'(390);
			43637: out = 16'(-77);
			43638: out = 16'(162);
			43639: out = 16'(37);
			43640: out = 16'(-4);
			43641: out = 16'(112);
			43642: out = 16'(237);
			43643: out = 16'(334);
			43644: out = 16'(452);
			43645: out = 16'(558);
			43646: out = 16'(644);
			43647: out = 16'(427);
			43648: out = 16'(190);
			43649: out = 16'(99);
			43650: out = 16'(-434);
			43651: out = 16'(-782);
			43652: out = 16'(-897);
			43653: out = 16'(-604);
			43654: out = 16'(-187);
			43655: out = 16'(-95);
			43656: out = 16'(100);
			43657: out = 16'(120);
			43658: out = 16'(179);
			43659: out = 16'(46);
			43660: out = 16'(-90);
			43661: out = 16'(-262);
			43662: out = 16'(-199);
			43663: out = 16'(-15);
			43664: out = 16'(-35);
			43665: out = 16'(-258);
			43666: out = 16'(-878);
			43667: out = 16'(-702);
			43668: out = 16'(-484);
			43669: out = 16'(152);
			43670: out = 16'(121);
			43671: out = 16'(162);
			43672: out = 16'(-19);
			43673: out = 16'(369);
			43674: out = 16'(764);
			43675: out = 16'(832);
			43676: out = 16'(787);
			43677: out = 16'(604);
			43678: out = 16'(233);
			43679: out = 16'(29);
			43680: out = 16'(-76);
			43681: out = 16'(-53);
			43682: out = 16'(-128);
			43683: out = 16'(-309);
			43684: out = 16'(-307);
			43685: out = 16'(-200);
			43686: out = 16'(130);
			43687: out = 16'(139);
			43688: out = 16'(116);
			43689: out = 16'(88);
			43690: out = 16'(-32);
			43691: out = 16'(-227);
			43692: out = 16'(-1035);
			43693: out = 16'(-1084);
			43694: out = 16'(-1002);
			43695: out = 16'(-169);
			43696: out = 16'(-184);
			43697: out = 16'(-452);
			43698: out = 16'(-442);
			43699: out = 16'(-193);
			43700: out = 16'(249);
			43701: out = 16'(552);
			43702: out = 16'(814);
			43703: out = 16'(840);
			43704: out = 16'(560);
			43705: out = 16'(86);
			43706: out = 16'(-638);
			43707: out = 16'(-459);
			43708: out = 16'(-162);
			43709: out = 16'(-71);
			43710: out = 16'(1);
			43711: out = 16'(-87);
			43712: out = 16'(141);
			43713: out = 16'(109);
			43714: out = 16'(197);
			43715: out = 16'(113);
			43716: out = 16'(380);
			43717: out = 16'(660);
			43718: out = 16'(692);
			43719: out = 16'(453);
			43720: out = 16'(59);
			43721: out = 16'(-498);
			43722: out = 16'(-651);
			43723: out = 16'(-286);
			43724: out = 16'(-61);
			43725: out = 16'(54);
			43726: out = 16'(-308);
			43727: out = 16'(-281);
			43728: out = 16'(-267);
			43729: out = 16'(-101);
			43730: out = 16'(-61);
			43731: out = 16'(24);
			43732: out = 16'(594);
			43733: out = 16'(539);
			43734: out = 16'(251);
			43735: out = 16'(-11);
			43736: out = 16'(-154);
			43737: out = 16'(-103);
			43738: out = 16'(-258);
			43739: out = 16'(-304);
			43740: out = 16'(-295);
			43741: out = 16'(-181);
			43742: out = 16'(-46);
			43743: out = 16'(-69);
			43744: out = 16'(410);
			43745: out = 16'(694);
			43746: out = 16'(626);
			43747: out = 16'(352);
			43748: out = 16'(-23);
			43749: out = 16'(85);
			43750: out = 16'(-10);
			43751: out = 16'(41);
			43752: out = 16'(-496);
			43753: out = 16'(-380);
			43754: out = 16'(-110);
			43755: out = 16'(208);
			43756: out = 16'(301);
			43757: out = 16'(274);
			43758: out = 16'(0);
			43759: out = 16'(-71);
			43760: out = 16'(44);
			43761: out = 16'(44);
			43762: out = 16'(-51);
			43763: out = 16'(-309);
			43764: out = 16'(-793);
			43765: out = 16'(-1220);
			43766: out = 16'(-1255);
			43767: out = 16'(-1237);
			43768: out = 16'(-891);
			43769: out = 16'(-50);
			43770: out = 16'(524);
			43771: out = 16'(898);
			43772: out = 16'(866);
			43773: out = 16'(664);
			43774: out = 16'(255);
			43775: out = 16'(227);
			43776: out = 16'(27);
			43777: out = 16'(-31);
			43778: out = 16'(-522);
			43779: out = 16'(-706);
			43780: out = 16'(-679);
			43781: out = 16'(-181);
			43782: out = 16'(203);
			43783: out = 16'(312);
			43784: out = 16'(334);
			43785: out = 16'(316);
			43786: out = 16'(132);
			43787: out = 16'(232);
			43788: out = 16'(292);
			43789: out = 16'(348);
			43790: out = 16'(88);
			43791: out = 16'(-144);
			43792: out = 16'(-971);
			43793: out = 16'(-761);
			43794: out = 16'(179);
			43795: out = 16'(486);
			43796: out = 16'(600);
			43797: out = 16'(55);
			43798: out = 16'(48);
			43799: out = 16'(-139);
			43800: out = 16'(0);
			43801: out = 16'(-259);
			43802: out = 16'(-230);
			43803: out = 16'(12);
			43804: out = 16'(320);
			43805: out = 16'(435);
			43806: out = 16'(-10);
			43807: out = 16'(-286);
			43808: out = 16'(-548);
			43809: out = 16'(-669);
			43810: out = 16'(-556);
			43811: out = 16'(-213);
			43812: out = 16'(151);
			43813: out = 16'(539);
			43814: out = 16'(814);
			43815: out = 16'(705);
			43816: out = 16'(556);
			43817: out = 16'(468);
			43818: out = 16'(168);
			43819: out = 16'(-130);
			43820: out = 16'(-738);
			43821: out = 16'(-502);
			43822: out = 16'(-266);
			43823: out = 16'(-110);
			43824: out = 16'(8);
			43825: out = 16'(53);
			43826: out = 16'(-127);
			43827: out = 16'(-52);
			43828: out = 16'(58);
			43829: out = 16'(-58);
			43830: out = 16'(-36);
			43831: out = 16'(72);
			43832: out = 16'(-273);
			43833: out = 16'(-248);
			43834: out = 16'(-73);
			43835: out = 16'(39);
			43836: out = 16'(-143);
			43837: out = 16'(-917);
			43838: out = 16'(-795);
			43839: out = 16'(-440);
			43840: out = 16'(621);
			43841: out = 16'(857);
			43842: out = 16'(952);
			43843: out = 16'(491);
			43844: out = 16'(206);
			43845: out = 16'(-131);
			43846: out = 16'(453);
			43847: out = 16'(240);
			43848: out = 16'(-7);
			43849: out = 16'(-783);
			43850: out = 16'(-891);
			43851: out = 16'(-692);
			43852: out = 16'(-278);
			43853: out = 16'(-41);
			43854: out = 16'(71);
			43855: out = 16'(-69);
			43856: out = 16'(-32);
			43857: out = 16'(289);
			43858: out = 16'(417);
			43859: out = 16'(357);
			43860: out = 16'(-269);
			43861: out = 16'(-635);
			43862: out = 16'(-921);
			43863: out = 16'(-511);
			43864: out = 16'(-327);
			43865: out = 16'(-38);
			43866: out = 16'(33);
			43867: out = 16'(129);
			43868: out = 16'(53);
			43869: out = 16'(-49);
			43870: out = 16'(-50);
			43871: out = 16'(192);
			43872: out = 16'(211);
			43873: out = 16'(342);
			43874: out = 16'(42);
			43875: out = 16'(529);
			43876: out = 16'(508);
			43877: out = 16'(130);
			43878: out = 16'(-662);
			43879: out = 16'(-1045);
			43880: out = 16'(-6);
			43881: out = 16'(451);
			43882: out = 16'(852);
			43883: out = 16'(615);
			43884: out = 16'(562);
			43885: out = 16'(400);
			43886: out = 16'(148);
			43887: out = 16'(20);
			43888: out = 16'(10);
			43889: out = 16'(-257);
			43890: out = 16'(-545);
			43891: out = 16'(-947);
			43892: out = 16'(-1097);
			43893: out = 16'(-909);
			43894: out = 16'(-94);
			43895: out = 16'(3);
			43896: out = 16'(70);
			43897: out = 16'(-103);
			43898: out = 16'(-102);
			43899: out = 16'(-87);
			43900: out = 16'(69);
			43901: out = 16'(38);
			43902: out = 16'(-53);
			43903: out = 16'(320);
			43904: out = 16'(46);
			43905: out = 16'(-326);
			43906: out = 16'(-627);
			43907: out = 16'(-464);
			43908: out = 16'(154);
			43909: out = 16'(356);
			43910: out = 16'(594);
			43911: out = 16'(603);
			43912: out = 16'(785);
			43913: out = 16'(740);
			43914: out = 16'(611);
			43915: out = 16'(400);
			43916: out = 16'(193);
			43917: out = 16'(268);
			43918: out = 16'(18);
			43919: out = 16'(-167);
			43920: out = 16'(-366);
			43921: out = 16'(-292);
			43922: out = 16'(-149);
			43923: out = 16'(175);
			43924: out = 16'(253);
			43925: out = 16'(234);
			43926: out = 16'(-43);
			43927: out = 16'(-152);
			43928: out = 16'(-173);
			43929: out = 16'(-169);
			43930: out = 16'(-231);
			43931: out = 16'(-336);
			43932: out = 16'(-615);
			43933: out = 16'(-690);
			43934: out = 16'(-325);
			43935: out = 16'(-216);
			43936: out = 16'(-152);
			43937: out = 16'(-325);
			43938: out = 16'(-287);
			43939: out = 16'(-300);
			43940: out = 16'(-123);
			43941: out = 16'(-50);
			43942: out = 16'(116);
			43943: out = 16'(508);
			43944: out = 16'(851);
			43945: out = 16'(1093);
			43946: out = 16'(633);
			43947: out = 16'(163);
			43948: out = 16'(-373);
			43949: out = 16'(-249);
			43950: out = 16'(-101);
			43951: out = 16'(-6);
			43952: out = 16'(160);
			43953: out = 16'(331);
			43954: out = 16'(914);
			43955: out = 16'(712);
			43956: out = 16'(481);
			43957: out = 16'(46);
			43958: out = 16'(32);
			43959: out = 16'(-44);
			43960: out = 16'(-462);
			43961: out = 16'(-1017);
			43962: out = 16'(-1618);
			43963: out = 16'(-1574);
			43964: out = 16'(-1520);
			43965: out = 16'(-1516);
			43966: out = 16'(-469);
			43967: out = 16'(113);
			43968: out = 16'(341);
			43969: out = 16'(85);
			43970: out = 16'(-34);
			43971: out = 16'(-42);
			43972: out = 16'(215);
			43973: out = 16'(245);
			43974: out = 16'(-198);
			43975: out = 16'(-795);
			43976: out = 16'(-1298);
			43977: out = 16'(-897);
			43978: out = 16'(-461);
			43979: out = 16'(131);
			43980: out = 16'(864);
			43981: out = 16'(993);
			43982: out = 16'(619);
			43983: out = 16'(457);
			43984: out = 16'(314);
			43985: out = 16'(544);
			43986: out = 16'(86);
			43987: out = 16'(-124);
			43988: out = 16'(-294);
			43989: out = 16'(-182);
			43990: out = 16'(-69);
			43991: out = 16'(-77);
			43992: out = 16'(168);
			43993: out = 16'(379);
			43994: out = 16'(938);
			43995: out = 16'(741);
			43996: out = 16'(360);
			43997: out = 16'(-197);
			43998: out = 16'(-468);
			43999: out = 16'(-520);
			44000: out = 16'(-512);
			44001: out = 16'(-515);
			44002: out = 16'(-492);
			44003: out = 16'(-502);
			44004: out = 16'(-453);
			44005: out = 16'(-508);
			44006: out = 16'(-60);
			44007: out = 16'(97);
			44008: out = 16'(8);
			44009: out = 16'(-197);
			44010: out = 16'(-251);
			44011: out = 16'(-143);
			44012: out = 16'(492);
			44013: out = 16'(1078);
			44014: out = 16'(1108);
			44015: out = 16'(930);
			44016: out = 16'(513);
			44017: out = 16'(36);
			44018: out = 16'(-191);
			44019: out = 16'(-123);
			44020: out = 16'(108);
			44021: out = 16'(394);
			44022: out = 16'(565);
			44023: out = 16'(243);
			44024: out = 16'(-114);
			44025: out = 16'(-341);
			44026: out = 16'(-548);
			44027: out = 16'(-471);
			44028: out = 16'(-136);
			44029: out = 16'(-103);
			44030: out = 16'(-190);
			44031: out = 16'(-661);
			44032: out = 16'(-871);
			44033: out = 16'(-839);
			44034: out = 16'(-84);
			44035: out = 16'(280);
			44036: out = 16'(463);
			44037: out = 16'(188);
			44038: out = 16'(5);
			44039: out = 16'(-64);
			44040: out = 16'(37);
			44041: out = 16'(222);
			44042: out = 16'(429);
			44043: out = 16'(367);
			44044: out = 16'(87);
			44045: out = 16'(-290);
			44046: out = 16'(-993);
			44047: out = 16'(-1309);
			44048: out = 16'(-724);
			44049: out = 16'(-267);
			44050: out = 16'(222);
			44051: out = 16'(-75);
			44052: out = 16'(-12);
			44053: out = 16'(-35);
			44054: out = 16'(760);
			44055: out = 16'(627);
			44056: out = 16'(233);
			44057: out = 16'(17);
			44058: out = 16'(-114);
			44059: out = 16'(-63);
			44060: out = 16'(-266);
			44061: out = 16'(-373);
			44062: out = 16'(-528);
			44063: out = 16'(-125);
			44064: out = 16'(124);
			44065: out = 16'(109);
			44066: out = 16'(122);
			44067: out = 16'(108);
			44068: out = 16'(93);
			44069: out = 16'(-322);
			44070: out = 16'(-788);
			44071: out = 16'(-623);
			44072: out = 16'(-825);
			44073: out = 16'(-823);
			44074: out = 16'(-1300);
			44075: out = 16'(-851);
			44076: out = 16'(-154);
			44077: out = 16'(669);
			44078: out = 16'(812);
			44079: out = 16'(330);
			44080: out = 16'(207);
			44081: out = 16'(152);
			44082: out = 16'(366);
			44083: out = 16'(566);
			44084: out = 16'(584);
			44085: out = 16'(-35);
			44086: out = 16'(-256);
			44087: out = 16'(-591);
			44088: out = 16'(-808);
			44089: out = 16'(-722);
			44090: out = 16'(-326);
			44091: out = 16'(0);
			44092: out = 16'(302);
			44093: out = 16'(347);
			44094: out = 16'(829);
			44095: out = 16'(603);
			44096: out = 16'(128);
			44097: out = 16'(-42);
			44098: out = 16'(1);
			44099: out = 16'(342);
			44100: out = 16'(190);
			44101: out = 16'(-34);
			44102: out = 16'(-685);
			44103: out = 16'(-581);
			44104: out = 16'(-342);
			44105: out = 16'(114);
			44106: out = 16'(366);
			44107: out = 16'(486);
			44108: out = 16'(175);
			44109: out = 16'(101);
			44110: out = 16'(97);
			44111: out = 16'(106);
			44112: out = 16'(287);
			44113: out = 16'(466);
			44114: out = 16'(198);
			44115: out = 16'(-325);
			44116: out = 16'(-1143);
			44117: out = 16'(-529);
			44118: out = 16'(46);
			44119: out = 16'(848);
			44120: out = 16'(828);
			44121: out = 16'(715);
			44122: out = 16'(274);
			44123: out = 16'(152);
			44124: out = 16'(20);
			44125: out = 16'(117);
			44126: out = 16'(45);
			44127: out = 16'(17);
			44128: out = 16'(-338);
			44129: out = 16'(-187);
			44130: out = 16'(73);
			44131: out = 16'(-88);
			44132: out = 16'(-99);
			44133: out = 16'(-156);
			44134: out = 16'(-274);
			44135: out = 16'(-405);
			44136: out = 16'(-510);
			44137: out = 16'(-377);
			44138: out = 16'(-208);
			44139: out = 16'(65);
			44140: out = 16'(8);
			44141: out = 16'(-62);
			44142: out = 16'(106);
			44143: out = 16'(-140);
			44144: out = 16'(-378);
			44145: out = 16'(-627);
			44146: out = 16'(-788);
			44147: out = 16'(-824);
			44148: out = 16'(-172);
			44149: out = 16'(123);
			44150: out = 16'(409);
			44151: out = 16'(415);
			44152: out = 16'(729);
			44153: out = 16'(972);
			44154: out = 16'(1148);
			44155: out = 16'(815);
			44156: out = 16'(81);
			44157: out = 16'(-570);
			44158: out = 16'(-1060);
			44159: out = 16'(-1079);
			44160: out = 16'(-1030);
			44161: out = 16'(-728);
			44162: out = 16'(-347);
			44163: out = 16'(-5);
			44164: out = 16'(194);
			44165: out = 16'(104);
			44166: out = 16'(112);
			44167: out = 16'(121);
			44168: out = 16'(465);
			44169: out = 16'(381);
			44170: out = 16'(106);
			44171: out = 16'(-44);
			44172: out = 16'(-113);
			44173: out = 16'(-23);
			44174: out = 16'(-71);
			44175: out = 16'(21);
			44176: out = 16'(108);
			44177: out = 16'(372);
			44178: out = 16'(411);
			44179: out = 16'(-122);
			44180: out = 16'(-117);
			44181: out = 16'(-113);
			44182: out = 16'(157);
			44183: out = 16'(-98);
			44184: out = 16'(-344);
			44185: out = 16'(-673);
			44186: out = 16'(-388);
			44187: out = 16'(157);
			44188: out = 16'(83);
			44189: out = 16'(247);
			44190: out = 16'(290);
			44191: out = 16'(582);
			44192: out = 16'(634);
			44193: out = 16'(636);
			44194: out = 16'(365);
			44195: out = 16'(219);
			44196: out = 16'(273);
			44197: out = 16'(-1);
			44198: out = 16'(-302);
			44199: out = 16'(-724);
			44200: out = 16'(-753);
			44201: out = 16'(-670);
			44202: out = 16'(-180);
			44203: out = 16'(-110);
			44204: out = 16'(-153);
			44205: out = 16'(-547);
			44206: out = 16'(-643);
			44207: out = 16'(-571);
			44208: out = 16'(-211);
			44209: out = 16'(40);
			44210: out = 16'(96);
			44211: out = 16'(164);
			44212: out = 16'(-26);
			44213: out = 16'(-415);
			44214: out = 16'(-440);
			44215: out = 16'(-290);
			44216: out = 16'(137);
			44217: out = 16'(144);
			44218: out = 16'(89);
			44219: out = 16'(-219);
			44220: out = 16'(-99);
			44221: out = 16'(139);
			44222: out = 16'(-63);
			44223: out = 16'(158);
			44224: out = 16'(288);
			44225: out = 16'(719);
			44226: out = 16'(422);
			44227: out = 16'(-109);
			44228: out = 16'(-615);
			44229: out = 16'(-764);
			44230: out = 16'(-561);
			44231: out = 16'(-252);
			44232: out = 16'(20);
			44233: out = 16'(146);
			44234: out = 16'(28);
			44235: out = 16'(-45);
			44236: out = 16'(-255);
			44237: out = 16'(78);
			44238: out = 16'(374);
			44239: out = 16'(867);
			44240: out = 16'(510);
			44241: out = 16'(21);
			44242: out = 16'(-369);
			44243: out = 16'(-335);
			44244: out = 16'(-50);
			44245: out = 16'(203);
			44246: out = 16'(178);
			44247: out = 16'(-78);
			44248: out = 16'(-344);
			44249: out = 16'(-349);
			44250: out = 16'(-20);
			44251: out = 16'(461);
			44252: out = 16'(772);
			44253: out = 16'(675);
			44254: out = 16'(365);
			44255: out = 16'(-85);
			44256: out = 16'(-385);
			44257: out = 16'(-608);
			44258: out = 16'(-547);
			44259: out = 16'(-32);
			44260: out = 16'(185);
			44261: out = 16'(267);
			44262: out = 16'(498);
			44263: out = 16'(606);
			44264: out = 16'(679);
			44265: out = 16'(431);
			44266: out = 16'(244);
			44267: out = 16'(29);
			44268: out = 16'(58);
			44269: out = 16'(-56);
			44270: out = 16'(-340);
			44271: out = 16'(-459);
			44272: out = 16'(-431);
			44273: out = 16'(28);
			44274: out = 16'(-192);
			44275: out = 16'(-353);
			44276: out = 16'(-657);
			44277: out = 16'(-321);
			44278: out = 16'(92);
			44279: out = 16'(-95);
			44280: out = 16'(0);
			44281: out = 16'(18);
			44282: out = 16'(-51);
			44283: out = 16'(-109);
			44284: out = 16'(-115);
			44285: out = 16'(-415);
			44286: out = 16'(-383);
			44287: out = 16'(-96);
			44288: out = 16'(-128);
			44289: out = 16'(-61);
			44290: out = 16'(57);
			44291: out = 16'(-60);
			44292: out = 16'(-99);
			44293: out = 16'(61);
			44294: out = 16'(0);
			44295: out = 16'(-83);
			44296: out = 16'(-44);
			44297: out = 16'(-162);
			44298: out = 16'(-284);
			44299: out = 16'(-276);
			44300: out = 16'(-262);
			44301: out = 16'(-252);
			44302: out = 16'(-116);
			44303: out = 16'(-31);
			44304: out = 16'(71);
			44305: out = 16'(-22);
			44306: out = 16'(47);
			44307: out = 16'(282);
			44308: out = 16'(386);
			44309: out = 16'(321);
			44310: out = 16'(-69);
			44311: out = 16'(-50);
			44312: out = 16'(-4);
			44313: out = 16'(396);
			44314: out = 16'(241);
			44315: out = 16'(42);
			44316: out = 16'(-36);
			44317: out = 16'(-121);
			44318: out = 16'(-97);
			44319: out = 16'(-4);
			44320: out = 16'(183);
			44321: out = 16'(403);
			44322: out = 16'(512);
			44323: out = 16'(348);
			44324: out = 16'(-147);
			44325: out = 16'(-109);
			44326: out = 16'(-216);
			44327: out = 16'(-291);
			44328: out = 16'(-454);
			44329: out = 16'(-382);
			44330: out = 16'(69);
			44331: out = 16'(91);
			44332: out = 16'(50);
			44333: out = 16'(-130);
			44334: out = 16'(-51);
			44335: out = 16'(34);
			44336: out = 16'(-85);
			44337: out = 16'(-83);
			44338: out = 16'(-74);
			44339: out = 16'(26);
			44340: out = 16'(-71);
			44341: out = 16'(-342);
			44342: out = 16'(-13);
			44343: out = 16'(39);
			44344: out = 16'(92);
			44345: out = 16'(-192);
			44346: out = 16'(-302);
			44347: out = 16'(-313);
			44348: out = 16'(148);
			44349: out = 16'(470);
			44350: out = 16'(511);
			44351: out = 16'(377);
			44352: out = 16'(145);
			44353: out = 16'(-55);
			44354: out = 16'(-55);
			44355: out = 16'(93);
			44356: out = 16'(168);
			44357: out = 16'(162);
			44358: out = 16'(-67);
			44359: out = 16'(-353);
			44360: out = 16'(-667);
			44361: out = 16'(-802);
			44362: out = 16'(-601);
			44363: out = 16'(-300);
			44364: out = 16'(-92);
			44365: out = 16'(185);
			44366: out = 16'(204);
			44367: out = 16'(78);
			44368: out = 16'(-480);
			44369: out = 16'(-857);
			44370: out = 16'(-776);
			44371: out = 16'(-539);
			44372: out = 16'(-144);
			44373: out = 16'(70);
			44374: out = 16'(239);
			44375: out = 16'(266);
			44376: out = 16'(28);
			44377: out = 16'(0);
			44378: out = 16'(90);
			44379: out = 16'(109);
			44380: out = 16'(138);
			44381: out = 16'(119);
			44382: out = 16'(113);
			44383: out = 16'(131);
			44384: out = 16'(282);
			44385: out = 16'(156);
			44386: out = 16'(67);
			44387: out = 16'(-67);
			44388: out = 16'(97);
			44389: out = 16'(298);
			44390: out = 16'(213);
			44391: out = 16'(342);
			44392: out = 16'(360);
			44393: out = 16'(414);
			44394: out = 16'(148);
			44395: out = 16'(-186);
			44396: out = 16'(-437);
			44397: out = 16'(-331);
			44398: out = 16'(69);
			44399: out = 16'(3);
			44400: out = 16'(-34);
			44401: out = 16'(-341);
			44402: out = 16'(-280);
			44403: out = 16'(-316);
			44404: out = 16'(-258);
			44405: out = 16'(-406);
			44406: out = 16'(-463);
			44407: out = 16'(-629);
			44408: out = 16'(-230);
			44409: out = 16'(111);
			44410: out = 16'(-36);
			44411: out = 16'(-122);
			44412: out = 16'(-270);
			44413: out = 16'(-95);
			44414: out = 16'(-58);
			44415: out = 16'(-16);
			44416: out = 16'(210);
			44417: out = 16'(301);
			44418: out = 16'(260);
			44419: out = 16'(157);
			44420: out = 16'(120);
			44421: out = 16'(282);
			44422: out = 16'(315);
			44423: out = 16'(470);
			44424: out = 16'(491);
			44425: out = 16'(658);
			44426: out = 16'(524);
			44427: out = 16'(-24);
			44428: out = 16'(-498);
			44429: out = 16'(-863);
			44430: out = 16'(-665);
			44431: out = 16'(-451);
			44432: out = 16'(-57);
			44433: out = 16'(-33);
			44434: out = 16'(218);
			44435: out = 16'(367);
			44436: out = 16'(66);
			44437: out = 16'(-366);
			44438: out = 16'(-1003);
			44439: out = 16'(-857);
			44440: out = 16'(-695);
			44441: out = 16'(-411);
			44442: out = 16'(-510);
			44443: out = 16'(-580);
			44444: out = 16'(-542);
			44445: out = 16'(-568);
			44446: out = 16'(-443);
			44447: out = 16'(59);
			44448: out = 16'(394);
			44449: out = 16'(643);
			44450: out = 16'(201);
			44451: out = 16'(163);
			44452: out = 16'(156);
			44453: out = 16'(539);
			44454: out = 16'(474);
			44455: out = 16'(75);
			44456: out = 16'(259);
			44457: out = 16'(371);
			44458: out = 16'(753);
			44459: out = 16'(258);
			44460: out = 16'(44);
			44461: out = 16'(-109);
			44462: out = 16'(304);
			44463: out = 16'(557);
			44464: out = 16'(523);
			44465: out = 16'(247);
			44466: out = 16'(-49);
			44467: out = 16'(-142);
			44468: out = 16'(-78);
			44469: out = 16'(55);
			44470: out = 16'(-78);
			44471: out = 16'(-194);
			44472: out = 16'(-342);
			44473: out = 16'(-459);
			44474: out = 16'(-375);
			44475: out = 16'(-64);
			44476: out = 16'(-100);
			44477: out = 16'(-117);
			44478: out = 16'(-300);
			44479: out = 16'(-300);
			44480: out = 16'(-244);
			44481: out = 16'(-91);
			44482: out = 16'(109);
			44483: out = 16'(252);
			44484: out = 16'(-88);
			44485: out = 16'(6);
			44486: out = 16'(27);
			44487: out = 16'(49);
			44488: out = 16'(5);
			44489: out = 16'(55);
			44490: out = 16'(-85);
			44491: out = 16'(46);
			44492: out = 16'(233);
			44493: out = 16'(698);
			44494: out = 16'(790);
			44495: out = 16'(642);
			44496: out = 16'(110);
			44497: out = 16'(-165);
			44498: out = 16'(62);
			44499: out = 16'(-7);
			44500: out = 16'(-138);
			44501: out = 16'(-880);
			44502: out = 16'(-658);
			44503: out = 16'(-428);
			44504: out = 16'(-17);
			44505: out = 16'(-120);
			44506: out = 16'(-365);
			44507: out = 16'(-260);
			44508: out = 16'(-404);
			44509: out = 16'(-436);
			44510: out = 16'(-630);
			44511: out = 16'(-414);
			44512: out = 16'(98);
			44513: out = 16'(-18);
			44514: out = 16'(-106);
			44515: out = 16'(-263);
			44516: out = 16'(-378);
			44517: out = 16'(-410);
			44518: out = 16'(-240);
			44519: out = 16'(-131);
			44520: out = 16'(50);
			44521: out = 16'(241);
			44522: out = 16'(314);
			44523: out = 16'(245);
			44524: out = 16'(155);
			44525: out = 16'(15);
			44526: out = 16'(-46);
			44527: out = 16'(-110);
			44528: out = 16'(-65);
			44529: out = 16'(-39);
			44530: out = 16'(670);
			44531: out = 16'(853);
			44532: out = 16'(650);
			44533: out = 16'(358);
			44534: out = 16'(168);
			44535: out = 16'(247);
			44536: out = 16'(82);
			44537: out = 16'(39);
			44538: out = 16'(-11);
			44539: out = 16'(7);
			44540: out = 16'(-76);
			44541: out = 16'(-274);
			44542: out = 16'(-606);
			44543: out = 16'(-872);
			44544: out = 16'(-825);
			44545: out = 16'(-681);
			44546: out = 16'(-379);
			44547: out = 16'(-351);
			44548: out = 16'(-77);
			44549: out = 16'(110);
			44550: out = 16'(617);
			44551: out = 16'(639);
			44552: out = 16'(406);
			44553: out = 16'(-75);
			44554: out = 16'(-378);
			44555: out = 16'(-445);
			44556: out = 16'(-223);
			44557: out = 16'(47);
			44558: out = 16'(394);
			44559: out = 16'(161);
			44560: out = 16'(-132);
			44561: out = 16'(-234);
			44562: out = 16'(-199);
			44563: out = 16'(-17);
			44564: out = 16'(54);
			44565: out = 16'(71);
			44566: out = 16'(-98);
			44567: out = 16'(-44);
			44568: out = 16'(-34);
			44569: out = 16'(143);
			44570: out = 16'(42);
			44571: out = 16'(179);
			44572: out = 16'(202);
			44573: out = 16'(586);
			44574: out = 16'(578);
			44575: out = 16'(265);
			44576: out = 16'(-314);
			44577: out = 16'(-706);
			44578: out = 16'(-637);
			44579: out = 16'(-309);
			44580: out = 16'(77);
			44581: out = 16'(-129);
			44582: out = 16'(-227);
			44583: out = 16'(-494);
			44584: out = 16'(-117);
			44585: out = 16'(-181);
			44586: out = 16'(-251);
			44587: out = 16'(-289);
			44588: out = 16'(-172);
			44589: out = 16'(-37);
			44590: out = 16'(267);
			44591: out = 16'(540);
			44592: out = 16'(673);
			44593: out = 16'(637);
			44594: out = 16'(411);
			44595: out = 16'(133);
			44596: out = 16'(-189);
			44597: out = 16'(-289);
			44598: out = 16'(-179);
			44599: out = 16'(67);
			44600: out = 16'(244);
			44601: out = 16'(218);
			44602: out = 16'(128);
			44603: out = 16'(5);
			44604: out = 16'(-428);
			44605: out = 16'(-426);
			44606: out = 16'(-307);
			44607: out = 16'(8);
			44608: out = 16'(57);
			44609: out = 16'(51);
			44610: out = 16'(-685);
			44611: out = 16'(-908);
			44612: out = 16'(-262);
			44613: out = 16'(-58);
			44614: out = 16'(119);
			44615: out = 16'(-106);
			44616: out = 16'(-264);
			44617: out = 16'(-483);
			44618: out = 16'(-571);
			44619: out = 16'(-455);
			44620: out = 16'(-160);
			44621: out = 16'(472);
			44622: out = 16'(576);
			44623: out = 16'(382);
			44624: out = 16'(163);
			44625: out = 16'(32);
			44626: out = 16'(73);
			44627: out = 16'(49);
			44628: out = 16'(14);
			44629: out = 16'(-116);
			44630: out = 16'(-114);
			44631: out = 16'(-56);
			44632: out = 16'(79);
			44633: out = 16'(461);
			44634: out = 16'(702);
			44635: out = 16'(401);
			44636: out = 16'(137);
			44637: out = 16'(-201);
			44638: out = 16'(-104);
			44639: out = 16'(-190);
			44640: out = 16'(-95);
			44641: out = 16'(-184);
			44642: out = 16'(29);
			44643: out = 16'(230);
			44644: out = 16'(471);
			44645: out = 16'(355);
			44646: out = 16'(-143);
			44647: out = 16'(-94);
			44648: out = 16'(-104);
			44649: out = 16'(23);
			44650: out = 16'(-211);
			44651: out = 16'(-373);
			44652: out = 16'(-479);
			44653: out = 16'(-483);
			44654: out = 16'(-461);
			44655: out = 16'(-473);
			44656: out = 16'(-309);
			44657: out = 16'(-58);
			44658: out = 16'(-106);
			44659: out = 16'(155);
			44660: out = 16'(441);
			44661: out = 16'(631);
			44662: out = 16'(653);
			44663: out = 16'(495);
			44664: out = 16'(330);
			44665: out = 16'(113);
			44666: out = 16'(23);
			44667: out = 16'(-115);
			44668: out = 16'(6);
			44669: out = 16'(319);
			44670: out = 16'(382);
			44671: out = 16'(256);
			44672: out = 16'(61);
			44673: out = 16'(-580);
			44674: out = 16'(-1126);
			44675: out = 16'(-1190);
			44676: out = 16'(-909);
			44677: out = 16'(-359);
			44678: out = 16'(-221);
			44679: out = 16'(-3);
			44680: out = 16'(43);
			44681: out = 16'(228);
			44682: out = 16'(335);
			44683: out = 16'(557);
			44684: out = 16'(222);
			44685: out = 16'(-110);
			44686: out = 16'(-639);
			44687: out = 16'(-763);
			44688: out = 16'(-687);
			44689: out = 16'(70);
			44690: out = 16'(-30);
			44691: out = 16'(0);
			44692: out = 16'(58);
			44693: out = 16'(351);
			44694: out = 16'(528);
			44695: out = 16'(327);
			44696: out = 16'(-71);
			44697: out = 16'(-496);
			44698: out = 16'(-600);
			44699: out = 16'(-424);
			44700: out = 16'(122);
			44701: out = 16'(295);
			44702: out = 16'(468);
			44703: out = 16'(359);
			44704: out = 16'(430);
			44705: out = 16'(345);
			44706: out = 16'(421);
			44707: out = 16'(46);
			44708: out = 16'(-88);
			44709: out = 16'(44);
			44710: out = 16'(-6);
			44711: out = 16'(-180);
			44712: out = 16'(-236);
			44713: out = 16'(-664);
			44714: out = 16'(-1038);
			44715: out = 16'(-1189);
			44716: out = 16'(-878);
			44717: out = 16'(-360);
			44718: out = 16'(-16);
			44719: out = 16'(-30);
			44720: out = 16'(-450);
			44721: out = 16'(-497);
			44722: out = 16'(-525);
			44723: out = 16'(-164);
			44724: out = 16'(-374);
			44725: out = 16'(-273);
			44726: out = 16'(108);
			44727: out = 16'(249);
			44728: out = 16'(382);
			44729: out = 16'(429);
			44730: out = 16'(698);
			44731: out = 16'(894);
			44732: out = 16'(890);
			44733: out = 16'(594);
			44734: out = 16'(188);
			44735: out = 16'(139);
			44736: out = 16'(38);
			44737: out = 16'(39);
			44738: out = 16'(-61);
			44739: out = 16'(-87);
			44740: out = 16'(-87);
			44741: out = 16'(-225);
			44742: out = 16'(-346);
			44743: out = 16'(-461);
			44744: out = 16'(-347);
			44745: out = 16'(-239);
			44746: out = 16'(-118);
			44747: out = 16'(-112);
			44748: out = 16'(-112);
			44749: out = 16'(-257);
			44750: out = 16'(-120);
			44751: out = 16'(144);
			44752: out = 16'(634);
			44753: out = 16'(725);
			44754: out = 16'(629);
			44755: out = 16'(-223);
			44756: out = 16'(-660);
			44757: out = 16'(-772);
			44758: out = 16'(-443);
			44759: out = 16'(-151);
			44760: out = 16'(-72);
			44761: out = 16'(193);
			44762: out = 16'(237);
			44763: out = 16'(72);
			44764: out = 16'(-148);
			44765: out = 16'(-304);
			44766: out = 16'(-233);
			44767: out = 16'(-291);
			44768: out = 16'(-204);
			44769: out = 16'(-156);
			44770: out = 16'(181);
			44771: out = 16'(468);
			44772: out = 16'(691);
			44773: out = 16'(547);
			44774: out = 16'(188);
			44775: out = 16'(148);
			44776: out = 16'(0);
			44777: out = 16'(-59);
			44778: out = 16'(-13);
			44779: out = 16'(33);
			44780: out = 16'(17);
			44781: out = 16'(-21);
			44782: out = 16'(-169);
			44783: out = 16'(-441);
			44784: out = 16'(-579);
			44785: out = 16'(-616);
			44786: out = 16'(-443);
			44787: out = 16'(-443);
			44788: out = 16'(-417);
			44789: out = 16'(-431);
			44790: out = 16'(-275);
			44791: out = 16'(-22);
			44792: out = 16'(205);
			44793: out = 16'(488);
			44794: out = 16'(727);
			44795: out = 16'(392);
			44796: out = 16'(133);
			44797: out = 16'(-106);
			44798: out = 16'(-131);
			44799: out = 16'(-53);
			44800: out = 16'(43);
			44801: out = 16'(193);
			44802: out = 16'(294);
			44803: out = 16'(561);
			44804: out = 16'(276);
			44805: out = 16'(-51);
			44806: out = 16'(-260);
			44807: out = 16'(-171);
			44808: out = 16'(70);
			44809: out = 16'(-102);
			44810: out = 16'(-35);
			44811: out = 16'(-122);
			44812: out = 16'(-40);
			44813: out = 16'(-170);
			44814: out = 16'(-273);
			44815: out = 16'(-576);
			44816: out = 16'(-480);
			44817: out = 16'(-40);
			44818: out = 16'(358);
			44819: out = 16'(543);
			44820: out = 16'(38);
			44821: out = 16'(114);
			44822: out = 16'(-39);
			44823: out = 16'(-35);
			44824: out = 16'(-523);
			44825: out = 16'(-785);
			44826: out = 16'(-637);
			44827: out = 16'(-334);
			44828: out = 16'(28);
			44829: out = 16'(373);
			44830: out = 16'(395);
			44831: out = 16'(233);
			44832: out = 16'(-121);
			44833: out = 16'(-351);
			44834: out = 16'(-418);
			44835: out = 16'(-72);
			44836: out = 16'(115);
			44837: out = 16'(66);
			44838: out = 16'(-123);
			44839: out = 16'(-245);
			44840: out = 16'(109);
			44841: out = 16'(49);
			44842: out = 16'(140);
			44843: out = 16'(213);
			44844: out = 16'(532);
			44845: out = 16'(684);
			44846: out = 16'(305);
			44847: out = 16'(147);
			44848: out = 16'(9);
			44849: out = 16'(-242);
			44850: out = 16'(-299);
			44851: out = 16'(-289);
			44852: out = 16'(-104);
			44853: out = 16'(-41);
			44854: out = 16'(70);
			44855: out = 16'(-327);
			44856: out = 16'(-349);
			44857: out = 16'(108);
			44858: out = 16'(192);
			44859: out = 16'(220);
			44860: out = 16'(-125);
			44861: out = 16'(-78);
			44862: out = 16'(-37);
			44863: out = 16'(236);
			44864: out = 16'(175);
			44865: out = 16'(69);
			44866: out = 16'(241);
			44867: out = 16'(165);
			44868: out = 16'(75);
			44869: out = 16'(24);
			44870: out = 16'(53);
			44871: out = 16'(52);
			44872: out = 16'(116);
			44873: out = 16'(-140);
			44874: out = 16'(-632);
			44875: out = 16'(-767);
			44876: out = 16'(-762);
			44877: out = 16'(-648);
			44878: out = 16'(-254);
			44879: out = 16'(41);
			44880: out = 16'(448);
			44881: out = 16'(0);
			44882: out = 16'(-550);
			44883: out = 16'(-1057);
			44884: out = 16'(-861);
			44885: out = 16'(-275);
			44886: out = 16'(-24);
			44887: out = 16'(204);
			44888: out = 16'(120);
			44889: out = 16'(431);
			44890: out = 16'(446);
			44891: out = 16'(453);
			44892: out = 16'(338);
			44893: out = 16'(218);
			44894: out = 16'(124);
			44895: out = 16'(-16);
			44896: out = 16'(-178);
			44897: out = 16'(-619);
			44898: out = 16'(-196);
			44899: out = 16'(255);
			44900: out = 16'(790);
			44901: out = 16'(814);
			44902: out = 16'(621);
			44903: out = 16'(161);
			44904: out = 16'(-18);
			44905: out = 16'(-101);
			44906: out = 16'(-244);
			44907: out = 16'(-427);
			44908: out = 16'(-650);
			44909: out = 16'(-669);
			44910: out = 16'(-478);
			44911: out = 16'(-103);
			44912: out = 16'(176);
			44913: out = 16'(171);
			44914: out = 16'(-268);
			44915: out = 16'(-462);
			44916: out = 16'(-548);
			44917: out = 16'(64);
			44918: out = 16'(13);
			44919: out = 16'(-36);
			44920: out = 16'(-85);
			44921: out = 16'(-88);
			44922: out = 16'(-107);
			44923: out = 16'(-374);
			44924: out = 16'(-372);
			44925: out = 16'(-214);
			44926: out = 16'(43);
			44927: out = 16'(222);
			44928: out = 16'(275);
			44929: out = 16'(404);
			44930: out = 16'(475);
			44931: out = 16'(573);
			44932: out = 16'(465);
			44933: out = 16'(348);
			44934: out = 16'(256);
			44935: out = 16'(43);
			44936: out = 16'(-101);
			44937: out = 16'(38);
			44938: out = 16'(-46);
			44939: out = 16'(-80);
			44940: out = 16'(-96);
			44941: out = 16'(-27);
			44942: out = 16'(5);
			44943: out = 16'(-370);
			44944: out = 16'(-562);
			44945: out = 16'(-615);
			44946: out = 16'(-646);
			44947: out = 16'(-424);
			44948: out = 16'(105);
			44949: out = 16'(-16);
			44950: out = 16'(-108);
			44951: out = 16'(-442);
			44952: out = 16'(-207);
			44953: out = 16'(-54);
			44954: out = 16'(-17);
			44955: out = 16'(-59);
			44956: out = 16'(-56);
			44957: out = 16'(64);
			44958: out = 16'(116);
			44959: out = 16'(152);
			44960: out = 16'(404);
			44961: out = 16'(375);
			44962: out = 16'(230);
			44963: out = 16'(-13);
			44964: out = 16'(-184);
			44965: out = 16'(-264);
			44966: out = 16'(-32);
			44967: out = 16'(58);
			44968: out = 16'(-74);
			44969: out = 16'(-34);
			44970: out = 16'(-14);
			44971: out = 16'(296);
			44972: out = 16'(137);
			44973: out = 16'(95);
			44974: out = 16'(-96);
			44975: out = 16'(285);
			44976: out = 16'(577);
			44977: out = 16'(689);
			44978: out = 16'(343);
			44979: out = 16'(-217);
			44980: out = 16'(-510);
			44981: out = 16'(-905);
			44982: out = 16'(-1190);
			44983: out = 16'(-881);
			44984: out = 16'(-599);
			44985: out = 16'(-204);
			44986: out = 16'(-403);
			44987: out = 16'(-288);
			44988: out = 16'(-19);
			44989: out = 16'(336);
			44990: out = 16'(382);
			44991: out = 16'(-56);
			44992: out = 16'(-307);
			44993: out = 16'(-487);
			44994: out = 16'(-55);
			44995: out = 16'(-27);
			44996: out = 16'(6);
			44997: out = 16'(-16);
			44998: out = 16'(0);
			44999: out = 16'(9);
			45000: out = 16'(87);
			45001: out = 16'(217);
			45002: out = 16'(403);
			45003: out = 16'(463);
			45004: out = 16'(441);
			45005: out = 16'(196);
			45006: out = 16'(139);
			45007: out = 16'(68);
			45008: out = 16'(104);
			45009: out = 16'(63);
			45010: out = 16'(125);
			45011: out = 16'(177);
			45012: out = 16'(242);
			45013: out = 16'(140);
			45014: out = 16'(-39);
			45015: out = 16'(-407);
			45016: out = 16'(-692);
			45017: out = 16'(-537);
			45018: out = 16'(-322);
			45019: out = 16'(-74);
			45020: out = 16'(-167);
			45021: out = 16'(-357);
			45022: out = 16'(-663);
			45023: out = 16'(-1070);
			45024: out = 16'(-1204);
			45025: out = 16'(-842);
			45026: out = 16'(-434);
			45027: out = 16'(39);
			45028: out = 16'(63);
			45029: out = 16'(455);
			45030: out = 16'(604);
			45031: out = 16'(1060);
			45032: out = 16'(467);
			45033: out = 16'(-122);
			45034: out = 16'(-676);
			45035: out = 16'(-654);
			45036: out = 16'(-380);
			45037: out = 16'(-48);
			45038: out = 16'(61);
			45039: out = 16'(18);
			45040: out = 16'(105);
			45041: out = 16'(195);
			45042: out = 16'(276);
			45043: out = 16'(644);
			45044: out = 16'(795);
			45045: out = 16'(741);
			45046: out = 16'(262);
			45047: out = 16'(-141);
			45048: out = 16'(-161);
			45049: out = 16'(-143);
			45050: out = 16'(27);
			45051: out = 16'(34);
			45052: out = 16'(86);
			45053: out = 16'(29);
			45054: out = 16'(7);
			45055: out = 16'(-119);
			45056: out = 16'(-200);
			45057: out = 16'(-218);
			45058: out = 16'(-127);
			45059: out = 16'(83);
			45060: out = 16'(-23);
			45061: out = 16'(-181);
			45062: out = 16'(-502);
			45063: out = 16'(-202);
			45064: out = 16'(72);
			45065: out = 16'(388);
			45066: out = 16'(222);
			45067: out = 16'(64);
			45068: out = 16'(-53);
			45069: out = 16'(-7);
			45070: out = 16'(135);
			45071: out = 16'(441);
			45072: out = 16'(549);
			45073: out = 16'(569);
			45074: out = 16'(146);
			45075: out = 16'(25);
			45076: out = 16'(43);
			45077: out = 16'(-98);
			45078: out = 16'(-134);
			45079: out = 16'(-277);
			45080: out = 16'(-11);
			45081: out = 16'(-33);
			45082: out = 16'(-237);
			45083: out = 16'(-535);
			45084: out = 16'(-636);
			45085: out = 16'(-354);
			45086: out = 16'(-188);
			45087: out = 16'(72);
			45088: out = 16'(318);
			45089: out = 16'(409);
			45090: out = 16'(258);
			45091: out = 16'(-120);
			45092: out = 16'(-579);
			45093: out = 16'(-1018);
			45094: out = 16'(-939);
			45095: out = 16'(-950);
			45096: out = 16'(-893);
			45097: out = 16'(-135);
			45098: out = 16'(354);
			45099: out = 16'(655);
			45100: out = 16'(503);
			45101: out = 16'(305);
			45102: out = 16'(158);
			45103: out = 16'(-2);
			45104: out = 16'(-49);
			45105: out = 16'(-59);
			45106: out = 16'(-12);
			45107: out = 16'(3);
			45108: out = 16'(263);
			45109: out = 16'(115);
			45110: out = 16'(-17);
			45111: out = 16'(65);
			45112: out = 16'(147);
			45113: out = 16'(264);
			45114: out = 16'(437);
			45115: out = 16'(498);
			45116: out = 16'(449);
			45117: out = 16'(91);
			45118: out = 16'(-146);
			45119: out = 16'(-230);
			45120: out = 16'(-158);
			45121: out = 16'(-65);
			45122: out = 16'(-62);
			45123: out = 16'(38);
			45124: out = 16'(78);
			45125: out = 16'(39);
			45126: out = 16'(31);
			45127: out = 16'(60);
			45128: out = 16'(317);
			45129: out = 16'(283);
			45130: out = 16'(155);
			45131: out = 16'(-28);
			45132: out = 16'(-98);
			45133: out = 16'(-123);
			45134: out = 16'(-234);
			45135: out = 16'(-222);
			45136: out = 16'(-95);
			45137: out = 16'(-325);
			45138: out = 16'(-378);
			45139: out = 16'(-393);
			45140: out = 16'(-78);
			45141: out = 16'(144);
			45142: out = 16'(205);
			45143: out = 16'(84);
			45144: out = 16'(-82);
			45145: out = 16'(61);
			45146: out = 16'(-57);
			45147: out = 16'(-61);
			45148: out = 16'(0);
			45149: out = 16'(137);
			45150: out = 16'(180);
			45151: out = 16'(-23);
			45152: out = 16'(-277);
			45153: out = 16'(-528);
			45154: out = 16'(-546);
			45155: out = 16'(-425);
			45156: out = 16'(-204);
			45157: out = 16'(17);
			45158: out = 16'(125);
			45159: out = 16'(99);
			45160: out = 16'(-171);
			45161: out = 16'(-416);
			45162: out = 16'(-470);
			45163: out = 16'(-423);
			45164: out = 16'(-290);
			45165: out = 16'(-85);
			45166: out = 16'(31);
			45167: out = 16'(102);
			45168: out = 16'(105);
			45169: out = 16'(233);
			45170: out = 16'(398);
			45171: out = 16'(469);
			45172: out = 16'(487);
			45173: out = 16'(475);
			45174: out = 16'(179);
			45175: out = 16'(52);
			45176: out = 16'(35);
			45177: out = 16'(148);
			45178: out = 16'(176);
			45179: out = 16'(78);
			45180: out = 16'(-52);
			45181: out = 16'(-119);
			45182: out = 16'(-88);
			45183: out = 16'(148);
			45184: out = 16'(329);
			45185: out = 16'(210);
			45186: out = 16'(46);
			45187: out = 16'(-184);
			45188: out = 16'(-625);
			45189: out = 16'(-649);
			45190: out = 16'(-500);
			45191: out = 16'(-196);
			45192: out = 16'(-24);
			45193: out = 16'(34);
			45194: out = 16'(-359);
			45195: out = 16'(-508);
			45196: out = 16'(-342);
			45197: out = 16'(2);
			45198: out = 16'(369);
			45199: out = 16'(568);
			45200: out = 16'(488);
			45201: out = 16'(271);
			45202: out = 16'(253);
			45203: out = 16'(105);
			45204: out = 16'(73);
			45205: out = 16'(-115);
			45206: out = 16'(-65);
			45207: out = 16'(32);
			45208: out = 16'(73);
			45209: out = 16'(-5);
			45210: out = 16'(-80);
			45211: out = 16'(-73);
			45212: out = 16'(-64);
			45213: out = 16'(-80);
			45214: out = 16'(0);
			45215: out = 16'(27);
			45216: out = 16'(13);
			45217: out = 16'(-143);
			45218: out = 16'(-345);
			45219: out = 16'(-655);
			45220: out = 16'(-608);
			45221: out = 16'(-449);
			45222: out = 16'(-143);
			45223: out = 16'(15);
			45224: out = 16'(62);
			45225: out = 16'(217);
			45226: out = 16'(158);
			45227: out = 16'(90);
			45228: out = 16'(-54);
			45229: out = 16'(-130);
			45230: out = 16'(-254);
			45231: out = 16'(-201);
			45232: out = 16'(-272);
			45233: out = 16'(-347);
			45234: out = 16'(-573);
			45235: out = 16'(-580);
			45236: out = 16'(-348);
			45237: out = 16'(97);
			45238: out = 16'(494);
			45239: out = 16'(717);
			45240: out = 16'(642);
			45241: out = 16'(410);
			45242: out = 16'(136);
			45243: out = 16'(106);
			45244: out = 16'(242);
			45245: out = 16'(67);
			45246: out = 16'(52);
			45247: out = 16'(-112);
			45248: out = 16'(197);
			45249: out = 16'(91);
			45250: out = 16'(-46);
			45251: out = 16'(-426);
			45252: out = 16'(-468);
			45253: out = 16'(-250);
			45254: out = 16'(155);
			45255: out = 16'(346);
			45256: out = 16'(208);
			45257: out = 16'(-29);
			45258: out = 16'(-338);
			45259: out = 16'(-643);
			45260: out = 16'(-474);
			45261: out = 16'(-173);
			45262: out = 16'(-74);
			45263: out = 16'(24);
			45264: out = 16'(59);
			45265: out = 16'(33);
			45266: out = 16'(132);
			45267: out = 16'(214);
			45268: out = 16'(345);
			45269: out = 16'(209);
			45270: out = 16'(-47);
			45271: out = 16'(-194);
			45272: out = 16'(-128);
			45273: out = 16'(185);
			45274: out = 16'(538);
			45275: out = 16'(622);
			45276: out = 16'(97);
			45277: out = 16'(-341);
			45278: out = 16'(-742);
			45279: out = 16'(-670);
			45280: out = 16'(-363);
			45281: out = 16'(161);
			45282: out = 16'(353);
			45283: out = 16'(561);
			45284: out = 16'(544);
			45285: out = 16'(295);
			45286: out = 16'(108);
			45287: out = 16'(67);
			45288: out = 16'(28);
			45289: out = 16'(60);
			45290: out = 16'(-9);
			45291: out = 16'(-51);
			45292: out = 16'(-232);
			45293: out = 16'(-373);
			45294: out = 16'(-597);
			45295: out = 16'(-606);
			45296: out = 16'(-146);
			45297: out = 16'(64);
			45298: out = 16'(203);
			45299: out = 16'(-18);
			45300: out = 16'(-194);
			45301: out = 16'(-425);
			45302: out = 16'(-457);
			45303: out = 16'(-552);
			45304: out = 16'(-467);
			45305: out = 16'(-767);
			45306: out = 16'(-578);
			45307: out = 16'(-13);
			45308: out = 16'(327);
			45309: out = 16'(621);
			45310: out = 16'(706);
			45311: out = 16'(754);
			45312: out = 16'(593);
			45313: out = 16'(118);
			45314: out = 16'(-121);
			45315: out = 16'(-239);
			45316: out = 16'(-65);
			45317: out = 16'(-61);
			45318: out = 16'(-94);
			45319: out = 16'(-436);
			45320: out = 16'(-609);
			45321: out = 16'(-612);
			45322: out = 16'(-189);
			45323: out = 16'(238);
			45324: out = 16'(610);
			45325: out = 16'(433);
			45326: out = 16'(208);
			45327: out = 16'(-76);
			45328: out = 16'(-307);
			45329: out = 16'(-317);
			45330: out = 16'(-54);
			45331: out = 16'(40);
			45332: out = 16'(95);
			45333: out = 16'(59);
			45334: out = 16'(-48);
			45335: out = 16'(-65);
			45336: out = 16'(47);
			45337: out = 16'(267);
			45338: out = 16'(480);
			45339: out = 16'(459);
			45340: out = 16'(258);
			45341: out = 16'(-122);
			45342: out = 16'(-191);
			45343: out = 16'(-363);
			45344: out = 16'(-532);
			45345: out = 16'(-433);
			45346: out = 16'(-335);
			45347: out = 16'(-241);
			45348: out = 16'(-59);
			45349: out = 16'(98);
			45350: out = 16'(59);
			45351: out = 16'(325);
			45352: out = 16'(473);
			45353: out = 16'(594);
			45354: out = 16'(321);
			45355: out = 16'(15);
			45356: out = 16'(-76);
			45357: out = 16'(0);
			45358: out = 16'(185);
			45359: out = 16'(-44);
			45360: out = 16'(-209);
			45361: out = 16'(-426);
			45362: out = 16'(-531);
			45363: out = 16'(-478);
			45364: out = 16'(-234);
			45365: out = 16'(-42);
			45366: out = 16'(133);
			45367: out = 16'(189);
			45368: out = 16'(104);
			45369: out = 16'(-17);
			45370: out = 16'(34);
			45371: out = 16'(4);
			45372: out = 16'(2);
			45373: out = 16'(-264);
			45374: out = 16'(-128);
			45375: out = 16'(24);
			45376: out = 16'(-99);
			45377: out = 16'(-170);
			45378: out = 16'(-231);
			45379: out = 16'(297);
			45380: out = 16'(587);
			45381: out = 16'(800);
			45382: out = 16'(443);
			45383: out = 16'(172);
			45384: out = 16'(0);
			45385: out = 16'(-408);
			45386: out = 16'(-642);
			45387: out = 16'(-707);
			45388: out = 16'(-616);
			45389: out = 16'(-560);
			45390: out = 16'(-838);
			45391: out = 16'(-685);
			45392: out = 16'(-372);
			45393: out = 16'(496);
			45394: out = 16'(693);
			45395: out = 16'(682);
			45396: out = 16'(426);
			45397: out = 16'(137);
			45398: out = 16'(-75);
			45399: out = 16'(-87);
			45400: out = 16'(-34);
			45401: out = 16'(61);
			45402: out = 16'(54);
			45403: out = 16'(-1);
			45404: out = 16'(-265);
			45405: out = 16'(-190);
			45406: out = 16'(-6);
			45407: out = 16'(427);
			45408: out = 16'(515);
			45409: out = 16'(490);
			45410: out = 16'(73);
			45411: out = 16'(-57);
			45412: out = 16'(-176);
			45413: out = 16'(-255);
			45414: out = 16'(-306);
			45415: out = 16'(-282);
			45416: out = 16'(-393);
			45417: out = 16'(-416);
			45418: out = 16'(-396);
			45419: out = 16'(-298);
			45420: out = 16'(-159);
			45421: out = 16'(34);
			45422: out = 16'(48);
			45423: out = 16'(132);
			45424: out = 16'(326);
			45425: out = 16'(332);
			45426: out = 16'(255);
			45427: out = 16'(-119);
			45428: out = 16'(-192);
			45429: out = 16'(-279);
			45430: out = 16'(-91);
			45431: out = 16'(-336);
			45432: out = 16'(-554);
			45433: out = 16'(-690);
			45434: out = 16'(-446);
			45435: out = 16'(-39);
			45436: out = 16'(149);
			45437: out = 16'(257);
			45438: out = 16'(192);
			45439: out = 16'(129);
			45440: out = 16'(93);
			45441: out = 16'(232);
			45442: out = 16'(108);
			45443: out = 16'(53);
			45444: out = 16'(28);
			45445: out = 16'(41);
			45446: out = 16'(73);
			45447: out = 16'(46);
			45448: out = 16'(123);
			45449: out = 16'(232);
			45450: out = 16'(660);
			45451: out = 16'(510);
			45452: out = 16'(212);
			45453: out = 16'(-295);
			45454: out = 16'(-570);
			45455: out = 16'(-717);
			45456: out = 16'(-261);
			45457: out = 16'(-67);
			45458: out = 16'(-76);
			45459: out = 16'(-283);
			45460: out = 16'(-455);
			45461: out = 16'(-523);
			45462: out = 16'(-235);
			45463: out = 16'(31);
			45464: out = 16'(62);
			45465: out = 16'(101);
			45466: out = 16'(62);
			45467: out = 16'(101);
			45468: out = 16'(8);
			45469: out = 16'(-38);
			45470: out = 16'(293);
			45471: out = 16'(342);
			45472: out = 16'(312);
			45473: out = 16'(-37);
			45474: out = 16'(-156);
			45475: out = 16'(-87);
			45476: out = 16'(-98);
			45477: out = 16'(-32);
			45478: out = 16'(20);
			45479: out = 16'(-45);
			45480: out = 16'(-33);
			45481: out = 16'(209);
			45482: out = 16'(78);
			45483: out = 16'(121);
			45484: out = 16'(418);
			45485: out = 16'(304);
			45486: out = 16'(96);
			45487: out = 16'(-213);
			45488: out = 16'(-381);
			45489: out = 16'(-391);
			45490: out = 16'(-316);
			45491: out = 16'(-130);
			45492: out = 16'(13);
			45493: out = 16'(171);
			45494: out = 16'(97);
			45495: out = 16'(-130);
			45496: out = 16'(-552);
			45497: out = 16'(-673);
			45498: out = 16'(-335);
			45499: out = 16'(-481);
			45500: out = 16'(-582);
			45501: out = 16'(-985);
			45502: out = 16'(-668);
			45503: out = 16'(-393);
			45504: out = 16'(-218);
			45505: out = 16'(-36);
			45506: out = 16'(138);
			45507: out = 16'(246);
			45508: out = 16'(274);
			45509: out = 16'(263);
			45510: out = 16'(574);
			45511: out = 16'(637);
			45512: out = 16'(566);
			45513: out = 16'(119);
			45514: out = 16'(-183);
			45515: out = 16'(-342);
			45516: out = 16'(-127);
			45517: out = 16'(178);
			45518: out = 16'(295);
			45519: out = 16'(680);
			45520: out = 16'(789);
			45521: out = 16'(709);
			45522: out = 16'(298);
			45523: out = 16'(-127);
			45524: out = 16'(-663);
			45525: out = 16'(-594);
			45526: out = 16'(-335);
			45527: out = 16'(93);
			45528: out = 16'(213);
			45529: out = 16'(159);
			45530: out = 16'(-279);
			45531: out = 16'(-438);
			45532: out = 16'(-382);
			45533: out = 16'(31);
			45534: out = 16'(297);
			45535: out = 16'(442);
			45536: out = 16'(85);
			45537: out = 16'(-277);
			45538: out = 16'(-686);
			45539: out = 16'(-435);
			45540: out = 16'(-171);
			45541: out = 16'(1);
			45542: out = 16'(10);
			45543: out = 16'(-79);
			45544: out = 16'(53);
			45545: out = 16'(189);
			45546: out = 16'(336);
			45547: out = 16'(321);
			45548: out = 16'(262);
			45549: out = 16'(173);
			45550: out = 16'(184);
			45551: out = 16'(194);
			45552: out = 16'(300);
			45553: out = 16'(292);
			45554: out = 16'(232);
			45555: out = 16'(3);
			45556: out = 16'(0);
			45557: out = 16'(-106);
			45558: out = 16'(-427);
			45559: out = 16'(-369);
			45560: out = 16'(-248);
			45561: out = 16'(10);
			45562: out = 16'(-20);
			45563: out = 16'(-145);
			45564: out = 16'(-368);
			45565: out = 16'(-448);
			45566: out = 16'(-390);
			45567: out = 16'(-438);
			45568: out = 16'(-316);
			45569: out = 16'(-269);
			45570: out = 16'(-11);
			45571: out = 16'(-8);
			45572: out = 16'(-102);
			45573: out = 16'(-502);
			45574: out = 16'(-703);
			45575: out = 16'(-649);
			45576: out = 16'(-405);
			45577: out = 16'(-126);
			45578: out = 16'(-47);
			45579: out = 16'(134);
			45580: out = 16'(237);
			45581: out = 16'(-6);
			45582: out = 16'(12);
			45583: out = 16'(73);
			45584: out = 16'(106);
			45585: out = 16'(84);
			45586: out = 16'(72);
			45587: out = 16'(-39);
			45588: out = 16'(117);
			45589: out = 16'(488);
			45590: out = 16'(478);
			45591: out = 16'(369);
			45592: out = 16'(7);
			45593: out = 16'(30);
			45594: out = 16'(4);
			45595: out = 16'(34);
			45596: out = 16'(-138);
			45597: out = 16'(-279);
			45598: out = 16'(-79);
			45599: out = 16'(-265);
			45600: out = 16'(-412);
			45601: out = 16'(-528);
			45602: out = 16'(-302);
			45603: out = 16'(-13);
			45604: out = 16'(167);
			45605: out = 16'(203);
			45606: out = 16'(64);
			45607: out = 16'(-12);
			45608: out = 16'(-46);
			45609: out = 16'(68);
			45610: out = 16'(-81);
			45611: out = 16'(-75);
			45612: out = 16'(-60);
			45613: out = 16'(-53);
			45614: out = 16'(-70);
			45615: out = 16'(-225);
			45616: out = 16'(-320);
			45617: out = 16'(-324);
			45618: out = 16'(38);
			45619: out = 16'(1);
			45620: out = 16'(-22);
			45621: out = 16'(69);
			45622: out = 16'(218);
			45623: out = 16'(361);
			45624: out = 16'(340);
			45625: out = 16'(288);
			45626: out = 16'(192);
			45627: out = 16'(-32);
			45628: out = 16'(-144);
			45629: out = 16'(-107);
			45630: out = 16'(-86);
			45631: out = 16'(-69);
			45632: out = 16'(-65);
			45633: out = 16'(-88);
			45634: out = 16'(-127);
			45635: out = 16'(-269);
			45636: out = 16'(-56);
			45637: out = 16'(80);
			45638: out = 16'(98);
			45639: out = 16'(-142);
			45640: out = 16'(-420);
			45641: out = 16'(-253);
			45642: out = 16'(-111);
			45643: out = 16'(123);
			45644: out = 16'(55);
			45645: out = 16'(54);
			45646: out = 16'(-71);
			45647: out = 16'(-46);
			45648: out = 16'(-43);
			45649: out = 16'(95);
			45650: out = 16'(-19);
			45651: out = 16'(-60);
			45652: out = 16'(-94);
			45653: out = 16'(-180);
			45654: out = 16'(-258);
			45655: out = 16'(-209);
			45656: out = 16'(-242);
			45657: out = 16'(-189);
			45658: out = 16'(-95);
			45659: out = 16'(154);
			45660: out = 16'(376);
			45661: out = 16'(352);
			45662: out = 16'(239);
			45663: out = 16'(10);
			45664: out = 16'(-165);
			45665: out = 16'(-180);
			45666: out = 16'(103);
			45667: out = 16'(-33);
			45668: out = 16'(-58);
			45669: out = 16'(-124);
			45670: out = 16'(-1);
			45671: out = 16'(35);
			45672: out = 16'(39);
			45673: out = 16'(-55);
			45674: out = 16'(-99);
			45675: out = 16'(-119);
			45676: out = 16'(-10);
			45677: out = 16'(101);
			45678: out = 16'(174);
			45679: out = 16'(207);
			45680: out = 16'(186);
			45681: out = 16'(67);
			45682: out = 16'(-8);
			45683: out = 16'(40);
			45684: out = 16'(-66);
			45685: out = 16'(-61);
			45686: out = 16'(31);
			45687: out = 16'(-83);
			45688: out = 16'(-133);
			45689: out = 16'(-111);
			45690: out = 16'(-124);
			45691: out = 16'(-90);
			45692: out = 16'(12);
			45693: out = 16'(-10);
			45694: out = 16'(-96);
			45695: out = 16'(-82);
			45696: out = 16'(-255);
			45697: out = 16'(-391);
			45698: out = 16'(-140);
			45699: out = 16'(-76);
			45700: out = 16'(-50);
			45701: out = 16'(54);
			45702: out = 16'(86);
			45703: out = 16'(63);
			45704: out = 16'(-16);
			45705: out = 16'(-80);
			45706: out = 16'(-42);
			45707: out = 16'(-78);
			45708: out = 16'(-40);
			45709: out = 16'(32);
			45710: out = 16'(38);
			45711: out = 16'(4);
			45712: out = 16'(-59);
			45713: out = 16'(-11);
			45714: out = 16'(24);
			45715: out = 16'(-249);
			45716: out = 16'(-143);
			45717: out = 16'(-52);
			45718: out = 16'(270);
			45719: out = 16'(258);
			45720: out = 16'(39);
			45721: out = 16'(-157);
			45722: out = 16'(-288);
			45723: out = 16'(-244);
			45724: out = 16'(-264);
			45725: out = 16'(-245);
			45726: out = 16'(-417);
			45727: out = 16'(-176);
			45728: out = 16'(-8);
			45729: out = 16'(369);
			45730: out = 16'(136);
			45731: out = 16'(-122);
			45732: out = 16'(-450);
			45733: out = 16'(-524);
			45734: out = 16'(-458);
			45735: out = 16'(-127);
			45736: out = 16'(-8);
			45737: out = 16'(-37);
			45738: out = 16'(101);
			45739: out = 16'(101);
			45740: out = 16'(89);
			45741: out = 16'(43);
			45742: out = 16'(81);
			45743: out = 16'(112);
			45744: out = 16'(104);
			45745: out = 16'(92);
			45746: out = 16'(101);
			45747: out = 16'(68);
			45748: out = 16'(-3);
			45749: out = 16'(-513);
			45750: out = 16'(-220);
			45751: out = 16'(143);
			45752: out = 16'(299);
			45753: out = 16'(389);
			45754: out = 16'(313);
			45755: out = 16'(252);
			45756: out = 16'(130);
			45757: out = 16'(74);
			45758: out = 16'(-48);
			45759: out = 16'(-29);
			45760: out = 16'(28);
			45761: out = 16'(59);
			45762: out = 16'(56);
			45763: out = 16'(64);
			45764: out = 16'(-46);
			45765: out = 16'(-125);
			45766: out = 16'(-109);
			45767: out = 16'(-83);
			45768: out = 16'(-62);
			45769: out = 16'(26);
			45770: out = 16'(-39);
			45771: out = 16'(-139);
			45772: out = 16'(-343);
			45773: out = 16'(-456);
			45774: out = 16'(-503);
			45775: out = 16'(-59);
			45776: out = 16'(134);
			45777: out = 16'(219);
			45778: out = 16'(116);
			45779: out = 16'(79);
			45780: out = 16'(72);
			45781: out = 16'(37);
			45782: out = 16'(-15);
			45783: out = 16'(-214);
			45784: out = 16'(-149);
			45785: out = 16'(-61);
			45786: out = 16'(4);
			45787: out = 16'(58);
			45788: out = 16'(59);
			45789: out = 16'(251);
			45790: out = 16'(155);
			45791: out = 16'(-19);
			45792: out = 16'(-181);
			45793: out = 16'(-191);
			45794: out = 16'(-76);
			45795: out = 16'(-206);
			45796: out = 16'(-168);
			45797: out = 16'(-91);
			45798: out = 16'(-91);
			45799: out = 16'(-110);
			45800: out = 16'(-200);
			45801: out = 16'(-130);
			45802: out = 16'(-60);
			45803: out = 16'(-56);
			45804: out = 16'(-49);
			45805: out = 16'(-91);
			45806: out = 16'(39);
			45807: out = 16'(-35);
			45808: out = 16'(-88);
			45809: out = 16'(-292);
			45810: out = 16'(-223);
			45811: out = 16'(-52);
			45812: out = 16'(-38);
			45813: out = 16'(-74);
			45814: out = 16'(-204);
			45815: out = 16'(-280);
			45816: out = 16'(-267);
			45817: out = 16'(-169);
			45818: out = 16'(-106);
			45819: out = 16'(-46);
			45820: out = 16'(-34);
			45821: out = 16'(40);
			45822: out = 16'(147);
			45823: out = 16'(363);
			45824: out = 16'(448);
			45825: out = 16'(437);
			45826: out = 16'(205);
			45827: out = 16'(-14);
			45828: out = 16'(-236);
			45829: out = 16'(-104);
			45830: out = 16'(-72);
			45831: out = 16'(-47);
			45832: out = 16'(13);
			45833: out = 16'(10);
			45834: out = 16'(30);
			45835: out = 16'(-48);
			45836: out = 16'(0);
			45837: out = 16'(151);
			45838: out = 16'(252);
			45839: out = 16'(174);
			45840: out = 16'(-93);
			45841: out = 16'(-310);
			45842: out = 16'(-421);
			45843: out = 16'(0);
			45844: out = 16'(81);
			45845: out = 16'(161);
			45846: out = 16'(-71);
			45847: out = 16'(-60);
			45848: out = 16'(-62);
			45849: out = 16'(33);
			45850: out = 16'(-2);
			45851: out = 16'(-73);
			45852: out = 16'(17);
			45853: out = 16'(-69);
			45854: out = 16'(-227);
			45855: out = 16'(-121);
			45856: out = 16'(-83);
			45857: out = 16'(-62);
			45858: out = 16'(-75);
			45859: out = 16'(-107);
			45860: out = 16'(-90);
			45861: out = 16'(-67);
			45862: out = 16'(-42);
			45863: out = 16'(-73);
			45864: out = 16'(51);
			45865: out = 16'(202);
			45866: out = 16'(437);
			45867: out = 16'(457);
			45868: out = 16'(431);
			45869: out = 16'(65);
			45870: out = 16'(-112);
			45871: out = 16'(-241);
			45872: out = 16'(-132);
			45873: out = 16'(-181);
			45874: out = 16'(-349);
			45875: out = 16'(-345);
			45876: out = 16'(-274);
			45877: out = 16'(-93);
			45878: out = 16'(-1);
			45879: out = 16'(63);
			45880: out = 16'(151);
			45881: out = 16'(98);
			45882: out = 16'(-72);
			45883: out = 16'(-525);
			45884: out = 16'(-527);
			45885: out = 16'(-411);
			45886: out = 16'(-448);
			45887: out = 16'(-405);
			45888: out = 16'(-406);
			45889: out = 16'(-9);
			45890: out = 16'(37);
			45891: out = 16'(-36);
			45892: out = 16'(50);
			45893: out = 16'(177);
			45894: out = 16'(389);
			45895: out = 16'(203);
			45896: out = 16'(-40);
			45897: out = 16'(-286);
			45898: out = 16'(-388);
			45899: out = 16'(-381);
			45900: out = 16'(-322);
			45901: out = 16'(-128);
			45902: out = 16'(-7);
			45903: out = 16'(-10);
			45904: out = 16'(-82);
			45905: out = 16'(-145);
			45906: out = 16'(-2);
			45907: out = 16'(186);
			45908: out = 16'(303);
			45909: out = 16'(404);
			45910: out = 16'(252);
			45911: out = 16'(-39);
			45912: out = 16'(-140);
			45913: out = 16'(-153);
			45914: out = 16'(-36);
			45915: out = 16'(312);
			45916: out = 16'(469);
			45917: out = 16'(163);
			45918: out = 16'(-11);
			45919: out = 16'(-230);
			45920: out = 16'(60);
			45921: out = 16'(-36);
			45922: out = 16'(-26);
			45923: out = 16'(-104);
			45924: out = 16'(-9);
			45925: out = 16'(14);
			45926: out = 16'(55);
			45927: out = 16'(-151);
			45928: out = 16'(-436);
			45929: out = 16'(-429);
			45930: out = 16'(-294);
			45931: out = 16'(66);
			45932: out = 16'(33);
			45933: out = 16'(70);
			45934: out = 16'(20);
			45935: out = 16'(133);
			45936: out = 16'(234);
			45937: out = 16'(457);
			45938: out = 16'(475);
			45939: out = 16'(418);
			45940: out = 16'(33);
			45941: out = 16'(-83);
			45942: out = 16'(-269);
			45943: out = 16'(-271);
			45944: out = 16'(-551);
			45945: out = 16'(-791);
			45946: out = 16'(-844);
			45947: out = 16'(-449);
			45948: out = 16'(248);
			45949: out = 16'(478);
			45950: out = 16'(575);
			45951: out = 16'(359);
			45952: out = 16'(198);
			45953: out = 16'(-22);
			45954: out = 16'(-42);
			45955: out = 16'(-255);
			45956: out = 16'(-260);
			45957: out = 16'(7);
			45958: out = 16'(41);
			45959: out = 16'(10);
			45960: out = 16'(-179);
			45961: out = 16'(-107);
			45962: out = 16'(60);
			45963: out = 16'(50);
			45964: out = 16'(39);
			45965: out = 16'(-77);
			45966: out = 16'(-224);
			45967: out = 16'(-430);
			45968: out = 16'(-652);
			45969: out = 16'(-676);
			45970: out = 16'(-515);
			45971: out = 16'(-14);
			45972: out = 16'(-59);
			45973: out = 16'(-13);
			45974: out = 16'(-69);
			45975: out = 16'(171);
			45976: out = 16'(333);
			45977: out = 16'(419);
			45978: out = 16'(251);
			45979: out = 16'(44);
			45980: out = 16'(-29);
			45981: out = 16'(-60);
			45982: out = 16'(-13);
			45983: out = 16'(398);
			45984: out = 16'(506);
			45985: out = 16'(457);
			45986: out = 16'(254);
			45987: out = 16'(83);
			45988: out = 16'(52);
			45989: out = 16'(102);
			45990: out = 16'(169);
			45991: out = 16'(130);
			45992: out = 16'(81);
			45993: out = 16'(-85);
			45994: out = 16'(-288);
			45995: out = 16'(-490);
			45996: out = 16'(-550);
			45997: out = 16'(-465);
			45998: out = 16'(-271);
			45999: out = 16'(-65);
			46000: out = 16'(-172);
			46001: out = 16'(-234);
			46002: out = 16'(-311);
			46003: out = 16'(-117);
			46004: out = 16'(-38);
			46005: out = 16'(-30);
			46006: out = 16'(126);
			46007: out = 16'(190);
			46008: out = 16'(171);
			46009: out = 16'(105);
			46010: out = 16'(-17);
			46011: out = 16'(-52);
			46012: out = 16'(-145);
			46013: out = 16'(-222);
			46014: out = 16'(-301);
			46015: out = 16'(-234);
			46016: out = 16'(-154);
			46017: out = 16'(-90);
			46018: out = 16'(-7);
			46019: out = 16'(63);
			46020: out = 16'(267);
			46021: out = 16'(283);
			46022: out = 16'(280);
			46023: out = 16'(184);
			46024: out = 16'(220);
			46025: out = 16'(372);
			46026: out = 16'(217);
			46027: out = 16'(112);
			46028: out = 16'(12);
			46029: out = 16'(-3);
			46030: out = 16'(-8);
			46031: out = 16'(-119);
			46032: out = 16'(-75);
			46033: out = 16'(-72);
			46034: out = 16'(41);
			46035: out = 16'(-63);
			46036: out = 16'(-277);
			46037: out = 16'(-622);
			46038: out = 16'(-714);
			46039: out = 16'(-635);
			46040: out = 16'(-598);
			46041: out = 16'(-342);
			46042: out = 16'(-45);
			46043: out = 16'(-46);
			46044: out = 16'(-43);
			46045: out = 16'(-47);
			46046: out = 16'(42);
			46047: out = 16'(207);
			46048: out = 16'(597);
			46049: out = 16'(539);
			46050: out = 16'(418);
			46051: out = 16'(196);
			46052: out = 16'(40);
			46053: out = 16'(-66);
			46054: out = 16'(27);
			46055: out = 16'(-36);
			46056: out = 16'(-105);
			46057: out = 16'(-88);
			46058: out = 16'(-77);
			46059: out = 16'(-32);
			46060: out = 16'(102);
			46061: out = 16'(232);
			46062: out = 16'(352);
			46063: out = 16'(505);
			46064: out = 16'(493);
			46065: out = 16'(318);
			46066: out = 16'(138);
			46067: out = 16'(-54);
			46068: out = 16'(-93);
			46069: out = 16'(-352);
			46070: out = 16'(-461);
			46071: out = 16'(-255);
			46072: out = 16'(-115);
			46073: out = 16'(14);
			46074: out = 16'(-10);
			46075: out = 16'(-45);
			46076: out = 16'(-150);
			46077: out = 16'(-280);
			46078: out = 16'(-430);
			46079: out = 16'(-566);
			46080: out = 16'(-473);
			46081: out = 16'(-393);
			46082: out = 16'(-300);
			46083: out = 16'(-209);
			46084: out = 16'(-143);
			46085: out = 16'(55);
			46086: out = 16'(57);
			46087: out = 16'(104);
			46088: out = 16'(147);
			46089: out = 16'(265);
			46090: out = 16'(261);
			46091: out = 16'(286);
			46092: out = 16'(111);
			46093: out = 16'(-99);
			46094: out = 16'(-276);
			46095: out = 16'(-338);
			46096: out = 16'(-301);
			46097: out = 16'(-26);
			46098: out = 16'(29);
			46099: out = 16'(-60);
			46100: out = 16'(-69);
			46101: out = 16'(-31);
			46102: out = 16'(61);
			46103: out = 16'(136);
			46104: out = 16'(153);
			46105: out = 16'(28);
			46106: out = 16'(-96);
			46107: out = 16'(-253);
			46108: out = 16'(-293);
			46109: out = 16'(-324);
			46110: out = 16'(-278);
			46111: out = 16'(-208);
			46112: out = 16'(-126);
			46113: out = 16'(-44);
			46114: out = 16'(0);
			46115: out = 16'(150);
			46116: out = 16'(304);
			46117: out = 16'(281);
			46118: out = 16'(216);
			46119: out = 16'(47);
			46120: out = 16'(54);
			46121: out = 16'(79);
			46122: out = 16'(160);
			46123: out = 16'(100);
			46124: out = 16'(34);
			46125: out = 16'(15);
			46126: out = 16'(-5);
			46127: out = 16'(34);
			46128: out = 16'(27);
			46129: out = 16'(146);
			46130: out = 16'(259);
			46131: out = 16'(251);
			46132: out = 16'(152);
			46133: out = 16'(-2);
			46134: out = 16'(-57);
			46135: out = 16'(-148);
			46136: out = 16'(-231);
			46137: out = 16'(-159);
			46138: out = 16'(-87);
			46139: out = 16'(-86);
			46140: out = 16'(-5);
			46141: out = 16'(-17);
			46142: out = 16'(-90);
			46143: out = 16'(-73);
			46144: out = 16'(-56);
			46145: out = 16'(-4);
			46146: out = 16'(-38);
			46147: out = 16'(-77);
			46148: out = 16'(-106);
			46149: out = 16'(-150);
			46150: out = 16'(-244);
			46151: out = 16'(-191);
			46152: out = 16'(-364);
			46153: out = 16'(-568);
			46154: out = 16'(-570);
			46155: out = 16'(-365);
			46156: out = 16'(89);
			46157: out = 16'(96);
			46158: out = 16'(302);
			46159: out = 16'(459);
			46160: out = 16'(543);
			46161: out = 16'(535);
			46162: out = 16'(458);
			46163: out = 16'(212);
			46164: out = 16'(-111);
			46165: out = 16'(-647);
			46166: out = 16'(-845);
			46167: out = 16'(-895);
			46168: out = 16'(-375);
			46169: out = 16'(-262);
			46170: out = 16'(-126);
			46171: out = 16'(-13);
			46172: out = 16'(358);
			46173: out = 16'(763);
			46174: out = 16'(634);
			46175: out = 16'(350);
			46176: out = 16'(-124);
			46177: out = 16'(-426);
			46178: out = 16'(-539);
			46179: out = 16'(-297);
			46180: out = 16'(-160);
			46181: out = 16'(21);
			46182: out = 16'(147);
			46183: out = 16'(180);
			46184: out = 16'(166);
			46185: out = 16'(264);
			46186: out = 16'(257);
			46187: out = 16'(236);
			46188: out = 16'(63);
			46189: out = 16'(14);
			46190: out = 16'(-8);
			46191: out = 16'(-373);
			46192: out = 16'(-465);
			46193: out = 16'(-420);
			46194: out = 16'(-366);
			46195: out = 16'(-299);
			46196: out = 16'(-300);
			46197: out = 16'(-151);
			46198: out = 16'(-14);
			46199: out = 16'(52);
			46200: out = 16'(217);
			46201: out = 16'(279);
			46202: out = 16'(282);
			46203: out = 16'(105);
			46204: out = 16'(-79);
			46205: out = 16'(-175);
			46206: out = 16'(-148);
			46207: out = 16'(-96);
			46208: out = 16'(-73);
			46209: out = 16'(-201);
			46210: out = 16'(-436);
			46211: out = 16'(-401);
			46212: out = 16'(-362);
			46213: out = 16'(-140);
			46214: out = 16'(-99);
			46215: out = 16'(131);
			46216: out = 16'(495);
			46217: out = 16'(426);
			46218: out = 16'(319);
			46219: out = 16'(72);
			46220: out = 16'(-2);
			46221: out = 16'(-68);
			46222: out = 16'(-46);
			46223: out = 16'(-273);
			46224: out = 16'(-442);
			46225: out = 16'(-311);
			46226: out = 16'(-187);
			46227: out = 16'(10);
			46228: out = 16'(203);
			46229: out = 16'(407);
			46230: out = 16'(558);
			46231: out = 16'(589);
			46232: out = 16'(383);
			46233: out = 16'(-97);
			46234: out = 16'(1);
			46235: out = 16'(-28);
			46236: out = 16'(21);
			46237: out = 16'(-270);
			46238: out = 16'(-481);
			46239: out = 16'(-452);
			46240: out = 16'(-275);
			46241: out = 16'(5);
			46242: out = 16'(287);
			46243: out = 16'(479);
			46244: out = 16'(504);
			46245: out = 16'(115);
			46246: out = 16'(-205);
			46247: out = 16'(-451);
			46248: out = 16'(-463);
			46249: out = 16'(-439);
			46250: out = 16'(-439);
			46251: out = 16'(-160);
			46252: out = 16'(-89);
			46253: out = 16'(-201);
			46254: out = 16'(-182);
			46255: out = 16'(-143);
			46256: out = 16'(78);
			46257: out = 16'(114);
			46258: out = 16'(225);
			46259: out = 16'(352);
			46260: out = 16'(419);
			46261: out = 16'(425);
			46262: out = 16'(189);
			46263: out = 16'(73);
			46264: out = 16'(-22);
			46265: out = 16'(-101);
			46266: out = 16'(-151);
			46267: out = 16'(-235);
			46268: out = 16'(-68);
			46269: out = 16'(29);
			46270: out = 16'(18);
			46271: out = 16'(36);
			46272: out = 16'(-8);
			46273: out = 16'(-68);
			46274: out = 16'(-117);
			46275: out = 16'(-121);
			46276: out = 16'(-237);
			46277: out = 16'(-139);
			46278: out = 16'(-61);
			46279: out = 16'(1);
			46280: out = 16'(-150);
			46281: out = 16'(-356);
			46282: out = 16'(-225);
			46283: out = 16'(-116);
			46284: out = 16'(80);
			46285: out = 16'(102);
			46286: out = 16'(215);
			46287: out = 16'(233);
			46288: out = 16'(188);
			46289: out = 16'(61);
			46290: out = 16'(-113);
			46291: out = 16'(-191);
			46292: out = 16'(-228);
			46293: out = 16'(-235);
			46294: out = 16'(-134);
			46295: out = 16'(-15);
			46296: out = 16'(241);
			46297: out = 16'(190);
			46298: out = 16'(147);
			46299: out = 16'(226);
			46300: out = 16'(275);
			46301: out = 16'(310);
			46302: out = 16'(177);
			46303: out = 16'(-67);
			46304: out = 16'(-419);
			46305: out = 16'(-516);
			46306: out = 16'(-630);
			46307: out = 16'(-557);
			46308: out = 16'(-522);
			46309: out = 16'(-295);
			46310: out = 16'(-8);
			46311: out = 16'(212);
			46312: out = 16'(247);
			46313: out = 16'(165);
			46314: out = 16'(-40);
			46315: out = 16'(-269);
			46316: out = 16'(-409);
			46317: out = 16'(-410);
			46318: out = 16'(-259);
			46319: out = 16'(-11);
			46320: out = 16'(72);
			46321: out = 16'(39);
			46322: out = 16'(-37);
			46323: out = 16'(-90);
			46324: out = 16'(-72);
			46325: out = 16'(-73);
			46326: out = 16'(-109);
			46327: out = 16'(-209);
			46328: out = 16'(69);
			46329: out = 16'(268);
			46330: out = 16'(473);
			46331: out = 16'(353);
			46332: out = 16'(193);
			46333: out = 16'(-49);
			46334: out = 16'(-30);
			46335: out = 16'(79);
			46336: out = 16'(105);
			46337: out = 16'(256);
			46338: out = 16'(350);
			46339: out = 16'(431);
			46340: out = 16'(351);
			46341: out = 16'(192);
			46342: out = 16'(-49);
			46343: out = 16'(-84);
			46344: out = 16'(-29);
			46345: out = 16'(-75);
			46346: out = 16'(-125);
			46347: out = 16'(-90);
			46348: out = 16'(-282);
			46349: out = 16'(-386);
			46350: out = 16'(-490);
			46351: out = 16'(-260);
			46352: out = 16'(-73);
			46353: out = 16'(-4);
			46354: out = 16'(-173);
			46355: out = 16'(-352);
			46356: out = 16'(-111);
			46357: out = 16'(-41);
			46358: out = 16'(55);
			46359: out = 16'(22);
			46360: out = 16'(-76);
			46361: out = 16'(-248);
			46362: out = 16'(-464);
			46363: out = 16'(-620);
			46364: out = 16'(-639);
			46365: out = 16'(-441);
			46366: out = 16'(-151);
			46367: out = 16'(25);
			46368: out = 16'(358);
			46369: out = 16'(532);
			46370: out = 16'(569);
			46371: out = 16'(473);
			46372: out = 16'(307);
			46373: out = 16'(52);
			46374: out = 16'(-54);
			46375: out = 16'(-82);
			46376: out = 16'(-403);
			46377: out = 16'(-496);
			46378: out = 16'(-536);
			46379: out = 16'(-43);
			46380: out = 16'(159);
			46381: out = 16'(274);
			46382: out = 16'(30);
			46383: out = 16'(-79);
			46384: out = 16'(-74);
			46385: out = 16'(-22);
			46386: out = 16'(17);
			46387: out = 16'(-53);
			46388: out = 16'(6);
			46389: out = 16'(-1);
			46390: out = 16'(-78);
			46391: out = 16'(-89);
			46392: out = 16'(-74);
			46393: out = 16'(-61);
			46394: out = 16'(-42);
			46395: out = 16'(-44);
			46396: out = 16'(132);
			46397: out = 16'(160);
			46398: out = 16'(164);
			46399: out = 16'(47);
			46400: out = 16'(-22);
			46401: out = 16'(-106);
			46402: out = 16'(-70);
			46403: out = 16'(-37);
			46404: out = 16'(58);
			46405: out = 16'(-35);
			46406: out = 16'(-37);
			46407: out = 16'(23);
			46408: out = 16'(116);
			46409: out = 16'(152);
			46410: out = 16'(264);
			46411: out = 16'(70);
			46412: out = 16'(-93);
			46413: out = 16'(-101);
			46414: out = 16'(-75);
			46415: out = 16'(0);
			46416: out = 16'(-62);
			46417: out = 16'(-125);
			46418: out = 16'(-219);
			46419: out = 16'(-411);
			46420: out = 16'(-368);
			46421: out = 16'(-69);
			46422: out = 16'(0);
			46423: out = 16'(79);
			46424: out = 16'(34);
			46425: out = 16'(-15);
			46426: out = 16'(-54);
			46427: out = 16'(64);
			46428: out = 16'(29);
			46429: out = 16'(44);
			46430: out = 16'(32);
			46431: out = 16'(-206);
			46432: out = 16'(-485);
			46433: out = 16'(-304);
			46434: out = 16'(-340);
			46435: out = 16'(-296);
			46436: out = 16'(-425);
			46437: out = 16'(-278);
			46438: out = 16'(-11);
			46439: out = 16'(129);
			46440: out = 16'(161);
			46441: out = 16'(18);
			46442: out = 16'(55);
			46443: out = 16'(15);
			46444: out = 16'(-25);
			46445: out = 16'(-61);
			46446: out = 16'(-67);
			46447: out = 16'(36);
			46448: out = 16'(-11);
			46449: out = 16'(-19);
			46450: out = 16'(121);
			46451: out = 16'(316);
			46452: out = 16'(479);
			46453: out = 16'(197);
			46454: out = 16'(88);
			46455: out = 16'(0);
			46456: out = 16'(15);
			46457: out = 16'(-12);
			46458: out = 16'(-87);
			46459: out = 16'(28);
			46460: out = 16'(8);
			46461: out = 16'(-63);
			46462: out = 16'(-171);
			46463: out = 16'(-227);
			46464: out = 16'(-217);
			46465: out = 16'(-67);
			46466: out = 16'(91);
			46467: out = 16'(249);
			46468: out = 16'(165);
			46469: out = 16'(0);
			46470: out = 16'(47);
			46471: out = 16'(25);
			46472: out = 16'(12);
			46473: out = 16'(-350);
			46474: out = 16'(-569);
			46475: out = 16'(-685);
			46476: out = 16'(-442);
			46477: out = 16'(-95);
			46478: out = 16'(275);
			46479: out = 16'(425);
			46480: out = 16'(388);
			46481: out = 16'(39);
			46482: out = 16'(-37);
			46483: out = 16'(-93);
			46484: out = 16'(13);
			46485: out = 16'(-51);
			46486: out = 16'(-104);
			46487: out = 16'(-100);
			46488: out = 16'(-73);
			46489: out = 16'(-62);
			46490: out = 16'(-71);
			46491: out = 16'(-54);
			46492: out = 16'(-54);
			46493: out = 16'(117);
			46494: out = 16'(200);
			46495: out = 16'(257);
			46496: out = 16'(327);
			46497: out = 16'(334);
			46498: out = 16'(223);
			46499: out = 16'(170);
			46500: out = 16'(75);
			46501: out = 16'(12);
			46502: out = 16'(-296);
			46503: out = 16'(-508);
			46504: out = 16'(-458);
			46505: out = 16'(-412);
			46506: out = 16'(-290);
			46507: out = 16'(-27);
			46508: out = 16'(-12);
			46509: out = 16'(-68);
			46510: out = 16'(-59);
			46511: out = 16'(-59);
			46512: out = 16'(-62);
			46513: out = 16'(-73);
			46514: out = 16'(-208);
			46515: out = 16'(-439);
			46516: out = 16'(-446);
			46517: out = 16'(-338);
			46518: out = 16'(-72);
			46519: out = 16'(83);
			46520: out = 16'(219);
			46521: out = 16'(276);
			46522: out = 16'(221);
			46523: out = 16'(125);
			46524: out = 16'(75);
			46525: out = 16'(37);
			46526: out = 16'(28);
			46527: out = 16'(50);
			46528: out = 16'(-8);
			46529: out = 16'(-90);
			46530: out = 16'(-256);
			46531: out = 16'(-351);
			46532: out = 16'(-289);
			46533: out = 16'(-75);
			46534: out = 16'(72);
			46535: out = 16'(23);
			46536: out = 16'(447);
			46537: out = 16'(566);
			46538: out = 16'(571);
			46539: out = 16'(143);
			46540: out = 16'(-126);
			46541: out = 16'(-111);
			46542: out = 16'(28);
			46543: out = 16'(108);
			46544: out = 16'(-210);
			46545: out = 16'(-446);
			46546: out = 16'(-706);
			46547: out = 16'(-162);
			46548: out = 16'(-30);
			46549: out = 16'(36);
			46550: out = 16'(-244);
			46551: out = 16'(-443);
			46552: out = 16'(-682);
			46553: out = 16'(-327);
			46554: out = 16'(-69);
			46555: out = 16'(59);
			46556: out = 16'(232);
			46557: out = 16'(233);
			46558: out = 16'(-71);
			46559: out = 16'(-230);
			46560: out = 16'(-273);
			46561: out = 16'(31);
			46562: out = 16'(8);
			46563: out = 16'(-22);
			46564: out = 16'(151);
			46565: out = 16'(269);
			46566: out = 16'(394);
			46567: out = 16'(354);
			46568: out = 16'(371);
			46569: out = 16'(300);
			46570: out = 16'(178);
			46571: out = 16'(-38);
			46572: out = 16'(-291);
			46573: out = 16'(-479);
			46574: out = 16'(-570);
			46575: out = 16'(-550);
			46576: out = 16'(-321);
			46577: out = 16'(-49);
			46578: out = 16'(83);
			46579: out = 16'(230);
			46580: out = 16'(271);
			46581: out = 16'(197);
			46582: out = 16'(143);
			46583: out = 16'(90);
			46584: out = 16'(29);
			46585: out = 16'(-124);
			46586: out = 16'(-274);
			46587: out = 16'(-279);
			46588: out = 16'(-171);
			46589: out = 16'(17);
			46590: out = 16'(19);
			46591: out = 16'(11);
			46592: out = 16'(-61);
			46593: out = 16'(-6);
			46594: out = 16'(-39);
			46595: out = 16'(-158);
			46596: out = 16'(-174);
			46597: out = 16'(-138);
			46598: out = 16'(-59);
			46599: out = 16'(-1);
			46600: out = 16'(44);
			46601: out = 16'(7);
			46602: out = 16'(-12);
			46603: out = 16'(-39);
			46604: out = 16'(245);
			46605: out = 16'(266);
			46606: out = 16'(259);
			46607: out = 16'(50);
			46608: out = 16'(-21);
			46609: out = 16'(-20);
			46610: out = 16'(77);
			46611: out = 16'(59);
			46612: out = 16'(-75);
			46613: out = 16'(-204);
			46614: out = 16'(-296);
			46615: out = 16'(-372);
			46616: out = 16'(-195);
			46617: out = 16'(-51);
			46618: out = 16'(21);
			46619: out = 16'(-24);
			46620: out = 16'(-111);
			46621: out = 16'(-329);
			46622: out = 16'(-245);
			46623: out = 16'(-39);
			46624: out = 16'(68);
			46625: out = 16'(138);
			46626: out = 16'(102);
			46627: out = 16'(70);
			46628: out = 16'(-6);
			46629: out = 16'(-59);
			46630: out = 16'(0);
			46631: out = 16'(6);
			46632: out = 16'(9);
			46633: out = 16'(-166);
			46634: out = 16'(-290);
			46635: out = 16'(-431);
			46636: out = 16'(-186);
			46637: out = 16'(89);
			46638: out = 16'(89);
			46639: out = 16'(144);
			46640: out = 16'(107);
			46641: out = 16'(225);
			46642: out = 16'(74);
			46643: out = 16'(-49);
			46644: out = 16'(-156);
			46645: out = 16'(-133);
			46646: out = 16'(-47);
			46647: out = 16'(267);
			46648: out = 16'(306);
			46649: out = 16'(86);
			46650: out = 16'(38);
			46651: out = 16'(-8);
			46652: out = 16'(122);
			46653: out = 16'(36);
			46654: out = 16'(18);
			46655: out = 16'(-13);
			46656: out = 16'(-43);
			46657: out = 16'(-73);
			46658: out = 16'(-92);
			46659: out = 16'(-138);
			46660: out = 16'(-192);
			46661: out = 16'(-175);
			46662: out = 16'(-202);
			46663: out = 16'(-270);
			46664: out = 16'(-110);
			46665: out = 16'(-50);
			46666: out = 16'(16);
			46667: out = 16'(-190);
			46668: out = 16'(-256);
			46669: out = 16'(-246);
			46670: out = 16'(-85);
			46671: out = 16'(47);
			46672: out = 16'(0);
			46673: out = 16'(29);
			46674: out = 16'(65);
			46675: out = 16'(264);
			46676: out = 16'(197);
			46677: out = 16'(82);
			46678: out = 16'(-60);
			46679: out = 16'(-96);
			46680: out = 16'(-70);
			46681: out = 16'(1);
			46682: out = 16'(57);
			46683: out = 16'(111);
			46684: out = 16'(14);
			46685: out = 16'(-33);
			46686: out = 16'(-89);
			46687: out = 16'(-64);
			46688: out = 16'(-45);
			46689: out = 16'(-4);
			46690: out = 16'(-104);
			46691: out = 16'(-206);
			46692: out = 16'(-336);
			46693: out = 16'(-312);
			46694: out = 16'(-203);
			46695: out = 16'(88);
			46696: out = 16'(190);
			46697: out = 16'(287);
			46698: out = 16'(113);
			46699: out = 16'(149);
			46700: out = 16'(169);
			46701: out = 16'(141);
			46702: out = 16'(-29);
			46703: out = 16'(-261);
			46704: out = 16'(-490);
			46705: out = 16'(-443);
			46706: out = 16'(-62);
			46707: out = 16'(-23);
			46708: out = 16'(-1);
			46709: out = 16'(-171);
			46710: out = 16'(-272);
			46711: out = 16'(-331);
			46712: out = 16'(-156);
			46713: out = 16'(-118);
			46714: out = 16'(7);
			46715: out = 16'(236);
			46716: out = 16'(321);
			46717: out = 16'(326);
			46718: out = 16'(301);
			46719: out = 16'(160);
			46720: out = 16'(17);
			46721: out = 16'(-76);
			46722: out = 16'(-93);
			46723: out = 16'(-11);
			46724: out = 16'(-131);
			46725: out = 16'(-243);
			46726: out = 16'(-448);
			46727: out = 16'(-353);
			46728: out = 16'(-185);
			46729: out = 16'(24);
			46730: out = 16'(46);
			46731: out = 16'(27);
			46732: out = 16'(41);
			46733: out = 16'(-19);
			46734: out = 16'(-49);
			46735: out = 16'(0);
			46736: out = 16'(-20);
			46737: out = 16'(-44);
			46738: out = 16'(15);
			46739: out = 16'(7);
			46740: out = 16'(10);
			46741: out = 16'(1);
			46742: out = 16'(-2);
			46743: out = 16'(-74);
			46744: out = 16'(-54);
			46745: out = 16'(-170);
			46746: out = 16'(-432);
			46747: out = 16'(-448);
			46748: out = 16'(-364);
			46749: out = 16'(-97);
			46750: out = 16'(59);
			46751: out = 16'(117);
			46752: out = 16'(71);
			46753: out = 16'(-189);
			46754: out = 16'(-419);
			46755: out = 16'(-41);
			46756: out = 16'(173);
			46757: out = 16'(390);
			46758: out = 16'(364);
			46759: out = 16'(288);
			46760: out = 16'(88);
			46761: out = 16'(64);
			46762: out = 16'(-122);
			46763: out = 16'(-448);
			46764: out = 16'(-265);
			46765: out = 16'(-74);
			46766: out = 16'(191);
			46767: out = 16'(117);
			46768: out = 16'(-1);
			46769: out = 16'(-57);
			46770: out = 16'(-96);
			46771: out = 16'(-50);
			46772: out = 16'(-21);
			46773: out = 16'(24);
			46774: out = 16'(36);
			46775: out = 16'(105);
			46776: out = 16'(67);
			46777: out = 16'(-79);
			46778: out = 16'(-69);
			46779: out = 16'(-109);
			46780: out = 16'(-158);
			46781: out = 16'(-236);
			46782: out = 16'(-230);
			46783: out = 16'(-163);
			46784: out = 16'(-36);
			46785: out = 16'(21);
			46786: out = 16'(-55);
			46787: out = 16'(2);
			46788: out = 16'(14);
			46789: out = 16'(16);
			46790: out = 16'(21);
			46791: out = 16'(38);
			46792: out = 16'(-35);
			46793: out = 16'(-90);
			46794: out = 16'(-165);
			46795: out = 16'(-83);
			46796: out = 16'(-31);
			46797: out = 16'(53);
			46798: out = 16'(-38);
			46799: out = 16'(-25);
			46800: out = 16'(9);
			46801: out = 16'(96);
			46802: out = 16'(96);
			46803: out = 16'(31);
			46804: out = 16'(-32);
			46805: out = 16'(-75);
			46806: out = 16'(9);
			46807: out = 16'(18);
			46808: out = 16'(46);
			46809: out = 16'(182);
			46810: out = 16'(115);
			46811: out = 16'(19);
			46812: out = 16'(1);
			46813: out = 16'(12);
			46814: out = 16'(22);
			46815: out = 16'(35);
			46816: out = 16'(-69);
			46817: out = 16'(-269);
			46818: out = 16'(-315);
			46819: out = 16'(-321);
			46820: out = 16'(-153);
			46821: out = 16'(-101);
			46822: out = 16'(-80);
			46823: out = 16'(-251);
			46824: out = 16'(-133);
			46825: out = 16'(-56);
			46826: out = 16'(-29);
			46827: out = 16'(-45);
			46828: out = 16'(-49);
			46829: out = 16'(10);
			46830: out = 16'(27);
			46831: out = 16'(11);
			46832: out = 16'(-52);
			46833: out = 16'(-51);
			46834: out = 16'(-38);
			46835: out = 16'(-44);
			46836: out = 16'(-28);
			46837: out = 16'(-32);
			46838: out = 16'(-3);
			46839: out = 16'(7);
			46840: out = 16'(-76);
			46841: out = 16'(11);
			46842: out = 16'(69);
			46843: out = 16'(208);
			46844: out = 16'(68);
			46845: out = 16'(-63);
			46846: out = 16'(-72);
			46847: out = 16'(-60);
			46848: out = 16'(-38);
			46849: out = 16'(-48);
			46850: out = 16'(-78);
			46851: out = 16'(-169);
			46852: out = 16'(-86);
			46853: out = 16'(-36);
			46854: out = 16'(19);
			46855: out = 16'(-52);
			46856: out = 16'(-94);
			46857: out = 16'(-156);
			46858: out = 16'(-93);
			46859: out = 16'(-23);
			46860: out = 16'(124);
			46861: out = 16'(78);
			46862: out = 16'(37);
			46863: out = 16'(19);
			46864: out = 16'(-21);
			46865: out = 16'(-22);
			46866: out = 16'(189);
			46867: out = 16'(131);
			46868: out = 16'(20);
			46869: out = 16'(98);
			46870: out = 16'(99);
			46871: out = 16'(113);
			46872: out = 16'(23);
			46873: out = 16'(-4);
			46874: out = 16'(0);
			46875: out = 16'(-50);
			46876: out = 16'(-57);
			46877: out = 16'(35);
			46878: out = 16'(-36);
			46879: out = 16'(-69);
			46880: out = 16'(-92);
			46881: out = 16'(-31);
			46882: out = 16'(-9);
			46883: out = 16'(28);
			46884: out = 16'(-21);
			46885: out = 16'(-75);
			46886: out = 16'(-93);
			46887: out = 16'(-38);
			46888: out = 16'(18);
			46889: out = 16'(-63);
			46890: out = 16'(-151);
			46891: out = 16'(-290);
			46892: out = 16'(-116);
			46893: out = 16'(-74);
			46894: out = 16'(-77);
			46895: out = 16'(-8);
			46896: out = 16'(57);
			46897: out = 16'(196);
			46898: out = 16'(43);
			46899: out = 16'(-93);
			46900: out = 16'(-174);
			46901: out = 16'(-175);
			46902: out = 16'(-181);
			46903: out = 16'(-252);
			46904: out = 16'(-288);
			46905: out = 16'(-338);
			46906: out = 16'(-111);
			46907: out = 16'(0);
			46908: out = 16'(39);
			46909: out = 16'(54);
			46910: out = 16'(-47);
			46911: out = 16'(-245);
			46912: out = 16'(-312);
			46913: out = 16'(-280);
			46914: out = 16'(-35);
			46915: out = 16'(-46);
			46916: out = 16'(-17);
			46917: out = 16'(-32);
			46918: out = 16'(-29);
			46919: out = 16'(-12);
			46920: out = 16'(52);
			46921: out = 16'(35);
			46922: out = 16'(30);
			46923: out = 16'(48);
			46924: out = 16'(84);
			46925: out = 16'(123);
			46926: out = 16'(42);
			46927: out = 16'(-16);
			46928: out = 16'(-67);
			46929: out = 16'(81);
			46930: out = 16'(159);
			46931: out = 16'(190);
			46932: out = 16'(79);
			46933: out = 16'(23);
			46934: out = 16'(38);
			46935: out = 16'(26);
			46936: out = 16'(5);
			46937: out = 16'(-60);
			46938: out = 16'(41);
			46939: out = 16'(121);
			46940: out = 16'(5);
			46941: out = 16'(-10);
			46942: out = 16'(-73);
			46943: out = 16'(21);
			46944: out = 16'(-145);
			46945: out = 16'(-383);
			46946: out = 16'(-429);
			46947: out = 16'(-350);
			46948: out = 16'(-129);
			46949: out = 16'(-87);
			46950: out = 16'(6);
			46951: out = 16'(25);
			46952: out = 16'(115);
			46953: out = 16'(88);
			46954: out = 16'(39);
			46955: out = 16'(-206);
			46956: out = 16'(-331);
			46957: out = 16'(-151);
			46958: out = 16'(-120);
			46959: out = 16'(-45);
			46960: out = 16'(-78);
			46961: out = 16'(-11);
			46962: out = 16'(20);
			46963: out = 16'(-34);
			46964: out = 16'(3);
			46965: out = 16'(57);
			46966: out = 16'(102);
			46967: out = 16'(130);
			46968: out = 16'(122);
			46969: out = 16'(85);
			46970: out = 16'(-28);
			46971: out = 16'(-157);
			46972: out = 16'(-269);
			46973: out = 16'(-304);
			46974: out = 16'(-65);
			46975: out = 16'(-50);
			46976: out = 16'(-22);
			46977: out = 16'(-60);
			46978: out = 16'(62);
			46979: out = 16'(122);
			46980: out = 16'(71);
			46981: out = 16'(-56);
			46982: out = 16'(-161);
			46983: out = 16'(-247);
			46984: out = 16'(-175);
			46985: out = 16'(-59);
			46986: out = 16'(6);
			46987: out = 16'(-14);
			46988: out = 16'(-151);
			46989: out = 16'(-228);
			46990: out = 16'(-161);
			46991: out = 16'(53);
			46992: out = 16'(255);
			46993: out = 16'(374);
			46994: out = 16'(270);
			46995: out = 16'(125);
			46996: out = 16'(-82);
			46997: out = 16'(135);
			46998: out = 16'(30);
			46999: out = 16'(-61);
			47000: out = 16'(-78);
			47001: out = 16'(-43);
			47002: out = 16'(7);
			47003: out = 16'(-142);
			47004: out = 16'(-116);
			47005: out = 16'(23);
			47006: out = 16'(143);
			47007: out = 16'(225);
			47008: out = 16'(244);
			47009: out = 16'(278);
			47010: out = 16'(212);
			47011: out = 16'(105);
			47012: out = 16'(-74);
			47013: out = 16'(-227);
			47014: out = 16'(-354);
			47015: out = 16'(-364);
			47016: out = 16'(-373);
			47017: out = 16'(-431);
			47018: out = 16'(-393);
			47019: out = 16'(-319);
			47020: out = 16'(-265);
			47021: out = 16'(-160);
			47022: out = 16'(-45);
			47023: out = 16'(10);
			47024: out = 16'(17);
			47025: out = 16'(-66);
			47026: out = 16'(-17);
			47027: out = 16'(-24);
			47028: out = 16'(78);
			47029: out = 16'(-80);
			47030: out = 16'(-195);
			47031: out = 16'(-412);
			47032: out = 16'(-164);
			47033: out = 16'(115);
			47034: out = 16'(346);
			47035: out = 16'(388);
			47036: out = 16'(349);
			47037: out = 16'(365);
			47038: out = 16'(314);
			47039: out = 16'(254);
			47040: out = 16'(133);
			47041: out = 16'(58);
			47042: out = 16'(-25);
			47043: out = 16'(2);
			47044: out = 16'(-8);
			47045: out = 16'(20);
			47046: out = 16'(8);
			47047: out = 16'(9);
			47048: out = 16'(4);
			47049: out = 16'(26);
			47050: out = 16'(-7);
			47051: out = 16'(21);
			47052: out = 16'(-228);
			47053: out = 16'(-384);
			47054: out = 16'(-355);
			47055: out = 16'(-307);
			47056: out = 16'(-264);
			47057: out = 16'(-239);
			47058: out = 16'(-324);
			47059: out = 16'(-420);
			47060: out = 16'(-431);
			47061: out = 16'(-289);
			47062: out = 16'(-6);
			47063: out = 16'(32);
			47064: out = 16'(51);
			47065: out = 16'(-61);
			47066: out = 16'(-19);
			47067: out = 16'(17);
			47068: out = 16'(306);
			47069: out = 16'(208);
			47070: out = 16'(72);
			47071: out = 16'(-214);
			47072: out = 16'(-249);
			47073: out = 16'(-229);
			47074: out = 16'(-309);
			47075: out = 16'(-236);
			47076: out = 16'(-93);
			47077: out = 16'(176);
			47078: out = 16'(281);
			47079: out = 16'(291);
			47080: out = 16'(170);
			47081: out = 16'(123);
			47082: out = 16'(151);
			47083: out = 16'(4);
			47084: out = 16'(-44);
			47085: out = 16'(-70);
			47086: out = 16'(-117);
			47087: out = 16'(-159);
			47088: out = 16'(-137);
			47089: out = 16'(-141);
			47090: out = 16'(-125);
			47091: out = 16'(17);
			47092: out = 16'(13);
			47093: out = 16'(-37);
			47094: out = 16'(-29);
			47095: out = 16'(-41);
			47096: out = 16'(-21);
			47097: out = 16'(35);
			47098: out = 16'(-22);
			47099: out = 16'(-171);
			47100: out = 16'(12);
			47101: out = 16'(36);
			47102: out = 16'(61);
			47103: out = 16'(-11);
			47104: out = 16'(-12);
			47105: out = 16'(28);
			47106: out = 16'(204);
			47107: out = 16'(250);
			47108: out = 16'(-28);
			47109: out = 16'(-98);
			47110: out = 16'(-163);
			47111: out = 16'(-29);
			47112: out = 16'(-50);
			47113: out = 16'(-37);
			47114: out = 16'(-60);
			47115: out = 16'(-52);
			47116: out = 16'(-22);
			47117: out = 16'(141);
			47118: out = 16'(282);
			47119: out = 16'(425);
			47120: out = 16'(431);
			47121: out = 16'(307);
			47122: out = 16'(8);
			47123: out = 16'(-107);
			47124: out = 16'(-226);
			47125: out = 16'(-252);
			47126: out = 16'(-326);
			47127: out = 16'(-365);
			47128: out = 16'(-425);
			47129: out = 16'(-475);
			47130: out = 16'(-499);
			47131: out = 16'(-356);
			47132: out = 16'(-237);
			47133: out = 16'(-126);
			47134: out = 16'(-208);
			47135: out = 16'(-155);
			47136: out = 16'(-24);
			47137: out = 16'(96);
			47138: out = 16'(213);
			47139: out = 16'(306);
			47140: out = 16'(143);
			47141: out = 16'(21);
			47142: out = 16'(59);
			47143: out = 16'(-99);
			47144: out = 16'(-103);
			47145: out = 16'(28);
			47146: out = 16'(186);
			47147: out = 16'(305);
			47148: out = 16'(288);
			47149: out = 16'(203);
			47150: out = 16'(88);
			47151: out = 16'(-29);
			47152: out = 16'(-163);
			47153: out = 16'(-254);
			47154: out = 16'(-37);
			47155: out = 16'(31);
			47156: out = 16'(30);
			47157: out = 16'(23);
			47158: out = 16'(-7);
			47159: out = 16'(-9);
			47160: out = 16'(-31);
			47161: out = 16'(-54);
			47162: out = 16'(9);
			47163: out = 16'(-112);
			47164: out = 16'(-175);
			47165: out = 16'(-178);
			47166: out = 16'(-134);
			47167: out = 16'(-75);
			47168: out = 16'(-158);
			47169: out = 16'(-205);
			47170: out = 16'(-263);
			47171: out = 16'(-248);
			47172: out = 16'(-184);
			47173: out = 16'(-41);
			47174: out = 16'(-62);
			47175: out = 16'(1);
			47176: out = 16'(43);
			47177: out = 16'(165);
			47178: out = 16'(186);
			47179: out = 16'(31);
			47180: out = 16'(-21);
			47181: out = 16'(-86);
			47182: out = 16'(-57);
			47183: out = 16'(-90);
			47184: out = 16'(-70);
			47185: out = 16'(-253);
			47186: out = 16'(-131);
			47187: out = 16'(-9);
			47188: out = 16'(247);
			47189: out = 16'(210);
			47190: out = 16'(0);
			47191: out = 16'(59);
			47192: out = 16'(-4);
			47193: out = 16'(-39);
			47194: out = 16'(-76);
			47195: out = 16'(34);
			47196: out = 16'(291);
			47197: out = 16'(50);
			47198: out = 16'(-140);
			47199: out = 16'(-322);
			47200: out = 16'(-361);
			47201: out = 16'(-306);
			47202: out = 16'(-177);
			47203: out = 16'(-83);
			47204: out = 16'(-24);
			47205: out = 16'(37);
			47206: out = 16'(11);
			47207: out = 16'(-38);
			47208: out = 16'(110);
			47209: out = 16'(167);
			47210: out = 16'(180);
			47211: out = 16'(74);
			47212: out = 16'(22);
			47213: out = 16'(12);
			47214: out = 16'(-126);
			47215: out = 16'(-137);
			47216: out = 16'(10);
			47217: out = 16'(21);
			47218: out = 16'(44);
			47219: out = 16'(15);
			47220: out = 16'(-9);
			47221: out = 16'(-73);
			47222: out = 16'(-59);
			47223: out = 16'(-225);
			47224: out = 16'(-358);
			47225: out = 16'(-334);
			47226: out = 16'(-272);
			47227: out = 16'(-124);
			47228: out = 16'(-75);
			47229: out = 16'(100);
			47230: out = 16'(297);
			47231: out = 16'(164);
			47232: out = 16'(81);
			47233: out = 16'(18);
			47234: out = 16'(-34);
			47235: out = 16'(-26);
			47236: out = 16'(35);
			47237: out = 16'(-20);
			47238: out = 16'(-63);
			47239: out = 16'(-64);
			47240: out = 16'(-130);
			47241: out = 16'(-176);
			47242: out = 16'(-258);
			47243: out = 16'(-158);
			47244: out = 16'(-26);
			47245: out = 16'(245);
			47246: out = 16'(318);
			47247: out = 16'(343);
			47248: out = 16'(59);
			47249: out = 16'(-24);
			47250: out = 16'(-64);
			47251: out = 16'(139);
			47252: out = 16'(124);
			47253: out = 16'(-61);
			47254: out = 16'(-207);
			47255: out = 16'(-220);
			47256: out = 16'(0);
			47257: out = 16'(167);
			47258: out = 16'(252);
			47259: out = 16'(113);
			47260: out = 16'(4);
			47261: out = 16'(-138);
			47262: out = 16'(-321);
			47263: out = 16'(-316);
			47264: out = 16'(-247);
			47265: out = 16'(-104);
			47266: out = 16'(-136);
			47267: out = 16'(-258);
			47268: out = 16'(-389);
			47269: out = 16'(-326);
			47270: out = 16'(-34);
			47271: out = 16'(52);
			47272: out = 16'(190);
			47273: out = 16'(195);
			47274: out = 16'(159);
			47275: out = 16'(84);
			47276: out = 16'(-51);
			47277: out = 16'(0);
			47278: out = 16'(82);
			47279: out = 16'(253);
			47280: out = 16'(206);
			47281: out = 16'(54);
			47282: out = 16'(-104);
			47283: out = 16'(-305);
			47284: out = 16'(-430);
			47285: out = 16'(-226);
			47286: out = 16'(-23);
			47287: out = 16'(111);
			47288: out = 16'(257);
			47289: out = 16'(183);
			47290: out = 16'(-90);
			47291: out = 16'(-207);
			47292: out = 16'(-213);
			47293: out = 16'(18);
			47294: out = 16'(-46);
			47295: out = 16'(-78);
			47296: out = 16'(-66);
			47297: out = 16'(-124);
			47298: out = 16'(-172);
			47299: out = 16'(-324);
			47300: out = 16'(-176);
			47301: out = 16'(55);
			47302: out = 16'(29);
			47303: out = 16'(25);
			47304: out = 16'(-54);
			47305: out = 16'(116);
			47306: out = 16'(81);
			47307: out = 16'(19);
			47308: out = 16'(-313);
			47309: out = 16'(-449);
			47310: out = 16'(-386);
			47311: out = 16'(-385);
			47312: out = 16'(-225);
			47313: out = 16'(-52);
			47314: out = 16'(330);
			47315: out = 16'(568);
			47316: out = 16'(567);
			47317: out = 16'(505);
			47318: out = 16'(386);
			47319: out = 16'(226);
			47320: out = 16'(58);
			47321: out = 16'(-90);
			47322: out = 16'(-71);
			47323: out = 16'(-177);
			47324: out = 16'(-257);
			47325: out = 16'(-345);
			47326: out = 16'(-272);
			47327: out = 16'(-79);
			47328: out = 16'(128);
			47329: out = 16'(174);
			47330: out = 16'(34);
			47331: out = 16'(-209);
			47332: out = 16'(-404);
			47333: out = 16'(-509);
			47334: out = 16'(-334);
			47335: out = 16'(-77);
			47336: out = 16'(14);
			47337: out = 16'(79);
			47338: out = 16'(38);
			47339: out = 16'(38);
			47340: out = 16'(9);
			47341: out = 16'(32);
			47342: out = 16'(19);
			47343: out = 16'(108);
			47344: out = 16'(200);
			47345: out = 16'(310);
			47346: out = 16'(361);
			47347: out = 16'(411);
			47348: out = 16'(252);
			47349: out = 16'(89);
			47350: out = 16'(-65);
			47351: out = 16'(-102);
			47352: out = 16'(-128);
			47353: out = 16'(-289);
			47354: out = 16'(-193);
			47355: out = 16'(-50);
			47356: out = 16'(66);
			47357: out = 16'(140);
			47358: out = 16'(145);
			47359: out = 16'(91);
			47360: out = 16'(7);
			47361: out = 16'(-86);
			47362: out = 16'(-44);
			47363: out = 16'(-70);
			47364: out = 16'(-169);
			47365: out = 16'(-144);
			47366: out = 16'(-186);
			47367: out = 16'(-276);
			47368: out = 16'(-336);
			47369: out = 16'(-281);
			47370: out = 16'(-82);
			47371: out = 16'(-47);
			47372: out = 16'(-43);
			47373: out = 16'(-21);
			47374: out = 16'(-44);
			47375: out = 16'(-73);
			47376: out = 16'(-69);
			47377: out = 16'(-41);
			47378: out = 16'(-28);
			47379: out = 16'(-100);
			47380: out = 16'(-203);
			47381: out = 16'(-324);
			47382: out = 16'(-331);
			47383: out = 16'(-226);
			47384: out = 16'(26);
			47385: out = 16'(1);
			47386: out = 16'(50);
			47387: out = 16'(67);
			47388: out = 16'(129);
			47389: out = 16'(142);
			47390: out = 16'(118);
			47391: out = 16'(100);
			47392: out = 16'(48);
			47393: out = 16'(11);
			47394: out = 16'(-33);
			47395: out = 16'(-77);
			47396: out = 16'(-60);
			47397: out = 16'(-81);
			47398: out = 16'(-54);
			47399: out = 16'(-43);
			47400: out = 16'(-31);
			47401: out = 16'(-5);
			47402: out = 16'(-9);
			47403: out = 16'(45);
			47404: out = 16'(121);
			47405: out = 16'(155);
			47406: out = 16'(141);
			47407: out = 16'(-4);
			47408: out = 16'(-120);
			47409: out = 16'(-226);
			47410: out = 16'(-199);
			47411: out = 16'(-140);
			47412: out = 16'(-53);
			47413: out = 16'(-41);
			47414: out = 16'(82);
			47415: out = 16'(182);
			47416: out = 16'(176);
			47417: out = 16'(89);
			47418: out = 16'(-32);
			47419: out = 16'(-64);
			47420: out = 16'(-102);
			47421: out = 16'(-78);
			47422: out = 16'(-126);
			47423: out = 16'(-151);
			47424: out = 16'(-146);
			47425: out = 16'(-104);
			47426: out = 16'(-38);
			47427: out = 16'(46);
			47428: out = 16'(121);
			47429: out = 16'(182);
			47430: out = 16'(92);
			47431: out = 16'(162);
			47432: out = 16'(203);
			47433: out = 16'(177);
			47434: out = 16'(21);
			47435: out = 16'(-202);
			47436: out = 16'(-309);
			47437: out = 16'(-343);
			47438: out = 16'(-268);
			47439: out = 16'(-391);
			47440: out = 16'(-368);
			47441: out = 16'(-327);
			47442: out = 16'(-133);
			47443: out = 16'(-8);
			47444: out = 16'(80);
			47445: out = 16'(36);
			47446: out = 16'(4);
			47447: out = 16'(-46);
			47448: out = 16'(-62);
			47449: out = 16'(-51);
			47450: out = 16'(-106);
			47451: out = 16'(-167);
			47452: out = 16'(-173);
			47453: out = 16'(-86);
			47454: out = 16'(99);
			47455: out = 16'(246);
			47456: out = 16'(238);
			47457: out = 16'(160);
			47458: out = 16'(-28);
			47459: out = 16'(-101);
			47460: out = 16'(-140);
			47461: out = 16'(-61);
			47462: out = 16'(-85);
			47463: out = 16'(-54);
			47464: out = 16'(-92);
			47465: out = 16'(13);
			47466: out = 16'(84);
			47467: out = 16'(171);
			47468: out = 16'(113);
			47469: out = 16'(23);
			47470: out = 16'(-57);
			47471: out = 16'(-120);
			47472: out = 16'(-123);
			47473: out = 16'(-60);
			47474: out = 16'(16);
			47475: out = 16'(55);
			47476: out = 16'(67);
			47477: out = 16'(16);
			47478: out = 16'(-12);
			47479: out = 16'(-255);
			47480: out = 16'(-354);
			47481: out = 16'(-334);
			47482: out = 16'(-155);
			47483: out = 16'(-40);
			47484: out = 16'(-11);
			47485: out = 16'(-73);
			47486: out = 16'(-125);
			47487: out = 16'(-73);
			47488: out = 16'(0);
			47489: out = 16'(77);
			47490: out = 16'(-33);
			47491: out = 16'(-100);
			47492: out = 16'(-203);
			47493: out = 16'(-239);
			47494: out = 16'(-209);
			47495: out = 16'(-97);
			47496: out = 16'(-22);
			47497: out = 16'(14);
			47498: out = 16'(10);
			47499: out = 16'(71);
			47500: out = 16'(82);
			47501: out = 16'(87);
			47502: out = 16'(34);
			47503: out = 16'(-6);
			47504: out = 16'(-36);
			47505: out = 16'(-10);
			47506: out = 16'(30);
			47507: out = 16'(122);
			47508: out = 16'(96);
			47509: out = 16'(46);
			47510: out = 16'(31);
			47511: out = 16'(-39);
			47512: out = 16'(-70);
			47513: out = 16'(-29);
			47514: out = 16'(-10);
			47515: out = 16'(1);
			47516: out = 16'(43);
			47517: out = 16'(77);
			47518: out = 16'(106);
			47519: out = 16'(-2);
			47520: out = 16'(-101);
			47521: out = 16'(-188);
			47522: out = 16'(-227);
			47523: out = 16'(-155);
			47524: out = 16'(47);
			47525: out = 16'(109);
			47526: out = 16'(114);
			47527: out = 16'(-6);
			47528: out = 16'(-41);
			47529: out = 16'(-79);
			47530: out = 16'(-66);
			47531: out = 16'(-97);
			47532: out = 16'(-138);
			47533: out = 16'(-134);
			47534: out = 16'(-87);
			47535: out = 16'(-5);
			47536: out = 16'(7);
			47537: out = 16'(0);
			47538: out = 16'(0);
			47539: out = 16'(-128);
			47540: out = 16'(-165);
			47541: out = 16'(9);
			47542: out = 16'(90);
			47543: out = 16'(183);
			47544: out = 16'(9);
			47545: out = 16'(-24);
			47546: out = 16'(-96);
			47547: out = 16'(-106);
			47548: out = 16'(-199);
			47549: out = 16'(-251);
			47550: out = 16'(-101);
			47551: out = 16'(-33);
			47552: out = 16'(16);
			47553: out = 16'(-33);
			47554: out = 16'(-52);
			47555: out = 16'(-55);
			47556: out = 16'(38);
			47557: out = 16'(97);
			47558: out = 16'(181);
			47559: out = 16'(73);
			47560: out = 16'(-25);
			47561: out = 16'(-109);
			47562: out = 16'(-186);
			47563: out = 16'(-186);
			47564: out = 16'(-195);
			47565: out = 16'(-152);
			47566: out = 16'(-115);
			47567: out = 16'(-76);
			47568: out = 16'(-38);
			47569: out = 16'(14);
			47570: out = 16'(-35);
			47571: out = 16'(-28);
			47572: out = 16'(29);
			47573: out = 16'(-36);
			47574: out = 16'(-86);
			47575: out = 16'(-119);
			47576: out = 16'(-61);
			47577: out = 16'(-32);
			47578: out = 16'(-44);
			47579: out = 16'(-29);
			47580: out = 16'(-47);
			47581: out = 16'(-39);
			47582: out = 16'(-17);
			47583: out = 16'(33);
			47584: out = 16'(65);
			47585: out = 16'(107);
			47586: out = 16'(114);
			47587: out = 16'(36);
			47588: out = 16'(-39);
			47589: out = 16'(-130);
			47590: out = 16'(-179);
			47591: out = 16'(-137);
			47592: out = 16'(-1);
			47593: out = 16'(41);
			47594: out = 16'(94);
			47595: out = 16'(131);
			47596: out = 16'(46);
			47597: out = 16'(-16);
			47598: out = 16'(-57);
			47599: out = 16'(-70);
			47600: out = 16'(-74);
			47601: out = 16'(-42);
			47602: out = 16'(-112);
			47603: out = 16'(-196);
			47604: out = 16'(-245);
			47605: out = 16'(-206);
			47606: out = 16'(-105);
			47607: out = 16'(-135);
			47608: out = 16'(-95);
			47609: out = 16'(-58);
			47610: out = 16'(-19);
			47611: out = 16'(5);
			47612: out = 16'(2);
			47613: out = 16'(42);
			47614: out = 16'(102);
			47615: out = 16'(242);
			47616: out = 16'(135);
			47617: out = 16'(44);
			47618: out = 16'(-9);
			47619: out = 16'(-59);
			47620: out = 16'(-67);
			47621: out = 16'(-79);
			47622: out = 16'(-55);
			47623: out = 16'(-10);
			47624: out = 16'(-61);
			47625: out = 16'(-1);
			47626: out = 16'(65);
			47627: out = 16'(241);
			47628: out = 16'(227);
			47629: out = 16'(36);
			47630: out = 16'(-33);
			47631: out = 16'(-82);
			47632: out = 16'(-22);
			47633: out = 16'(-26);
			47634: out = 16'(-57);
			47635: out = 16'(-213);
			47636: out = 16'(-236);
			47637: out = 16'(-259);
			47638: out = 16'(-76);
			47639: out = 16'(-79);
			47640: out = 16'(-49);
			47641: out = 16'(-44);
			47642: out = 16'(-72);
			47643: out = 16'(-73);
			47644: out = 16'(-178);
			47645: out = 16'(-179);
			47646: out = 16'(-122);
			47647: out = 16'(-90);
			47648: out = 16'(-49);
			47649: out = 16'(-70);
			47650: out = 16'(-9);
			47651: out = 16'(0);
			47652: out = 16'(6);
			47653: out = 16'(84);
			47654: out = 16'(155);
			47655: out = 16'(220);
			47656: out = 16'(232);
			47657: out = 16'(192);
			47658: out = 16'(2);
			47659: out = 16'(-119);
			47660: out = 16'(-216);
			47661: out = 16'(-91);
			47662: out = 16'(-64);
			47663: out = 16'(-62);
			47664: out = 16'(-27);
			47665: out = 16'(29);
			47666: out = 16'(38);
			47667: out = 16'(115);
			47668: out = 16'(75);
			47669: out = 16'(-23);
			47670: out = 16'(-192);
			47671: out = 16'(-284);
			47672: out = 16'(-205);
			47673: out = 16'(-127);
			47674: out = 16'(-25);
			47675: out = 16'(0);
			47676: out = 16'(-28);
			47677: out = 16'(-73);
			47678: out = 16'(-60);
			47679: out = 16'(-106);
			47680: out = 16'(-120);
			47681: out = 16'(-78);
			47682: out = 16'(-21);
			47683: out = 16'(10);
			47684: out = 16'(10);
			47685: out = 16'(-21);
			47686: out = 16'(-35);
			47687: out = 16'(-126);
			47688: out = 16'(-134);
			47689: out = 16'(-133);
			47690: out = 16'(-46);
			47691: out = 16'(-13);
			47692: out = 16'(-70);
			47693: out = 16'(-129);
			47694: out = 16'(-189);
			47695: out = 16'(-125);
			47696: out = 16'(-59);
			47697: out = 16'(27);
			47698: out = 16'(2);
			47699: out = 16'(56);
			47700: out = 16'(71);
			47701: out = 16'(122);
			47702: out = 16'(82);
			47703: out = 16'(-15);
			47704: out = 16'(-255);
			47705: out = 16'(-317);
			47706: out = 16'(-237);
			47707: out = 16'(-188);
			47708: out = 16'(-57);
			47709: out = 16'(12);
			47710: out = 16'(134);
			47711: out = 16'(179);
			47712: out = 16'(21);
			47713: out = 16'(-28);
			47714: out = 16'(-54);
			47715: out = 16'(14);
			47716: out = 16'(-18);
			47717: out = 16'(-66);
			47718: out = 16'(-220);
			47719: out = 16'(-231);
			47720: out = 16'(-170);
			47721: out = 16'(-87);
			47722: out = 16'(-12);
			47723: out = 16'(30);
			47724: out = 16'(119);
			47725: out = 16'(122);
			47726: out = 16'(75);
			47727: out = 16'(1);
			47728: out = 16'(-39);
			47729: out = 16'(12);
			47730: out = 16'(-70);
			47731: out = 16'(-118);
			47732: out = 16'(-78);
			47733: out = 16'(-16);
			47734: out = 16'(5);
			47735: out = 16'(0);
			47736: out = 16'(-16);
			47737: out = 16'(-48);
			47738: out = 16'(-47);
			47739: out = 16'(-31);
			47740: out = 16'(-41);
			47741: out = 16'(93);
			47742: out = 16'(137);
			47743: out = 16'(130);
			47744: out = 16'(0);
			47745: out = 16'(-114);
			47746: out = 16'(-188);
			47747: out = 16'(-116);
			47748: out = 16'(-54);
			47749: out = 16'(-72);
			47750: out = 16'(-47);
			47751: out = 16'(-12);
			47752: out = 16'(162);
			47753: out = 16'(187);
			47754: out = 16'(176);
			47755: out = 16'(17);
			47756: out = 16'(-26);
			47757: out = 16'(-57);
			47758: out = 16'(-10);
			47759: out = 16'(-10);
			47760: out = 16'(-62);
			47761: out = 16'(-209);
			47762: out = 16'(-287);
			47763: out = 16'(-321);
			47764: out = 16'(-162);
			47765: out = 16'(7);
			47766: out = 16'(116);
			47767: out = 16'(108);
			47768: out = 16'(46);
			47769: out = 16'(13);
			47770: out = 16'(-110);
			47771: out = 16'(-196);
			47772: out = 16'(-74);
			47773: out = 16'(-26);
			47774: out = 16'(24);
			47775: out = 16'(-57);
			47776: out = 16'(-93);
			47777: out = 16'(-113);
			47778: out = 16'(-73);
			47779: out = 16'(-17);
			47780: out = 16'(18);
			47781: out = 16'(19);
			47782: out = 16'(12);
			47783: out = 16'(-2);
			47784: out = 16'(-8);
			47785: out = 16'(19);
			47786: out = 16'(115);
			47787: out = 16'(127);
			47788: out = 16'(110);
			47789: out = 16'(3);
			47790: out = 16'(-32);
			47791: out = 16'(-20);
			47792: out = 16'(-45);
			47793: out = 16'(-44);
			47794: out = 16'(2);
			47795: out = 16'(-48);
			47796: out = 16'(-60);
			47797: out = 16'(-11);
			47798: out = 16'(-165);
			47799: out = 16'(-226);
			47800: out = 16'(-339);
			47801: out = 16'(-157);
			47802: out = 16'(-29);
			47803: out = 16'(0);
			47804: out = 16'(-122);
			47805: out = 16'(-188);
			47806: out = 16'(-128);
			47807: out = 16'(-56);
			47808: out = 16'(6);
			47809: out = 16'(-44);
			47810: out = 16'(-2);
			47811: out = 16'(33);
			47812: out = 16'(45);
			47813: out = 16'(134);
			47814: out = 16'(248);
			47815: out = 16'(282);
			47816: out = 16'(217);
			47817: out = 16'(41);
			47818: out = 16'(-80);
			47819: out = 16'(-179);
			47820: out = 16'(-112);
			47821: out = 16'(-236);
			47822: out = 16'(-257);
			47823: out = 16'(-272);
			47824: out = 16'(-149);
			47825: out = 16'(-38);
			47826: out = 16'(-7);
			47827: out = 16'(1);
			47828: out = 16'(-14);
			47829: out = 16'(14);
			47830: out = 16'(19);
			47831: out = 16'(-2);
			47832: out = 16'(-41);
			47833: out = 16'(-138);
			47834: out = 16'(-263);
			47835: out = 16'(-205);
			47836: out = 16'(-127);
			47837: out = 16'(-44);
			47838: out = 16'(-51);
			47839: out = 16'(-37);
			47840: out = 16'(-121);
			47841: out = 16'(-108);
			47842: out = 16'(-117);
			47843: out = 16'(-56);
			47844: out = 16'(-90);
			47845: out = 16'(-106);
			47846: out = 16'(-185);
			47847: out = 16'(-75);
			47848: out = 16'(35);
			47849: out = 16'(64);
			47850: out = 16'(141);
			47851: out = 16'(202);
			47852: out = 16'(49);
			47853: out = 16'(-9);
			47854: out = 16'(-37);
			47855: out = 16'(5);
			47856: out = 16'(13);
			47857: out = 16'(-43);
			47858: out = 16'(-48);
			47859: out = 16'(-49);
			47860: out = 16'(-26);
			47861: out = 16'(-11);
			47862: out = 16'(43);
			47863: out = 16'(122);
			47864: out = 16'(92);
			47865: out = 16'(58);
			47866: out = 16'(14);
			47867: out = 16'(-22);
			47868: out = 16'(-16);
			47869: out = 16'(-46);
			47870: out = 16'(-46);
			47871: out = 16'(-42);
			47872: out = 16'(28);
			47873: out = 16'(112);
			47874: out = 16'(226);
			47875: out = 16'(114);
			47876: out = 16'(-21);
			47877: out = 16'(-201);
			47878: out = 16'(-165);
			47879: out = 16'(-142);
			47880: out = 16'(-130);
			47881: out = 16'(-136);
			47882: out = 16'(-132);
			47883: out = 16'(-21);
			47884: out = 16'(9);
			47885: out = 16'(23);
			47886: out = 16'(119);
			47887: out = 16'(64);
			47888: out = 16'(-9);
			47889: out = 16'(-102);
			47890: out = 16'(-186);
			47891: out = 16'(-262);
			47892: out = 16'(-65);
			47893: out = 16'(-11);
			47894: out = 16'(-51);
			47895: out = 16'(-67);
			47896: out = 16'(-45);
			47897: out = 16'(7);
			47898: out = 16'(15);
			47899: out = 16'(8);
			47900: out = 16'(0);
			47901: out = 16'(-123);
			47902: out = 16'(-204);
			47903: out = 16'(-254);
			47904: out = 16'(-127);
			47905: out = 16'(22);
			47906: out = 16'(110);
			47907: out = 16'(94);
			47908: out = 16'(-13);
			47909: out = 16'(-169);
			47910: out = 16'(-136);
			47911: out = 16'(14);
			47912: out = 16'(-47);
			47913: out = 16'(-122);
			47914: out = 16'(-328);
			47915: out = 16'(-304);
			47916: out = 16'(-277);
			47917: out = 16'(-174);
			47918: out = 16'(-78);
			47919: out = 16'(19);
			47920: out = 16'(122);
			47921: out = 16'(128);
			47922: out = 16'(72);
			47923: out = 16'(-5);
			47924: out = 16'(-23);
			47925: out = 16'(27);
			47926: out = 16'(76);
			47927: out = 16'(71);
			47928: out = 16'(24);
			47929: out = 16'(21);
			47930: out = 16'(-38);
			47931: out = 16'(-114);
			47932: out = 16'(-164);
			47933: out = 16'(-151);
			47934: out = 16'(-49);
			47935: out = 16'(-61);
			47936: out = 16'(-26);
			47937: out = 16'(0);
			47938: out = 16'(12);
			47939: out = 16'(5);
			47940: out = 16'(6);
			47941: out = 16'(2);
			47942: out = 16'(-6);
			47943: out = 16'(-104);
			47944: out = 16'(-65);
			47945: out = 16'(43);
			47946: out = 16'(105);
			47947: out = 16'(145);
			47948: out = 16'(113);
			47949: out = 16'(-5);
			47950: out = 16'(-115);
			47951: out = 16'(-177);
			47952: out = 16'(-206);
			47953: out = 16'(-155);
			47954: out = 16'(-126);
			47955: out = 16'(-27);
			47956: out = 16'(12);
			47957: out = 16'(-27);
			47958: out = 16'(-77);
			47959: out = 16'(-133);
			47960: out = 16'(-122);
			47961: out = 16'(-75);
			47962: out = 16'(-52);
			47963: out = 16'(30);
			47964: out = 16'(0);
			47965: out = 16'(-35);
			47966: out = 16'(-51);
			47967: out = 16'(-44);
			47968: out = 16'(-21);
			47969: out = 16'(47);
			47970: out = 16'(71);
			47971: out = 16'(15);
			47972: out = 16'(31);
			47973: out = 16'(13);
			47974: out = 16'(14);
			47975: out = 16'(17);
			47976: out = 16'(-8);
			47977: out = 16'(0);
			47978: out = 16'(-6);
			47979: out = 16'(-1);
			47980: out = 16'(-52);
			47981: out = 16'(-35);
			47982: out = 16'(-43);
			47983: out = 16'(-30);
			47984: out = 16'(-39);
			47985: out = 16'(-75);
			47986: out = 16'(-62);
			47987: out = 16'(-19);
			47988: out = 16'(19);
			47989: out = 16'(102);
			47990: out = 16'(129);
			47991: out = 16'(136);
			47992: out = 16'(20);
			47993: out = 16'(-66);
			47994: out = 16'(7);
			47995: out = 16'(-38);
			47996: out = 16'(-48);
			47997: out = 16'(0);
			47998: out = 16'(15);
			47999: out = 16'(-27);
			48000: out = 16'(-110);
			48001: out = 16'(-147);
			48002: out = 16'(-121);
			48003: out = 16'(-194);
			48004: out = 16'(-160);
			48005: out = 16'(-123);
			48006: out = 16'(-54);
			48007: out = 16'(-48);
			48008: out = 16'(-47);
			48009: out = 16'(-148);
			48010: out = 16'(-161);
			48011: out = 16'(-19);
			48012: out = 16'(-19);
			48013: out = 16'(41);
			48014: out = 16'(11);
			48015: out = 16'(31);
			48016: out = 16'(10);
			48017: out = 16'(14);
			48018: out = 16'(-84);
			48019: out = 16'(-181);
			48020: out = 16'(-4);
			48021: out = 16'(-7);
			48022: out = 16'(8);
			48023: out = 16'(-50);
			48024: out = 16'(-41);
			48025: out = 16'(28);
			48026: out = 16'(105);
			48027: out = 16'(109);
			48028: out = 16'(20);
			48029: out = 16'(-45);
			48030: out = 16'(-46);
			48031: out = 16'(-9);
			48032: out = 16'(3);
			48033: out = 16'(11);
			48034: out = 16'(-47);
			48035: out = 16'(-50);
			48036: out = 16'(-64);
			48037: out = 16'(14);
			48038: out = 16'(1);
			48039: out = 16'(14);
			48040: out = 16'(-204);
			48041: out = 16'(-293);
			48042: out = 16'(-304);
			48043: out = 16'(-313);
			48044: out = 16'(-254);
			48045: out = 16'(-28);
			48046: out = 16'(0);
			48047: out = 16'(3);
			48048: out = 16'(-124);
			48049: out = 16'(-24);
			48050: out = 16'(33);
			48051: out = 16'(145);
			48052: out = 16'(40);
			48053: out = 16'(-39);
			48054: out = 16'(-24);
			48055: out = 16'(29);
			48056: out = 16'(151);
			48057: out = 16'(77);
			48058: out = 16'(88);
			48059: out = 16'(70);
			48060: out = 16'(170);
			48061: out = 16'(143);
			48062: out = 16'(61);
			48063: out = 16'(25);
			48064: out = 16'(-14);
			48065: out = 16'(-58);
			48066: out = 16'(-74);
			48067: out = 16'(-57);
			48068: out = 16'(-12);
			48069: out = 16'(-26);
			48070: out = 16'(-21);
			48071: out = 16'(-150);
			48072: out = 16'(-68);
			48073: out = 16'(-3);
			48074: out = 16'(-14);
			48075: out = 16'(-91);
			48076: out = 16'(-223);
			48077: out = 16'(-177);
			48078: out = 16'(-182);
			48079: out = 16'(-116);
			48080: out = 16'(-188);
			48081: out = 16'(-150);
			48082: out = 16'(-51);
			48083: out = 16'(-24);
			48084: out = 16'(0);
			default: out = 0;
		endcase
	end
endmodule
