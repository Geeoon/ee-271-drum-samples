module open_hihat_lookup(index, out);
	input logic unsigned [12:0] index;
	output logic signed [15:0] out;
	always_comb begin
		case(index)
			0: out = 16'(0);
			1: out = 16'(210);
			2: out = 16'(426);
			3: out = 16'(775);
			4: out = 16'(-680);
			5: out = 16'(-24513);
			6: out = 16'(-7222);
			7: out = 16'(16446);
			8: out = 16'(11029);
			9: out = 16'(-14513);
			10: out = 16'(-7655);
			11: out = 16'(-7438);
			12: out = 16'(-7514);
			13: out = 16'(-4116);
			14: out = 16'(3581);
			15: out = 16'(-14156);
			16: out = 16'(-13716);
			17: out = 16'(-11132);
			18: out = 16'(-4441);
			19: out = 16'(-16318);
			20: out = 16'(-4714);
			21: out = 16'(898);
			22: out = 16'(3404);
			23: out = 16'(3352);
			24: out = 16'(-3418);
			25: out = 16'(-12889);
			26: out = 16'(4873);
			27: out = 16'(-3071);
			28: out = 16'(9156);
			29: out = 16'(25125);
			30: out = 16'(-17429);
			31: out = 16'(4691);
			32: out = 16'(4042);
			33: out = 16'(-5393);
			34: out = 16'(70);
			35: out = 16'(-8951);
			36: out = 16'(18295);
			37: out = 16'(-4335);
			38: out = 16'(-3027);
			39: out = 16'(16170);
			40: out = 16'(14447);
			41: out = 16'(-20155);
			42: out = 16'(710);
			43: out = 16'(-38);
			44: out = 16'(4186);
			45: out = 16'(7281);
			46: out = 16'(-19716);
			47: out = 16'(-17731);
			48: out = 16'(-16072);
			49: out = 16'(3013);
			50: out = 16'(1801);
			51: out = 16'(7567);
			52: out = 16'(-6729);
			53: out = 16'(577);
			54: out = 16'(-6227);
			55: out = 16'(29435);
			56: out = 16'(8913);
			57: out = 16'(24668);
			58: out = 16'(10903);
			59: out = 16'(-4099);
			60: out = 16'(-28925);
			61: out = 16'(-16457);
			62: out = 16'(-7727);
			63: out = 16'(-10172);
			64: out = 16'(18398);
			65: out = 16'(-8283);
			66: out = 16'(15586);
			67: out = 16'(12797);
			68: out = 16'(-7303);
			69: out = 16'(7744);
			70: out = 16'(-12778);
			71: out = 16'(1551);
			72: out = 16'(8020);
			73: out = 16'(-12665);
			74: out = 16'(-1501);
			75: out = 16'(-24511);
			76: out = 16'(-5456);
			77: out = 16'(11607);
			78: out = 16'(2132);
			79: out = 16'(-1479);
			80: out = 16'(9800);
			81: out = 16'(16486);
			82: out = 16'(-3931);
			83: out = 16'(74);
			84: out = 16'(10295);
			85: out = 16'(11521);
			86: out = 16'(21437);
			87: out = 16'(-29852);
			88: out = 16'(-27513);
			89: out = 16'(8790);
			90: out = 16'(-12426);
			91: out = 16'(-15958);
			92: out = 16'(8038);
			93: out = 16'(-14820);
			94: out = 16'(6424);
			95: out = 16'(-13523);
			96: out = 16'(25268);
			97: out = 16'(-15338);
			98: out = 16'(21207);
			99: out = 16'(16454);
			100: out = 16'(-9599);
			101: out = 16'(1759);
			102: out = 16'(9228);
			103: out = 16'(6351);
			104: out = 16'(-24674);
			105: out = 16'(21353);
			106: out = 16'(-3217);
			107: out = 16'(28842);
			108: out = 16'(-26367);
			109: out = 16'(684);
			110: out = 16'(10265);
			111: out = 16'(-7898);
			112: out = 16'(-6829);
			113: out = 16'(6221);
			114: out = 16'(-19207);
			115: out = 16'(12328);
			116: out = 16'(-18359);
			117: out = 16'(19903);
			118: out = 16'(5124);
			119: out = 16'(1451);
			120: out = 16'(-807);
			121: out = 16'(12310);
			122: out = 16'(1725);
			123: out = 16'(-2630);
			124: out = 16'(-4205);
			125: out = 16'(4279);
			126: out = 16'(-17281);
			127: out = 16'(6235);
			128: out = 16'(-3291);
			129: out = 16'(-7193);
			130: out = 16'(23886);
			131: out = 16'(870);
			132: out = 16'(26057);
			133: out = 16'(1512);
			134: out = 16'(4963);
			135: out = 16'(913);
			136: out = 16'(-1094);
			137: out = 16'(-12028);
			138: out = 16'(21427);
			139: out = 16'(5095);
			140: out = 16'(32173);
			141: out = 16'(28374);
			142: out = 16'(-15415);
			143: out = 16'(-5522);
			144: out = 16'(-12471);
			145: out = 16'(-26122);
			146: out = 16'(-23193);
			147: out = 16'(14769);
			148: out = 16'(-7209);
			149: out = 16'(20223);
			150: out = 16'(-4583);
			151: out = 16'(14177);
			152: out = 16'(-7334);
			153: out = 16'(12918);
			154: out = 16'(29059);
			155: out = 16'(9338);
			156: out = 16'(3394);
			157: out = 16'(-7337);
			158: out = 16'(-9398);
			159: out = 16'(2267);
			160: out = 16'(22873);
			161: out = 16'(-3467);
			162: out = 16'(-148);
			163: out = 16'(951);
			164: out = 16'(-8225);
			165: out = 16'(-6423);
			166: out = 16'(1917);
			167: out = 16'(6747);
			168: out = 16'(15440);
			169: out = 16'(13573);
			170: out = 16'(18141);
			171: out = 16'(4901);
			172: out = 16'(11765);
			173: out = 16'(11811);
			174: out = 16'(14070);
			175: out = 16'(14921);
			176: out = 16'(-17025);
			177: out = 16'(-20857);
			178: out = 16'(29888);
			179: out = 16'(-17411);
			180: out = 16'(-31351);
			181: out = 16'(28195);
			182: out = 16'(-4414);
			183: out = 16'(12041);
			184: out = 16'(2804);
			185: out = 16'(16826);
			186: out = 16'(-1995);
			187: out = 16'(-172);
			188: out = 16'(-1553);
			189: out = 16'(29449);
			190: out = 16'(-1254);
			191: out = 16'(-12404);
			192: out = 16'(-2375);
			193: out = 16'(-7274);
			194: out = 16'(-14352);
			195: out = 16'(13059);
			196: out = 16'(-1908);
			197: out = 16'(25263);
			198: out = 16'(-2490);
			199: out = 16'(-21087);
			200: out = 16'(30659);
			201: out = 16'(12929);
			202: out = 16'(2612);
			203: out = 16'(356);
			204: out = 16'(-4177);
			205: out = 16'(7376);
			206: out = 16'(13273);
			207: out = 16'(-4246);
			208: out = 16'(3368);
			209: out = 16'(-1412);
			210: out = 16'(-7941);
			211: out = 16'(2332);
			212: out = 16'(11594);
			213: out = 16'(-31725);
			214: out = 16'(-19816);
			215: out = 16'(-6235);
			216: out = 16'(-4099);
			217: out = 16'(-4754);
			218: out = 16'(11471);
			219: out = 16'(-3431);
			220: out = 16'(-4929);
			221: out = 16'(-24123);
			222: out = 16'(20163);
			223: out = 16'(2125);
			224: out = 16'(-1192);
			225: out = 16'(4874);
			226: out = 16'(8776);
			227: out = 16'(-27683);
			228: out = 16'(-15844);
			229: out = 16'(21236);
			230: out = 16'(-20626);
			231: out = 16'(-10957);
			232: out = 16'(-25393);
			233: out = 16'(17964);
			234: out = 16'(-5523);
			235: out = 16'(-3556);
			236: out = 16'(-28510);
			237: out = 16'(19292);
			238: out = 16'(-12510);
			239: out = 16'(-686);
			240: out = 16'(-1942);
			241: out = 16'(16958);
			242: out = 16'(-8239);
			243: out = 16'(-27104);
			244: out = 16'(5882);
			245: out = 16'(-9722);
			246: out = 16'(18748);
			247: out = 16'(3163);
			248: out = 16'(-11210);
			249: out = 16'(-12784);
			250: out = 16'(-3384);
			251: out = 16'(-20597);
			252: out = 16'(4142);
			253: out = 16'(-29415);
			254: out = 16'(20647);
			255: out = 16'(-14210);
			256: out = 16'(10004);
			257: out = 16'(-7222);
			258: out = 16'(13437);
			259: out = 16'(-11660);
			260: out = 16'(-5348);
			261: out = 16'(-9815);
			262: out = 16'(-31509);
			263: out = 16'(4775);
			264: out = 16'(-5904);
			265: out = 16'(-23802);
			266: out = 16'(-530);
			267: out = 16'(14737);
			268: out = 16'(-14229);
			269: out = 16'(4204);
			270: out = 16'(4505);
			271: out = 16'(-6542);
			272: out = 16'(18136);
			273: out = 16'(-13637);
			274: out = 16'(-14312);
			275: out = 16'(-847);
			276: out = 16'(9010);
			277: out = 16'(12095);
			278: out = 16'(-13980);
			279: out = 16'(-15425);
			280: out = 16'(-2914);
			281: out = 16'(8984);
			282: out = 16'(14196);
			283: out = 16'(-19114);
			284: out = 16'(-7798);
			285: out = 16'(20352);
			286: out = 16'(-12930);
			287: out = 16'(-24592);
			288: out = 16'(18046);
			289: out = 16'(4874);
			290: out = 16'(-181);
			291: out = 16'(21946);
			292: out = 16'(22324);
			293: out = 16'(-20009);
			294: out = 16'(19388);
			295: out = 16'(1981);
			296: out = 16'(-7643);
			297: out = 16'(17710);
			298: out = 16'(7770);
			299: out = 16'(8267);
			300: out = 16'(18802);
			301: out = 16'(17446);
			302: out = 16'(20988);
			303: out = 16'(11212);
			304: out = 16'(8298);
			305: out = 16'(-11131);
			306: out = 16'(4944);
			307: out = 16'(25905);
			308: out = 16'(-26644);
			309: out = 16'(-4637);
			310: out = 16'(-25741);
			311: out = 16'(17658);
			312: out = 16'(-3815);
			313: out = 16'(13834);
			314: out = 16'(15756);
			315: out = 16'(-26547);
			316: out = 16'(-12169);
			317: out = 16'(-22301);
			318: out = 16'(456);
			319: out = 16'(9708);
			320: out = 16'(-18977);
			321: out = 16'(-15235);
			322: out = 16'(9123);
			323: out = 16'(-11038);
			324: out = 16'(-9469);
			325: out = 16'(10682);
			326: out = 16'(6527);
			327: out = 16'(18229);
			328: out = 16'(-25509);
			329: out = 16'(-11001);
			330: out = 16'(11488);
			331: out = 16'(-26102);
			332: out = 16'(1909);
			333: out = 16'(24865);
			334: out = 16'(17402);
			335: out = 16'(3079);
			336: out = 16'(11222);
			337: out = 16'(11203);
			338: out = 16'(8750);
			339: out = 16'(22023);
			340: out = 16'(8340);
			341: out = 16'(0);
			342: out = 16'(-11556);
			343: out = 16'(-2160);
			344: out = 16'(-5740);
			345: out = 16'(-935);
			346: out = 16'(-21060);
			347: out = 16'(1955);
			348: out = 16'(-9653);
			349: out = 16'(16246);
			350: out = 16'(-25230);
			351: out = 16'(4166);
			352: out = 16'(-17731);
			353: out = 16'(3550);
			354: out = 16'(-5161);
			355: out = 16'(16080);
			356: out = 16'(1292);
			357: out = 16'(-14510);
			358: out = 16'(-21649);
			359: out = 16'(-1742);
			360: out = 16'(-538);
			361: out = 16'(-19150);
			362: out = 16'(21162);
			363: out = 16'(5161);
			364: out = 16'(-9890);
			365: out = 16'(855);
			366: out = 16'(17570);
			367: out = 16'(-4324);
			368: out = 16'(8311);
			369: out = 16'(-4925);
			370: out = 16'(-2984);
			371: out = 16'(12265);
			372: out = 16'(-8754);
			373: out = 16'(2330);
			374: out = 16'(4887);
			375: out = 16'(-6384);
			376: out = 16'(18476);
			377: out = 16'(-8015);
			378: out = 16'(-18963);
			379: out = 16'(12998);
			380: out = 16'(3354);
			381: out = 16'(-23322);
			382: out = 16'(5712);
			383: out = 16'(-2071);
			384: out = 16'(-6747);
			385: out = 16'(18313);
			386: out = 16'(-12305);
			387: out = 16'(1943);
			388: out = 16'(6542);
			389: out = 16'(11792);
			390: out = 16'(-11872);
			391: out = 16'(4853);
			392: out = 16'(6177);
			393: out = 16'(-4158);
			394: out = 16'(-28945);
			395: out = 16'(-10018);
			396: out = 16'(-512);
			397: out = 16'(-10507);
			398: out = 16'(7317);
			399: out = 16'(1003);
			400: out = 16'(-3576);
			401: out = 16'(-14400);
			402: out = 16'(-4465);
			403: out = 16'(6550);
			404: out = 16'(11030);
			405: out = 16'(-12802);
			406: out = 16'(18119);
			407: out = 16'(-2277);
			408: out = 16'(-9468);
			409: out = 16'(1509);
			410: out = 16'(7673);
			411: out = 16'(6476);
			412: out = 16'(16828);
			413: out = 16'(-7630);
			414: out = 16'(-25080);
			415: out = 16'(-9192);
			416: out = 16'(-11255);
			417: out = 16'(20469);
			418: out = 16'(-21803);
			419: out = 16'(-18225);
			420: out = 16'(1000);
			421: out = 16'(-7691);
			422: out = 16'(9521);
			423: out = 16'(-8553);
			424: out = 16'(-14483);
			425: out = 16'(3076);
			426: out = 16'(21950);
			427: out = 16'(-23585);
			428: out = 16'(6533);
			429: out = 16'(13959);
			430: out = 16'(-19812);
			431: out = 16'(10793);
			432: out = 16'(20276);
			433: out = 16'(-18702);
			434: out = 16'(342);
			435: out = 16'(5817);
			436: out = 16'(1106);
			437: out = 16'(7954);
			438: out = 16'(-22749);
			439: out = 16'(15651);
			440: out = 16'(28386);
			441: out = 16'(-20168);
			442: out = 16'(8702);
			443: out = 16'(-9273);
			444: out = 16'(-9490);
			445: out = 16'(-21634);
			446: out = 16'(25285);
			447: out = 16'(6440);
			448: out = 16'(-532);
			449: out = 16'(-5569);
			450: out = 16'(2619);
			451: out = 16'(10592);
			452: out = 16'(10873);
			453: out = 16'(-8966);
			454: out = 16'(17137);
			455: out = 16'(-10177);
			456: out = 16'(-2672);
			457: out = 16'(-1429);
			458: out = 16'(-8572);
			459: out = 16'(10880);
			460: out = 16'(7290);
			461: out = 16'(14553);
			462: out = 16'(15907);
			463: out = 16'(18352);
			464: out = 16'(-4118);
			465: out = 16'(5704);
			466: out = 16'(5521);
			467: out = 16'(1097);
			468: out = 16'(10752);
			469: out = 16'(25178);
			470: out = 16'(-3456);
			471: out = 16'(-17870);
			472: out = 16'(13389);
			473: out = 16'(6504);
			474: out = 16'(637);
			475: out = 16'(7934);
			476: out = 16'(23162);
			477: out = 16'(18141);
			478: out = 16'(-21631);
			479: out = 16'(-6805);
			480: out = 16'(1606);
			481: out = 16'(-1581);
			482: out = 16'(3321);
			483: out = 16'(16750);
			484: out = 16'(-2318);
			485: out = 16'(9271);
			486: out = 16'(-9968);
			487: out = 16'(-10785);
			488: out = 16'(12515);
			489: out = 16'(7089);
			490: out = 16'(7278);
			491: out = 16'(895);
			492: out = 16'(9144);
			493: out = 16'(894);
			494: out = 16'(3637);
			495: out = 16'(15496);
			496: out = 16'(-7057);
			497: out = 16'(-5316);
			498: out = 16'(-15510);
			499: out = 16'(1050);
			500: out = 16'(-11891);
			501: out = 16'(-11401);
			502: out = 16'(12050);
			503: out = 16'(2731);
			504: out = 16'(7109);
			505: out = 16'(-2561);
			506: out = 16'(-27315);
			507: out = 16'(-13546);
			508: out = 16'(2993);
			509: out = 16'(-2477);
			510: out = 16'(10049);
			511: out = 16'(-475);
			512: out = 16'(3916);
			513: out = 16'(14925);
			514: out = 16'(-2970);
			515: out = 16'(937);
			516: out = 16'(-2006);
			517: out = 16'(7107);
			518: out = 16'(21596);
			519: out = 16'(5185);
			520: out = 16'(-16039);
			521: out = 16'(2341);
			522: out = 16'(-316);
			523: out = 16'(-5022);
			524: out = 16'(11883);
			525: out = 16'(-8600);
			526: out = 16'(-6399);
			527: out = 16'(-2339);
			528: out = 16'(-11069);
			529: out = 16'(-32246);
			530: out = 16'(213);
			531: out = 16'(246);
			532: out = 16'(3076);
			533: out = 16'(11189);
			534: out = 16'(-1575);
			535: out = 16'(-8157);
			536: out = 16'(9965);
			537: out = 16'(7415);
			538: out = 16'(9355);
			539: out = 16'(16862);
			540: out = 16'(-14668);
			541: out = 16'(-13360);
			542: out = 16'(-30867);
			543: out = 16'(3604);
			544: out = 16'(-15132);
			545: out = 16'(20757);
			546: out = 16'(2749);
			547: out = 16'(-2090);
			548: out = 16'(-4489);
			549: out = 16'(-1304);
			550: out = 16'(-9144);
			551: out = 16'(-12295);
			552: out = 16'(-18355);
			553: out = 16'(-8791);
			554: out = 16'(2558);
			555: out = 16'(-7713);
			556: out = 16'(-12950);
			557: out = 16'(2596);
			558: out = 16'(3828);
			559: out = 16'(6203);
			560: out = 16'(19421);
			561: out = 16'(-1545);
			562: out = 16'(2853);
			563: out = 16'(-7625);
			564: out = 16'(-21376);
			565: out = 16'(-5846);
			566: out = 16'(3963);
			567: out = 16'(-11589);
			568: out = 16'(13797);
			569: out = 16'(-340);
			570: out = 16'(15505);
			571: out = 16'(331);
			572: out = 16'(-28590);
			573: out = 16'(4047);
			574: out = 16'(296);
			575: out = 16'(-1474);
			576: out = 16'(4771);
			577: out = 16'(-2067);
			578: out = 16'(1665);
			579: out = 16'(9779);
			580: out = 16'(6094);
			581: out = 16'(3337);
			582: out = 16'(7699);
			583: out = 16'(-9841);
			584: out = 16'(-5377);
			585: out = 16'(-1225);
			586: out = 16'(-20612);
			587: out = 16'(1557);
			588: out = 16'(10331);
			589: out = 16'(3249);
			590: out = 16'(21039);
			591: out = 16'(3134);
			592: out = 16'(10598);
			593: out = 16'(3785);
			594: out = 16'(13144);
			595: out = 16'(-5030);
			596: out = 16'(5287);
			597: out = 16'(-9452);
			598: out = 16'(5310);
			599: out = 16'(-12402);
			600: out = 16'(4857);
			601: out = 16'(2599);
			602: out = 16'(2747);
			603: out = 16'(6912);
			604: out = 16'(10752);
			605: out = 16'(11116);
			606: out = 16'(-1394);
			607: out = 16'(-3821);
			608: out = 16'(-23402);
			609: out = 16'(2449);
			610: out = 16'(12542);
			611: out = 16'(16004);
			612: out = 16'(-5467);
			613: out = 16'(-4988);
			614: out = 16'(3012);
			615: out = 16'(-13446);
			616: out = 16'(6143);
			617: out = 16'(-2203);
			618: out = 16'(975);
			619: out = 16'(2907);
			620: out = 16'(-13020);
			621: out = 16'(8863);
			622: out = 16'(3575);
			623: out = 16'(-29733);
			624: out = 16'(13823);
			625: out = 16'(5801);
			626: out = 16'(393);
			627: out = 16'(-10491);
			628: out = 16'(10892);
			629: out = 16'(-10333);
			630: out = 16'(-12795);
			631: out = 16'(-6513);
			632: out = 16'(4978);
			633: out = 16'(3642);
			634: out = 16'(-4348);
			635: out = 16'(-4492);
			636: out = 16'(7177);
			637: out = 16'(-1782);
			638: out = 16'(8023);
			639: out = 16'(13445);
			640: out = 16'(676);
			641: out = 16'(3011);
			642: out = 16'(6053);
			643: out = 16'(1878);
			644: out = 16'(6239);
			645: out = 16'(-13009);
			646: out = 16'(11609);
			647: out = 16'(11217);
			648: out = 16'(-2752);
			649: out = 16'(-4095);
			650: out = 16'(-268);
			651: out = 16'(7514);
			652: out = 16'(1807);
			653: out = 16'(5361);
			654: out = 16'(6681);
			655: out = 16'(12459);
			656: out = 16'(-238);
			657: out = 16'(-8114);
			658: out = 16'(10268);
			659: out = 16'(-2014);
			660: out = 16'(-9472);
			661: out = 16'(5084);
			662: out = 16'(7039);
			663: out = 16'(804);
			664: out = 16'(1693);
			665: out = 16'(-1416);
			666: out = 16'(7370);
			667: out = 16'(-648);
			668: out = 16'(8091);
			669: out = 16'(1536);
			670: out = 16'(-8978);
			671: out = 16'(-4657);
			672: out = 16'(-3887);
			673: out = 16'(-4634);
			674: out = 16'(-3539);
			675: out = 16'(-12207);
			676: out = 16'(-4176);
			677: out = 16'(2612);
			678: out = 16'(-10488);
			679: out = 16'(4795);
			680: out = 16'(-7617);
			681: out = 16'(186);
			682: out = 16'(-9047);
			683: out = 16'(16302);
			684: out = 16'(-10967);
			685: out = 16'(-3297);
			686: out = 16'(2873);
			687: out = 16'(205);
			688: out = 16'(-2102);
			689: out = 16'(-8083);
			690: out = 16'(-6052);
			691: out = 16'(-6480);
			692: out = 16'(-10897);
			693: out = 16'(-4095);
			694: out = 16'(-4168);
			695: out = 16'(11203);
			696: out = 16'(10349);
			697: out = 16'(-6117);
			698: out = 16'(-1555);
			699: out = 16'(-2201);
			700: out = 16'(-15289);
			701: out = 16'(-4757);
			702: out = 16'(-3080);
			703: out = 16'(-991);
			704: out = 16'(6034);
			705: out = 16'(-2611);
			706: out = 16'(-1819);
			707: out = 16'(1375);
			708: out = 16'(-5694);
			709: out = 16'(2702);
			710: out = 16'(8691);
			711: out = 16'(1485);
			712: out = 16'(-12063);
			713: out = 16'(-9082);
			714: out = 16'(2307);
			715: out = 16'(2660);
			716: out = 16'(8205);
			717: out = 16'(22088);
			718: out = 16'(-6762);
			719: out = 16'(2710);
			720: out = 16'(4490);
			721: out = 16'(-4086);
			722: out = 16'(-7428);
			723: out = 16'(-3362);
			724: out = 16'(-3316);
			725: out = 16'(11561);
			726: out = 16'(-4657);
			727: out = 16'(1695);
			728: out = 16'(-2255);
			729: out = 16'(-3905);
			730: out = 16'(1358);
			731: out = 16'(18396);
			732: out = 16'(11184);
			733: out = 16'(-1987);
			734: out = 16'(7915);
			735: out = 16'(859);
			736: out = 16'(9630);
			737: out = 16'(-8290);
			738: out = 16'(-9539);
			739: out = 16'(17399);
			740: out = 16'(5152);
			741: out = 16'(1401);
			742: out = 16'(-4513);
			743: out = 16'(294);
			744: out = 16'(-15417);
			745: out = 16'(9099);
			746: out = 16'(2022);
			747: out = 16'(12654);
			748: out = 16'(2520);
			749: out = 16'(-4783);
			750: out = 16'(9958);
			751: out = 16'(-137);
			752: out = 16'(5578);
			753: out = 16'(1045);
			754: out = 16'(11547);
			755: out = 16'(-2251);
			756: out = 16'(1474);
			757: out = 16'(-1439);
			758: out = 16'(5058);
			759: out = 16'(-718);
			760: out = 16'(2285);
			761: out = 16'(-439);
			762: out = 16'(-4282);
			763: out = 16'(-11483);
			764: out = 16'(-2468);
			765: out = 16'(12425);
			766: out = 16'(-8203);
			767: out = 16'(-3079);
			768: out = 16'(2584);
			769: out = 16'(16467);
			770: out = 16'(-2097);
			771: out = 16'(-5334);
			772: out = 16'(2836);
			773: out = 16'(9646);
			774: out = 16'(-1404);
			775: out = 16'(7228);
			776: out = 16'(6744);
			777: out = 16'(-12022);
			778: out = 16'(5428);
			779: out = 16'(-2858);
			780: out = 16'(9984);
			781: out = 16'(-5047);
			782: out = 16'(12607);
			783: out = 16'(1692);
			784: out = 16'(7686);
			785: out = 16'(-1375);
			786: out = 16'(4246);
			787: out = 16'(6541);
			788: out = 16'(-491);
			789: out = 16'(-1266);
			790: out = 16'(4755);
			791: out = 16'(-3605);
			792: out = 16'(1934);
			793: out = 16'(5336);
			794: out = 16'(-12380);
			795: out = 16'(5905);
			796: out = 16'(-9656);
			797: out = 16'(9686);
			798: out = 16'(2628);
			799: out = 16'(-6766);
			800: out = 16'(-9193);
			801: out = 16'(11599);
			802: out = 16'(-1938);
			803: out = 16'(10395);
			804: out = 16'(-12908);
			805: out = 16'(3255);
			806: out = 16'(-3017);
			807: out = 16'(-3284);
			808: out = 16'(-7519);
			809: out = 16'(5601);
			810: out = 16'(-703);
			811: out = 16'(3259);
			812: out = 16'(-4789);
			813: out = 16'(-10980);
			814: out = 16'(8719);
			815: out = 16'(-6025);
			816: out = 16'(50);
			817: out = 16'(-1422);
			818: out = 16'(2750);
			819: out = 16'(-8720);
			820: out = 16'(6126);
			821: out = 16'(-11075);
			822: out = 16'(-1067);
			823: out = 16'(-8261);
			824: out = 16'(4320);
			825: out = 16'(-6728);
			826: out = 16'(-7690);
			827: out = 16'(-5222);
			828: out = 16'(9536);
			829: out = 16'(-642);
			830: out = 16'(8699);
			831: out = 16'(-6253);
			832: out = 16'(741);
			833: out = 16'(3348);
			834: out = 16'(-7083);
			835: out = 16'(-2274);
			836: out = 16'(9950);
			837: out = 16'(4037);
			838: out = 16'(2816);
			839: out = 16'(-754);
			840: out = 16'(3131);
			841: out = 16'(-9565);
			842: out = 16'(7664);
			843: out = 16'(1684);
			844: out = 16'(9617);
			845: out = 16'(-2674);
			846: out = 16'(-6884);
			847: out = 16'(1358);
			848: out = 16'(-13763);
			849: out = 16'(1211);
			850: out = 16'(5225);
			851: out = 16'(11451);
			852: out = 16'(-3899);
			853: out = 16'(6201);
			854: out = 16'(-7774);
			855: out = 16'(-1894);
			856: out = 16'(-9685);
			857: out = 16'(3217);
			858: out = 16'(-6388);
			859: out = 16'(5825);
			860: out = 16'(-11690);
			861: out = 16'(9435);
			862: out = 16'(-6377);
			863: out = 16'(596);
			864: out = 16'(-1281);
			865: out = 16'(5104);
			866: out = 16'(-7364);
			867: out = 16'(2867);
			868: out = 16'(-1504);
			869: out = 16'(-4881);
			870: out = 16'(950);
			871: out = 16'(-2470);
			872: out = 16'(-5519);
			873: out = 16'(7819);
			874: out = 16'(6931);
			875: out = 16'(-2999);
			876: out = 16'(2929);
			877: out = 16'(-1319);
			878: out = 16'(-13315);
			879: out = 16'(5206);
			880: out = 16'(-503);
			881: out = 16'(423);
			882: out = 16'(603);
			883: out = 16'(-10272);
			884: out = 16'(-6841);
			885: out = 16'(-3485);
			886: out = 16'(1402);
			887: out = 16'(3741);
			888: out = 16'(983);
			889: out = 16'(-9765);
			890: out = 16'(7805);
			891: out = 16'(5751);
			892: out = 16'(-1958);
			893: out = 16'(-290);
			894: out = 16'(11159);
			895: out = 16'(-822);
			896: out = 16'(5421);
			897: out = 16'(1963);
			898: out = 16'(-3693);
			899: out = 16'(-946);
			900: out = 16'(-15250);
			901: out = 16'(736);
			902: out = 16'(7463);
			903: out = 16'(-5906);
			904: out = 16'(410);
			905: out = 16'(8546);
			906: out = 16'(-10802);
			907: out = 16'(3734);
			908: out = 16'(-322);
			909: out = 16'(4041);
			910: out = 16'(7871);
			911: out = 16'(-7785);
			912: out = 16'(-5045);
			913: out = 16'(4179);
			914: out = 16'(-4545);
			915: out = 16'(-3340);
			916: out = 16'(6197);
			917: out = 16'(49);
			918: out = 16'(4399);
			919: out = 16'(161);
			920: out = 16'(6576);
			921: out = 16'(-1374);
			922: out = 16'(225);
			923: out = 16'(-1038);
			924: out = 16'(14405);
			925: out = 16'(-310);
			926: out = 16'(-4137);
			927: out = 16'(2618);
			928: out = 16'(1465);
			929: out = 16'(1556);
			930: out = 16'(9217);
			931: out = 16'(10886);
			932: out = 16'(-8618);
			933: out = 16'(959);
			934: out = 16'(3266);
			935: out = 16'(2262);
			936: out = 16'(-4429);
			937: out = 16'(141);
			938: out = 16'(-7458);
			939: out = 16'(8506);
			940: out = 16'(-1073);
			941: out = 16'(-3692);
			942: out = 16'(-1766);
			943: out = 16'(6959);
			944: out = 16'(-658);
			945: out = 16'(6028);
			946: out = 16'(1280);
			947: out = 16'(-1831);
			948: out = 16'(4005);
			949: out = 16'(-7520);
			950: out = 16'(835);
			951: out = 16'(-188);
			952: out = 16'(-4742);
			953: out = 16'(-10535);
			954: out = 16'(7946);
			955: out = 16'(-6426);
			956: out = 16'(334);
			957: out = 16'(-57);
			958: out = 16'(1351);
			959: out = 16'(-10519);
			960: out = 16'(1806);
			961: out = 16'(-5481);
			962: out = 16'(289);
			963: out = 16'(-781);
			964: out = 16'(-2151);
			965: out = 16'(6291);
			966: out = 16'(-2127);
			967: out = 16'(-6345);
			968: out = 16'(1717);
			969: out = 16'(-3934);
			970: out = 16'(-3189);
			971: out = 16'(9267);
			972: out = 16'(1729);
			973: out = 16'(-8583);
			974: out = 16'(-5518);
			975: out = 16'(-9379);
			976: out = 16'(-165);
			977: out = 16'(13143);
			978: out = 16'(-12152);
			979: out = 16'(2208);
			980: out = 16'(3117);
			981: out = 16'(872);
			982: out = 16'(-802);
			983: out = 16'(3826);
			984: out = 16'(-10234);
			985: out = 16'(-199);
			986: out = 16'(-1009);
			987: out = 16'(1554);
			988: out = 16'(-3352);
			989: out = 16'(-5603);
			990: out = 16'(5817);
			991: out = 16'(7396);
			992: out = 16'(-3303);
			993: out = 16'(3007);
			994: out = 16'(-2402);
			995: out = 16'(3167);
			996: out = 16'(942);
			997: out = 16'(-12587);
			998: out = 16'(2715);
			999: out = 16'(3819);
			1000: out = 16'(1925);
			1001: out = 16'(2024);
			1002: out = 16'(2109);
			1003: out = 16'(-4825);
			1004: out = 16'(-2679);
			1005: out = 16'(-8596);
			1006: out = 16'(1800);
			1007: out = 16'(-8689);
			1008: out = 16'(2102);
			1009: out = 16'(-5858);
			1010: out = 16'(-1997);
			1011: out = 16'(-1685);
			1012: out = 16'(-5582);
			1013: out = 16'(4068);
			1014: out = 16'(3648);
			1015: out = 16'(6160);
			1016: out = 16'(4245);
			1017: out = 16'(149);
			1018: out = 16'(-1012);
			1019: out = 16'(1970);
			1020: out = 16'(-9782);
			1021: out = 16'(7051);
			1022: out = 16'(-7604);
			1023: out = 16'(8196);
			1024: out = 16'(-9434);
			1025: out = 16'(1762);
			1026: out = 16'(-19619);
			1027: out = 16'(2637);
			1028: out = 16'(-5111);
			1029: out = 16'(-1672);
			1030: out = 16'(5266);
			1031: out = 16'(-1985);
			1032: out = 16'(2148);
			1033: out = 16'(2639);
			1034: out = 16'(5962);
			1035: out = 16'(5027);
			1036: out = 16'(4879);
			1037: out = 16'(-5203);
			1038: out = 16'(5668);
			1039: out = 16'(-282);
			1040: out = 16'(-6097);
			1041: out = 16'(2988);
			1042: out = 16'(-8177);
			1043: out = 16'(-1069);
			1044: out = 16'(2387);
			1045: out = 16'(8679);
			1046: out = 16'(-5765);
			1047: out = 16'(6935);
			1048: out = 16'(7168);
			1049: out = 16'(8556);
			1050: out = 16'(2750);
			1051: out = 16'(6590);
			1052: out = 16'(4435);
			1053: out = 16'(10451);
			1054: out = 16'(-7469);
			1055: out = 16'(-6173);
			1056: out = 16'(14);
			1057: out = 16'(7923);
			1058: out = 16'(229);
			1059: out = 16'(-6782);
			1060: out = 16'(-3889);
			1061: out = 16'(-2373);
			1062: out = 16'(1136);
			1063: out = 16'(-2904);
			1064: out = 16'(708);
			1065: out = 16'(-374);
			1066: out = 16'(2982);
			1067: out = 16'(870);
			1068: out = 16'(2920);
			1069: out = 16'(-12074);
			1070: out = 16'(375);
			1071: out = 16'(3598);
			1072: out = 16'(2265);
			1073: out = 16'(3120);
			1074: out = 16'(5532);
			1075: out = 16'(827);
			1076: out = 16'(714);
			1077: out = 16'(-4575);
			1078: out = 16'(1648);
			1079: out = 16'(1580);
			1080: out = 16'(2632);
			1081: out = 16'(3050);
			1082: out = 16'(-2304);
			1083: out = 16'(-9335);
			1084: out = 16'(6971);
			1085: out = 16'(-973);
			1086: out = 16'(-5871);
			1087: out = 16'(2226);
			1088: out = 16'(2113);
			1089: out = 16'(-1387);
			1090: out = 16'(3226);
			1091: out = 16'(-157);
			1092: out = 16'(-7544);
			1093: out = 16'(6148);
			1094: out = 16'(420);
			1095: out = 16'(768);
			1096: out = 16'(-73);
			1097: out = 16'(-5060);
			1098: out = 16'(1922);
			1099: out = 16'(8912);
			1100: out = 16'(-9030);
			1101: out = 16'(9380);
			1102: out = 16'(1345);
			1103: out = 16'(1054);
			1104: out = 16'(-6272);
			1105: out = 16'(5648);
			1106: out = 16'(-3925);
			1107: out = 16'(2230);
			1108: out = 16'(739);
			1109: out = 16'(466);
			1110: out = 16'(-3474);
			1111: out = 16'(-7879);
			1112: out = 16'(2819);
			1113: out = 16'(-2455);
			1114: out = 16'(3217);
			1115: out = 16'(-407);
			1116: out = 16'(12164);
			1117: out = 16'(-3430);
			1118: out = 16'(-415);
			1119: out = 16'(1550);
			1120: out = 16'(-1924);
			1121: out = 16'(-597);
			1122: out = 16'(2623);
			1123: out = 16'(-12655);
			1124: out = 16'(4785);
			1125: out = 16'(282);
			1126: out = 16'(-422);
			1127: out = 16'(-1097);
			1128: out = 16'(-1817);
			1129: out = 16'(-751);
			1130: out = 16'(-789);
			1131: out = 16'(2425);
			1132: out = 16'(-12007);
			1133: out = 16'(3736);
			1134: out = 16'(2273);
			1135: out = 16'(2475);
			1136: out = 16'(-651);
			1137: out = 16'(-3932);
			1138: out = 16'(51);
			1139: out = 16'(2951);
			1140: out = 16'(86);
			1141: out = 16'(-1594);
			1142: out = 16'(11632);
			1143: out = 16'(-7671);
			1144: out = 16'(287);
			1145: out = 16'(-2138);
			1146: out = 16'(-6675);
			1147: out = 16'(-1197);
			1148: out = 16'(5365);
			1149: out = 16'(-3563);
			1150: out = 16'(5845);
			1151: out = 16'(-7258);
			1152: out = 16'(-4182);
			1153: out = 16'(387);
			1154: out = 16'(182);
			1155: out = 16'(-6636);
			1156: out = 16'(2078);
			1157: out = 16'(-1967);
			1158: out = 16'(877);
			1159: out = 16'(-553);
			1160: out = 16'(-3179);
			1161: out = 16'(-2736);
			1162: out = 16'(-3649);
			1163: out = 16'(1125);
			1164: out = 16'(21);
			1165: out = 16'(4236);
			1166: out = 16'(944);
			1167: out = 16'(9067);
			1168: out = 16'(-4645);
			1169: out = 16'(-3122);
			1170: out = 16'(1237);
			1171: out = 16'(-1282);
			1172: out = 16'(1001);
			1173: out = 16'(-1367);
			1174: out = 16'(-777);
			1175: out = 16'(1724);
			1176: out = 16'(250);
			1177: out = 16'(-3434);
			1178: out = 16'(-450);
			1179: out = 16'(-575);
			1180: out = 16'(-1497);
			1181: out = 16'(-345);
			1182: out = 16'(-3241);
			1183: out = 16'(-6694);
			1184: out = 16'(170);
			1185: out = 16'(9768);
			1186: out = 16'(8917);
			1187: out = 16'(-10645);
			1188: out = 16'(63);
			1189: out = 16'(1815);
			1190: out = 16'(4814);
			1191: out = 16'(2432);
			1192: out = 16'(-3514);
			1193: out = 16'(-1330);
			1194: out = 16'(10576);
			1195: out = 16'(4178);
			1196: out = 16'(-3429);
			1197: out = 16'(2947);
			1198: out = 16'(2911);
			1199: out = 16'(606);
			1200: out = 16'(10583);
			1201: out = 16'(-9852);
			1202: out = 16'(-4577);
			1203: out = 16'(2127);
			1204: out = 16'(1745);
			1205: out = 16'(-1596);
			1206: out = 16'(-3346);
			1207: out = 16'(2705);
			1208: out = 16'(-1900);
			1209: out = 16'(-117);
			1210: out = 16'(-877);
			1211: out = 16'(3183);
			1212: out = 16'(-4279);
			1213: out = 16'(4981);
			1214: out = 16'(-6170);
			1215: out = 16'(602);
			1216: out = 16'(3182);
			1217: out = 16'(32);
			1218: out = 16'(-550);
			1219: out = 16'(4671);
			1220: out = 16'(-7901);
			1221: out = 16'(-385);
			1222: out = 16'(10504);
			1223: out = 16'(71);
			1224: out = 16'(-8703);
			1225: out = 16'(138);
			1226: out = 16'(-7447);
			1227: out = 16'(5515);
			1228: out = 16'(6394);
			1229: out = 16'(-9105);
			1230: out = 16'(5317);
			1231: out = 16'(606);
			1232: out = 16'(-2996);
			1233: out = 16'(-375);
			1234: out = 16'(-228);
			1235: out = 16'(945);
			1236: out = 16'(1368);
			1237: out = 16'(-384);
			1238: out = 16'(3669);
			1239: out = 16'(2505);
			1240: out = 16'(-3297);
			1241: out = 16'(4067);
			1242: out = 16'(729);
			1243: out = 16'(2791);
			1244: out = 16'(3668);
			1245: out = 16'(8173);
			1246: out = 16'(-2030);
			1247: out = 16'(-1077);
			1248: out = 16'(-1149);
			1249: out = 16'(2051);
			1250: out = 16'(3070);
			1251: out = 16'(-426);
			1252: out = 16'(-1484);
			1253: out = 16'(-402);
			1254: out = 16'(-1525);
			1255: out = 16'(-8600);
			1256: out = 16'(6125);
			1257: out = 16'(285);
			1258: out = 16'(5826);
			1259: out = 16'(5596);
			1260: out = 16'(3534);
			1261: out = 16'(1467);
			1262: out = 16'(774);
			1263: out = 16'(-1134);
			1264: out = 16'(3233);
			1265: out = 16'(-6622);
			1266: out = 16'(-485);
			1267: out = 16'(-7195);
			1268: out = 16'(-1371);
			1269: out = 16'(-7565);
			1270: out = 16'(53);
			1271: out = 16'(-714);
			1272: out = 16'(-891);
			1273: out = 16'(-383);
			1274: out = 16'(-4561);
			1275: out = 16'(-6976);
			1276: out = 16'(-204);
			1277: out = 16'(-1428);
			1278: out = 16'(-1923);
			1279: out = 16'(781);
			1280: out = 16'(-4549);
			1281: out = 16'(-3259);
			1282: out = 16'(314);
			1283: out = 16'(1116);
			1284: out = 16'(1527);
			1285: out = 16'(1965);
			1286: out = 16'(560);
			1287: out = 16'(-4869);
			1288: out = 16'(544);
			1289: out = 16'(6864);
			1290: out = 16'(3409);
			1291: out = 16'(629);
			1292: out = 16'(1284);
			1293: out = 16'(-4003);
			1294: out = 16'(-6793);
			1295: out = 16'(-1644);
			1296: out = 16'(3308);
			1297: out = 16'(-9384);
			1298: out = 16'(-445);
			1299: out = 16'(-5568);
			1300: out = 16'(1608);
			1301: out = 16'(6737);
			1302: out = 16'(1218);
			1303: out = 16'(-9162);
			1304: out = 16'(2893);
			1305: out = 16'(998);
			1306: out = 16'(4188);
			1307: out = 16'(3881);
			1308: out = 16'(582);
			1309: out = 16'(4591);
			1310: out = 16'(-2679);
			1311: out = 16'(1215);
			1312: out = 16'(4724);
			1313: out = 16'(1152);
			1314: out = 16'(-2214);
			1315: out = 16'(-5724);
			1316: out = 16'(3351);
			1317: out = 16'(-1490);
			1318: out = 16'(43);
			1319: out = 16'(-5353);
			1320: out = 16'(-3622);
			1321: out = 16'(-5456);
			1322: out = 16'(1661);
			1323: out = 16'(101);
			1324: out = 16'(5395);
			1325: out = 16'(7945);
			1326: out = 16'(10455);
			1327: out = 16'(788);
			1328: out = 16'(-613);
			1329: out = 16'(-653);
			1330: out = 16'(-3595);
			1331: out = 16'(-5336);
			1332: out = 16'(4774);
			1333: out = 16'(-6965);
			1334: out = 16'(-8245);
			1335: out = 16'(2174);
			1336: out = 16'(-619);
			1337: out = 16'(-529);
			1338: out = 16'(2111);
			1339: out = 16'(3203);
			1340: out = 16'(1115);
			1341: out = 16'(7781);
			1342: out = 16'(-1810);
			1343: out = 16'(-1356);
			1344: out = 16'(3277);
			1345: out = 16'(-4665);
			1346: out = 16'(-4155);
			1347: out = 16'(-8383);
			1348: out = 16'(6474);
			1349: out = 16'(3717);
			1350: out = 16'(-267);
			1351: out = 16'(6260);
			1352: out = 16'(-11651);
			1353: out = 16'(1472);
			1354: out = 16'(3782);
			1355: out = 16'(1355);
			1356: out = 16'(-5393);
			1357: out = 16'(1600);
			1358: out = 16'(-2459);
			1359: out = 16'(7847);
			1360: out = 16'(80);
			1361: out = 16'(5802);
			1362: out = 16'(2446);
			1363: out = 16'(5994);
			1364: out = 16'(4839);
			1365: out = 16'(-2299);
			1366: out = 16'(36);
			1367: out = 16'(-134);
			1368: out = 16'(1242);
			1369: out = 16'(-3023);
			1370: out = 16'(5363);
			1371: out = 16'(-275);
			1372: out = 16'(-346);
			1373: out = 16'(-1561);
			1374: out = 16'(-7645);
			1375: out = 16'(-887);
			1376: out = 16'(-1959);
			1377: out = 16'(-218);
			1378: out = 16'(8240);
			1379: out = 16'(3374);
			1380: out = 16'(-6133);
			1381: out = 16'(4474);
			1382: out = 16'(-592);
			1383: out = 16'(-10874);
			1384: out = 16'(-431);
			1385: out = 16'(55);
			1386: out = 16'(-4187);
			1387: out = 16'(-923);
			1388: out = 16'(1994);
			1389: out = 16'(-3272);
			1390: out = 16'(6680);
			1391: out = 16'(1955);
			1392: out = 16'(10626);
			1393: out = 16'(-4501);
			1394: out = 16'(3485);
			1395: out = 16'(-6064);
			1396: out = 16'(-4694);
			1397: out = 16'(839);
			1398: out = 16'(-13773);
			1399: out = 16'(5002);
			1400: out = 16'(9523);
			1401: out = 16'(764);
			1402: out = 16'(1008);
			1403: out = 16'(2174);
			1404: out = 16'(6830);
			1405: out = 16'(3957);
			1406: out = 16'(-7585);
			1407: out = 16'(11698);
			1408: out = 16'(-4239);
			1409: out = 16'(-7258);
			1410: out = 16'(8881);
			1411: out = 16'(-173);
			1412: out = 16'(-4593);
			1413: out = 16'(3802);
			1414: out = 16'(6264);
			1415: out = 16'(-390);
			1416: out = 16'(6745);
			1417: out = 16'(-4704);
			1418: out = 16'(3948);
			1419: out = 16'(1551);
			1420: out = 16'(-11338);
			1421: out = 16'(449);
			1422: out = 16'(816);
			1423: out = 16'(-2073);
			1424: out = 16'(3369);
			1425: out = 16'(-2183);
			1426: out = 16'(-866);
			1427: out = 16'(9345);
			1428: out = 16'(-6579);
			1429: out = 16'(-193);
			1430: out = 16'(2000);
			1431: out = 16'(228);
			1432: out = 16'(-1197);
			1433: out = 16'(9203);
			1434: out = 16'(-7623);
			1435: out = 16'(1237);
			1436: out = 16'(1497);
			1437: out = 16'(-1750);
			1438: out = 16'(-1699);
			1439: out = 16'(-299);
			1440: out = 16'(656);
			1441: out = 16'(998);
			1442: out = 16'(-231);
			1443: out = 16'(-624);
			1444: out = 16'(-2071);
			1445: out = 16'(4283);
			1446: out = 16'(4539);
			1447: out = 16'(-427);
			1448: out = 16'(-1212);
			1449: out = 16'(-7799);
			1450: out = 16'(4754);
			1451: out = 16'(5027);
			1452: out = 16'(3737);
			1453: out = 16'(-5691);
			1454: out = 16'(7284);
			1455: out = 16'(-1877);
			1456: out = 16'(-681);
			1457: out = 16'(-6763);
			1458: out = 16'(-9663);
			1459: out = 16'(-4061);
			1460: out = 16'(5769);
			1461: out = 16'(-2151);
			1462: out = 16'(686);
			1463: out = 16'(-1681);
			1464: out = 16'(1461);
			1465: out = 16'(1145);
			1466: out = 16'(-5306);
			1467: out = 16'(8705);
			1468: out = 16'(-681);
			1469: out = 16'(-2718);
			1470: out = 16'(2082);
			1471: out = 16'(-9945);
			1472: out = 16'(-144);
			1473: out = 16'(5384);
			1474: out = 16'(-4735);
			1475: out = 16'(3838);
			1476: out = 16'(-743);
			1477: out = 16'(2026);
			1478: out = 16'(832);
			1479: out = 16'(-5135);
			1480: out = 16'(5532);
			1481: out = 16'(1701);
			1482: out = 16'(-7315);
			1483: out = 16'(-917);
			1484: out = 16'(-1836);
			1485: out = 16'(-6793);
			1486: out = 16'(3280);
			1487: out = 16'(5509);
			1488: out = 16'(-5588);
			1489: out = 16'(-2062);
			1490: out = 16'(-2018);
			1491: out = 16'(2309);
			1492: out = 16'(2840);
			1493: out = 16'(-10733);
			1494: out = 16'(251);
			1495: out = 16'(4512);
			1496: out = 16'(1630);
			1497: out = 16'(2936);
			1498: out = 16'(-251);
			1499: out = 16'(3499);
			1500: out = 16'(6806);
			1501: out = 16'(241);
			1502: out = 16'(-4673);
			1503: out = 16'(8132);
			1504: out = 16'(-4411);
			1505: out = 16'(-666);
			1506: out = 16'(5709);
			1507: out = 16'(-2345);
			1508: out = 16'(3551);
			1509: out = 16'(3209);
			1510: out = 16'(-70);
			1511: out = 16'(-2834);
			1512: out = 16'(-3152);
			1513: out = 16'(-3822);
			1514: out = 16'(2737);
			1515: out = 16'(-7309);
			1516: out = 16'(1399);
			1517: out = 16'(519);
			1518: out = 16'(4167);
			1519: out = 16'(4540);
			1520: out = 16'(-2990);
			1521: out = 16'(-3156);
			1522: out = 16'(-2842);
			1523: out = 16'(-6928);
			1524: out = 16'(144);
			1525: out = 16'(-5349);
			1526: out = 16'(-1649);
			1527: out = 16'(-2647);
			1528: out = 16'(1518);
			1529: out = 16'(-2410);
			1530: out = 16'(7682);
			1531: out = 16'(-8241);
			1532: out = 16'(3064);
			1533: out = 16'(-358);
			1534: out = 16'(-6981);
			1535: out = 16'(2953);
			1536: out = 16'(4215);
			1537: out = 16'(-1896);
			1538: out = 16'(-10098);
			1539: out = 16'(-1082);
			1540: out = 16'(-2750);
			1541: out = 16'(2660);
			1542: out = 16'(1137);
			1543: out = 16'(2842);
			1544: out = 16'(2781);
			1545: out = 16'(1176);
			1546: out = 16'(731);
			1547: out = 16'(2654);
			1548: out = 16'(-889);
			1549: out = 16'(5811);
			1550: out = 16'(666);
			1551: out = 16'(-2678);
			1552: out = 16'(-2117);
			1553: out = 16'(-66);
			1554: out = 16'(1500);
			1555: out = 16'(3079);
			1556: out = 16'(-592);
			1557: out = 16'(-1756);
			1558: out = 16'(2352);
			1559: out = 16'(-288);
			1560: out = 16'(8566);
			1561: out = 16'(5428);
			1562: out = 16'(-8339);
			1563: out = 16'(4568);
			1564: out = 16'(-3156);
			1565: out = 16'(326);
			1566: out = 16'(-5338);
			1567: out = 16'(932);
			1568: out = 16'(-7316);
			1569: out = 16'(234);
			1570: out = 16'(1419);
			1571: out = 16'(-2120);
			1572: out = 16'(6318);
			1573: out = 16'(-7133);
			1574: out = 16'(445);
			1575: out = 16'(2841);
			1576: out = 16'(1784);
			1577: out = 16'(5642);
			1578: out = 16'(-1516);
			1579: out = 16'(801);
			1580: out = 16'(9404);
			1581: out = 16'(287);
			1582: out = 16'(-6453);
			1583: out = 16'(1422);
			1584: out = 16'(-2212);
			1585: out = 16'(2391);
			1586: out = 16'(-4776);
			1587: out = 16'(-346);
			1588: out = 16'(-10936);
			1589: out = 16'(-556);
			1590: out = 16'(-662);
			1591: out = 16'(-1901);
			1592: out = 16'(3982);
			1593: out = 16'(-2965);
			1594: out = 16'(7431);
			1595: out = 16'(-5053);
			1596: out = 16'(5006);
			1597: out = 16'(-2267);
			1598: out = 16'(3350);
			1599: out = 16'(-1005);
			1600: out = 16'(2626);
			1601: out = 16'(-669);
			1602: out = 16'(3069);
			1603: out = 16'(4866);
			1604: out = 16'(-169);
			1605: out = 16'(349);
			1606: out = 16'(196);
			1607: out = 16'(5559);
			1608: out = 16'(-3953);
			1609: out = 16'(-64);
			1610: out = 16'(5029);
			1611: out = 16'(-7188);
			1612: out = 16'(-1789);
			1613: out = 16'(5749);
			1614: out = 16'(-1869);
			1615: out = 16'(1388);
			1616: out = 16'(-863);
			1617: out = 16'(-7933);
			1618: out = 16'(-2750);
			1619: out = 16'(3823);
			1620: out = 16'(-7809);
			1621: out = 16'(-5539);
			1622: out = 16'(-4715);
			1623: out = 16'(6935);
			1624: out = 16'(1235);
			1625: out = 16'(1411);
			1626: out = 16'(1211);
			1627: out = 16'(7682);
			1628: out = 16'(1316);
			1629: out = 16'(6137);
			1630: out = 16'(-2669);
			1631: out = 16'(803);
			1632: out = 16'(-789);
			1633: out = 16'(-636);
			1634: out = 16'(-3324);
			1635: out = 16'(-4009);
			1636: out = 16'(-4144);
			1637: out = 16'(-984);
			1638: out = 16'(790);
			1639: out = 16'(148);
			1640: out = 16'(2561);
			1641: out = 16'(-6756);
			1642: out = 16'(-85);
			1643: out = 16'(-9494);
			1644: out = 16'(-4017);
			1645: out = 16'(5076);
			1646: out = 16'(-935);
			1647: out = 16'(262);
			1648: out = 16'(4773);
			1649: out = 16'(1799);
			1650: out = 16'(658);
			1651: out = 16'(4102);
			1652: out = 16'(-5201);
			1653: out = 16'(814);
			1654: out = 16'(3954);
			1655: out = 16'(1573);
			1656: out = 16'(1682);
			1657: out = 16'(860);
			1658: out = 16'(-4235);
			1659: out = 16'(-2573);
			1660: out = 16'(-1638);
			1661: out = 16'(-89);
			1662: out = 16'(3799);
			1663: out = 16'(7286);
			1664: out = 16'(639);
			1665: out = 16'(644);
			1666: out = 16'(-8204);
			1667: out = 16'(2458);
			1668: out = 16'(-7220);
			1669: out = 16'(-308);
			1670: out = 16'(1581);
			1671: out = 16'(-2963);
			1672: out = 16'(-9);
			1673: out = 16'(-6514);
			1674: out = 16'(927);
			1675: out = 16'(882);
			1676: out = 16'(7383);
			1677: out = 16'(-1569);
			1678: out = 16'(5747);
			1679: out = 16'(-1947);
			1680: out = 16'(8319);
			1681: out = 16'(-1395);
			1682: out = 16'(4626);
			1683: out = 16'(-399);
			1684: out = 16'(1658);
			1685: out = 16'(-7779);
			1686: out = 16'(-5609);
			1687: out = 16'(-3508);
			1688: out = 16'(-6709);
			1689: out = 16'(1458);
			1690: out = 16'(5158);
			1691: out = 16'(1074);
			1692: out = 16'(824);
			1693: out = 16'(3774);
			1694: out = 16'(-2009);
			1695: out = 16'(6821);
			1696: out = 16'(-426);
			1697: out = 16'(-112);
			1698: out = 16'(-6580);
			1699: out = 16'(-123);
			1700: out = 16'(1882);
			1701: out = 16'(1520);
			1702: out = 16'(-3114);
			1703: out = 16'(-1822);
			1704: out = 16'(3958);
			1705: out = 16'(1395);
			1706: out = 16'(-5277);
			1707: out = 16'(5931);
			1708: out = 16'(3327);
			1709: out = 16'(-2340);
			1710: out = 16'(-3646);
			1711: out = 16'(98);
			1712: out = 16'(-297);
			1713: out = 16'(7442);
			1714: out = 16'(2980);
			1715: out = 16'(-492);
			1716: out = 16'(-3180);
			1717: out = 16'(-1451);
			1718: out = 16'(3608);
			1719: out = 16'(-197);
			1720: out = 16'(3859);
			1721: out = 16'(-51);
			1722: out = 16'(923);
			1723: out = 16'(2444);
			1724: out = 16'(2204);
			1725: out = 16'(-498);
			1726: out = 16'(6253);
			1727: out = 16'(738);
			1728: out = 16'(622);
			1729: out = 16'(4647);
			1730: out = 16'(3644);
			1731: out = 16'(-938);
			1732: out = 16'(5627);
			1733: out = 16'(-456);
			1734: out = 16'(-1022);
			1735: out = 16'(-6015);
			1736: out = 16'(-10734);
			1737: out = 16'(476);
			1738: out = 16'(319);
			1739: out = 16'(-3438);
			1740: out = 16'(1574);
			1741: out = 16'(983);
			1742: out = 16'(-2868);
			1743: out = 16'(5097);
			1744: out = 16'(-7761);
			1745: out = 16'(-3870);
			1746: out = 16'(4455);
			1747: out = 16'(-1144);
			1748: out = 16'(3399);
			1749: out = 16'(2930);
			1750: out = 16'(-8021);
			1751: out = 16'(-4072);
			1752: out = 16'(1938);
			1753: out = 16'(-5993);
			1754: out = 16'(7214);
			1755: out = 16'(3056);
			1756: out = 16'(4750);
			1757: out = 16'(6727);
			1758: out = 16'(-3020);
			1759: out = 16'(-4978);
			1760: out = 16'(498);
			1761: out = 16'(-11402);
			1762: out = 16'(2938);
			1763: out = 16'(758);
			1764: out = 16'(-1757);
			1765: out = 16'(3261);
			1766: out = 16'(370);
			1767: out = 16'(-1671);
			1768: out = 16'(-1733);
			1769: out = 16'(2464);
			1770: out = 16'(-609);
			1771: out = 16'(3006);
			1772: out = 16'(-1653);
			1773: out = 16'(4740);
			1774: out = 16'(-4579);
			1775: out = 16'(-63);
			1776: out = 16'(-2199);
			1777: out = 16'(2433);
			1778: out = 16'(-1436);
			1779: out = 16'(6809);
			1780: out = 16'(441);
			1781: out = 16'(513);
			1782: out = 16'(5495);
			1783: out = 16'(-4144);
			1784: out = 16'(-1835);
			1785: out = 16'(4697);
			1786: out = 16'(-7707);
			1787: out = 16'(4456);
			1788: out = 16'(-6673);
			1789: out = 16'(3401);
			1790: out = 16'(-1912);
			1791: out = 16'(-814);
			1792: out = 16'(-2706);
			1793: out = 16'(-3063);
			1794: out = 16'(-91);
			1795: out = 16'(-5815);
			1796: out = 16'(1086);
			1797: out = 16'(2146);
			1798: out = 16'(1078);
			1799: out = 16'(2918);
			1800: out = 16'(-4536);
			1801: out = 16'(141);
			1802: out = 16'(7114);
			1803: out = 16'(1617);
			1804: out = 16'(-3099);
			1805: out = 16'(1676);
			1806: out = 16'(-2584);
			1807: out = 16'(5320);
			1808: out = 16'(-2667);
			1809: out = 16'(54);
			1810: out = 16'(-4713);
			1811: out = 16'(-40);
			1812: out = 16'(-2912);
			1813: out = 16'(831);
			1814: out = 16'(1677);
			1815: out = 16'(348);
			1816: out = 16'(671);
			1817: out = 16'(-668);
			1818: out = 16'(-5167);
			1819: out = 16'(-7443);
			1820: out = 16'(2014);
			1821: out = 16'(-1910);
			1822: out = 16'(7572);
			1823: out = 16'(-5449);
			1824: out = 16'(2073);
			1825: out = 16'(-852);
			1826: out = 16'(4723);
			1827: out = 16'(-5105);
			1828: out = 16'(-3708);
			1829: out = 16'(712);
			1830: out = 16'(-5295);
			1831: out = 16'(945);
			1832: out = 16'(-45);
			1833: out = 16'(-1437);
			1834: out = 16'(-795);
			1835: out = 16'(-1867);
			1836: out = 16'(-4674);
			1837: out = 16'(4416);
			1838: out = 16'(2882);
			1839: out = 16'(2078);
			1840: out = 16'(8175);
			1841: out = 16'(-329);
			1842: out = 16'(3084);
			1843: out = 16'(-7972);
			1844: out = 16'(-1636);
			1845: out = 16'(-4786);
			1846: out = 16'(-4248);
			1847: out = 16'(755);
			1848: out = 16'(361);
			1849: out = 16'(-1064);
			1850: out = 16'(-702);
			1851: out = 16'(-141);
			1852: out = 16'(-1783);
			1853: out = 16'(4879);
			1854: out = 16'(-2164);
			1855: out = 16'(4225);
			1856: out = 16'(-3287);
			1857: out = 16'(-1100);
			1858: out = 16'(3468);
			1859: out = 16'(-777);
			1860: out = 16'(41);
			1861: out = 16'(1970);
			1862: out = 16'(-1989);
			1863: out = 16'(-3539);
			1864: out = 16'(-1533);
			1865: out = 16'(-581);
			1866: out = 16'(2216);
			1867: out = 16'(2889);
			1868: out = 16'(1915);
			1869: out = 16'(4458);
			1870: out = 16'(2404);
			1871: out = 16'(-1210);
			1872: out = 16'(4576);
			1873: out = 16'(242);
			1874: out = 16'(-393);
			1875: out = 16'(7927);
			1876: out = 16'(-5378);
			1877: out = 16'(-3156);
			1878: out = 16'(2831);
			1879: out = 16'(-3494);
			1880: out = 16'(-180);
			1881: out = 16'(2353);
			1882: out = 16'(208);
			1883: out = 16'(3235);
			1884: out = 16'(1240);
			1885: out = 16'(59);
			1886: out = 16'(5147);
			1887: out = 16'(-8936);
			1888: out = 16'(1438);
			1889: out = 16'(-2118);
			1890: out = 16'(1472);
			1891: out = 16'(941);
			1892: out = 16'(3486);
			1893: out = 16'(-3002);
			1894: out = 16'(-2753);
			1895: out = 16'(600);
			1896: out = 16'(1013);
			1897: out = 16'(4631);
			1898: out = 16'(-1256);
			1899: out = 16'(1611);
			1900: out = 16'(-4355);
			1901: out = 16'(1691);
			1902: out = 16'(3179);
			1903: out = 16'(2238);
			1904: out = 16'(838);
			1905: out = 16'(409);
			1906: out = 16'(279);
			1907: out = 16'(-182);
			1908: out = 16'(2594);
			1909: out = 16'(-2568);
			1910: out = 16'(2081);
			1911: out = 16'(-2578);
			1912: out = 16'(-2264);
			1913: out = 16'(342);
			1914: out = 16'(2609);
			1915: out = 16'(-3996);
			1916: out = 16'(1256);
			1917: out = 16'(917);
			1918: out = 16'(1423);
			1919: out = 16'(7246);
			1920: out = 16'(-1721);
			1921: out = 16'(3134);
			1922: out = 16'(3896);
			1923: out = 16'(-3052);
			1924: out = 16'(-2750);
			1925: out = 16'(4019);
			1926: out = 16'(546);
			1927: out = 16'(9);
			1928: out = 16'(4797);
			1929: out = 16'(-5986);
			1930: out = 16'(4957);
			1931: out = 16'(2776);
			1932: out = 16'(-1762);
			1933: out = 16'(628);
			1934: out = 16'(-226);
			1935: out = 16'(-2845);
			1936: out = 16'(-618);
			1937: out = 16'(360);
			1938: out = 16'(-791);
			1939: out = 16'(5138);
			1940: out = 16'(-3675);
			1941: out = 16'(6093);
			1942: out = 16'(-142);
			1943: out = 16'(1672);
			1944: out = 16'(1074);
			1945: out = 16'(1861);
			1946: out = 16'(-3108);
			1947: out = 16'(-7306);
			1948: out = 16'(-183);
			1949: out = 16'(-2173);
			1950: out = 16'(5349);
			1951: out = 16'(-5078);
			1952: out = 16'(4062);
			1953: out = 16'(-6659);
			1954: out = 16'(2277);
			1955: out = 16'(-4091);
			1956: out = 16'(2136);
			1957: out = 16'(525);
			1958: out = 16'(3644);
			1959: out = 16'(2384);
			1960: out = 16'(-6126);
			1961: out = 16'(1642);
			1962: out = 16'(-8338);
			1963: out = 16'(216);
			1964: out = 16'(-5723);
			1965: out = 16'(1710);
			1966: out = 16'(-1271);
			1967: out = 16'(4433);
			1968: out = 16'(1299);
			1969: out = 16'(2194);
			1970: out = 16'(98);
			1971: out = 16'(1925);
			1972: out = 16'(-602);
			1973: out = 16'(-774);
			1974: out = 16'(3070);
			1975: out = 16'(-699);
			1976: out = 16'(-2250);
			1977: out = 16'(-3541);
			1978: out = 16'(-86);
			1979: out = 16'(1432);
			1980: out = 16'(-189);
			1981: out = 16'(2515);
			1982: out = 16'(-1206);
			1983: out = 16'(-1190);
			1984: out = 16'(2160);
			1985: out = 16'(936);
			1986: out = 16'(-1404);
			1987: out = 16'(3059);
			1988: out = 16'(-1255);
			1989: out = 16'(-2501);
			1990: out = 16'(-5394);
			1991: out = 16'(2057);
			1992: out = 16'(-1663);
			1993: out = 16'(1242);
			1994: out = 16'(2505);
			1995: out = 16'(-408);
			1996: out = 16'(-165);
			1997: out = 16'(-2660);
			1998: out = 16'(836);
			1999: out = 16'(2933);
			2000: out = 16'(997);
			2001: out = 16'(2549);
			2002: out = 16'(-482);
			2003: out = 16'(-429);
			2004: out = 16'(-292);
			2005: out = 16'(-1272);
			2006: out = 16'(-7122);
			2007: out = 16'(8398);
			2008: out = 16'(1661);
			2009: out = 16'(226);
			2010: out = 16'(1135);
			2011: out = 16'(-592);
			2012: out = 16'(2525);
			2013: out = 16'(-3800);
			2014: out = 16'(4233);
			2015: out = 16'(-900);
			2016: out = 16'(530);
			2017: out = 16'(-4207);
			2018: out = 16'(843);
			2019: out = 16'(-5055);
			2020: out = 16'(59);
			2021: out = 16'(225);
			2022: out = 16'(139);
			2023: out = 16'(-1373);
			2024: out = 16'(-450);
			2025: out = 16'(3381);
			2026: out = 16'(-8989);
			2027: out = 16'(-742);
			2028: out = 16'(-4819);
			2029: out = 16'(4461);
			2030: out = 16'(-1478);
			2031: out = 16'(3273);
			2032: out = 16'(556);
			2033: out = 16'(-2565);
			2034: out = 16'(1631);
			2035: out = 16'(-905);
			2036: out = 16'(7587);
			2037: out = 16'(1264);
			2038: out = 16'(4450);
			2039: out = 16'(-2526);
			2040: out = 16'(3203);
			2041: out = 16'(2109);
			2042: out = 16'(944);
			2043: out = 16'(-391);
			2044: out = 16'(306);
			2045: out = 16'(-779);
			2046: out = 16'(3656);
			2047: out = 16'(299);
			2048: out = 16'(-1129);
			2049: out = 16'(794);
			2050: out = 16'(-8157);
			2051: out = 16'(4819);
			2052: out = 16'(-789);
			2053: out = 16'(-909);
			2054: out = 16'(-898);
			2055: out = 16'(-2527);
			2056: out = 16'(-3259);
			2057: out = 16'(-640);
			2058: out = 16'(899);
			2059: out = 16'(1750);
			2060: out = 16'(2097);
			2061: out = 16'(23);
			2062: out = 16'(1916);
			2063: out = 16'(-1687);
			2064: out = 16'(5267);
			2065: out = 16'(-1083);
			2066: out = 16'(641);
			2067: out = 16'(-2978);
			2068: out = 16'(-4457);
			2069: out = 16'(2714);
			2070: out = 16'(4795);
			2071: out = 16'(-4531);
			2072: out = 16'(191);
			2073: out = 16'(3069);
			2074: out = 16'(-3496);
			2075: out = 16'(-3890);
			2076: out = 16'(-270);
			2077: out = 16'(-2611);
			2078: out = 16'(-4397);
			2079: out = 16'(-1221);
			2080: out = 16'(-4538);
			2081: out = 16'(2787);
			2082: out = 16'(516);
			2083: out = 16'(1098);
			2084: out = 16'(5798);
			2085: out = 16'(-2369);
			2086: out = 16'(5419);
			2087: out = 16'(5427);
			2088: out = 16'(1381);
			2089: out = 16'(4656);
			2090: out = 16'(1985);
			2091: out = 16'(-1891);
			2092: out = 16'(-971);
			2093: out = 16'(-370);
			2094: out = 16'(-4336);
			2095: out = 16'(-2263);
			2096: out = 16'(152);
			2097: out = 16'(-1037);
			2098: out = 16'(496);
			2099: out = 16'(-1768);
			2100: out = 16'(-1223);
			2101: out = 16'(1259);
			2102: out = 16'(-7719);
			2103: out = 16'(278);
			2104: out = 16'(-821);
			2105: out = 16'(-824);
			2106: out = 16'(1038);
			2107: out = 16'(101);
			2108: out = 16'(-580);
			2109: out = 16'(-1127);
			2110: out = 16'(1163);
			2111: out = 16'(-563);
			2112: out = 16'(-2988);
			2113: out = 16'(2971);
			2114: out = 16'(4996);
			2115: out = 16'(1916);
			2116: out = 16'(3461);
			2117: out = 16'(2186);
			2118: out = 16'(678);
			2119: out = 16'(2787);
			2120: out = 16'(-2021);
			2121: out = 16'(3069);
			2122: out = 16'(-2373);
			2123: out = 16'(-1389);
			2124: out = 16'(-209);
			2125: out = 16'(-3449);
			2126: out = 16'(25);
			2127: out = 16'(-832);
			2128: out = 16'(-1282);
			2129: out = 16'(1074);
			2130: out = 16'(4525);
			2131: out = 16'(652);
			2132: out = 16'(6245);
			2133: out = 16'(-569);
			2134: out = 16'(-1782);
			2135: out = 16'(-2507);
			2136: out = 16'(1609);
			2137: out = 16'(-3809);
			2138: out = 16'(1166);
			2139: out = 16'(-47);
			2140: out = 16'(-1690);
			2141: out = 16'(1776);
			2142: out = 16'(2668);
			2143: out = 16'(1101);
			2144: out = 16'(-2402);
			2145: out = 16'(-5154);
			2146: out = 16'(-14);
			2147: out = 16'(-3127);
			2148: out = 16'(-4455);
			2149: out = 16'(2085);
			2150: out = 16'(-2070);
			2151: out = 16'(-5120);
			2152: out = 16'(691);
			2153: out = 16'(-7394);
			2154: out = 16'(1078);
			2155: out = 16'(1411);
			2156: out = 16'(-4892);
			2157: out = 16'(-2645);
			2158: out = 16'(3042);
			2159: out = 16'(-5274);
			2160: out = 16'(-1376);
			2161: out = 16'(3871);
			2162: out = 16'(-347);
			2163: out = 16'(2652);
			2164: out = 16'(-860);
			2165: out = 16'(3436);
			2166: out = 16'(2111);
			2167: out = 16'(880);
			2168: out = 16'(339);
			2169: out = 16'(-481);
			2170: out = 16'(-6512);
			2171: out = 16'(414);
			2172: out = 16'(4755);
			2173: out = 16'(-928);
			2174: out = 16'(5278);
			2175: out = 16'(375);
			2176: out = 16'(67);
			2177: out = 16'(-8831);
			2178: out = 16'(2392);
			2179: out = 16'(-1543);
			2180: out = 16'(200);
			2181: out = 16'(-4704);
			2182: out = 16'(1719);
			2183: out = 16'(5586);
			2184: out = 16'(-2458);
			2185: out = 16'(-647);
			2186: out = 16'(-79);
			2187: out = 16'(-1767);
			2188: out = 16'(-3942);
			2189: out = 16'(2122);
			2190: out = 16'(-642);
			2191: out = 16'(1756);
			2192: out = 16'(974);
			2193: out = 16'(1104);
			2194: out = 16'(217);
			2195: out = 16'(48);
			2196: out = 16'(302);
			2197: out = 16'(1414);
			2198: out = 16'(3963);
			2199: out = 16'(-602);
			2200: out = 16'(-3557);
			2201: out = 16'(-2673);
			2202: out = 16'(1960);
			2203: out = 16'(-3410);
			2204: out = 16'(-1851);
			2205: out = 16'(3964);
			2206: out = 16'(-3565);
			2207: out = 16'(442);
			2208: out = 16'(1317);
			2209: out = 16'(-2361);
			2210: out = 16'(-5530);
			2211: out = 16'(2127);
			2212: out = 16'(-2465);
			2213: out = 16'(-2679);
			2214: out = 16'(3537);
			2215: out = 16'(458);
			2216: out = 16'(2474);
			2217: out = 16'(-2314);
			2218: out = 16'(-2442);
			2219: out = 16'(3974);
			2220: out = 16'(1155);
			2221: out = 16'(-788);
			2222: out = 16'(-89);
			2223: out = 16'(-1395);
			2224: out = 16'(363);
			2225: out = 16'(824);
			2226: out = 16'(-3580);
			2227: out = 16'(-516);
			2228: out = 16'(-346);
			2229: out = 16'(554);
			2230: out = 16'(771);
			2231: out = 16'(4483);
			2232: out = 16'(-1159);
			2233: out = 16'(1203);
			2234: out = 16'(879);
			2235: out = 16'(-165);
			2236: out = 16'(5031);
			2237: out = 16'(-5193);
			2238: out = 16'(1605);
			2239: out = 16'(-940);
			2240: out = 16'(2556);
			2241: out = 16'(-94);
			2242: out = 16'(4041);
			2243: out = 16'(-829);
			2244: out = 16'(-211);
			2245: out = 16'(-231);
			2246: out = 16'(907);
			2247: out = 16'(289);
			2248: out = 16'(-466);
			2249: out = 16'(2472);
			2250: out = 16'(-367);
			2251: out = 16'(348);
			2252: out = 16'(-874);
			2253: out = 16'(-1840);
			2254: out = 16'(-1525);
			2255: out = 16'(3461);
			2256: out = 16'(-7245);
			2257: out = 16'(709);
			2258: out = 16'(3398);
			2259: out = 16'(-4633);
			2260: out = 16'(2738);
			2261: out = 16'(-1341);
			2262: out = 16'(445);
			2263: out = 16'(-1883);
			2264: out = 16'(4189);
			2265: out = 16'(-3903);
			2266: out = 16'(1665);
			2267: out = 16'(-1037);
			2268: out = 16'(-1619);
			2269: out = 16'(2524);
			2270: out = 16'(-144);
			2271: out = 16'(-2770);
			2272: out = 16'(-2851);
			2273: out = 16'(1149);
			2274: out = 16'(-4374);
			2275: out = 16'(3011);
			2276: out = 16'(-604);
			2277: out = 16'(1583);
			2278: out = 16'(-3042);
			2279: out = 16'(-663);
			2280: out = 16'(3389);
			2281: out = 16'(-467);
			2282: out = 16'(-180);
			2283: out = 16'(2222);
			2284: out = 16'(866);
			2285: out = 16'(-8127);
			2286: out = 16'(2068);
			2287: out = 16'(-2759);
			2288: out = 16'(713);
			2289: out = 16'(-752);
			2290: out = 16'(1072);
			2291: out = 16'(-919);
			2292: out = 16'(2100);
			2293: out = 16'(986);
			2294: out = 16'(2821);
			2295: out = 16'(1761);
			2296: out = 16'(-171);
			2297: out = 16'(-490);
			2298: out = 16'(2831);
			2299: out = 16'(638);
			2300: out = 16'(3028);
			2301: out = 16'(2660);
			2302: out = 16'(292);
			2303: out = 16'(-1993);
			2304: out = 16'(-172);
			2305: out = 16'(3294);
			2306: out = 16'(517);
			2307: out = 16'(-176);
			2308: out = 16'(1951);
			2309: out = 16'(-269);
			2310: out = 16'(695);
			2311: out = 16'(600);
			2312: out = 16'(305);
			2313: out = 16'(3645);
			2314: out = 16'(2212);
			2315: out = 16'(-1339);
			2316: out = 16'(-418);
			2317: out = 16'(156);
			2318: out = 16'(-4322);
			2319: out = 16'(873);
			2320: out = 16'(1424);
			2321: out = 16'(1161);
			2322: out = 16'(-99);
			2323: out = 16'(130);
			2324: out = 16'(1023);
			2325: out = 16'(1815);
			2326: out = 16'(101);
			2327: out = 16'(-981);
			2328: out = 16'(429);
			2329: out = 16'(-5995);
			2330: out = 16'(-991);
			2331: out = 16'(-578);
			2332: out = 16'(768);
			2333: out = 16'(1671);
			2334: out = 16'(-1132);
			2335: out = 16'(3531);
			2336: out = 16'(-1321);
			2337: out = 16'(-155);
			2338: out = 16'(-589);
			2339: out = 16'(-589);
			2340: out = 16'(643);
			2341: out = 16'(1325);
			2342: out = 16'(2094);
			2343: out = 16'(493);
			2344: out = 16'(-4929);
			2345: out = 16'(-26);
			2346: out = 16'(2895);
			2347: out = 16'(-1928);
			2348: out = 16'(1625);
			2349: out = 16'(-2781);
			2350: out = 16'(150);
			2351: out = 16'(2238);
			2352: out = 16'(-1249);
			2353: out = 16'(-836);
			2354: out = 16'(1507);
			2355: out = 16'(306);
			2356: out = 16'(-3887);
			2357: out = 16'(-1028);
			2358: out = 16'(817);
			2359: out = 16'(-1820);
			2360: out = 16'(-3303);
			2361: out = 16'(585);
			2362: out = 16'(-1157);
			2363: out = 16'(1812);
			2364: out = 16'(933);
			2365: out = 16'(3267);
			2366: out = 16'(4213);
			2367: out = 16'(614);
			2368: out = 16'(3488);
			2369: out = 16'(-332);
			2370: out = 16'(-1518);
			2371: out = 16'(-421);
			2372: out = 16'(-960);
			2373: out = 16'(473);
			2374: out = 16'(-1022);
			2375: out = 16'(-4363);
			2376: out = 16'(3345);
			2377: out = 16'(-2370);
			2378: out = 16'(-184);
			2379: out = 16'(1769);
			2380: out = 16'(677);
			2381: out = 16'(-4023);
			2382: out = 16'(4022);
			2383: out = 16'(1143);
			2384: out = 16'(-1252);
			2385: out = 16'(-1958);
			2386: out = 16'(-1217);
			2387: out = 16'(-19);
			2388: out = 16'(-3455);
			2389: out = 16'(610);
			2390: out = 16'(2147);
			2391: out = 16'(-2968);
			2392: out = 16'(777);
			2393: out = 16'(-807);
			2394: out = 16'(-3204);
			2395: out = 16'(4135);
			2396: out = 16'(-993);
			2397: out = 16'(618);
			2398: out = 16'(729);
			2399: out = 16'(-605);
			2400: out = 16'(-5649);
			2401: out = 16'(2311);
			2402: out = 16'(-3094);
			2403: out = 16'(462);
			2404: out = 16'(139);
			2405: out = 16'(-3753);
			2406: out = 16'(120);
			2407: out = 16'(-1178);
			2408: out = 16'(-83);
			2409: out = 16'(1880);
			2410: out = 16'(-1081);
			2411: out = 16'(-1344);
			2412: out = 16'(2809);
			2413: out = 16'(-417);
			2414: out = 16'(-1858);
			2415: out = 16'(2393);
			2416: out = 16'(-2);
			2417: out = 16'(-3962);
			2418: out = 16'(-854);
			2419: out = 16'(473);
			2420: out = 16'(294);
			2421: out = 16'(178);
			2422: out = 16'(-3693);
			2423: out = 16'(3929);
			2424: out = 16'(-1820);
			2425: out = 16'(-3595);
			2426: out = 16'(795);
			2427: out = 16'(752);
			2428: out = 16'(-727);
			2429: out = 16'(-444);
			2430: out = 16'(-2091);
			2431: out = 16'(2032);
			2432: out = 16'(624);
			2433: out = 16'(374);
			2434: out = 16'(-984);
			2435: out = 16'(1065);
			2436: out = 16'(-3331);
			2437: out = 16'(-401);
			2438: out = 16'(-312);
			2439: out = 16'(1298);
			2440: out = 16'(-1620);
			2441: out = 16'(611);
			2442: out = 16'(2096);
			2443: out = 16'(-524);
			2444: out = 16'(1606);
			2445: out = 16'(182);
			2446: out = 16'(1199);
			2447: out = 16'(-5244);
			2448: out = 16'(-265);
			2449: out = 16'(-620);
			2450: out = 16'(-1916);
			2451: out = 16'(-51);
			2452: out = 16'(4);
			2453: out = 16'(562);
			2454: out = 16'(543);
			2455: out = 16'(-217);
			2456: out = 16'(131);
			2457: out = 16'(3415);
			2458: out = 16'(-5120);
			2459: out = 16'(1392);
			2460: out = 16'(210);
			2461: out = 16'(-4429);
			2462: out = 16'(-378);
			2463: out = 16'(-730);
			2464: out = 16'(1544);
			2465: out = 16'(1156);
			2466: out = 16'(-674);
			2467: out = 16'(295);
			2468: out = 16'(4735);
			2469: out = 16'(-194);
			2470: out = 16'(2219);
			2471: out = 16'(2770);
			2472: out = 16'(-3164);
			2473: out = 16'(-139);
			2474: out = 16'(-93);
			2475: out = 16'(-226);
			2476: out = 16'(-1923);
			2477: out = 16'(-1636);
			2478: out = 16'(74);
			2479: out = 16'(2449);
			2480: out = 16'(508);
			2481: out = 16'(2331);
			2482: out = 16'(1711);
			2483: out = 16'(-73);
			2484: out = 16'(263);
			2485: out = 16'(-2);
			2486: out = 16'(1511);
			2487: out = 16'(3693);
			2488: out = 16'(747);
			2489: out = 16'(-3017);
			2490: out = 16'(1201);
			2491: out = 16'(-3270);
			2492: out = 16'(-320);
			2493: out = 16'(-475);
			2494: out = 16'(1412);
			2495: out = 16'(2980);
			2496: out = 16'(1806);
			2497: out = 16'(1986);
			2498: out = 16'(2018);
			2499: out = 16'(1692);
			2500: out = 16'(-1011);
			2501: out = 16'(1515);
			2502: out = 16'(-2556);
			2503: out = 16'(-439);
			2504: out = 16'(-3889);
			2505: out = 16'(799);
			2506: out = 16'(1052);
			2507: out = 16'(-904);
			2508: out = 16'(1571);
			2509: out = 16'(-1846);
			2510: out = 16'(1817);
			2511: out = 16'(1072);
			2512: out = 16'(223);
			2513: out = 16'(1812);
			2514: out = 16'(32);
			2515: out = 16'(-803);
			2516: out = 16'(622);
			2517: out = 16'(-985);
			2518: out = 16'(-3985);
			2519: out = 16'(2930);
			2520: out = 16'(121);
			2521: out = 16'(-16);
			2522: out = 16'(1311);
			2523: out = 16'(-1334);
			2524: out = 16'(-1626);
			2525: out = 16'(-1296);
			2526: out = 16'(-5274);
			2527: out = 16'(1748);
			2528: out = 16'(-2020);
			2529: out = 16'(847);
			2530: out = 16'(-692);
			2531: out = 16'(1268);
			2532: out = 16'(-2338);
			2533: out = 16'(637);
			2534: out = 16'(932);
			2535: out = 16'(-2409);
			2536: out = 16'(-539);
			2537: out = 16'(-3022);
			2538: out = 16'(1211);
			2539: out = 16'(-1366);
			2540: out = 16'(-772);
			2541: out = 16'(229);
			2542: out = 16'(2646);
			2543: out = 16'(753);
			2544: out = 16'(1553);
			2545: out = 16'(1907);
			2546: out = 16'(267);
			2547: out = 16'(219);
			2548: out = 16'(684);
			2549: out = 16'(3760);
			2550: out = 16'(-1092);
			2551: out = 16'(-2023);
			2552: out = 16'(1584);
			2553: out = 16'(-2214);
			2554: out = 16'(992);
			2555: out = 16'(-1663);
			2556: out = 16'(554);
			2557: out = 16'(-2004);
			2558: out = 16'(-434);
			2559: out = 16'(-1548);
			2560: out = 16'(1405);
			2561: out = 16'(787);
			2562: out = 16'(-2007);
			2563: out = 16'(216);
			2564: out = 16'(-2291);
			2565: out = 16'(1423);
			2566: out = 16'(-220);
			2567: out = 16'(584);
			2568: out = 16'(686);
			2569: out = 16'(-458);
			2570: out = 16'(-1728);
			2571: out = 16'(-1529);
			2572: out = 16'(752);
			2573: out = 16'(-22);
			2574: out = 16'(421);
			2575: out = 16'(-1388);
			2576: out = 16'(141);
			2577: out = 16'(1387);
			2578: out = 16'(-3519);
			2579: out = 16'(-72);
			2580: out = 16'(-1346);
			2581: out = 16'(-3156);
			2582: out = 16'(372);
			2583: out = 16'(-466);
			2584: out = 16'(-1516);
			2585: out = 16'(1764);
			2586: out = 16'(948);
			2587: out = 16'(-574);
			2588: out = 16'(-4);
			2589: out = 16'(-455);
			2590: out = 16'(1853);
			2591: out = 16'(2942);
			2592: out = 16'(-619);
			2593: out = 16'(977);
			2594: out = 16'(-4080);
			2595: out = 16'(-1675);
			2596: out = 16'(1168);
			2597: out = 16'(1439);
			2598: out = 16'(2916);
			2599: out = 16'(-3448);
			2600: out = 16'(2311);
			2601: out = 16'(936);
			2602: out = 16'(1578);
			2603: out = 16'(822);
			2604: out = 16'(1494);
			2605: out = 16'(2428);
			2606: out = 16'(1732);
			2607: out = 16'(-214);
			2608: out = 16'(-3898);
			2609: out = 16'(2657);
			2610: out = 16'(-718);
			2611: out = 16'(614);
			2612: out = 16'(-4203);
			2613: out = 16'(1918);
			2614: out = 16'(-614);
			2615: out = 16'(984);
			2616: out = 16'(2895);
			2617: out = 16'(-1063);
			2618: out = 16'(-2197);
			2619: out = 16'(1600);
			2620: out = 16'(-1151);
			2621: out = 16'(-2747);
			2622: out = 16'(4377);
			2623: out = 16'(-166);
			2624: out = 16'(2292);
			2625: out = 16'(472);
			2626: out = 16'(-665);
			2627: out = 16'(-595);
			2628: out = 16'(1418);
			2629: out = 16'(-1843);
			2630: out = 16'(1840);
			2631: out = 16'(-570);
			2632: out = 16'(1346);
			2633: out = 16'(-1006);
			2634: out = 16'(885);
			2635: out = 16'(0);
			2636: out = 16'(-2773);
			2637: out = 16'(-1357);
			2638: out = 16'(860);
			2639: out = 16'(3222);
			2640: out = 16'(-3296);
			2641: out = 16'(551);
			2642: out = 16'(157);
			2643: out = 16'(-3730);
			2644: out = 16'(-115);
			2645: out = 16'(-72);
			2646: out = 16'(287);
			2647: out = 16'(947);
			2648: out = 16'(232);
			2649: out = 16'(-2158);
			2650: out = 16'(-600);
			2651: out = 16'(-2940);
			2652: out = 16'(-40);
			2653: out = 16'(1116);
			2654: out = 16'(-825);
			2655: out = 16'(192);
			2656: out = 16'(375);
			2657: out = 16'(1849);
			2658: out = 16'(1748);
			2659: out = 16'(406);
			2660: out = 16'(-235);
			2661: out = 16'(0);
			2662: out = 16'(520);
			2663: out = 16'(-454);
			2664: out = 16'(2460);
			2665: out = 16'(2030);
			2666: out = 16'(345);
			2667: out = 16'(-1428);
			2668: out = 16'(2495);
			2669: out = 16'(-921);
			2670: out = 16'(-998);
			2671: out = 16'(-655);
			2672: out = 16'(179);
			2673: out = 16'(-764);
			2674: out = 16'(-176);
			2675: out = 16'(-122);
			2676: out = 16'(130);
			2677: out = 16'(-657);
			2678: out = 16'(-253);
			2679: out = 16'(-1276);
			2680: out = 16'(-3141);
			2681: out = 16'(2467);
			2682: out = 16'(1151);
			2683: out = 16'(32);
			2684: out = 16'(-822);
			2685: out = 16'(-1601);
			2686: out = 16'(-4571);
			2687: out = 16'(2809);
			2688: out = 16'(-988);
			2689: out = 16'(-2214);
			2690: out = 16'(143);
			2691: out = 16'(684);
			2692: out = 16'(-163);
			2693: out = 16'(1492);
			2694: out = 16'(2942);
			2695: out = 16'(1173);
			2696: out = 16'(-242);
			2697: out = 16'(-2522);
			2698: out = 16'(-56);
			2699: out = 16'(-454);
			2700: out = 16'(-532);
			2701: out = 16'(296);
			2702: out = 16'(-1935);
			2703: out = 16'(-1825);
			2704: out = 16'(332);
			2705: out = 16'(2059);
			2706: out = 16'(31);
			2707: out = 16'(490);
			2708: out = 16'(1347);
			2709: out = 16'(-39);
			2710: out = 16'(-101);
			2711: out = 16'(-1378);
			2712: out = 16'(1203);
			2713: out = 16'(-109);
			2714: out = 16'(7);
			2715: out = 16'(-36);
			2716: out = 16'(17);
			2717: out = 16'(-4142);
			2718: out = 16'(-1715);
			2719: out = 16'(648);
			2720: out = 16'(-196);
			2721: out = 16'(-155);
			2722: out = 16'(-187);
			2723: out = 16'(-291);
			2724: out = 16'(-1676);
			2725: out = 16'(319);
			2726: out = 16'(84);
			2727: out = 16'(-1015);
			2728: out = 16'(144);
			2729: out = 16'(-1864);
			2730: out = 16'(-1175);
			2731: out = 16'(-1282);
			2732: out = 16'(392);
			2733: out = 16'(964);
			2734: out = 16'(1477);
			2735: out = 16'(-510);
			2736: out = 16'(417);
			2737: out = 16'(-1393);
			2738: out = 16'(3161);
			2739: out = 16'(2492);
			2740: out = 16'(-294);
			2741: out = 16'(-398);
			2742: out = 16'(-26);
			2743: out = 16'(-669);
			2744: out = 16'(-169);
			2745: out = 16'(2372);
			2746: out = 16'(-1794);
			2747: out = 16'(-229);
			2748: out = 16'(-1304);
			2749: out = 16'(1288);
			2750: out = 16'(18);
			2751: out = 16'(259);
			2752: out = 16'(-3024);
			2753: out = 16'(208);
			2754: out = 16'(-2731);
			2755: out = 16'(-1143);
			2756: out = 16'(2465);
			2757: out = 16'(1433);
			2758: out = 16'(1206);
			2759: out = 16'(-2192);
			2760: out = 16'(774);
			2761: out = 16'(-2166);
			2762: out = 16'(3880);
			2763: out = 16'(198);
			2764: out = 16'(341);
			2765: out = 16'(1077);
			2766: out = 16'(-1454);
			2767: out = 16'(-262);
			2768: out = 16'(275);
			2769: out = 16'(1818);
			2770: out = 16'(-1734);
			2771: out = 16'(1917);
			2772: out = 16'(-2384);
			2773: out = 16'(310);
			2774: out = 16'(-2529);
			2775: out = 16'(471);
			2776: out = 16'(1369);
			2777: out = 16'(-429);
			2778: out = 16'(-940);
			2779: out = 16'(309);
			2780: out = 16'(-1435);
			2781: out = 16'(-721);
			2782: out = 16'(-1117);
			2783: out = 16'(-3822);
			2784: out = 16'(92);
			2785: out = 16'(269);
			2786: out = 16'(1110);
			2787: out = 16'(940);
			2788: out = 16'(-154);
			2789: out = 16'(-63);
			2790: out = 16'(2010);
			2791: out = 16'(708);
			2792: out = 16'(-2205);
			2793: out = 16'(2079);
			2794: out = 16'(-311);
			2795: out = 16'(379);
			2796: out = 16'(5);
			2797: out = 16'(-1395);
			2798: out = 16'(2003);
			2799: out = 16'(-2029);
			2800: out = 16'(-353);
			2801: out = 16'(-568);
			2802: out = 16'(-972);
			2803: out = 16'(-919);
			2804: out = 16'(3622);
			2805: out = 16'(-319);
			2806: out = 16'(1333);
			2807: out = 16'(-2938);
			2808: out = 16'(-1902);
			2809: out = 16'(2472);
			2810: out = 16'(-624);
			2811: out = 16'(2598);
			2812: out = 16'(2240);
			2813: out = 16'(743);
			2814: out = 16'(-750);
			2815: out = 16'(408);
			2816: out = 16'(-102);
			2817: out = 16'(263);
			2818: out = 16'(1163);
			2819: out = 16'(-1312);
			2820: out = 16'(-550);
			2821: out = 16'(-1528);
			2822: out = 16'(898);
			2823: out = 16'(-1810);
			2824: out = 16'(2290);
			2825: out = 16'(-1409);
			2826: out = 16'(376);
			2827: out = 16'(-323);
			2828: out = 16'(918);
			2829: out = 16'(-555);
			2830: out = 16'(-2014);
			2831: out = 16'(315);
			2832: out = 16'(-1404);
			2833: out = 16'(2337);
			2834: out = 16'(-615);
			2835: out = 16'(1151);
			2836: out = 16'(-1668);
			2837: out = 16'(5);
			2838: out = 16'(-1019);
			2839: out = 16'(206);
			2840: out = 16'(4);
			2841: out = 16'(3087);
			2842: out = 16'(-220);
			2843: out = 16'(291);
			2844: out = 16'(-189);
			2845: out = 16'(-2298);
			2846: out = 16'(1920);
			2847: out = 16'(166);
			2848: out = 16'(704);
			2849: out = 16'(-2372);
			2850: out = 16'(-18);
			2851: out = 16'(-1831);
			2852: out = 16'(1954);
			2853: out = 16'(-1582);
			2854: out = 16'(266);
			2855: out = 16'(883);
			2856: out = 16'(-1105);
			2857: out = 16'(181);
			2858: out = 16'(-293);
			2859: out = 16'(746);
			2860: out = 16'(-972);
			2861: out = 16'(3338);
			2862: out = 16'(-167);
			2863: out = 16'(452);
			2864: out = 16'(-835);
			2865: out = 16'(-249);
			2866: out = 16'(-450);
			2867: out = 16'(16);
			2868: out = 16'(1732);
			2869: out = 16'(719);
			2870: out = 16'(-677);
			2871: out = 16'(-207);
			2872: out = 16'(-1469);
			2873: out = 16'(-1009);
			2874: out = 16'(736);
			2875: out = 16'(5);
			2876: out = 16'(403);
			2877: out = 16'(572);
			2878: out = 16'(-393);
			2879: out = 16'(2520);
			2880: out = 16'(-2762);
			2881: out = 16'(675);
			2882: out = 16'(472);
			2883: out = 16'(-731);
			2884: out = 16'(1479);
			2885: out = 16'(-474);
			2886: out = 16'(1124);
			2887: out = 16'(340);
			2888: out = 16'(-69);
			2889: out = 16'(-51);
			2890: out = 16'(203);
			2891: out = 16'(-2017);
			2892: out = 16'(739);
			2893: out = 16'(-469);
			2894: out = 16'(-204);
			2895: out = 16'(-1877);
			2896: out = 16'(1337);
			2897: out = 16'(-337);
			2898: out = 16'(-681);
			2899: out = 16'(-67);
			2900: out = 16'(-4599);
			2901: out = 16'(1858);
			2902: out = 16'(-267);
			2903: out = 16'(683);
			2904: out = 16'(527);
			2905: out = 16'(1165);
			2906: out = 16'(-942);
			2907: out = 16'(188);
			2908: out = 16'(569);
			2909: out = 16'(89);
			2910: out = 16'(251);
			2911: out = 16'(-312);
			2912: out = 16'(277);
			2913: out = 16'(-2648);
			2914: out = 16'(-239);
			2915: out = 16'(-1191);
			2916: out = 16'(2632);
			2917: out = 16'(-2367);
			2918: out = 16'(240);
			2919: out = 16'(689);
			2920: out = 16'(458);
			2921: out = 16'(756);
			2922: out = 16'(-779);
			2923: out = 16'(1339);
			2924: out = 16'(-275);
			2925: out = 16'(-1090);
			2926: out = 16'(-353);
			2927: out = 16'(340);
			2928: out = 16'(-164);
			2929: out = 16'(-351);
			2930: out = 16'(383);
			2931: out = 16'(-285);
			2932: out = 16'(-635);
			2933: out = 16'(709);
			2934: out = 16'(1030);
			2935: out = 16'(1892);
			2936: out = 16'(-336);
			2937: out = 16'(470);
			2938: out = 16'(136);
			2939: out = 16'(95);
			2940: out = 16'(-250);
			2941: out = 16'(1966);
			2942: out = 16'(-1688);
			2943: out = 16'(-540);
			2944: out = 16'(724);
			2945: out = 16'(309);
			2946: out = 16'(-1266);
			2947: out = 16'(1066);
			2948: out = 16'(-1548);
			2949: out = 16'(3285);
			2950: out = 16'(-49);
			2951: out = 16'(-1356);
			2952: out = 16'(-1031);
			2953: out = 16'(425);
			2954: out = 16'(403);
			2955: out = 16'(-1685);
			2956: out = 16'(-143);
			2957: out = 16'(-362);
			2958: out = 16'(2094);
			2959: out = 16'(197);
			2960: out = 16'(226);
			2961: out = 16'(-628);
			2962: out = 16'(-179);
			2963: out = 16'(136);
			2964: out = 16'(1725);
			2965: out = 16'(359);
			2966: out = 16'(327);
			2967: out = 16'(1340);
			2968: out = 16'(-670);
			2969: out = 16'(902);
			2970: out = 16'(-850);
			2971: out = 16'(3630);
			2972: out = 16'(689);
			2973: out = 16'(-104);
			2974: out = 16'(-117);
			2975: out = 16'(293);
			2976: out = 16'(1281);
			2977: out = 16'(-436);
			2978: out = 16'(-548);
			2979: out = 16'(-2056);
			2980: out = 16'(1849);
			2981: out = 16'(210);
			2982: out = 16'(1121);
			2983: out = 16'(-1319);
			2984: out = 16'(117);
			2985: out = 16'(-1333);
			2986: out = 16'(1621);
			2987: out = 16'(280);
			2988: out = 16'(-1844);
			2989: out = 16'(-862);
			2990: out = 16'(371);
			2991: out = 16'(57);
			2992: out = 16'(-1296);
			2993: out = 16'(1302);
			2994: out = 16'(-952);
			2995: out = 16'(427);
			2996: out = 16'(331);
			2997: out = 16'(1955);
			2998: out = 16'(-1143);
			2999: out = 16'(1200);
			3000: out = 16'(-660);
			3001: out = 16'(-74);
			3002: out = 16'(-1373);
			3003: out = 16'(-1464);
			3004: out = 16'(1793);
			3005: out = 16'(-1495);
			3006: out = 16'(2101);
			3007: out = 16'(881);
			3008: out = 16'(-348);
			3009: out = 16'(-675);
			3010: out = 16'(-1433);
			3011: out = 16'(-2036);
			3012: out = 16'(569);
			3013: out = 16'(-1207);
			3014: out = 16'(696);
			3015: out = 16'(1581);
			3016: out = 16'(-4356);
			3017: out = 16'(1836);
			3018: out = 16'(-592);
			3019: out = 16'(174);
			3020: out = 16'(108);
			3021: out = 16'(-17);
			3022: out = 16'(1006);
			3023: out = 16'(694);
			3024: out = 16'(1051);
			3025: out = 16'(-85);
			3026: out = 16'(-737);
			3027: out = 16'(896);
			3028: out = 16'(528);
			3029: out = 16'(-784);
			3030: out = 16'(-229);
			3031: out = 16'(924);
			3032: out = 16'(-156);
			3033: out = 16'(119);
			3034: out = 16'(-1538);
			3035: out = 16'(-459);
			3036: out = 16'(1101);
			3037: out = 16'(-310);
			3038: out = 16'(-650);
			3039: out = 16'(483);
			3040: out = 16'(-1385);
			3041: out = 16'(170);
			3042: out = 16'(478);
			3043: out = 16'(-1916);
			3044: out = 16'(1573);
			3045: out = 16'(-406);
			3046: out = 16'(333);
			3047: out = 16'(-489);
			3048: out = 16'(1550);
			3049: out = 16'(282);
			3050: out = 16'(1016);
			3051: out = 16'(143);
			3052: out = 16'(2415);
			3053: out = 16'(-429);
			3054: out = 16'(-119);
			3055: out = 16'(-253);
			3056: out = 16'(-1034);
			3057: out = 16'(714);
			3058: out = 16'(-3153);
			3059: out = 16'(1124);
			3060: out = 16'(-621);
			3061: out = 16'(1148);
			3062: out = 16'(-2014);
			3063: out = 16'(416);
			3064: out = 16'(-1038);
			3065: out = 16'(921);
			3066: out = 16'(-1512);
			3067: out = 16'(-1182);
			3068: out = 16'(704);
			3069: out = 16'(1073);
			3070: out = 16'(1111);
			3071: out = 16'(-717);
			3072: out = 16'(612);
			3073: out = 16'(-2025);
			3074: out = 16'(1776);
			3075: out = 16'(1309);
			3076: out = 16'(213);
			3077: out = 16'(-454);
			3078: out = 16'(681);
			3079: out = 16'(572);
			3080: out = 16'(-708);
			3081: out = 16'(-140);
			3082: out = 16'(168);
			3083: out = 16'(288);
			3084: out = 16'(-190);
			3085: out = 16'(-1217);
			3086: out = 16'(-1617);
			3087: out = 16'(1328);
			3088: out = 16'(426);
			3089: out = 16'(472);
			3090: out = 16'(644);
			3091: out = 16'(-718);
			3092: out = 16'(1277);
			3093: out = 16'(975);
			3094: out = 16'(-686);
			3095: out = 16'(-158);
			3096: out = 16'(-749);
			3097: out = 16'(-354);
			3098: out = 16'(1635);
			3099: out = 16'(-1583);
			3100: out = 16'(-2);
			3101: out = 16'(709);
			3102: out = 16'(-2233);
			3103: out = 16'(2588);
			3104: out = 16'(1655);
			3105: out = 16'(1886);
			3106: out = 16'(911);
			3107: out = 16'(68);
			3108: out = 16'(-730);
			3109: out = 16'(-539);
			3110: out = 16'(-1201);
			3111: out = 16'(7);
			3112: out = 16'(-321);
			3113: out = 16'(-3356);
			3114: out = 16'(43);
			3115: out = 16'(-227);
			3116: out = 16'(1828);
			3117: out = 16'(-3112);
			3118: out = 16'(638);
			3119: out = 16'(-102);
			3120: out = 16'(-1167);
			3121: out = 16'(340);
			3122: out = 16'(209);
			3123: out = 16'(116);
			3124: out = 16'(540);
			3125: out = 16'(2157);
			3126: out = 16'(-967);
			3127: out = 16'(2030);
			3128: out = 16'(-1161);
			3129: out = 16'(433);
			3130: out = 16'(571);
			3131: out = 16'(-1274);
			3132: out = 16'(1049);
			3133: out = 16'(-1051);
			3134: out = 16'(1537);
			3135: out = 16'(-1258);
			3136: out = 16'(1748);
			3137: out = 16'(-2342);
			3138: out = 16'(386);
			3139: out = 16'(-240);
			3140: out = 16'(-386);
			3141: out = 16'(-1037);
			3142: out = 16'(84);
			3143: out = 16'(-251);
			3144: out = 16'(209);
			3145: out = 16'(-520);
			3146: out = 16'(-1099);
			3147: out = 16'(837);
			3148: out = 16'(1010);
			3149: out = 16'(2248);
			3150: out = 16'(239);
			3151: out = 16'(170);
			3152: out = 16'(-818);
			3153: out = 16'(863);
			3154: out = 16'(-417);
			3155: out = 16'(-602);
			3156: out = 16'(-1642);
			3157: out = 16'(-1655);
			3158: out = 16'(1574);
			3159: out = 16'(-156);
			3160: out = 16'(1122);
			3161: out = 16'(-1906);
			3162: out = 16'(200);
			3163: out = 16'(-905);
			3164: out = 16'(112);
			3165: out = 16'(-297);
			3166: out = 16'(94);
			3167: out = 16'(-813);
			3168: out = 16'(3);
			3169: out = 16'(-1564);
			3170: out = 16'(131);
			3171: out = 16'(1876);
			3172: out = 16'(633);
			3173: out = 16'(75);
			3174: out = 16'(668);
			3175: out = 16'(-1351);
			3176: out = 16'(-1352);
			3177: out = 16'(-420);
			3178: out = 16'(309);
			3179: out = 16'(-232);
			3180: out = 16'(523);
			3181: out = 16'(-437);
			3182: out = 16'(-168);
			3183: out = 16'(180);
			3184: out = 16'(-1246);
			3185: out = 16'(1203);
			3186: out = 16'(-758);
			3187: out = 16'(87);
			3188: out = 16'(-2452);
			3189: out = 16'(1071);
			3190: out = 16'(-408);
			3191: out = 16'(1703);
			3192: out = 16'(-852);
			3193: out = 16'(932);
			3194: out = 16'(-32);
			3195: out = 16'(415);
			3196: out = 16'(499);
			3197: out = 16'(-396);
			3198: out = 16'(1444);
			3199: out = 16'(-1);
			3200: out = 16'(-334);
			3201: out = 16'(1577);
			3202: out = 16'(258);
			3203: out = 16'(-1068);
			3204: out = 16'(1950);
			3205: out = 16'(-706);
			3206: out = 16'(-59);
			3207: out = 16'(775);
			3208: out = 16'(-865);
			3209: out = 16'(-479);
			3210: out = 16'(117);
			3211: out = 16'(214);
			3212: out = 16'(-1258);
			3213: out = 16'(-1317);
			3214: out = 16'(79);
			3215: out = 16'(28);
			3216: out = 16'(-101);
			3217: out = 16'(496);
			3218: out = 16'(303);
			3219: out = 16'(56);
			3220: out = 16'(1030);
			3221: out = 16'(-1333);
			3222: out = 16'(464);
			3223: out = 16'(786);
			3224: out = 16'(1322);
			3225: out = 16'(324);
			3226: out = 16'(858);
			3227: out = 16'(367);
			3228: out = 16'(25);
			3229: out = 16'(-2850);
			3230: out = 16'(-437);
			3231: out = 16'(-95);
			3232: out = 16'(-497);
			3233: out = 16'(1191);
			3234: out = 16'(217);
			3235: out = 16'(-1766);
			3236: out = 16'(1561);
			3237: out = 16'(1056);
			3238: out = 16'(1608);
			3239: out = 16'(455);
			3240: out = 16'(-573);
			3241: out = 16'(949);
			3242: out = 16'(1489);
			3243: out = 16'(-1767);
			3244: out = 16'(470);
			3245: out = 16'(751);
			3246: out = 16'(-1402);
			3247: out = 16'(840);
			3248: out = 16'(-224);
			3249: out = 16'(432);
			3250: out = 16'(519);
			3251: out = 16'(-93);
			3252: out = 16'(54);
			3253: out = 16'(1894);
			3254: out = 16'(324);
			3255: out = 16'(555);
			3256: out = 16'(-2790);
			3257: out = 16'(-2637);
			3258: out = 16'(-2599);
			3259: out = 16'(-436);
			3260: out = 16'(-52);
			3261: out = 16'(-259);
			3262: out = 16'(-1444);
			3263: out = 16'(856);
			3264: out = 16'(1298);
			3265: out = 16'(-72);
			3266: out = 16'(327);
			3267: out = 16'(46);
			3268: out = 16'(793);
			3269: out = 16'(1258);
			3270: out = 16'(-968);
			3271: out = 16'(416);
			3272: out = 16'(101);
			3273: out = 16'(7);
			3274: out = 16'(984);
			3275: out = 16'(-386);
			3276: out = 16'(-844);
			3277: out = 16'(1024);
			3278: out = 16'(-545);
			3279: out = 16'(-26);
			3280: out = 16'(-418);
			3281: out = 16'(347);
			3282: out = 16'(867);
			3283: out = 16'(1280);
			3284: out = 16'(-867);
			3285: out = 16'(-251);
			3286: out = 16'(903);
			3287: out = 16'(-1167);
			3288: out = 16'(-159);
			3289: out = 16'(-7);
			3290: out = 16'(555);
			3291: out = 16'(302);
			3292: out = 16'(152);
			3293: out = 16'(-414);
			3294: out = 16'(-241);
			3295: out = 16'(-1499);
			3296: out = 16'(320);
			3297: out = 16'(-528);
			3298: out = 16'(-320);
			3299: out = 16'(795);
			3300: out = 16'(1002);
			3301: out = 16'(-122);
			3302: out = 16'(94);
			3303: out = 16'(258);
			3304: out = 16'(123);
			3305: out = 16'(662);
			3306: out = 16'(59);
			3307: out = 16'(20);
			3308: out = 16'(-1008);
			3309: out = 16'(68);
			3310: out = 16'(-1848);
			3311: out = 16'(-487);
			3312: out = 16'(1078);
			3313: out = 16'(-316);
			3314: out = 16'(777);
			3315: out = 16'(397);
			3316: out = 16'(1025);
			3317: out = 16'(352);
			3318: out = 16'(245);
			3319: out = 16'(605);
			3320: out = 16'(147);
			3321: out = 16'(-1310);
			3322: out = 16'(380);
			3323: out = 16'(424);
			3324: out = 16'(278);
			3325: out = 16'(-754);
			3326: out = 16'(-28);
			3327: out = 16'(173);
			3328: out = 16'(-1029);
			3329: out = 16'(477);
			3330: out = 16'(886);
			3331: out = 16'(125);
			3332: out = 16'(7);
			3333: out = 16'(1315);
			3334: out = 16'(-1666);
			3335: out = 16'(-336);
			3336: out = 16'(662);
			3337: out = 16'(156);
			3338: out = 16'(710);
			3339: out = 16'(2288);
			3340: out = 16'(-958);
			3341: out = 16'(2200);
			3342: out = 16'(1267);
			3343: out = 16'(-24);
			3344: out = 16'(-698);
			3345: out = 16'(-1737);
			3346: out = 16'(-607);
			3347: out = 16'(-895);
			3348: out = 16'(177);
			3349: out = 16'(340);
			3350: out = 16'(398);
			3351: out = 16'(-296);
			3352: out = 16'(-49);
			3353: out = 16'(-112);
			3354: out = 16'(151);
			3355: out = 16'(214);
			3356: out = 16'(1362);
			3357: out = 16'(-278);
			3358: out = 16'(46);
			3359: out = 16'(-2262);
			3360: out = 16'(-267);
			3361: out = 16'(367);
			3362: out = 16'(-7);
			3363: out = 16'(-420);
			3364: out = 16'(303);
			3365: out = 16'(-367);
			3366: out = 16'(375);
			3367: out = 16'(-121);
			3368: out = 16'(-1361);
			3369: out = 16'(2087);
			3370: out = 16'(611);
			3371: out = 16'(571);
			3372: out = 16'(463);
			3373: out = 16'(419);
			3374: out = 16'(288);
			3375: out = 16'(-78);
			3376: out = 16'(-252);
			3377: out = 16'(-285);
			3378: out = 16'(-1638);
			3379: out = 16'(-198);
			3380: out = 16'(-99);
			3381: out = 16'(336);
			3382: out = 16'(948);
			3383: out = 16'(-195);
			3384: out = 16'(2356);
			3385: out = 16'(183);
			3386: out = 16'(141);
			3387: out = 16'(-373);
			3388: out = 16'(-825);
			3389: out = 16'(-812);
			3390: out = 16'(646);
			3391: out = 16'(-957);
			3392: out = 16'(1198);
			3393: out = 16'(78);
			3394: out = 16'(-891);
			3395: out = 16'(-801);
			3396: out = 16'(599);
			3397: out = 16'(1433);
			3398: out = 16'(890);
			3399: out = 16'(343);
			3400: out = 16'(-1195);
			3401: out = 16'(309);
			3402: out = 16'(-1658);
			3403: out = 16'(-141);
			3404: out = 16'(-1283);
			3405: out = 16'(-652);
			3406: out = 16'(-19);
			3407: out = 16'(8);
			3408: out = 16'(-442);
			3409: out = 16'(53);
			3410: out = 16'(-1463);
			3411: out = 16'(-1800);
			3412: out = 16'(-686);
			3413: out = 16'(89);
			3414: out = 16'(-16);
			3415: out = 16'(663);
			3416: out = 16'(-556);
			3417: out = 16'(604);
			3418: out = 16'(206);
			3419: out = 16'(2265);
			3420: out = 16'(-141);
			3421: out = 16'(-736);
			3422: out = 16'(398);
			3423: out = 16'(-1159);
			3424: out = 16'(-198);
			3425: out = 16'(284);
			3426: out = 16'(-1276);
			3427: out = 16'(319);
			3428: out = 16'(-57);
			3429: out = 16'(-785);
			3430: out = 16'(-421);
			3431: out = 16'(1080);
			3432: out = 16'(-842);
			3433: out = 16'(-52);
			3434: out = 16'(628);
			3435: out = 16'(-2290);
			3436: out = 16'(495);
			3437: out = 16'(353);
			3438: out = 16'(-450);
			3439: out = 16'(2063);
			3440: out = 16'(-1119);
			3441: out = 16'(-41);
			3442: out = 16'(809);
			3443: out = 16'(-2025);
			3444: out = 16'(-1467);
			3445: out = 16'(1003);
			3446: out = 16'(-1587);
			3447: out = 16'(-737);
			3448: out = 16'(656);
			3449: out = 16'(91);
			3450: out = 16'(1028);
			3451: out = 16'(407);
			3452: out = 16'(110);
			3453: out = 16'(-207);
			3454: out = 16'(-294);
			3455: out = 16'(-764);
			3456: out = 16'(-527);
			3457: out = 16'(-942);
			3458: out = 16'(261);
			3459: out = 16'(293);
			3460: out = 16'(-1063);
			3461: out = 16'(1598);
			3462: out = 16'(128);
			3463: out = 16'(-458);
			3464: out = 16'(160);
			3465: out = 16'(192);
			3466: out = 16'(-315);
			3467: out = 16'(54);
			3468: out = 16'(619);
			3469: out = 16'(259);
			3470: out = 16'(-120);
			3471: out = 16'(-431);
			3472: out = 16'(-538);
			3473: out = 16'(-1590);
			3474: out = 16'(709);
			3475: out = 16'(-692);
			3476: out = 16'(668);
			3477: out = 16'(-389);
			3478: out = 16'(-604);
			3479: out = 16'(-178);
			3480: out = 16'(-301);
			3481: out = 16'(-847);
			3482: out = 16'(675);
			3483: out = 16'(606);
			3484: out = 16'(580);
			3485: out = 16'(1154);
			3486: out = 16'(-673);
			3487: out = 16'(236);
			3488: out = 16'(-41);
			3489: out = 16'(599);
			3490: out = 16'(151);
			3491: out = 16'(1334);
			3492: out = 16'(-561);
			3493: out = 16'(165);
			3494: out = 16'(-56);
			3495: out = 16'(867);
			3496: out = 16'(109);
			3497: out = 16'(-26);
			3498: out = 16'(-494);
			3499: out = 16'(-854);
			3500: out = 16'(491);
			3501: out = 16'(86);
			3502: out = 16'(249);
			3503: out = 16'(-665);
			3504: out = 16'(1804);
			3505: out = 16'(-1035);
			3506: out = 16'(-418);
			3507: out = 16'(316);
			3508: out = 16'(-1374);
			3509: out = 16'(294);
			3510: out = 16'(83);
			3511: out = 16'(-1955);
			3512: out = 16'(824);
			3513: out = 16'(-394);
			3514: out = 16'(-944);
			3515: out = 16'(968);
			3516: out = 16'(547);
			3517: out = 16'(177);
			3518: out = 16'(-196);
			3519: out = 16'(1116);
			3520: out = 16'(-337);
			3521: out = 16'(-16);
			3522: out = 16'(-1120);
			3523: out = 16'(-904);
			3524: out = 16'(-1924);
			3525: out = 16'(-503);
			3526: out = 16'(402);
			3527: out = 16'(-651);
			3528: out = 16'(-117);
			3529: out = 16'(-350);
			3530: out = 16'(-199);
			3531: out = 16'(1113);
			3532: out = 16'(734);
			3533: out = 16'(365);
			3534: out = 16'(906);
			3535: out = 16'(-105);
			3536: out = 16'(471);
			3537: out = 16'(667);
			3538: out = 16'(-601);
			3539: out = 16'(477);
			3540: out = 16'(399);
			3541: out = 16'(516);
			3542: out = 16'(877);
			3543: out = 16'(-2019);
			3544: out = 16'(133);
			3545: out = 16'(-448);
			3546: out = 16'(142);
			3547: out = 16'(-930);
			3548: out = 16'(442);
			3549: out = 16'(-1426);
			3550: out = 16'(1863);
			3551: out = 16'(247);
			3552: out = 16'(328);
			3553: out = 16'(-1705);
			3554: out = 16'(-1149);
			3555: out = 16'(474);
			3556: out = 16'(262);
			3557: out = 16'(-252);
			3558: out = 16'(-2283);
			3559: out = 16'(4);
			3560: out = 16'(-284);
			3561: out = 16'(-1565);
			3562: out = 16'(174);
			3563: out = 16'(111);
			3564: out = 16'(-26);
			3565: out = 16'(499);
			3566: out = 16'(-324);
			3567: out = 16'(-295);
			3568: out = 16'(231);
			3569: out = 16'(-70);
			3570: out = 16'(-41);
			3571: out = 16'(-899);
			3572: out = 16'(-33);
			3573: out = 16'(-201);
			3574: out = 16'(983);
			3575: out = 16'(-64);
			3576: out = 16'(-164);
			3577: out = 16'(-453);
			3578: out = 16'(768);
			3579: out = 16'(374);
			3580: out = 16'(-957);
			3581: out = 16'(252);
			3582: out = 16'(1000);
			3583: out = 16'(-318);
			3584: out = 16'(-718);
			3585: out = 16'(1415);
			3586: out = 16'(121);
			3587: out = 16'(119);
			3588: out = 16'(591);
			3589: out = 16'(-194);
			3590: out = 16'(-464);
			3591: out = 16'(-1449);
			3592: out = 16'(-162);
			3593: out = 16'(137);
			3594: out = 16'(273);
			3595: out = 16'(-874);
			3596: out = 16'(-16);
			3597: out = 16'(466);
			3598: out = 16'(1271);
			3599: out = 16'(67);
			3600: out = 16'(-1756);
			3601: out = 16'(454);
			3602: out = 16'(-1731);
			3603: out = 16'(1188);
			3604: out = 16'(-141);
			3605: out = 16'(783);
			3606: out = 16'(-375);
			3607: out = 16'(-7);
			3608: out = 16'(-186);
			3609: out = 16'(1434);
			3610: out = 16'(153);
			3611: out = 16'(-133);
			3612: out = 16'(642);
			3613: out = 16'(-617);
			3614: out = 16'(-428);
			3615: out = 16'(-149);
			3616: out = 16'(-560);
			3617: out = 16'(219);
			3618: out = 16'(-601);
			3619: out = 16'(76);
			3620: out = 16'(-416);
			3621: out = 16'(51);
			3622: out = 16'(51);
			3623: out = 16'(663);
			3624: out = 16'(6);
			3625: out = 16'(155);
			3626: out = 16'(-294);
			3627: out = 16'(240);
			3628: out = 16'(-475);
			3629: out = 16'(200);
			3630: out = 16'(-8);
			3631: out = 16'(243);
			3632: out = 16'(2069);
			3633: out = 16'(1310);
			3634: out = 16'(932);
			3635: out = 16'(484);
			3636: out = 16'(171);
			3637: out = 16'(-2024);
			3638: out = 16'(23);
			3639: out = 16'(-289);
			3640: out = 16'(-341);
			3641: out = 16'(616);
			3642: out = 16'(157);
			3643: out = 16'(119);
			3644: out = 16'(-405);
			3645: out = 16'(-235);
			3646: out = 16'(-508);
			3647: out = 16'(1093);
			3648: out = 16'(-68);
			3649: out = 16'(1087);
			3650: out = 16'(-480);
			3651: out = 16'(-961);
			3652: out = 16'(-276);
			3653: out = 16'(31);
			3654: out = 16'(198);
			3655: out = 16'(-708);
			3656: out = 16'(792);
			3657: out = 16'(-542);
			3658: out = 16'(483);
			3659: out = 16'(25);
			3660: out = 16'(109);
			3661: out = 16'(-873);
			3662: out = 16'(608);
			3663: out = 16'(544);
			3664: out = 16'(-502);
			3665: out = 16'(229);
			3666: out = 16'(-123);
			3667: out = 16'(-634);
			3668: out = 16'(1195);
			3669: out = 16'(-221);
			3670: out = 16'(-207);
			3671: out = 16'(42);
			3672: out = 16'(117);
			3673: out = 16'(-944);
			3674: out = 16'(190);
			3675: out = 16'(948);
			3676: out = 16'(174);
			3677: out = 16'(119);
			3678: out = 16'(-383);
			3679: out = 16'(833);
			3680: out = 16'(-713);
			3681: out = 16'(97);
			3682: out = 16'(228);
			3683: out = 16'(-301);
			3684: out = 16'(25);
			3685: out = 16'(35);
			3686: out = 16'(-967);
			3687: out = 16'(865);
			3688: out = 16'(-1074);
			3689: out = 16'(-52);
			3690: out = 16'(-10);
			3691: out = 16'(1019);
			3692: out = 16'(-702);
			3693: out = 16'(66);
			3694: out = 16'(-134);
			3695: out = 16'(97);
			3696: out = 16'(470);
			3697: out = 16'(-472);
			3698: out = 16'(16);
			3699: out = 16'(-49);
			3700: out = 16'(39);
			3701: out = 16'(-672);
			3702: out = 16'(794);
			3703: out = 16'(-129);
			3704: out = 16'(1019);
			3705: out = 16'(-987);
			3706: out = 16'(-138);
			3707: out = 16'(-457);
			3708: out = 16'(-1630);
			3709: out = 16'(915);
			3710: out = 16'(28);
			3711: out = 16'(254);
			3712: out = 16'(-194);
			3713: out = 16'(203);
			3714: out = 16'(-744);
			3715: out = 16'(546);
			3716: out = 16'(-288);
			3717: out = 16'(-304);
			3718: out = 16'(89);
			3719: out = 16'(-83);
			3720: out = 16'(-476);
			3721: out = 16'(-320);
			3722: out = 16'(-746);
			3723: out = 16'(-602);
			3724: out = 16'(-42);
			3725: out = 16'(-135);
			3726: out = 16'(675);
			3727: out = 16'(1350);
			3728: out = 16'(272);
			3729: out = 16'(-1133);
			3730: out = 16'(718);
			3731: out = 16'(99);
			3732: out = 16'(268);
			3733: out = 16'(106);
			3734: out = 16'(331);
			3735: out = 16'(-660);
			3736: out = 16'(-93);
			3737: out = 16'(-115);
			3738: out = 16'(-743);
			3739: out = 16'(168);
			3740: out = 16'(403);
			3741: out = 16'(-46);
			3742: out = 16'(-1187);
			3743: out = 16'(-522);
			3744: out = 16'(910);
			3745: out = 16'(-251);
			3746: out = 16'(-575);
			3747: out = 16'(303);
			3748: out = 16'(-90);
			3749: out = 16'(519);
			3750: out = 16'(178);
			3751: out = 16'(-1019);
			3752: out = 16'(305);
			3753: out = 16'(267);
			3754: out = 16'(-1230);
			3755: out = 16'(-434);
			3756: out = 16'(-70);
			3757: out = 16'(-1211);
			3758: out = 16'(-1260);
			3759: out = 16'(-396);
			3760: out = 16'(178);
			3761: out = 16'(568);
			3762: out = 16'(205);
			3763: out = 16'(567);
			3764: out = 16'(332);
			3765: out = 16'(-2019);
			3766: out = 16'(174);
			3767: out = 16'(709);
			3768: out = 16'(48);
			3769: out = 16'(109);
			3770: out = 16'(-485);
			3771: out = 16'(352);
			3772: out = 16'(129);
			3773: out = 16'(42);
			3774: out = 16'(-587);
			3775: out = 16'(940);
			3776: out = 16'(-130);
			3777: out = 16'(12);
			3778: out = 16'(688);
			3779: out = 16'(-326);
			3780: out = 16'(74);
			3781: out = 16'(711);
			3782: out = 16'(-250);
			3783: out = 16'(-127);
			3784: out = 16'(-192);
			3785: out = 16'(-8);
			3786: out = 16'(958);
			3787: out = 16'(-115);
			3788: out = 16'(-442);
			3789: out = 16'(255);
			3790: out = 16'(-455);
			3791: out = 16'(-323);
			3792: out = 16'(628);
			3793: out = 16'(-552);
			3794: out = 16'(-357);
			3795: out = 16'(-46);
			3796: out = 16'(1012);
			3797: out = 16'(183);
			3798: out = 16'(138);
			3799: out = 16'(-1048);
			3800: out = 16'(478);
			3801: out = 16'(-85);
			3802: out = 16'(-166);
			3803: out = 16'(-1359);
			3804: out = 16'(-196);
			3805: out = 16'(257);
			3806: out = 16'(-360);
			3807: out = 16'(567);
			3808: out = 16'(114);
			3809: out = 16'(303);
			3810: out = 16'(-54);
			3811: out = 16'(198);
			3812: out = 16'(537);
			3813: out = 16'(-64);
			3814: out = 16'(-582);
			3815: out = 16'(933);
			3816: out = 16'(-298);
			3817: out = 16'(649);
			3818: out = 16'(520);
			3819: out = 16'(-332);
			3820: out = 16'(-13);
			3821: out = 16'(482);
			3822: out = 16'(-393);
			3823: out = 16'(516);
			3824: out = 16'(-438);
			3825: out = 16'(-1092);
			3826: out = 16'(-871);
			3827: out = 16'(-224);
			3828: out = 16'(947);
			3829: out = 16'(179);
			3830: out = 16'(97);
			3831: out = 16'(-997);
			3832: out = 16'(-143);
			3833: out = 16'(668);
			3834: out = 16'(-37);
			3835: out = 16'(-32);
			3836: out = 16'(-490);
			3837: out = 16'(-695);
			3838: out = 16'(-367);
			3839: out = 16'(-8);
			3840: out = 16'(49);
			3841: out = 16'(-176);
			3842: out = 16'(-337);
			3843: out = 16'(-312);
			3844: out = 16'(566);
			3845: out = 16'(76);
			3846: out = 16'(-120);
			3847: out = 16'(307);
			3848: out = 16'(-1035);
			3849: out = 16'(68);
			3850: out = 16'(-24);
			3851: out = 16'(-244);
			3852: out = 16'(-284);
			3853: out = 16'(514);
			3854: out = 16'(-377);
			3855: out = 16'(-100);
			3856: out = 16'(-313);
			3857: out = 16'(-102);
			3858: out = 16'(940);
			3859: out = 16'(50);
			3860: out = 16'(-25);
			3861: out = 16'(129);
			3862: out = 16'(61);
			3863: out = 16'(-500);
			3864: out = 16'(134);
			3865: out = 16'(-4);
			3866: out = 16'(-442);
			3867: out = 16'(-1409);
			3868: out = 16'(-2153);
			3869: out = 16'(523);
			3870: out = 16'(-200);
			3871: out = 16'(-462);
			3872: out = 16'(339);
			3873: out = 16'(-78);
			3874: out = 16'(121);
			3875: out = 16'(373);
			3876: out = 16'(-66);
			3877: out = 16'(20);
			3878: out = 16'(140);
			3879: out = 16'(-698);
			3880: out = 16'(263);
			3881: out = 16'(-509);
			3882: out = 16'(-487);
			3883: out = 16'(930);
			3884: out = 16'(242);
			3885: out = 16'(-589);
			3886: out = 16'(316);
			3887: out = 16'(90);
			3888: out = 16'(-315);
			3889: out = 16'(64);
			3890: out = 16'(13);
			3891: out = 16'(-531);
			3892: out = 16'(152);
			3893: out = 16'(-108);
			3894: out = 16'(-246);
			3895: out = 16'(1198);
			3896: out = 16'(-67);
			3897: out = 16'(45);
			3898: out = 16'(1141);
			3899: out = 16'(96);
			3900: out = 16'(-420);
			3901: out = 16'(-81);
			3902: out = 16'(168);
			3903: out = 16'(-57);
			3904: out = 16'(-873);
			3905: out = 16'(-586);
			3906: out = 16'(671);
			3907: out = 16'(-368);
			3908: out = 16'(-484);
			3909: out = 16'(259);
			3910: out = 16'(408);
			3911: out = 16'(314);
			3912: out = 16'(81);
			3913: out = 16'(-60);
			3914: out = 16'(-323);
			3915: out = 16'(835);
			3916: out = 16'(-1509);
			3917: out = 16'(-204);
			3918: out = 16'(36);
			3919: out = 16'(-977);
			3920: out = 16'(248);
			3921: out = 16'(-140);
			3922: out = 16'(-30);
			3923: out = 16'(-104);
			3924: out = 16'(492);
			3925: out = 16'(14);
			3926: out = 16'(1044);
			3927: out = 16'(-152);
			3928: out = 16'(336);
			3929: out = 16'(260);
			3930: out = 16'(-1583);
			3931: out = 16'(839);
			3932: out = 16'(-949);
			3933: out = 16'(-20);
			3934: out = 16'(177);
			3935: out = 16'(301);
			3936: out = 16'(-461);
			3937: out = 16'(707);
			3938: out = 16'(-387);
			3939: out = 16'(711);
			3940: out = 16'(559);
			3941: out = 16'(31);
			3942: out = 16'(-97);
			3943: out = 16'(-409);
			3944: out = 16'(-255);
			3945: out = 16'(141);
			3946: out = 16'(-134);
			3947: out = 16'(73);
			3948: out = 16'(214);
			3949: out = 16'(-876);
			3950: out = 16'(194);
			3951: out = 16'(-230);
			3952: out = 16'(-129);
			3953: out = 16'(70);
			3954: out = 16'(35);
			3955: out = 16'(535);
			3956: out = 16'(80);
			3957: out = 16'(-1065);
			3958: out = 16'(103);
			3959: out = 16'(185);
			3960: out = 16'(-89);
			3961: out = 16'(1304);
			3962: out = 16'(178);
			3963: out = 16'(328);
			3964: out = 16'(-44);
			3965: out = 16'(-63);
			3966: out = 16'(402);
			3967: out = 16'(62);
			3968: out = 16'(-41);
			3969: out = 16'(-129);
			3970: out = 16'(45);
			3971: out = 16'(103);
			3972: out = 16'(946);
			3973: out = 16'(-1369);
			3974: out = 16'(-397);
			3975: out = 16'(1080);
			3976: out = 16'(-165);
			3977: out = 16'(232);
			3978: out = 16'(829);
			3979: out = 16'(69);
			3980: out = 16'(312);
			3981: out = 16'(438);
			3982: out = 16'(-63);
			3983: out = 16'(284);
			3984: out = 16'(-9);
			3985: out = 16'(-1362);
			3986: out = 16'(243);
			3987: out = 16'(-357);
			3988: out = 16'(-117);
			3989: out = 16'(900);
			3990: out = 16'(15);
			3991: out = 16'(232);
			3992: out = 16'(574);
			3993: out = 16'(374);
			3994: out = 16'(865);
			3995: out = 16'(32);
			3996: out = 16'(-258);
			3997: out = 16'(224);
			3998: out = 16'(-696);
			3999: out = 16'(-52);
			4000: out = 16'(-104);
			4001: out = 16'(270);
			4002: out = 16'(-818);
			4003: out = 16'(499);
			4004: out = 16'(166);
			4005: out = 16'(-667);
			4006: out = 16'(-54);
			4007: out = 16'(-824);
			4008: out = 16'(-265);
			4009: out = 16'(4);
			4010: out = 16'(-95);
			4011: out = 16'(-281);
			4012: out = 16'(637);
			4013: out = 16'(-1164);
			4014: out = 16'(-1425);
			4015: out = 16'(-31);
			4016: out = 16'(190);
			4017: out = 16'(-20);
			4018: out = 16'(755);
			4019: out = 16'(-452);
			4020: out = 16'(-723);
			4021: out = 16'(-142);
			4022: out = 16'(-873);
			4023: out = 16'(436);
			4024: out = 16'(163);
			4025: out = 16'(-97);
			4026: out = 16'(561);
			4027: out = 16'(65);
			4028: out = 16'(-73);
			4029: out = 16'(-186);
			4030: out = 16'(371);
			4031: out = 16'(-263);
			4032: out = 16'(-8);
			4033: out = 16'(34);
			4034: out = 16'(-57);
			4035: out = 16'(749);
			4036: out = 16'(133);
			4037: out = 16'(-442);
			4038: out = 16'(201);
			4039: out = 16'(-157);
			4040: out = 16'(880);
			4041: out = 16'(333);
			4042: out = 16'(-61);
			4043: out = 16'(-15);
			4044: out = 16'(258);
			4045: out = 16'(461);
			4046: out = 16'(139);
			4047: out = 16'(183);
			4048: out = 16'(-628);
			4049: out = 16'(-558);
			4050: out = 16'(-332);
			4051: out = 16'(-57);
			4052: out = 16'(-151);
			4053: out = 16'(91);
			4054: out = 16'(258);
			4055: out = 16'(-240);
			4056: out = 16'(-1051);
			4057: out = 16'(-655);
			4058: out = 16'(630);
			4059: out = 16'(0);
			4060: out = 16'(141);
			4061: out = 16'(-269);
			4062: out = 16'(-28);
			4063: out = 16'(-304);
			4064: out = 16'(-325);
			4065: out = 16'(407);
			4066: out = 16'(-973);
			4067: out = 16'(-170);
			4068: out = 16'(352);
			4069: out = 16'(575);
			4070: out = 16'(468);
			4071: out = 16'(99);
			4072: out = 16'(-44);
			4073: out = 16'(-9);
			4074: out = 16'(727);
			4075: out = 16'(-555);
			4076: out = 16'(112);
			4077: out = 16'(670);
			4078: out = 16'(-4);
			4079: out = 16'(85);
			4080: out = 16'(532);
			4081: out = 16'(92);
			4082: out = 16'(-27);
			4083: out = 16'(-35);
			4084: out = 16'(1);
			4085: out = 16'(-206);
			4086: out = 16'(-974);
			4087: out = 16'(-69);
			4088: out = 16'(93);
			4089: out = 16'(189);
			4090: out = 16'(-78);
			4091: out = 16'(218);
			4092: out = 16'(-603);
			4093: out = 16'(-157);
			4094: out = 16'(88);
			4095: out = 16'(258);
			4096: out = 16'(84);
			4097: out = 16'(407);
			4098: out = 16'(-789);
			4099: out = 16'(-472);
			4100: out = 16'(246);
			4101: out = 16'(-109);
			4102: out = 16'(99);
			4103: out = 16'(-115);
			4104: out = 16'(76);
			4105: out = 16'(-504);
			4106: out = 16'(595);
			4107: out = 16'(6);
			4108: out = 16'(294);
			4109: out = 16'(-34);
			4110: out = 16'(-693);
			4111: out = 16'(-159);
			4112: out = 16'(323);
			4113: out = 16'(-155);
			4114: out = 16'(-211);
			4115: out = 16'(-470);
			4116: out = 16'(-438);
			4117: out = 16'(398);
			4118: out = 16'(-179);
			4119: out = 16'(-149);
			4120: out = 16'(140);
			4121: out = 16'(34);
			4122: out = 16'(-138);
			4123: out = 16'(55);
			4124: out = 16'(-101);
			4125: out = 16'(17);
			4126: out = 16'(642);
			4127: out = 16'(-43);
			4128: out = 16'(-217);
			4129: out = 16'(1010);
			4130: out = 16'(-701);
			4131: out = 16'(58);
			4132: out = 16'(207);
			4133: out = 16'(-254);
			4134: out = 16'(425);
			4135: out = 16'(-86);
			4136: out = 16'(303);
			4137: out = 16'(-98);
			4138: out = 16'(106);
			4139: out = 16'(-314);
			4140: out = 16'(139);
			4141: out = 16'(-523);
			4142: out = 16'(41);
			4143: out = 16'(744);
			4144: out = 16'(-404);
			4145: out = 16'(-717);
			4146: out = 16'(154);
			4147: out = 16'(25);
			4148: out = 16'(381);
			4149: out = 16'(-546);
			4150: out = 16'(15);
			4151: out = 16'(49);
			4152: out = 16'(-277);
			4153: out = 16'(-138);
			4154: out = 16'(-230);
			4155: out = 16'(59);
			4156: out = 16'(-992);
			4157: out = 16'(130);
			4158: out = 16'(-89);
			4159: out = 16'(-77);
			4160: out = 16'(-366);
			4161: out = 16'(-353);
			4162: out = 16'(-43);
			4163: out = 16'(-157);
			4164: out = 16'(-46);
			4165: out = 16'(-128);
			4166: out = 16'(268);
			4167: out = 16'(-134);
			4168: out = 16'(-792);
			4169: out = 16'(618);
			4170: out = 16'(-219);
			4171: out = 16'(-87);
			4172: out = 16'(661);
			4173: out = 16'(-689);
			4174: out = 16'(27);
			4175: out = 16'(344);
			4176: out = 16'(-1039);
			4177: out = 16'(226);
			4178: out = 16'(-20);
			4179: out = 16'(111);
			4180: out = 16'(90);
			4181: out = 16'(-709);
			4182: out = 16'(89);
			4183: out = 16'(209);
			4184: out = 16'(-424);
			4185: out = 16'(347);
			4186: out = 16'(-434);
			4187: out = 16'(-147);
			4188: out = 16'(420);
			4189: out = 16'(-69);
			4190: out = 16'(-10);
			4191: out = 16'(848);
			4192: out = 16'(-375);
			4193: out = 16'(-142);
			4194: out = 16'(157);
			4195: out = 16'(-38);
			4196: out = 16'(-441);
			4197: out = 16'(-91);
			4198: out = 16'(-74);
			4199: out = 16'(140);
			4200: out = 16'(-147);
			4201: out = 16'(294);
			4202: out = 16'(284);
			4203: out = 16'(-82);
			4204: out = 16'(-17);
			4205: out = 16'(541);
			4206: out = 16'(-343);
			4207: out = 16'(244);
			4208: out = 16'(-108);
			4209: out = 16'(-516);
			4210: out = 16'(178);
			4211: out = 16'(-295);
			4212: out = 16'(239);
			4213: out = 16'(4);
			4214: out = 16'(-295);
			4215: out = 16'(-607);
			4216: out = 16'(182);
			4217: out = 16'(29);
			4218: out = 16'(-40);
			4219: out = 16'(-196);
			4220: out = 16'(-28);
			4221: out = 16'(-50);
			4222: out = 16'(490);
			4223: out = 16'(-422);
			4224: out = 16'(-112);
			4225: out = 16'(-130);
			4226: out = 16'(-44);
			4227: out = 16'(61);
			4228: out = 16'(230);
			4229: out = 16'(-132);
			4230: out = 16'(117);
			4231: out = 16'(-104);
			4232: out = 16'(-50);
			4233: out = 16'(51);
			4234: out = 16'(-104);
			4235: out = 16'(-44);
			4236: out = 16'(36);
			4237: out = 16'(-120);
			4238: out = 16'(-139);
			4239: out = 16'(61);
			4240: out = 16'(-94);
			4241: out = 16'(405);
			4242: out = 16'(356);
			4243: out = 16'(-552);
			4244: out = 16'(361);
			4245: out = 16'(839);
			4246: out = 16'(-865);
			4247: out = 16'(-139);
			4248: out = 16'(85);
			4249: out = 16'(-17);
			4250: out = 16'(-49);
			4251: out = 16'(-88);
			4252: out = 16'(210);
			4253: out = 16'(118);
			4254: out = 16'(506);
			4255: out = 16'(205);
			4256: out = 16'(238);
			4257: out = 16'(55);
			4258: out = 16'(154);
			4259: out = 16'(146);
			4260: out = 16'(149);
			4261: out = 16'(-679);
			4262: out = 16'(-609);
			4263: out = 16'(55);
			4264: out = 16'(-261);
			4265: out = 16'(281);
			4266: out = 16'(-278);
			4267: out = 16'(290);
			4268: out = 16'(-674);
			4269: out = 16'(78);
			4270: out = 16'(-355);
			4271: out = 16'(591);
			4272: out = 16'(-160);
			4273: out = 16'(594);
			4274: out = 16'(-818);
			4275: out = 16'(-68);
			4276: out = 16'(-263);
			4277: out = 16'(-491);
			4278: out = 16'(-332);
			4279: out = 16'(183);
			4280: out = 16'(48);
			4281: out = 16'(-92);
			4282: out = 16'(284);
			4283: out = 16'(-868);
			4284: out = 16'(-248);
			4285: out = 16'(-269);
			4286: out = 16'(134);
			4287: out = 16'(32);
			4288: out = 16'(-15);
			4289: out = 16'(-224);
			4290: out = 16'(86);
			4291: out = 16'(-291);
			4292: out = 16'(439);
			4293: out = 16'(-447);
			4294: out = 16'(679);
			4295: out = 16'(35);
			4296: out = 16'(-226);
			4297: out = 16'(315);
			4298: out = 16'(-131);
			4299: out = 16'(-1113);
			4300: out = 16'(-19);
			4301: out = 16'(54);
			4302: out = 16'(138);
			4303: out = 16'(-647);
			4304: out = 16'(-137);
			4305: out = 16'(400);
			4306: out = 16'(619);
			4307: out = 16'(233);
			4308: out = 16'(168);
			4309: out = 16'(10);
			4310: out = 16'(-337);
			4311: out = 16'(108);
			4312: out = 16'(-599);
			4313: out = 16'(-1024);
			4314: out = 16'(-123);
			4315: out = 16'(31);
			4316: out = 16'(-323);
			4317: out = 16'(226);
			4318: out = 16'(-223);
			4319: out = 16'(455);
			4320: out = 16'(-125);
			4321: out = 16'(-302);
			4322: out = 16'(-425);
			4323: out = 16'(-9);
			4324: out = 16'(137);
			4325: out = 16'(-8);
			4326: out = 16'(-521);
			4327: out = 16'(-789);
			4328: out = 16'(83);
			4329: out = 16'(-861);
			4330: out = 16'(124);
			4331: out = 16'(293);
			4332: out = 16'(-83);
			4333: out = 16'(230);
			4334: out = 16'(96);
			4335: out = 16'(-593);
			4336: out = 16'(258);
			4337: out = 16'(114);
			4338: out = 16'(362);
			4339: out = 16'(-333);
			4340: out = 16'(-121);
			4341: out = 16'(364);
			4342: out = 16'(530);
			4343: out = 16'(63);
			4344: out = 16'(52);
			4345: out = 16'(125);
			4346: out = 16'(-160);
			4347: out = 16'(294);
			4348: out = 16'(-147);
			4349: out = 16'(65);
			4350: out = 16'(54);
			4351: out = 16'(-106);
			4352: out = 16'(-26);
			4353: out = 16'(351);
			4354: out = 16'(-640);
			4355: out = 16'(-292);
			4356: out = 16'(-318);
			4357: out = 16'(-171);
			4358: out = 16'(364);
			4359: out = 16'(-89);
			4360: out = 16'(-418);
			4361: out = 16'(-12);
			4362: out = 16'(-295);
			4363: out = 16'(-422);
			4364: out = 16'(-28);
			4365: out = 16'(-90);
			4366: out = 16'(297);
			4367: out = 16'(117);
			4368: out = 16'(-103);
			4369: out = 16'(-388);
			4370: out = 16'(-137);
			4371: out = 16'(-126);
			4372: out = 16'(25);
			4373: out = 16'(-82);
			4374: out = 16'(-85);
			4375: out = 16'(480);
			4376: out = 16'(-100);
			4377: out = 16'(-315);
			4378: out = 16'(475);
			4379: out = 16'(-42);
			4380: out = 16'(546);
			4381: out = 16'(-114);
			4382: out = 16'(22);
			4383: out = 16'(-2);
			4384: out = 16'(-199);
			4385: out = 16'(429);
			4386: out = 16'(67);
			4387: out = 16'(130);
			4388: out = 16'(204);
			4389: out = 16'(29);
			4390: out = 16'(-80);
			4391: out = 16'(74);
			4392: out = 16'(101);
			4393: out = 16'(55);
			4394: out = 16'(-420);
			4395: out = 16'(431);
			4396: out = 16'(19);
			4397: out = 16'(-3);
			4398: out = 16'(-99);
			4399: out = 16'(68);
			4400: out = 16'(45);
			4401: out = 16'(-40);
			4402: out = 16'(251);
			4403: out = 16'(5);
			4404: out = 16'(200);
			4405: out = 16'(-467);
			4406: out = 16'(-884);
			4407: out = 16'(95);
			4408: out = 16'(-395);
			4409: out = 16'(16);
			4410: out = 16'(-47);
			4411: out = 16'(-543);
			4412: out = 16'(45);
			4413: out = 16'(-307);
			4414: out = 16'(-245);
			4415: out = 16'(135);
			4416: out = 16'(-73);
			4417: out = 16'(-392);
			4418: out = 16'(215);
			4419: out = 16'(-100);
			4420: out = 16'(27);
			4421: out = 16'(457);
			4422: out = 16'(52);
			4423: out = 16'(40);
			4424: out = 16'(234);
			4425: out = 16'(-133);
			4426: out = 16'(185);
			4427: out = 16'(192);
			4428: out = 16'(-545);
			4429: out = 16'(35);
			4430: out = 16'(38);
			4431: out = 16'(321);
			4432: out = 16'(26);
			4433: out = 16'(-63);
			4434: out = 16'(-44);
			4435: out = 16'(54);
			4436: out = 16'(-270);
			4437: out = 16'(560);
			4438: out = 16'(-271);
			4439: out = 16'(29);
			4440: out = 16'(-30);
			4441: out = 16'(265);
			4442: out = 16'(-146);
			4443: out = 16'(-160);
			4444: out = 16'(-230);
			4445: out = 16'(-237);
			4446: out = 16'(-237);
			4447: out = 16'(-470);
			4448: out = 16'(-86);
			4449: out = 16'(-93);
			4450: out = 16'(212);
			4451: out = 16'(-319);
			4452: out = 16'(257);
			4453: out = 16'(266);
			4454: out = 16'(-478);
			4455: out = 16'(-60);
			4456: out = 16'(-14);
			4457: out = 16'(-444);
			4458: out = 16'(-55);
			4459: out = 16'(203);
			4460: out = 16'(-152);
			4461: out = 16'(-444);
			4462: out = 16'(-353);
			4463: out = 16'(118);
			4464: out = 16'(310);
			4465: out = 16'(100);
			4466: out = 16'(-48);
			4467: out = 16'(189);
			4468: out = 16'(-352);
			4469: out = 16'(427);
			4470: out = 16'(-274);
			4471: out = 16'(-53);
			4472: out = 16'(-100);
			4473: out = 16'(-431);
			4474: out = 16'(150);
			4475: out = 16'(-120);
			4476: out = 16'(-98);
			4477: out = 16'(172);
			4478: out = 16'(-171);
			4479: out = 16'(-425);
			4480: out = 16'(-173);
			4481: out = 16'(-251);
			4482: out = 16'(587);
			4483: out = 16'(-84);
			4484: out = 16'(-9);
			4485: out = 16'(162);
			4486: out = 16'(-9);
			4487: out = 16'(-269);
			4488: out = 16'(-603);
			4489: out = 16'(144);
			4490: out = 16'(5);
			4491: out = 16'(-85);
			4492: out = 16'(253);
			4493: out = 16'(82);
			4494: out = 16'(-430);
			4495: out = 16'(-151);
			4496: out = 16'(200);
			4497: out = 16'(183);
			4498: out = 16'(-393);
			4499: out = 16'(-322);
			4500: out = 16'(-236);
			4501: out = 16'(234);
			4502: out = 16'(-557);
			4503: out = 16'(-64);
			4504: out = 16'(-236);
			4505: out = 16'(-28);
			4506: out = 16'(-3);
			4507: out = 16'(-117);
			4508: out = 16'(179);
			4509: out = 16'(-14);
			4510: out = 16'(-266);
			4511: out = 16'(-55);
			4512: out = 16'(197);
			4513: out = 16'(-137);
			4514: out = 16'(-292);
			4515: out = 16'(351);
			4516: out = 16'(20);
			4517: out = 16'(-114);
			4518: out = 16'(367);
			4519: out = 16'(102);
			4520: out = 16'(-49);
			4521: out = 16'(87);
			4522: out = 16'(-57);
			4523: out = 16'(-72);
			4524: out = 16'(39);
			4525: out = 16'(95);
			4526: out = 16'(54);
			4527: out = 16'(-1);
			4528: out = 16'(-126);
			4529: out = 16'(217);
			4530: out = 16'(-4);
			4531: out = 16'(-327);
			4532: out = 16'(-36);
			4533: out = 16'(-7);
			4534: out = 16'(116);
			4535: out = 16'(432);
			4536: out = 16'(-341);
			4537: out = 16'(-84);
			4538: out = 16'(38);
			4539: out = 16'(-544);
			4540: out = 16'(180);
			4541: out = 16'(361);
			4542: out = 16'(-214);
			4543: out = 16'(26);
			4544: out = 16'(485);
			4545: out = 16'(-549);
			4546: out = 16'(-41);
			4547: out = 16'(204);
			4548: out = 16'(-318);
			4549: out = 16'(521);
			4550: out = 16'(27);
			4551: out = 16'(-232);
			4552: out = 16'(179);
			4553: out = 16'(-402);
			4554: out = 16'(-10);
			4555: out = 16'(198);
			4556: out = 16'(-68);
			4557: out = 16'(-145);
			4558: out = 16'(263);
			4559: out = 16'(166);
			4560: out = 16'(1);
			4561: out = 16'(-25);
			4562: out = 16'(84);
			4563: out = 16'(-362);
			4564: out = 16'(-298);
			4565: out = 16'(152);
			4566: out = 16'(280);
			4567: out = 16'(42);
			4568: out = 16'(175);
			4569: out = 16'(503);
			4570: out = 16'(565);
			4571: out = 16'(-223);
			4572: out = 16'(-204);
			4573: out = 16'(-321);
			4574: out = 16'(328);
			4575: out = 16'(-116);
			4576: out = 16'(364);
			4577: out = 16'(72);
			4578: out = 16'(391);
			4579: out = 16'(-464);
			4580: out = 16'(-30);
			4581: out = 16'(142);
			4582: out = 16'(-157);
			4583: out = 16'(330);
			4584: out = 16'(410);
			4585: out = 16'(61);
			4586: out = 16'(251);
			4587: out = 16'(-243);
			4588: out = 16'(-412);
			4589: out = 16'(-275);
			4590: out = 16'(-238);
			4591: out = 16'(471);
			4592: out = 16'(99);
			4593: out = 16'(435);
			4594: out = 16'(84);
			4595: out = 16'(-171);
			4596: out = 16'(240);
			4597: out = 16'(528);
			4598: out = 16'(-321);
			4599: out = 16'(25);
			4600: out = 16'(-292);
			4601: out = 16'(-551);
			4602: out = 16'(94);
			4603: out = 16'(240);
			4604: out = 16'(-118);
			4605: out = 16'(-830);
			4606: out = 16'(-75);
			4607: out = 16'(2);
			4608: out = 16'(185);
			4609: out = 16'(-187);
			4610: out = 16'(89);
			4611: out = 16'(-3);
			4612: out = 16'(-31);
			4613: out = 16'(-253);
			4614: out = 16'(-248);
			4615: out = 16'(105);
			4616: out = 16'(-633);
			4617: out = 16'(22);
			4618: out = 16'(-36);
			4619: out = 16'(-293);
			4620: out = 16'(-100);
			4621: out = 16'(-120);
			4622: out = 16'(37);
			4623: out = 16'(-44);
			4624: out = 16'(-49);
			4625: out = 16'(62);
			4626: out = 16'(-130);
			4627: out = 16'(-272);
			4628: out = 16'(-354);
			4629: out = 16'(-125);
			4630: out = 16'(-26);
			4631: out = 16'(107);
			4632: out = 16'(169);
			4633: out = 16'(121);
			4634: out = 16'(463);
			4635: out = 16'(-10);
			4636: out = 16'(-224);
			4637: out = 16'(-4);
			4638: out = 16'(-372);
			4639: out = 16'(-341);
			4640: out = 16'(316);
			4641: out = 16'(-70);
			4642: out = 16'(-22);
			4643: out = 16'(54);
			4644: out = 16'(-16);
			4645: out = 16'(-62);
			4646: out = 16'(-256);
			4647: out = 16'(110);
			4648: out = 16'(113);
			4649: out = 16'(-233);
			4650: out = 16'(99);
			4651: out = 16'(24);
			4652: out = 16'(-120);
			4653: out = 16'(-130);
			4654: out = 16'(74);
			4655: out = 16'(-479);
			4656: out = 16'(-429);
			4657: out = 16'(32);
			4658: out = 16'(-229);
			4659: out = 16'(59);
			4660: out = 16'(-99);
			4661: out = 16'(84);
			4662: out = 16'(-210);
			4663: out = 16'(-159);
			4664: out = 16'(-241);
			4665: out = 16'(-472);
			4666: out = 16'(68);
			4667: out = 16'(134);
			4668: out = 16'(-243);
			4669: out = 16'(82);
			4670: out = 16'(-64);
			4671: out = 16'(-128);
			4672: out = 16'(9);
			4673: out = 16'(-684);
			4674: out = 16'(121);
			4675: out = 16'(-70);
			4676: out = 16'(70);
			4677: out = 16'(287);
			4678: out = 16'(19);
			4679: out = 16'(-228);
			4680: out = 16'(48);
			4681: out = 16'(-96);
			4682: out = 16'(-644);
			4683: out = 16'(677);
			4684: out = 16'(-405);
			4685: out = 16'(178);
			4686: out = 16'(524);
			4687: out = 16'(-37);
			4688: out = 16'(-31);
			4689: out = 16'(-120);
			4690: out = 16'(-437);
			4691: out = 16'(93);
			4692: out = 16'(30);
			4693: out = 16'(43);
			4694: out = 16'(53);
			4695: out = 16'(294);
			4696: out = 16'(-55);
			4697: out = 16'(-148);
			4698: out = 16'(166);
			4699: out = 16'(-413);
			4700: out = 16'(575);
			4701: out = 16'(-20);
			4702: out = 16'(75);
			4703: out = 16'(175);
			4704: out = 16'(-143);
			4705: out = 16'(-424);
			4706: out = 16'(6);
			4707: out = 16'(-423);
			4708: out = 16'(40);
			4709: out = 16'(50);
			4710: out = 16'(0);
			4711: out = 16'(-398);
			4712: out = 16'(236);
			4713: out = 16'(-256);
			4714: out = 16'(-103);
			4715: out = 16'(53);
			4716: out = 16'(-101);
			4717: out = 16'(63);
			4718: out = 16'(-75);
			4719: out = 16'(-46);
			4720: out = 16'(271);
			4721: out = 16'(-118);
			4722: out = 16'(-39);
			4723: out = 16'(169);
			4724: out = 16'(-193);
			4725: out = 16'(144);
			4726: out = 16'(230);
			4727: out = 16'(19);
			4728: out = 16'(-65);
			4729: out = 16'(59);
			4730: out = 16'(-207);
			4731: out = 16'(390);
			4732: out = 16'(494);
			4733: out = 16'(-22);
			4734: out = 16'(-13);
			4735: out = 16'(-101);
			4736: out = 16'(92);
			4737: out = 16'(-113);
			4738: out = 16'(-61);
			4739: out = 16'(-55);
			4740: out = 16'(146);
			4741: out = 16'(-195);
			4742: out = 16'(150);
			4743: out = 16'(250);
			4744: out = 16'(-359);
			4745: out = 16'(36);
			4746: out = 16'(-435);
			4747: out = 16'(-242);
			4748: out = 16'(-13);
			4749: out = 16'(50);
			4750: out = 16'(-42);
			4751: out = 16'(145);
			4752: out = 16'(-238);
			4753: out = 16'(-366);
			4754: out = 16'(-519);
			4755: out = 16'(50);
			4756: out = 16'(17);
			4757: out = 16'(-261);
			4758: out = 16'(-4);
			4759: out = 16'(-313);
			4760: out = 16'(-159);
			4761: out = 16'(67);
			4762: out = 16'(60);
			4763: out = 16'(-8);
			4764: out = 16'(-79);
			4765: out = 16'(184);
			4766: out = 16'(317);
			4767: out = 16'(90);
			4768: out = 16'(6);
			4769: out = 16'(-20);
			4770: out = 16'(25);
			4771: out = 16'(-176);
			4772: out = 16'(-89);
			4773: out = 16'(165);
			4774: out = 16'(69);
			4775: out = 16'(-43);
			4776: out = 16'(238);
			4777: out = 16'(-74);
			4778: out = 16'(21);
			4779: out = 16'(3);
			4780: out = 16'(159);
			4781: out = 16'(-341);
			4782: out = 16'(76);
			4783: out = 16'(-281);
			4784: out = 16'(65);
			4785: out = 16'(-36);
			4786: out = 16'(143);
			4787: out = 16'(-105);
			4788: out = 16'(49);
			4789: out = 16'(201);
			4790: out = 16'(66);
			4791: out = 16'(116);
			4792: out = 16'(-33);
			4793: out = 16'(-169);
			4794: out = 16'(-219);
			4795: out = 16'(-504);
			4796: out = 16'(-189);
			4797: out = 16'(-430);
			4798: out = 16'(-55);
			4799: out = 16'(-41);
			4800: out = 16'(-140);
			4801: out = 16'(-329);
			4802: out = 16'(-242);
			4803: out = 16'(-384);
			4804: out = 16'(35);
			4805: out = 16'(11);
			4806: out = 16'(67);
			4807: out = 16'(-101);
			4808: out = 16'(-137);
			4809: out = 16'(-56);
			4810: out = 16'(-186);
			4811: out = 16'(-15);
			4812: out = 16'(-338);
			4813: out = 16'(-52);
			4814: out = 16'(-6);
			4815: out = 16'(218);
			4816: out = 16'(-88);
			4817: out = 16'(-28);
			4818: out = 16'(-472);
			4819: out = 16'(76);
			4820: out = 16'(200);
			4821: out = 16'(70);
			4822: out = 16'(261);
			4823: out = 16'(41);
			4824: out = 16'(28);
			4825: out = 16'(-75);
			4826: out = 16'(58);
			4827: out = 16'(-292);
			4828: out = 16'(452);
			4829: out = 16'(-37);
			4830: out = 16'(-410);
			default: out = 0;
		endcase
	end
endmodule
