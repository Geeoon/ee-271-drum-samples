module crash1_lookup(index, out);
	input logic unsigned [13:0] index;
	output logic signed [15:0] out;
	always_comb begin
		case(index)
			0: out = 16'(0);
			1: out = 16'(2);
			2: out = 16'(51);
			3: out = 16'(221);
			4: out = 16'(7393);
			5: out = 16'(-7947);
			6: out = 16'(-17672);
			7: out = 16'(1158);
			8: out = 16'(-3561);
			9: out = 16'(4337);
			10: out = 16'(5764);
			11: out = 16'(-6430);
			12: out = 16'(1002);
			13: out = 16'(-17884);
			14: out = 16'(4223);
			15: out = 16'(1278);
			16: out = 16'(-3472);
			17: out = 16'(-15365);
			18: out = 16'(7238);
			19: out = 16'(4586);
			20: out = 16'(8160);
			21: out = 16'(2571);
			22: out = 16'(-4257);
			23: out = 16'(1746);
			24: out = 16'(-2157);
			25: out = 16'(-1052);
			26: out = 16'(1123);
			27: out = 16'(5095);
			28: out = 16'(-1967);
			29: out = 16'(-7995);
			30: out = 16'(-19886);
			31: out = 16'(-774);
			32: out = 16'(1002);
			33: out = 16'(328);
			34: out = 16'(-2747);
			35: out = 16'(-8747);
			36: out = 16'(5024);
			37: out = 16'(-2132);
			38: out = 16'(-93);
			39: out = 16'(-4889);
			40: out = 16'(2324);
			41: out = 16'(3380);
			42: out = 16'(-6473);
			43: out = 16'(-15);
			44: out = 16'(10069);
			45: out = 16'(-4101);
			46: out = 16'(5284);
			47: out = 16'(-18236);
			48: out = 16'(4678);
			49: out = 16'(9490);
			50: out = 16'(1824);
			51: out = 16'(-19023);
			52: out = 16'(-7128);
			53: out = 16'(-3696);
			54: out = 16'(3813);
			55: out = 16'(12465);
			56: out = 16'(277);
			57: out = 16'(-11942);
			58: out = 16'(-6189);
			59: out = 16'(952);
			60: out = 16'(11610);
			61: out = 16'(-1676);
			62: out = 16'(-5131);
			63: out = 16'(-18131);
			64: out = 16'(-1421);
			65: out = 16'(-9221);
			66: out = 16'(-1311);
			67: out = 16'(1662);
			68: out = 16'(10664);
			69: out = 16'(17930);
			70: out = 16'(14586);
			71: out = 16'(19457);
			72: out = 16'(7105);
			73: out = 16'(-5882);
			74: out = 16'(-6544);
			75: out = 16'(-10904);
			76: out = 16'(-5890);
			77: out = 16'(7079);
			78: out = 16'(-3427);
			79: out = 16'(7874);
			80: out = 16'(26215);
			81: out = 16'(23310);
			82: out = 16'(13998);
			83: out = 16'(-8432);
			84: out = 16'(-12070);
			85: out = 16'(-11037);
			86: out = 16'(-26753);
			87: out = 16'(-32767);
			88: out = 16'(-18141);
			89: out = 16'(-21127);
			90: out = 16'(3286);
			91: out = 16'(-3470);
			92: out = 16'(799);
			93: out = 16'(25093);
			94: out = 16'(11789);
			95: out = 16'(13533);
			96: out = 16'(14706);
			97: out = 16'(10960);
			98: out = 16'(14511);
			99: out = 16'(8254);
			100: out = 16'(12531);
			101: out = 16'(11216);
			102: out = 16'(15009);
			103: out = 16'(3977);
			104: out = 16'(-14221);
			105: out = 16'(-22545);
			106: out = 16'(-19618);
			107: out = 16'(-21414);
			108: out = 16'(-27693);
			109: out = 16'(-24426);
			110: out = 16'(-11647);
			111: out = 16'(-20014);
			112: out = 16'(-9526);
			113: out = 16'(-14599);
			114: out = 16'(3090);
			115: out = 16'(6749);
			116: out = 16'(24628);
			117: out = 16'(24224);
			118: out = 16'(17326);
			119: out = 16'(-221);
			120: out = 16'(-2707);
			121: out = 16'(3994);
			122: out = 16'(14931);
			123: out = 16'(-5093);
			124: out = 16'(12536);
			125: out = 16'(137);
			126: out = 16'(2192);
			127: out = 16'(13298);
			128: out = 16'(-15771);
			129: out = 16'(12724);
			130: out = 16'(1337);
			131: out = 16'(-1993);
			132: out = 16'(-1422);
			133: out = 16'(-6330);
			134: out = 16'(-1587);
			135: out = 16'(-4005);
			136: out = 16'(-13910);
			137: out = 16'(-6615);
			138: out = 16'(4931);
			139: out = 16'(10872);
			140: out = 16'(-15854);
			141: out = 16'(2671);
			142: out = 16'(-148);
			143: out = 16'(5009);
			144: out = 16'(-5199);
			145: out = 16'(673);
			146: out = 16'(5693);
			147: out = 16'(-7553);
			148: out = 16'(2574);
			149: out = 16'(-11750);
			150: out = 16'(5113);
			151: out = 16'(12496);
			152: out = 16'(-16871);
			153: out = 16'(271);
			154: out = 16'(-3622);
			155: out = 16'(77);
			156: out = 16'(-2983);
			157: out = 16'(-26303);
			158: out = 16'(-9408);
			159: out = 16'(6907);
			160: out = 16'(12018);
			161: out = 16'(22072);
			162: out = 16'(4045);
			163: out = 16'(13512);
			164: out = 16'(13765);
			165: out = 16'(-3408);
			166: out = 16'(18258);
			167: out = 16'(-13912);
			168: out = 16'(-2011);
			169: out = 16'(-7978);
			170: out = 16'(-13154);
			171: out = 16'(-5501);
			172: out = 16'(-11745);
			173: out = 16'(-5953);
			174: out = 16'(422);
			175: out = 16'(7514);
			176: out = 16'(6878);
			177: out = 16'(21627);
			178: out = 16'(14613);
			179: out = 16'(13065);
			180: out = 16'(6047);
			181: out = 16'(2245);
			182: out = 16'(19977);
			183: out = 16'(-11133);
			184: out = 16'(-4249);
			185: out = 16'(-3572);
			186: out = 16'(-25717);
			187: out = 16'(-2156);
			188: out = 16'(-27933);
			189: out = 16'(-2498);
			190: out = 16'(-16482);
			191: out = 16'(9109);
			192: out = 16'(3692);
			193: out = 16'(1722);
			194: out = 16'(14163);
			195: out = 16'(6236);
			196: out = 16'(-8821);
			197: out = 16'(-1973);
			198: out = 16'(3884);
			199: out = 16'(7636);
			200: out = 16'(9802);
			201: out = 16'(4994);
			202: out = 16'(16544);
			203: out = 16'(-1286);
			204: out = 16'(4287);
			205: out = 16'(-9631);
			206: out = 16'(1387);
			207: out = 16'(-6432);
			208: out = 16'(3138);
			209: out = 16'(-3794);
			210: out = 16'(5442);
			211: out = 16'(-4987);
			212: out = 16'(2964);
			213: out = 16'(13205);
			214: out = 16'(21212);
			215: out = 16'(1927);
			216: out = 16'(-8510);
			217: out = 16'(14594);
			218: out = 16'(8113);
			219: out = 16'(-2632);
			220: out = 16'(-20192);
			221: out = 16'(-9895);
			222: out = 16'(-27961);
			223: out = 16'(-8170);
			224: out = 16'(-29960);
			225: out = 16'(-21383);
			226: out = 16'(14054);
			227: out = 16'(-17361);
			228: out = 16'(19201);
			229: out = 16'(-2415);
			230: out = 16'(28022);
			231: out = 16'(22157);
			232: out = 16'(11160);
			233: out = 16'(25390);
			234: out = 16'(566);
			235: out = 16'(-2854);
			236: out = 16'(-1266);
			237: out = 16'(-12704);
			238: out = 16'(-1768);
			239: out = 16'(-8200);
			240: out = 16'(9948);
			241: out = 16'(-2295);
			242: out = 16'(4576);
			243: out = 16'(-7556);
			244: out = 16'(369);
			245: out = 16'(-15972);
			246: out = 16'(-162);
			247: out = 16'(2925);
			248: out = 16'(-10333);
			249: out = 16'(19447);
			250: out = 16'(978);
			251: out = 16'(-5885);
			252: out = 16'(18576);
			253: out = 16'(-2129);
			254: out = 16'(25613);
			255: out = 16'(2284);
			256: out = 16'(9917);
			257: out = 16'(816);
			258: out = 16'(6528);
			259: out = 16'(-9055);
			260: out = 16'(-1910);
			261: out = 16'(-2983);
			262: out = 16'(-27792);
			263: out = 16'(-12221);
			264: out = 16'(-20419);
			265: out = 16'(2770);
			266: out = 16'(-23466);
			267: out = 16'(7132);
			268: out = 16'(-6367);
			269: out = 16'(23171);
			270: out = 16'(23630);
			271: out = 16'(8211);
			272: out = 16'(10043);
			273: out = 16'(-5970);
			274: out = 16'(-18143);
			275: out = 16'(-5625);
			276: out = 16'(17191);
			277: out = 16'(5233);
			278: out = 16'(-20997);
			279: out = 16'(5609);
			280: out = 16'(-10415);
			281: out = 16'(6630);
			282: out = 16'(11709);
			283: out = 16'(8179);
			284: out = 16'(-1174);
			285: out = 16'(-4527);
			286: out = 16'(-5854);
			287: out = 16'(-10680);
			288: out = 16'(24704);
			289: out = 16'(-9359);
			290: out = 16'(-5960);
			291: out = 16'(6126);
			292: out = 16'(13411);
			293: out = 16'(9150);
			294: out = 16'(-362);
			295: out = 16'(12437);
			296: out = 16'(-5198);
			297: out = 16'(29368);
			298: out = 16'(11433);
			299: out = 16'(13264);
			300: out = 16'(9859);
			301: out = 16'(-16045);
			302: out = 16'(-1901);
			303: out = 16'(-19354);
			304: out = 16'(24059);
			305: out = 16'(-7037);
			306: out = 16'(2463);
			307: out = 16'(13727);
			308: out = 16'(-16273);
			309: out = 16'(8613);
			310: out = 16'(-195);
			311: out = 16'(-7581);
			312: out = 16'(-2303);
			313: out = 16'(-853);
			314: out = 16'(816);
			315: out = 16'(-469);
			316: out = 16'(-7604);
			317: out = 16'(1666);
			318: out = 16'(-7854);
			319: out = 16'(-3010);
			320: out = 16'(-5735);
			321: out = 16'(19474);
			322: out = 16'(14989);
			323: out = 16'(-14437);
			324: out = 16'(-1812);
			325: out = 16'(-15772);
			326: out = 16'(-2851);
			327: out = 16'(5182);
			328: out = 16'(7556);
			329: out = 16'(-8330);
			330: out = 16'(3907);
			331: out = 16'(-8149);
			332: out = 16'(-2058);
			333: out = 16'(-8266);
			334: out = 16'(17227);
			335: out = 16'(3799);
			336: out = 16'(18826);
			337: out = 16'(6393);
			338: out = 16'(31091);
			339: out = 16'(3455);
			340: out = 16'(26760);
			341: out = 16'(7279);
			342: out = 16'(6783);
			343: out = 16'(13749);
			344: out = 16'(-11542);
			345: out = 16'(-13204);
			346: out = 16'(-1612);
			347: out = 16'(-19702);
			348: out = 16'(-15479);
			349: out = 16'(-8223);
			350: out = 16'(-5439);
			351: out = 16'(-2046);
			352: out = 16'(-12692);
			353: out = 16'(917);
			354: out = 16'(-444);
			355: out = 16'(5225);
			356: out = 16'(-8713);
			357: out = 16'(-11264);
			358: out = 16'(13522);
			359: out = 16'(2353);
			360: out = 16'(7055);
			361: out = 16'(5541);
			362: out = 16'(14327);
			363: out = 16'(-4301);
			364: out = 16'(-2273);
			365: out = 16'(-6596);
			366: out = 16'(-5132);
			367: out = 16'(-1048);
			368: out = 16'(-11244);
			369: out = 16'(14546);
			370: out = 16'(3906);
			371: out = 16'(-19413);
			372: out = 16'(-20609);
			373: out = 16'(-28061);
			374: out = 16'(14451);
			375: out = 16'(1539);
			376: out = 16'(841);
			377: out = 16'(12664);
			378: out = 16'(4469);
			379: out = 16'(6388);
			380: out = 16'(10826);
			381: out = 16'(554);
			382: out = 16'(15374);
			383: out = 16'(934);
			384: out = 16'(16537);
			385: out = 16'(17814);
			386: out = 16'(-445);
			387: out = 16'(17720);
			388: out = 16'(-3074);
			389: out = 16'(14372);
			390: out = 16'(-17036);
			391: out = 16'(-16407);
			392: out = 16'(-9386);
			393: out = 16'(-8155);
			394: out = 16'(2575);
			395: out = 16'(-29284);
			396: out = 16'(-8502);
			397: out = 16'(-26305);
			398: out = 16'(-2927);
			399: out = 16'(5757);
			400: out = 16'(5363);
			401: out = 16'(16618);
			402: out = 16'(-3316);
			403: out = 16'(12422);
			404: out = 16'(10184);
			405: out = 16'(-437);
			406: out = 16'(23168);
			407: out = 16'(-27639);
			408: out = 16'(29054);
			409: out = 16'(-24524);
			410: out = 16'(6092);
			411: out = 16'(-4616);
			412: out = 16'(-11861);
			413: out = 16'(7062);
			414: out = 16'(-1514);
			415: out = 16'(-15227);
			416: out = 16'(-22157);
			417: out = 16'(586);
			418: out = 16'(-3645);
			419: out = 16'(13052);
			420: out = 16'(13772);
			421: out = 16'(11196);
			422: out = 16'(13161);
			423: out = 16'(-742);
			424: out = 16'(9810);
			425: out = 16'(3686);
			426: out = 16'(13918);
			427: out = 16'(6942);
			428: out = 16'(-6164);
			429: out = 16'(-2202);
			430: out = 16'(4071);
			431: out = 16'(4424);
			432: out = 16'(9898);
			433: out = 16'(-9330);
			434: out = 16'(-21883);
			435: out = 16'(-11117);
			436: out = 16'(-11492);
			437: out = 16'(-1352);
			438: out = 16'(-2471);
			439: out = 16'(-3497);
			440: out = 16'(12287);
			441: out = 16'(-6746);
			442: out = 16'(463);
			443: out = 16'(-18660);
			444: out = 16'(11441);
			445: out = 16'(-26954);
			446: out = 16'(-7289);
			447: out = 16'(17035);
			448: out = 16'(3870);
			449: out = 16'(11913);
			450: out = 16'(21502);
			451: out = 16'(-3368);
			452: out = 16'(351);
			453: out = 16'(-26189);
			454: out = 16'(6527);
			455: out = 16'(-27999);
			456: out = 16'(25757);
			457: out = 16'(-14539);
			458: out = 16'(597);
			459: out = 16'(2798);
			460: out = 16'(-23380);
			461: out = 16'(-9950);
			462: out = 16'(-24961);
			463: out = 16'(29692);
			464: out = 16'(13742);
			465: out = 16'(15591);
			466: out = 16'(6914);
			467: out = 16'(-16246);
			468: out = 16'(110);
			469: out = 16'(-7322);
			470: out = 16'(-20276);
			471: out = 16'(-685);
			472: out = 16'(-5284);
			473: out = 16'(-16091);
			474: out = 16'(-11409);
			475: out = 16'(1100);
			476: out = 16'(-17523);
			477: out = 16'(-4188);
			478: out = 16'(-7498);
			479: out = 16'(15637);
			480: out = 16'(4620);
			481: out = 16'(7382);
			482: out = 16'(20376);
			483: out = 16'(-9280);
			484: out = 16'(23570);
			485: out = 16'(-1739);
			486: out = 16'(4277);
			487: out = 16'(5058);
			488: out = 16'(-607);
			489: out = 16'(4304);
			490: out = 16'(959);
			491: out = 16'(-2176);
			492: out = 16'(-1071);
			493: out = 16'(-27377);
			494: out = 16'(-6908);
			495: out = 16'(-6988);
			496: out = 16'(-4462);
			497: out = 16'(21647);
			498: out = 16'(-9548);
			499: out = 16'(-19029);
			500: out = 16'(-3824);
			501: out = 16'(11136);
			502: out = 16'(2846);
			503: out = 16'(11172);
			504: out = 16'(-2869);
			505: out = 16'(6701);
			506: out = 16'(3534);
			507: out = 16'(-12478);
			508: out = 16'(3820);
			509: out = 16'(528);
			510: out = 16'(4423);
			511: out = 16'(11248);
			512: out = 16'(-5585);
			513: out = 16'(25514);
			514: out = 16'(-4264);
			515: out = 16'(-156);
			516: out = 16'(19073);
			517: out = 16'(-14865);
			518: out = 16'(14289);
			519: out = 16'(754);
			520: out = 16'(-2894);
			521: out = 16'(20287);
			522: out = 16'(1339);
			523: out = 16'(-30297);
			524: out = 16'(-9101);
			525: out = 16'(-19274);
			526: out = 16'(3380);
			527: out = 16'(-8430);
			528: out = 16'(26137);
			529: out = 16'(-9917);
			530: out = 16'(-2676);
			531: out = 16'(-29676);
			532: out = 16'(-11215);
			533: out = 16'(-4748);
			534: out = 16'(12546);
			535: out = 16'(-3202);
			536: out = 16'(15266);
			537: out = 16'(6123);
			538: out = 16'(0);
			539: out = 16'(-10997);
			540: out = 16'(907);
			541: out = 16'(1036);
			542: out = 16'(1089);
			543: out = 16'(19887);
			544: out = 16'(-12990);
			545: out = 16'(13250);
			546: out = 16'(-17002);
			547: out = 16'(17223);
			548: out = 16'(-653);
			549: out = 16'(5659);
			550: out = 16'(8794);
			551: out = 16'(-29173);
			552: out = 16'(385);
			553: out = 16'(1498);
			554: out = 16'(-12309);
			555: out = 16'(29407);
			556: out = 16'(-10276);
			557: out = 16'(1685);
			558: out = 16'(6012);
			559: out = 16'(5025);
			560: out = 16'(18653);
			561: out = 16'(13314);
			562: out = 16'(-6792);
			563: out = 16'(-28151);
			564: out = 16'(3211);
			565: out = 16'(8164);
			566: out = 16'(1842);
			567: out = 16'(17481);
			568: out = 16'(-17872);
			569: out = 16'(7967);
			570: out = 16'(-30415);
			571: out = 16'(-4518);
			572: out = 16'(4611);
			573: out = 16'(-23344);
			574: out = 16'(10390);
			575: out = 16'(-3253);
			576: out = 16'(11127);
			577: out = 16'(-11029);
			578: out = 16'(-14452);
			579: out = 16'(211);
			580: out = 16'(-10776);
			581: out = 16'(12820);
			582: out = 16'(-3797);
			583: out = 16'(17099);
			584: out = 16'(-139);
			585: out = 16'(15360);
			586: out = 16'(6541);
			587: out = 16'(14074);
			588: out = 16'(4282);
			589: out = 16'(-2367);
			590: out = 16'(-24766);
			591: out = 16'(8291);
			592: out = 16'(1515);
			593: out = 16'(-8864);
			594: out = 16'(98);
			595: out = 16'(6482);
			596: out = 16'(-26963);
			597: out = 16'(110);
			598: out = 16'(-259);
			599: out = 16'(6676);
			600: out = 16'(24137);
			601: out = 16'(-24786);
			602: out = 16'(-3279);
			603: out = 16'(-330);
			604: out = 16'(8130);
			605: out = 16'(-18824);
			606: out = 16'(19549);
			607: out = 16'(-6383);
			608: out = 16'(6580);
			609: out = 16'(-2331);
			610: out = 16'(-10380);
			611: out = 16'(4818);
			612: out = 16'(10232);
			613: out = 16'(22005);
			614: out = 16'(-10772);
			615: out = 16'(7412);
			616: out = 16'(-19188);
			617: out = 16'(11188);
			618: out = 16'(-6403);
			619: out = 16'(2311);
			620: out = 16'(-8332);
			621: out = 16'(-22438);
			622: out = 16'(8270);
			623: out = 16'(-4197);
			624: out = 16'(4357);
			625: out = 16'(8545);
			626: out = 16'(12132);
			627: out = 16'(2611);
			628: out = 16'(19199);
			629: out = 16'(623);
			630: out = 16'(-22790);
			631: out = 16'(2674);
			632: out = 16'(-1555);
			633: out = 16'(8734);
			634: out = 16'(9523);
			635: out = 16'(-4419);
			636: out = 16'(906);
			637: out = 16'(7427);
			638: out = 16'(25343);
			639: out = 16'(-27201);
			640: out = 16'(18152);
			641: out = 16'(-23305);
			642: out = 16'(-29418);
			643: out = 16'(7836);
			644: out = 16'(12848);
			645: out = 16'(29887);
			646: out = 16'(15881);
			647: out = 16'(-24373);
			648: out = 16'(1630);
			649: out = 16'(633);
			650: out = 16'(-744);
			651: out = 16'(7789);
			652: out = 16'(15634);
			653: out = 16'(-11049);
			654: out = 16'(15370);
			655: out = 16'(134);
			656: out = 16'(3681);
			657: out = 16'(14913);
			658: out = 16'(-27812);
			659: out = 16'(-5927);
			660: out = 16'(-17779);
			661: out = 16'(-12281);
			662: out = 16'(-5674);
			663: out = 16'(2428);
			664: out = 16'(7395);
			665: out = 16'(3597);
			666: out = 16'(1707);
			667: out = 16'(-10544);
			668: out = 16'(-11885);
			669: out = 16'(8104);
			670: out = 16'(2729);
			671: out = 16'(16656);
			672: out = 16'(4296);
			673: out = 16'(-11664);
			674: out = 16'(-9509);
			675: out = 16'(-13403);
			676: out = 16'(494);
			677: out = 16'(-637);
			678: out = 16'(21103);
			679: out = 16'(-2184);
			680: out = 16'(12894);
			681: out = 16'(-108);
			682: out = 16'(-9309);
			683: out = 16'(1995);
			684: out = 16'(7010);
			685: out = 16'(1143);
			686: out = 16'(2433);
			687: out = 16'(398);
			688: out = 16'(-5577);
			689: out = 16'(11943);
			690: out = 16'(-4285);
			691: out = 16'(20560);
			692: out = 16'(-30932);
			693: out = 16'(1104);
			694: out = 16'(-15931);
			695: out = 16'(-11894);
			696: out = 16'(11008);
			697: out = 16'(-2208);
			698: out = 16'(2586);
			699: out = 16'(-550);
			700: out = 16'(-4094);
			701: out = 16'(-10215);
			702: out = 16'(-836);
			703: out = 16'(4113);
			704: out = 16'(-8944);
			705: out = 16'(-11862);
			706: out = 16'(2315);
			707: out = 16'(-17742);
			708: out = 16'(10714);
			709: out = 16'(9984);
			710: out = 16'(3025);
			711: out = 16'(414);
			712: out = 16'(5160);
			713: out = 16'(1139);
			714: out = 16'(8859);
			715: out = 16'(13722);
			716: out = 16'(-628);
			717: out = 16'(4670);
			718: out = 16'(-1470);
			719: out = 16'(-2388);
			720: out = 16'(5337);
			721: out = 16'(3524);
			722: out = 16'(15138);
			723: out = 16'(13605);
			724: out = 16'(-5971);
			725: out = 16'(11422);
			726: out = 16'(-7801);
			727: out = 16'(1152);
			728: out = 16'(2638);
			729: out = 16'(7557);
			730: out = 16'(-3797);
			731: out = 16'(14446);
			732: out = 16'(-11244);
			733: out = 16'(13809);
			734: out = 16'(-5930);
			735: out = 16'(15824);
			736: out = 16'(2448);
			737: out = 16'(-5948);
			738: out = 16'(7532);
			739: out = 16'(-20077);
			740: out = 16'(14045);
			741: out = 16'(-4064);
			742: out = 16'(14353);
			743: out = 16'(12689);
			744: out = 16'(-6853);
			745: out = 16'(-18009);
			746: out = 16'(-5844);
			747: out = 16'(5673);
			748: out = 16'(-4618);
			749: out = 16'(2708);
			750: out = 16'(-6999);
			751: out = 16'(9525);
			752: out = 16'(-17515);
			753: out = 16'(1724);
			754: out = 16'(14070);
			755: out = 16'(-17306);
			756: out = 16'(24754);
			757: out = 16'(-1169);
			758: out = 16'(-4215);
			759: out = 16'(19404);
			760: out = 16'(-3057);
			761: out = 16'(13544);
			762: out = 16'(11679);
			763: out = 16'(5331);
			764: out = 16'(-20917);
			765: out = 16'(5242);
			766: out = 16'(-12795);
			767: out = 16'(12835);
			768: out = 16'(-4491);
			769: out = 16'(14880);
			770: out = 16'(-7349);
			771: out = 16'(19339);
			772: out = 16'(-6531);
			773: out = 16'(13184);
			774: out = 16'(-12681);
			775: out = 16'(12455);
			776: out = 16'(-15727);
			777: out = 16'(5361);
			778: out = 16'(-832);
			779: out = 16'(-1825);
			780: out = 16'(7326);
			781: out = 16'(-9068);
			782: out = 16'(15193);
			783: out = 16'(-20607);
			784: out = 16'(-1949);
			785: out = 16'(-17045);
			786: out = 16'(-11471);
			787: out = 16'(1641);
			788: out = 16'(2028);
			789: out = 16'(-15928);
			790: out = 16'(4938);
			791: out = 16'(-28171);
			792: out = 16'(-176);
			793: out = 16'(874);
			794: out = 16'(2823);
			795: out = 16'(6535);
			796: out = 16'(4383);
			797: out = 16'(-10608);
			798: out = 16'(-3194);
			799: out = 16'(-5776);
			800: out = 16'(-1996);
			801: out = 16'(1063);
			802: out = 16'(-18779);
			803: out = 16'(12324);
			804: out = 16'(-15101);
			805: out = 16'(22883);
			806: out = 16'(-3375);
			807: out = 16'(5663);
			808: out = 16'(-27780);
			809: out = 16'(-19660);
			810: out = 16'(-6666);
			811: out = 16'(929);
			812: out = 16'(14156);
			813: out = 16'(9252);
			814: out = 16'(-1223);
			815: out = 16'(12599);
			816: out = 16'(-5269);
			817: out = 16'(-6303);
			818: out = 16'(22893);
			819: out = 16'(5928);
			820: out = 16'(-16456);
			821: out = 16'(8460);
			822: out = 16'(-8170);
			823: out = 16'(3210);
			824: out = 16'(4485);
			825: out = 16'(-13215);
			826: out = 16'(18236);
			827: out = 16'(-6215);
			828: out = 16'(11837);
			829: out = 16'(-2074);
			830: out = 16'(17317);
			831: out = 16'(-2532);
			832: out = 16'(-15896);
			833: out = 16'(5257);
			834: out = 16'(-6317);
			835: out = 16'(-65);
			836: out = 16'(-8583);
			837: out = 16'(17562);
			838: out = 16'(-16891);
			839: out = 16'(4025);
			840: out = 16'(12335);
			841: out = 16'(-3092);
			842: out = 16'(-65);
			843: out = 16'(-4628);
			844: out = 16'(436);
			845: out = 16'(6822);
			846: out = 16'(13412);
			847: out = 16'(9567);
			848: out = 16'(-2304);
			849: out = 16'(19526);
			850: out = 16'(-12558);
			851: out = 16'(5726);
			852: out = 16'(13084);
			853: out = 16'(-2607);
			854: out = 16'(-612);
			855: out = 16'(6167);
			856: out = 16'(-16965);
			857: out = 16'(8611);
			858: out = 16'(13808);
			859: out = 16'(-13067);
			860: out = 16'(18866);
			861: out = 16'(3137);
			862: out = 16'(-1849);
			863: out = 16'(-6755);
			864: out = 16'(-389);
			865: out = 16'(-24467);
			866: out = 16'(10502);
			867: out = 16'(3865);
			868: out = 16'(799);
			869: out = 16'(13289);
			870: out = 16'(-5645);
			871: out = 16'(-2932);
			872: out = 16'(-5582);
			873: out = 16'(10027);
			874: out = 16'(-9139);
			875: out = 16'(-1833);
			876: out = 16'(9375);
			877: out = 16'(2106);
			878: out = 16'(-13069);
			879: out = 16'(11694);
			880: out = 16'(-3590);
			881: out = 16'(-6334);
			882: out = 16'(7158);
			883: out = 16'(15300);
			884: out = 16'(-26833);
			885: out = 16'(26803);
			886: out = 16'(-12746);
			887: out = 16'(2762);
			888: out = 16'(-20501);
			889: out = 16'(2362);
			890: out = 16'(-9165);
			891: out = 16'(-2900);
			892: out = 16'(-529);
			893: out = 16'(-18356);
			894: out = 16'(23158);
			895: out = 16'(-11780);
			896: out = 16'(2785);
			897: out = 16'(5594);
			898: out = 16'(-1504);
			899: out = 16'(-4785);
			900: out = 16'(3825);
			901: out = 16'(2527);
			902: out = 16'(2635);
			903: out = 16'(1839);
			904: out = 16'(-2212);
			905: out = 16'(582);
			906: out = 16'(10010);
			907: out = 16'(3234);
			908: out = 16'(-11492);
			909: out = 16'(-3287);
			910: out = 16'(-4935);
			911: out = 16'(-952);
			912: out = 16'(-8451);
			913: out = 16'(3457);
			914: out = 16'(4049);
			915: out = 16'(-4047);
			916: out = 16'(148);
			917: out = 16'(-14189);
			918: out = 16'(5601);
			919: out = 16'(11250);
			920: out = 16'(-938);
			921: out = 16'(13659);
			922: out = 16'(-8410);
			923: out = 16'(1171);
			924: out = 16'(-7269);
			925: out = 16'(-12994);
			926: out = 16'(233);
			927: out = 16'(-7271);
			928: out = 16'(7810);
			929: out = 16'(-18457);
			930: out = 16'(-3317);
			931: out = 16'(-7967);
			932: out = 16'(1991);
			933: out = 16'(4437);
			934: out = 16'(-4003);
			935: out = 16'(1932);
			936: out = 16'(-3787);
			937: out = 16'(-4952);
			938: out = 16'(8153);
			939: out = 16'(1618);
			940: out = 16'(-9291);
			941: out = 16'(1800);
			942: out = 16'(11216);
			943: out = 16'(-27578);
			944: out = 16'(14522);
			945: out = 16'(-6003);
			946: out = 16'(-10307);
			947: out = 16'(4935);
			948: out = 16'(-15727);
			949: out = 16'(6678);
			950: out = 16'(-8461);
			951: out = 16'(7423);
			952: out = 16'(-6918);
			953: out = 16'(21216);
			954: out = 16'(-815);
			955: out = 16'(-938);
			956: out = 16'(-5995);
			957: out = 16'(6556);
			958: out = 16'(-9233);
			959: out = 16'(19038);
			960: out = 16'(14767);
			961: out = 16'(11959);
			962: out = 16'(5915);
			963: out = 16'(-4444);
			964: out = 16'(2979);
			965: out = 16'(2838);
			966: out = 16'(-1271);
			967: out = 16'(8111);
			968: out = 16'(-10426);
			969: out = 16'(-2139);
			970: out = 16'(-3653);
			971: out = 16'(-5866);
			972: out = 16'(17742);
			973: out = 16'(-7658);
			974: out = 16'(8644);
			975: out = 16'(-1314);
			976: out = 16'(4288);
			977: out = 16'(-6840);
			978: out = 16'(-7091);
			979: out = 16'(708);
			980: out = 16'(-1553);
			981: out = 16'(1258);
			982: out = 16'(-10468);
			983: out = 16'(1307);
			984: out = 16'(-1407);
			985: out = 16'(4990);
			986: out = 16'(-9854);
			987: out = 16'(4985);
			988: out = 16'(-1797);
			989: out = 16'(7808);
			990: out = 16'(9979);
			991: out = 16'(17742);
			992: out = 16'(6378);
			993: out = 16'(1179);
			994: out = 16'(-11756);
			995: out = 16'(-3376);
			996: out = 16'(14336);
			997: out = 16'(-20258);
			998: out = 16'(9209);
			999: out = 16'(15956);
			1000: out = 16'(-10928);
			1001: out = 16'(7924);
			1002: out = 16'(-11151);
			1003: out = 16'(9108);
			1004: out = 16'(334);
			1005: out = 16'(12182);
			1006: out = 16'(-8751);
			1007: out = 16'(8473);
			1008: out = 16'(-8098);
			1009: out = 16'(2019);
			1010: out = 16'(-297);
			1011: out = 16'(-2290);
			1012: out = 16'(-10718);
			1013: out = 16'(-14411);
			1014: out = 16'(14446);
			1015: out = 16'(-8601);
			1016: out = 16'(-2903);
			1017: out = 16'(9266);
			1018: out = 16'(664);
			1019: out = 16'(-8266);
			1020: out = 16'(-10224);
			1021: out = 16'(6943);
			1022: out = 16'(-3560);
			1023: out = 16'(8886);
			1024: out = 16'(2182);
			1025: out = 16'(-18223);
			1026: out = 16'(6599);
			1027: out = 16'(-6913);
			1028: out = 16'(-9187);
			1029: out = 16'(19529);
			1030: out = 16'(3586);
			1031: out = 16'(-9714);
			1032: out = 16'(571);
			1033: out = 16'(-2542);
			1034: out = 16'(-24682);
			1035: out = 16'(3353);
			1036: out = 16'(-4348);
			1037: out = 16'(-3370);
			1038: out = 16'(8307);
			1039: out = 16'(-6921);
			1040: out = 16'(-1554);
			1041: out = 16'(12368);
			1042: out = 16'(1166);
			1043: out = 16'(-11720);
			1044: out = 16'(21348);
			1045: out = 16'(-14274);
			1046: out = 16'(11076);
			1047: out = 16'(-11432);
			1048: out = 16'(-1943);
			1049: out = 16'(3467);
			1050: out = 16'(8672);
			1051: out = 16'(6723);
			1052: out = 16'(-15708);
			1053: out = 16'(-897);
			1054: out = 16'(-19158);
			1055: out = 16'(1098);
			1056: out = 16'(-11294);
			1057: out = 16'(9385);
			1058: out = 16'(979);
			1059: out = 16'(-13504);
			1060: out = 16'(-9151);
			1061: out = 16'(9486);
			1062: out = 16'(3722);
			1063: out = 16'(10980);
			1064: out = 16'(-4915);
			1065: out = 16'(3835);
			1066: out = 16'(-8739);
			1067: out = 16'(-3295);
			1068: out = 16'(3130);
			1069: out = 16'(19631);
			1070: out = 16'(11381);
			1071: out = 16'(-6495);
			1072: out = 16'(-4034);
			1073: out = 16'(-2136);
			1074: out = 16'(-14386);
			1075: out = 16'(-12495);
			1076: out = 16'(2236);
			1077: out = 16'(1584);
			1078: out = 16'(3218);
			1079: out = 16'(-754);
			1080: out = 16'(4114);
			1081: out = 16'(4760);
			1082: out = 16'(14175);
			1083: out = 16'(2870);
			1084: out = 16'(3059);
			1085: out = 16'(10592);
			1086: out = 16'(-2807);
			1087: out = 16'(221);
			1088: out = 16'(-9121);
			1089: out = 16'(11547);
			1090: out = 16'(-8844);
			1091: out = 16'(-3629);
			1092: out = 16'(-5007);
			1093: out = 16'(-25837);
			1094: out = 16'(5220);
			1095: out = 16'(12375);
			1096: out = 16'(-1249);
			1097: out = 16'(-6363);
			1098: out = 16'(13312);
			1099: out = 16'(-30504);
			1100: out = 16'(8188);
			1101: out = 16'(9115);
			1102: out = 16'(-5063);
			1103: out = 16'(16989);
			1104: out = 16'(-15620);
			1105: out = 16'(2716);
			1106: out = 16'(11999);
			1107: out = 16'(4721);
			1108: out = 16'(1397);
			1109: out = 16'(3515);
			1110: out = 16'(279);
			1111: out = 16'(-5220);
			1112: out = 16'(-8813);
			1113: out = 16'(3627);
			1114: out = 16'(8114);
			1115: out = 16'(4154);
			1116: out = 16'(9152);
			1117: out = 16'(-5569);
			1118: out = 16'(-6325);
			1119: out = 16'(11141);
			1120: out = 16'(-8669);
			1121: out = 16'(2980);
			1122: out = 16'(2967);
			1123: out = 16'(10190);
			1124: out = 16'(181);
			1125: out = 16'(3106);
			1126: out = 16'(2038);
			1127: out = 16'(-783);
			1128: out = 16'(-5443);
			1129: out = 16'(3521);
			1130: out = 16'(-25140);
			1131: out = 16'(10145);
			1132: out = 16'(1470);
			1133: out = 16'(2291);
			1134: out = 16'(16921);
			1135: out = 16'(-18916);
			1136: out = 16'(1087);
			1137: out = 16'(4672);
			1138: out = 16'(-25696);
			1139: out = 16'(8156);
			1140: out = 16'(-3788);
			1141: out = 16'(-739);
			1142: out = 16'(3606);
			1143: out = 16'(-15320);
			1144: out = 16'(14304);
			1145: out = 16'(3693);
			1146: out = 16'(-198);
			1147: out = 16'(-915);
			1148: out = 16'(9699);
			1149: out = 16'(-4387);
			1150: out = 16'(-9521);
			1151: out = 16'(1803);
			1152: out = 16'(5099);
			1153: out = 16'(7904);
			1154: out = 16'(-2504);
			1155: out = 16'(2066);
			1156: out = 16'(-11583);
			1157: out = 16'(8175);
			1158: out = 16'(-13163);
			1159: out = 16'(-436);
			1160: out = 16'(12246);
			1161: out = 16'(-10929);
			1162: out = 16'(1768);
			1163: out = 16'(6022);
			1164: out = 16'(-7583);
			1165: out = 16'(9384);
			1166: out = 16'(-7661);
			1167: out = 16'(-1281);
			1168: out = 16'(718);
			1169: out = 16'(-6920);
			1170: out = 16'(-6173);
			1171: out = 16'(7210);
			1172: out = 16'(87);
			1173: out = 16'(20084);
			1174: out = 16'(-16333);
			1175: out = 16'(-12594);
			1176: out = 16'(10961);
			1177: out = 16'(-15784);
			1178: out = 16'(4377);
			1179: out = 16'(14);
			1180: out = 16'(7517);
			1181: out = 16'(1906);
			1182: out = 16'(-3643);
			1183: out = 16'(-11551);
			1184: out = 16'(3541);
			1185: out = 16'(-1173);
			1186: out = 16'(13470);
			1187: out = 16'(16177);
			1188: out = 16'(-16355);
			1189: out = 16'(-9017);
			1190: out = 16'(1857);
			1191: out = 16'(12773);
			1192: out = 16'(3738);
			1193: out = 16'(5905);
			1194: out = 16'(-9336);
			1195: out = 16'(-19928);
			1196: out = 16'(16230);
			1197: out = 16'(-8373);
			1198: out = 16'(13899);
			1199: out = 16'(1341);
			1200: out = 16'(-11353);
			1201: out = 16'(17);
			1202: out = 16'(-3225);
			1203: out = 16'(667);
			1204: out = 16'(11114);
			1205: out = 16'(8766);
			1206: out = 16'(3548);
			1207: out = 16'(3241);
			1208: out = 16'(-23210);
			1209: out = 16'(-222);
			1210: out = 16'(3523);
			1211: out = 16'(698);
			1212: out = 16'(6054);
			1213: out = 16'(-16230);
			1214: out = 16'(3841);
			1215: out = 16'(-8923);
			1216: out = 16'(-2935);
			1217: out = 16'(-21722);
			1218: out = 16'(17476);
			1219: out = 16'(531);
			1220: out = 16'(-8259);
			1221: out = 16'(2088);
			1222: out = 16'(-16387);
			1223: out = 16'(-5834);
			1224: out = 16'(4689);
			1225: out = 16'(8573);
			1226: out = 16'(5688);
			1227: out = 16'(-6301);
			1228: out = 16'(1787);
			1229: out = 16'(-16911);
			1230: out = 16'(16151);
			1231: out = 16'(-21881);
			1232: out = 16'(16691);
			1233: out = 16'(-5517);
			1234: out = 16'(-13149);
			1235: out = 16'(7783);
			1236: out = 16'(-11851);
			1237: out = 16'(9905);
			1238: out = 16'(-2619);
			1239: out = 16'(19673);
			1240: out = 16'(-7048);
			1241: out = 16'(4945);
			1242: out = 16'(-12136);
			1243: out = 16'(-6745);
			1244: out = 16'(7068);
			1245: out = 16'(-17537);
			1246: out = 16'(3385);
			1247: out = 16'(-3796);
			1248: out = 16'(-6869);
			1249: out = 16'(11159);
			1250: out = 16'(13729);
			1251: out = 16'(-5733);
			1252: out = 16'(-11043);
			1253: out = 16'(4521);
			1254: out = 16'(-5318);
			1255: out = 16'(5663);
			1256: out = 16'(1600);
			1257: out = 16'(11384);
			1258: out = 16'(15723);
			1259: out = 16'(1297);
			1260: out = 16'(13308);
			1261: out = 16'(-13969);
			1262: out = 16'(-2742);
			1263: out = 16'(3024);
			1264: out = 16'(11090);
			1265: out = 16'(1203);
			1266: out = 16'(-3022);
			1267: out = 16'(-11075);
			1268: out = 16'(-8686);
			1269: out = 16'(14553);
			1270: out = 16'(-19954);
			1271: out = 16'(3367);
			1272: out = 16'(-2377);
			1273: out = 16'(-5500);
			1274: out = 16'(8940);
			1275: out = 16'(787);
			1276: out = 16'(284);
			1277: out = 16'(114);
			1278: out = 16'(8478);
			1279: out = 16'(-26897);
			1280: out = 16'(1807);
			1281: out = 16'(-11668);
			1282: out = 16'(-8385);
			1283: out = 16'(12592);
			1284: out = 16'(-2105);
			1285: out = 16'(1925);
			1286: out = 16'(-7575);
			1287: out = 16'(8614);
			1288: out = 16'(-6190);
			1289: out = 16'(5022);
			1290: out = 16'(-26129);
			1291: out = 16'(-2010);
			1292: out = 16'(2074);
			1293: out = 16'(-3653);
			1294: out = 16'(4751);
			1295: out = 16'(-1153);
			1296: out = 16'(1892);
			1297: out = 16'(-6727);
			1298: out = 16'(-551);
			1299: out = 16'(156);
			1300: out = 16'(3826);
			1301: out = 16'(17007);
			1302: out = 16'(6229);
			1303: out = 16'(10342);
			1304: out = 16'(-22146);
			1305: out = 16'(747);
			1306: out = 16'(-2063);
			1307: out = 16'(2563);
			1308: out = 16'(-2107);
			1309: out = 16'(8970);
			1310: out = 16'(-5361);
			1311: out = 16'(-22118);
			1312: out = 16'(8583);
			1313: out = 16'(-9702);
			1314: out = 16'(10448);
			1315: out = 16'(3505);
			1316: out = 16'(-2493);
			1317: out = 16'(7520);
			1318: out = 16'(-12737);
			1319: out = 16'(-458);
			1320: out = 16'(-3077);
			1321: out = 16'(23762);
			1322: out = 16'(-15935);
			1323: out = 16'(17220);
			1324: out = 16'(-21803);
			1325: out = 16'(5662);
			1326: out = 16'(6073);
			1327: out = 16'(-22711);
			1328: out = 16'(19156);
			1329: out = 16'(7260);
			1330: out = 16'(8);
			1331: out = 16'(-8991);
			1332: out = 16'(-5005);
			1333: out = 16'(1580);
			1334: out = 16'(7344);
			1335: out = 16'(-15320);
			1336: out = 16'(-5254);
			1337: out = 16'(17519);
			1338: out = 16'(-15302);
			1339: out = 16'(3810);
			1340: out = 16'(2400);
			1341: out = 16'(24109);
			1342: out = 16'(-12183);
			1343: out = 16'(-3707);
			1344: out = 16'(-954);
			1345: out = 16'(-12000);
			1346: out = 16'(21271);
			1347: out = 16'(-13822);
			1348: out = 16'(8395);
			1349: out = 16'(16987);
			1350: out = 16'(-1331);
			1351: out = 16'(-5883);
			1352: out = 16'(-8456);
			1353: out = 16'(11148);
			1354: out = 16'(-270);
			1355: out = 16'(18115);
			1356: out = 16'(2031);
			1357: out = 16'(9147);
			1358: out = 16'(17243);
			1359: out = 16'(-12632);
			1360: out = 16'(11651);
			1361: out = 16'(-10454);
			1362: out = 16'(10948);
			1363: out = 16'(-10894);
			1364: out = 16'(-4845);
			1365: out = 16'(11884);
			1366: out = 16'(-15946);
			1367: out = 16'(4375);
			1368: out = 16'(-22530);
			1369: out = 16'(4744);
			1370: out = 16'(-26284);
			1371: out = 16'(-511);
			1372: out = 16'(3870);
			1373: out = 16'(-9158);
			1374: out = 16'(-1060);
			1375: out = 16'(-1095);
			1376: out = 16'(5951);
			1377: out = 16'(390);
			1378: out = 16'(2186);
			1379: out = 16'(-8765);
			1380: out = 16'(13889);
			1381: out = 16'(-28005);
			1382: out = 16'(17224);
			1383: out = 16'(1075);
			1384: out = 16'(-694);
			1385: out = 16'(13208);
			1386: out = 16'(-10216);
			1387: out = 16'(1260);
			1388: out = 16'(12971);
			1389: out = 16'(-26722);
			1390: out = 16'(7405);
			1391: out = 16'(3459);
			1392: out = 16'(3976);
			1393: out = 16'(5115);
			1394: out = 16'(11064);
			1395: out = 16'(-24905);
			1396: out = 16'(14107);
			1397: out = 16'(-16641);
			1398: out = 16'(6358);
			1399: out = 16'(5594);
			1400: out = 16'(-26254);
			1401: out = 16'(4945);
			1402: out = 16'(-23842);
			1403: out = 16'(2284);
			1404: out = 16'(-21386);
			1405: out = 16'(1588);
			1406: out = 16'(-2430);
			1407: out = 16'(-14210);
			1408: out = 16'(-1287);
			1409: out = 16'(-19366);
			1410: out = 16'(13483);
			1411: out = 16'(-5450);
			1412: out = 16'(-9343);
			1413: out = 16'(4244);
			1414: out = 16'(-9947);
			1415: out = 16'(-5294);
			1416: out = 16'(-10259);
			1417: out = 16'(-8233);
			1418: out = 16'(-3810);
			1419: out = 16'(10818);
			1420: out = 16'(-13287);
			1421: out = 16'(18952);
			1422: out = 16'(-5855);
			1423: out = 16'(-21240);
			1424: out = 16'(15870);
			1425: out = 16'(-25462);
			1426: out = 16'(9258);
			1427: out = 16'(-3685);
			1428: out = 16'(3015);
			1429: out = 16'(40);
			1430: out = 16'(17841);
			1431: out = 16'(-12937);
			1432: out = 16'(7157);
			1433: out = 16'(-199);
			1434: out = 16'(-3261);
			1435: out = 16'(13569);
			1436: out = 16'(10880);
			1437: out = 16'(1569);
			1438: out = 16'(-9345);
			1439: out = 16'(-2169);
			1440: out = 16'(-19024);
			1441: out = 16'(-9317);
			1442: out = 16'(16130);
			1443: out = 16'(626);
			1444: out = 16'(15859);
			1445: out = 16'(-1176);
			1446: out = 16'(-4118);
			1447: out = 16'(-5148);
			1448: out = 16'(-19397);
			1449: out = 16'(8100);
			1450: out = 16'(-9859);
			1451: out = 16'(953);
			1452: out = 16'(-18486);
			1453: out = 16'(1342);
			1454: out = 16'(-18147);
			1455: out = 16'(24299);
			1456: out = 16'(-500);
			1457: out = 16'(-9956);
			1458: out = 16'(16331);
			1459: out = 16'(-27113);
			1460: out = 16'(3209);
			1461: out = 16'(-19710);
			1462: out = 16'(5017);
			1463: out = 16'(7237);
			1464: out = 16'(11320);
			1465: out = 16'(7616);
			1466: out = 16'(501);
			1467: out = 16'(1342);
			1468: out = 16'(-1529);
			1469: out = 16'(-10917);
			1470: out = 16'(9075);
			1471: out = 16'(-8429);
			1472: out = 16'(6332);
			1473: out = 16'(-7334);
			1474: out = 16'(6738);
			1475: out = 16'(5602);
			1476: out = 16'(-9590);
			1477: out = 16'(10144);
			1478: out = 16'(-15787);
			1479: out = 16'(-23430);
			1480: out = 16'(1416);
			1481: out = 16'(10024);
			1482: out = 16'(438);
			1483: out = 16'(12654);
			1484: out = 16'(-14676);
			1485: out = 16'(533);
			1486: out = 16'(-13975);
			1487: out = 16'(8863);
			1488: out = 16'(-24200);
			1489: out = 16'(19846);
			1490: out = 16'(-16447);
			1491: out = 16'(-3353);
			1492: out = 16'(-886);
			1493: out = 16'(-29225);
			1494: out = 16'(12651);
			1495: out = 16'(-2228);
			1496: out = 16'(-26623);
			1497: out = 16'(15552);
			1498: out = 16'(-3286);
			1499: out = 16'(-326);
			1500: out = 16'(10419);
			1501: out = 16'(-203);
			1502: out = 16'(11841);
			1503: out = 16'(3219);
			1504: out = 16'(2204);
			1505: out = 16'(-4127);
			1506: out = 16'(-7008);
			1507: out = 16'(-7319);
			1508: out = 16'(1683);
			1509: out = 16'(-13906);
			1510: out = 16'(2495);
			1511: out = 16'(-11183);
			1512: out = 16'(1994);
			1513: out = 16'(-3405);
			1514: out = 16'(1405);
			1515: out = 16'(1961);
			1516: out = 16'(-3777);
			1517: out = 16'(-4901);
			1518: out = 16'(-2122);
			1519: out = 16'(7352);
			1520: out = 16'(1709);
			1521: out = 16'(7116);
			1522: out = 16'(-3563);
			1523: out = 16'(6531);
			1524: out = 16'(-9651);
			1525: out = 16'(232);
			1526: out = 16'(4768);
			1527: out = 16'(-925);
			1528: out = 16'(2582);
			1529: out = 16'(4974);
			1530: out = 16'(-32118);
			1531: out = 16'(8796);
			1532: out = 16'(-13123);
			1533: out = 16'(-781);
			1534: out = 16'(1957);
			1535: out = 16'(3444);
			1536: out = 16'(3437);
			1537: out = 16'(18077);
			1538: out = 16'(4546);
			1539: out = 16'(7049);
			1540: out = 16'(2064);
			1541: out = 16'(-2458);
			1542: out = 16'(8840);
			1543: out = 16'(-18384);
			1544: out = 16'(19502);
			1545: out = 16'(-30390);
			1546: out = 16'(21062);
			1547: out = 16'(-5357);
			1548: out = 16'(456);
			1549: out = 16'(742);
			1550: out = 16'(-338);
			1551: out = 16'(2953);
			1552: out = 16'(5759);
			1553: out = 16'(20935);
			1554: out = 16'(9773);
			1555: out = 16'(-9862);
			1556: out = 16'(11843);
			1557: out = 16'(780);
			1558: out = 16'(2336);
			1559: out = 16'(2699);
			1560: out = 16'(9990);
			1561: out = 16'(-27095);
			1562: out = 16'(15490);
			1563: out = 16'(-7414);
			1564: out = 16'(-6560);
			1565: out = 16'(11469);
			1566: out = 16'(-27906);
			1567: out = 16'(17782);
			1568: out = 16'(-6462);
			1569: out = 16'(361);
			1570: out = 16'(-1880);
			1571: out = 16'(1705);
			1572: out = 16'(-107);
			1573: out = 16'(8128);
			1574: out = 16'(2507);
			1575: out = 16'(-3200);
			1576: out = 16'(94);
			1577: out = 16'(1455);
			1578: out = 16'(16142);
			1579: out = 16'(-26721);
			1580: out = 16'(12983);
			1581: out = 16'(-19682);
			1582: out = 16'(706);
			1583: out = 16'(-1282);
			1584: out = 16'(-13421);
			1585: out = 16'(3173);
			1586: out = 16'(-3389);
			1587: out = 16'(-13899);
			1588: out = 16'(13792);
			1589: out = 16'(-20179);
			1590: out = 16'(19159);
			1591: out = 16'(5419);
			1592: out = 16'(14816);
			1593: out = 16'(-26704);
			1594: out = 16'(2289);
			1595: out = 16'(-11176);
			1596: out = 16'(8253);
			1597: out = 16'(-14964);
			1598: out = 16'(10201);
			1599: out = 16'(-3510);
			1600: out = 16'(-14432);
			1601: out = 16'(-8653);
			1602: out = 16'(-16827);
			1603: out = 16'(11612);
			1604: out = 16'(1137);
			1605: out = 16'(18195);
			1606: out = 16'(-1237);
			1607: out = 16'(153);
			1608: out = 16'(1412);
			1609: out = 16'(13852);
			1610: out = 16'(6669);
			1611: out = 16'(3486);
			1612: out = 16'(14360);
			1613: out = 16'(-1722);
			1614: out = 16'(-9970);
			1615: out = 16'(11885);
			1616: out = 16'(-11234);
			1617: out = 16'(4664);
			1618: out = 16'(-298);
			1619: out = 16'(8178);
			1620: out = 16'(1064);
			1621: out = 16'(-9513);
			1622: out = 16'(6475);
			1623: out = 16'(-3922);
			1624: out = 16'(14701);
			1625: out = 16'(-1582);
			1626: out = 16'(-741);
			1627: out = 16'(16795);
			1628: out = 16'(-8038);
			1629: out = 16'(-7418);
			1630: out = 16'(25407);
			1631: out = 16'(-7992);
			1632: out = 16'(4914);
			1633: out = 16'(17751);
			1634: out = 16'(-1949);
			1635: out = 16'(3165);
			1636: out = 16'(3355);
			1637: out = 16'(6698);
			1638: out = 16'(5409);
			1639: out = 16'(-16156);
			1640: out = 16'(-3046);
			1641: out = 16'(3869);
			1642: out = 16'(12200);
			1643: out = 16'(10356);
			1644: out = 16'(9075);
			1645: out = 16'(-8167);
			1646: out = 16'(14138);
			1647: out = 16'(-4871);
			1648: out = 16'(-10864);
			1649: out = 16'(9033);
			1650: out = 16'(-17930);
			1651: out = 16'(12402);
			1652: out = 16'(-24143);
			1653: out = 16'(6379);
			1654: out = 16'(351);
			1655: out = 16'(-2828);
			1656: out = 16'(1559);
			1657: out = 16'(12908);
			1658: out = 16'(1080);
			1659: out = 16'(17916);
			1660: out = 16'(-5248);
			1661: out = 16'(7068);
			1662: out = 16'(16904);
			1663: out = 16'(-13674);
			1664: out = 16'(12917);
			1665: out = 16'(7307);
			1666: out = 16'(1703);
			1667: out = 16'(4333);
			1668: out = 16'(2835);
			1669: out = 16'(20021);
			1670: out = 16'(965);
			1671: out = 16'(-7938);
			1672: out = 16'(9511);
			1673: out = 16'(-30714);
			1674: out = 16'(8209);
			1675: out = 16'(1628);
			1676: out = 16'(-6320);
			1677: out = 16'(10859);
			1678: out = 16'(-5929);
			1679: out = 16'(10992);
			1680: out = 16'(-4236);
			1681: out = 16'(-22035);
			1682: out = 16'(2332);
			1683: out = 16'(-3944);
			1684: out = 16'(-8569);
			1685: out = 16'(1574);
			1686: out = 16'(-6731);
			1687: out = 16'(7898);
			1688: out = 16'(-24085);
			1689: out = 16'(6352);
			1690: out = 16'(-3906);
			1691: out = 16'(-4863);
			1692: out = 16'(-7602);
			1693: out = 16'(14320);
			1694: out = 16'(7519);
			1695: out = 16'(9900);
			1696: out = 16'(7509);
			1697: out = 16'(-18828);
			1698: out = 16'(17187);
			1699: out = 16'(-1275);
			1700: out = 16'(11659);
			1701: out = 16'(733);
			1702: out = 16'(-4002);
			1703: out = 16'(14265);
			1704: out = 16'(2620);
			1705: out = 16'(-409);
			1706: out = 16'(7802);
			1707: out = 16'(-16775);
			1708: out = 16'(14816);
			1709: out = 16'(-7081);
			1710: out = 16'(-991);
			1711: out = 16'(5367);
			1712: out = 16'(407);
			1713: out = 16'(-3722);
			1714: out = 16'(21708);
			1715: out = 16'(-18471);
			1716: out = 16'(-3672);
			1717: out = 16'(13069);
			1718: out = 16'(-5715);
			1719: out = 16'(146);
			1720: out = 16'(-6328);
			1721: out = 16'(13417);
			1722: out = 16'(202);
			1723: out = 16'(-599);
			1724: out = 16'(3359);
			1725: out = 16'(-8290);
			1726: out = 16'(-274);
			1727: out = 16'(11819);
			1728: out = 16'(-12625);
			1729: out = 16'(10712);
			1730: out = 16'(-11443);
			1731: out = 16'(-10404);
			1732: out = 16'(13679);
			1733: out = 16'(-411);
			1734: out = 16'(-300);
			1735: out = 16'(4699);
			1736: out = 16'(-10765);
			1737: out = 16'(10744);
			1738: out = 16'(796);
			1739: out = 16'(7187);
			1740: out = 16'(13917);
			1741: out = 16'(-6427);
			1742: out = 16'(13914);
			1743: out = 16'(-22166);
			1744: out = 16'(7107);
			1745: out = 16'(5866);
			1746: out = 16'(5197);
			1747: out = 16'(-5943);
			1748: out = 16'(9063);
			1749: out = 16'(-21264);
			1750: out = 16'(14646);
			1751: out = 16'(-837);
			1752: out = 16'(-5184);
			1753: out = 16'(10233);
			1754: out = 16'(-11950);
			1755: out = 16'(-22255);
			1756: out = 16'(9771);
			1757: out = 16'(-2105);
			1758: out = 16'(-871);
			1759: out = 16'(-1302);
			1760: out = 16'(5964);
			1761: out = 16'(-1018);
			1762: out = 16'(-16481);
			1763: out = 16'(10843);
			1764: out = 16'(-20284);
			1765: out = 16'(17109);
			1766: out = 16'(-745);
			1767: out = 16'(-16067);
			1768: out = 16'(-11281);
			1769: out = 16'(7951);
			1770: out = 16'(-26011);
			1771: out = 16'(14120);
			1772: out = 16'(1833);
			1773: out = 16'(49);
			1774: out = 16'(13175);
			1775: out = 16'(-18124);
			1776: out = 16'(-2984);
			1777: out = 16'(-15465);
			1778: out = 16'(8503);
			1779: out = 16'(4538);
			1780: out = 16'(3405);
			1781: out = 16'(-2311);
			1782: out = 16'(3743);
			1783: out = 16'(-215);
			1784: out = 16'(7946);
			1785: out = 16'(-29425);
			1786: out = 16'(11897);
			1787: out = 16'(-6756);
			1788: out = 16'(-14343);
			1789: out = 16'(17584);
			1790: out = 16'(4114);
			1791: out = 16'(-3265);
			1792: out = 16'(12294);
			1793: out = 16'(-17806);
			1794: out = 16'(3770);
			1795: out = 16'(-414);
			1796: out = 16'(-19479);
			1797: out = 16'(-4461);
			1798: out = 16'(7114);
			1799: out = 16'(12066);
			1800: out = 16'(12652);
			1801: out = 16'(10960);
			1802: out = 16'(-1606);
			1803: out = 16'(2493);
			1804: out = 16'(-28410);
			1805: out = 16'(6952);
			1806: out = 16'(399);
			1807: out = 16'(7017);
			1808: out = 16'(14006);
			1809: out = 16'(-3112);
			1810: out = 16'(-2750);
			1811: out = 16'(-5553);
			1812: out = 16'(-27117);
			1813: out = 16'(14631);
			1814: out = 16'(-12777);
			1815: out = 16'(16254);
			1816: out = 16'(9486);
			1817: out = 16'(-4858);
			1818: out = 16'(8039);
			1819: out = 16'(-25994);
			1820: out = 16'(-8027);
			1821: out = 16'(-3161);
			1822: out = 16'(-5042);
			1823: out = 16'(-5788);
			1824: out = 16'(11936);
			1825: out = 16'(2844);
			1826: out = 16'(9749);
			1827: out = 16'(-4750);
			1828: out = 16'(14084);
			1829: out = 16'(-17590);
			1830: out = 16'(7272);
			1831: out = 16'(6593);
			1832: out = 16'(114);
			1833: out = 16'(6499);
			1834: out = 16'(6741);
			1835: out = 16'(13259);
			1836: out = 16'(15818);
			1837: out = 16'(2935);
			1838: out = 16'(-25550);
			1839: out = 16'(753);
			1840: out = 16'(-11634);
			1841: out = 16'(-5481);
			1842: out = 16'(8300);
			1843: out = 16'(7299);
			1844: out = 16'(-13127);
			1845: out = 16'(4118);
			1846: out = 16'(-21692);
			1847: out = 16'(6738);
			1848: out = 16'(-12053);
			1849: out = 16'(150);
			1850: out = 16'(-1975);
			1851: out = 16'(-5);
			1852: out = 16'(12255);
			1853: out = 16'(9957);
			1854: out = 16'(-19458);
			1855: out = 16'(3142);
			1856: out = 16'(-26054);
			1857: out = 16'(-20052);
			1858: out = 16'(4284);
			1859: out = 16'(-26098);
			1860: out = 16'(12636);
			1861: out = 16'(-1048);
			1862: out = 16'(1045);
			1863: out = 16'(2346);
			1864: out = 16'(9652);
			1865: out = 16'(-15261);
			1866: out = 16'(7191);
			1867: out = 16'(-15154);
			1868: out = 16'(1454);
			1869: out = 16'(-12619);
			1870: out = 16'(13858);
			1871: out = 16'(-8789);
			1872: out = 16'(2431);
			1873: out = 16'(13109);
			1874: out = 16'(-9637);
			1875: out = 16'(-13831);
			1876: out = 16'(5452);
			1877: out = 16'(-7922);
			1878: out = 16'(-4204);
			1879: out = 16'(11016);
			1880: out = 16'(-2610);
			1881: out = 16'(787);
			1882: out = 16'(-327);
			1883: out = 16'(-2345);
			1884: out = 16'(-12037);
			1885: out = 16'(10397);
			1886: out = 16'(10273);
			1887: out = 16'(12596);
			1888: out = 16'(-4396);
			1889: out = 16'(8207);
			1890: out = 16'(-29392);
			1891: out = 16'(-298);
			1892: out = 16'(1988);
			1893: out = 16'(-2414);
			1894: out = 16'(-3128);
			1895: out = 16'(1877);
			1896: out = 16'(-6656);
			1897: out = 16'(7857);
			1898: out = 16'(-9850);
			1899: out = 16'(-888);
			1900: out = 16'(9705);
			1901: out = 16'(-6980);
			1902: out = 16'(18387);
			1903: out = 16'(-3005);
			1904: out = 16'(1099);
			1905: out = 16'(2605);
			1906: out = 16'(-4134);
			1907: out = 16'(940);
			1908: out = 16'(13101);
			1909: out = 16'(-4749);
			1910: out = 16'(1663);
			1911: out = 16'(-16638);
			1912: out = 16'(5808);
			1913: out = 16'(4520);
			1914: out = 16'(-1885);
			1915: out = 16'(5695);
			1916: out = 16'(9140);
			1917: out = 16'(-5813);
			1918: out = 16'(1236);
			1919: out = 16'(9645);
			1920: out = 16'(-5928);
			1921: out = 16'(24397);
			1922: out = 16'(-13554);
			1923: out = 16'(9571);
			1924: out = 16'(5228);
			1925: out = 16'(-9093);
			1926: out = 16'(750);
			1927: out = 16'(-16109);
			1928: out = 16'(-375);
			1929: out = 16'(6290);
			1930: out = 16'(-7225);
			1931: out = 16'(18378);
			1932: out = 16'(-13248);
			1933: out = 16'(13746);
			1934: out = 16'(5047);
			1935: out = 16'(-3844);
			1936: out = 16'(1242);
			1937: out = 16'(-4001);
			1938: out = 16'(-1378);
			1939: out = 16'(2813);
			1940: out = 16'(9165);
			1941: out = 16'(3096);
			1942: out = 16'(9016);
			1943: out = 16'(-6497);
			1944: out = 16'(16215);
			1945: out = 16'(-8018);
			1946: out = 16'(-17111);
			1947: out = 16'(-21521);
			1948: out = 16'(82);
			1949: out = 16'(-5997);
			1950: out = 16'(13783);
			1951: out = 16'(640);
			1952: out = 16'(-2546);
			1953: out = 16'(-1766);
			1954: out = 16'(14898);
			1955: out = 16'(-2117);
			1956: out = 16'(-3740);
			1957: out = 16'(14980);
			1958: out = 16'(-4838);
			1959: out = 16'(-9747);
			1960: out = 16'(10448);
			1961: out = 16'(-9162);
			1962: out = 16'(-7229);
			1963: out = 16'(13290);
			1964: out = 16'(-12686);
			1965: out = 16'(14971);
			1966: out = 16'(10045);
			1967: out = 16'(-3564);
			1968: out = 16'(13621);
			1969: out = 16'(11228);
			1970: out = 16'(-6489);
			1971: out = 16'(15314);
			1972: out = 16'(-7527);
			1973: out = 16'(10113);
			1974: out = 16'(2279);
			1975: out = 16'(-2947);
			1976: out = 16'(8837);
			1977: out = 16'(-17407);
			1978: out = 16'(7445);
			1979: out = 16'(-15568);
			1980: out = 16'(-19243);
			1981: out = 16'(-13088);
			1982: out = 16'(-2095);
			1983: out = 16'(-6002);
			1984: out = 16'(-11564);
			1985: out = 16'(-17605);
			1986: out = 16'(-2746);
			1987: out = 16'(-5457);
			1988: out = 16'(15523);
			1989: out = 16'(-3588);
			1990: out = 16'(1631);
			1991: out = 16'(-12195);
			1992: out = 16'(8382);
			1993: out = 16'(-10013);
			1994: out = 16'(9891);
			1995: out = 16'(5150);
			1996: out = 16'(2026);
			1997: out = 16'(761);
			1998: out = 16'(-8479);
			1999: out = 16'(3980);
			2000: out = 16'(-7611);
			2001: out = 16'(15103);
			2002: out = 16'(9520);
			2003: out = 16'(4484);
			2004: out = 16'(-3710);
			2005: out = 16'(20879);
			2006: out = 16'(-11631);
			2007: out = 16'(17779);
			2008: out = 16'(-532);
			2009: out = 16'(1549);
			2010: out = 16'(26780);
			2011: out = 16'(-11026);
			2012: out = 16'(3165);
			2013: out = 16'(2976);
			2014: out = 16'(-22742);
			2015: out = 16'(7784);
			2016: out = 16'(-4480);
			2017: out = 16'(16585);
			2018: out = 16'(238);
			2019: out = 16'(-918);
			2020: out = 16'(5938);
			2021: out = 16'(7100);
			2022: out = 16'(9269);
			2023: out = 16'(749);
			2024: out = 16'(14993);
			2025: out = 16'(2049);
			2026: out = 16'(14643);
			2027: out = 16'(-7145);
			2028: out = 16'(1570);
			2029: out = 16'(8173);
			2030: out = 16'(-7272);
			2031: out = 16'(2992);
			2032: out = 16'(-12876);
			2033: out = 16'(-174);
			2034: out = 16'(-830);
			2035: out = 16'(-2685);
			2036: out = 16'(7052);
			2037: out = 16'(-23475);
			2038: out = 16'(5280);
			2039: out = 16'(-10778);
			2040: out = 16'(3668);
			2041: out = 16'(-8648);
			2042: out = 16'(-14079);
			2043: out = 16'(-8171);
			2044: out = 16'(12437);
			2045: out = 16'(12070);
			2046: out = 16'(-13680);
			2047: out = 16'(13087);
			2048: out = 16'(-8333);
			2049: out = 16'(4194);
			2050: out = 16'(-13414);
			2051: out = 16'(6576);
			2052: out = 16'(399);
			2053: out = 16'(-2207);
			2054: out = 16'(4624);
			2055: out = 16'(-2492);
			2056: out = 16'(-117);
			2057: out = 16'(17791);
			2058: out = 16'(-18517);
			2059: out = 16'(5109);
			2060: out = 16'(-1896);
			2061: out = 16'(-10877);
			2062: out = 16'(16889);
			2063: out = 16'(6384);
			2064: out = 16'(6504);
			2065: out = 16'(-6175);
			2066: out = 16'(-2247);
			2067: out = 16'(5201);
			2068: out = 16'(-1263);
			2069: out = 16'(-7967);
			2070: out = 16'(4219);
			2071: out = 16'(-10980);
			2072: out = 16'(13731);
			2073: out = 16'(-6680);
			2074: out = 16'(3475);
			2075: out = 16'(1076);
			2076: out = 16'(5708);
			2077: out = 16'(-4521);
			2078: out = 16'(-8335);
			2079: out = 16'(7586);
			2080: out = 16'(-13170);
			2081: out = 16'(2524);
			2082: out = 16'(-1586);
			2083: out = 16'(14947);
			2084: out = 16'(-10669);
			2085: out = 16'(766);
			2086: out = 16'(-11628);
			2087: out = 16'(4926);
			2088: out = 16'(-5388);
			2089: out = 16'(3741);
			2090: out = 16'(1968);
			2091: out = 16'(10558);
			2092: out = 16'(12968);
			2093: out = 16'(5599);
			2094: out = 16'(-10688);
			2095: out = 16'(1482);
			2096: out = 16'(15141);
			2097: out = 16'(-6927);
			2098: out = 16'(7264);
			2099: out = 16'(1085);
			2100: out = 16'(5362);
			2101: out = 16'(12768);
			2102: out = 16'(-4014);
			2103: out = 16'(1485);
			2104: out = 16'(-1127);
			2105: out = 16'(-601);
			2106: out = 16'(3098);
			2107: out = 16'(-683);
			2108: out = 16'(946);
			2109: out = 16'(-4884);
			2110: out = 16'(4324);
			2111: out = 16'(-1207);
			2112: out = 16'(6389);
			2113: out = 16'(-2293);
			2114: out = 16'(898);
			2115: out = 16'(-4513);
			2116: out = 16'(-4371);
			2117: out = 16'(8924);
			2118: out = 16'(-23413);
			2119: out = 16'(11687);
			2120: out = 16'(-1610);
			2121: out = 16'(-4790);
			2122: out = 16'(1416);
			2123: out = 16'(-3761);
			2124: out = 16'(8494);
			2125: out = 16'(15757);
			2126: out = 16'(3086);
			2127: out = 16'(1548);
			2128: out = 16'(14805);
			2129: out = 16'(-4336);
			2130: out = 16'(4008);
			2131: out = 16'(708);
			2132: out = 16'(-17867);
			2133: out = 16'(15685);
			2134: out = 16'(8565);
			2135: out = 16'(23212);
			2136: out = 16'(-11680);
			2137: out = 16'(9023);
			2138: out = 16'(-12593);
			2139: out = 16'(-8928);
			2140: out = 16'(9232);
			2141: out = 16'(-7551);
			2142: out = 16'(2976);
			2143: out = 16'(-1285);
			2144: out = 16'(-13601);
			2145: out = 16'(13637);
			2146: out = 16'(9315);
			2147: out = 16'(-11946);
			2148: out = 16'(12637);
			2149: out = 16'(1635);
			2150: out = 16'(-23576);
			2151: out = 16'(970);
			2152: out = 16'(13569);
			2153: out = 16'(-3126);
			2154: out = 16'(885);
			2155: out = 16'(-18468);
			2156: out = 16'(-7878);
			2157: out = 16'(1720);
			2158: out = 16'(5470);
			2159: out = 16'(2598);
			2160: out = 16'(-9600);
			2161: out = 16'(12516);
			2162: out = 16'(-5271);
			2163: out = 16'(5446);
			2164: out = 16'(7655);
			2165: out = 16'(2229);
			2166: out = 16'(-22660);
			2167: out = 16'(12874);
			2168: out = 16'(-16282);
			2169: out = 16'(10433);
			2170: out = 16'(10968);
			2171: out = 16'(-5392);
			2172: out = 16'(6082);
			2173: out = 16'(-13732);
			2174: out = 16'(-3069);
			2175: out = 16'(-15460);
			2176: out = 16'(7580);
			2177: out = 16'(8106);
			2178: out = 16'(-23443);
			2179: out = 16'(1461);
			2180: out = 16'(10110);
			2181: out = 16'(-13212);
			2182: out = 16'(13718);
			2183: out = 16'(-5369);
			2184: out = 16'(-1675);
			2185: out = 16'(3184);
			2186: out = 16'(13038);
			2187: out = 16'(4756);
			2188: out = 16'(7568);
			2189: out = 16'(-7863);
			2190: out = 16'(-331);
			2191: out = 16'(-3113);
			2192: out = 16'(5064);
			2193: out = 16'(420);
			2194: out = 16'(-978);
			2195: out = 16'(7488);
			2196: out = 16'(9368);
			2197: out = 16'(-1403);
			2198: out = 16'(4679);
			2199: out = 16'(-10428);
			2200: out = 16'(875);
			2201: out = 16'(6871);
			2202: out = 16'(2110);
			2203: out = 16'(-3602);
			2204: out = 16'(453);
			2205: out = 16'(-2345);
			2206: out = 16'(-14628);
			2207: out = 16'(3758);
			2208: out = 16'(12261);
			2209: out = 16'(7459);
			2210: out = 16'(-3873);
			2211: out = 16'(-10472);
			2212: out = 16'(-7780);
			2213: out = 16'(414);
			2214: out = 16'(9326);
			2215: out = 16'(-2482);
			2216: out = 16'(8363);
			2217: out = 16'(2138);
			2218: out = 16'(-10113);
			2219: out = 16'(14042);
			2220: out = 16'(-17705);
			2221: out = 16'(-3444);
			2222: out = 16'(12533);
			2223: out = 16'(-1136);
			2224: out = 16'(20407);
			2225: out = 16'(10078);
			2226: out = 16'(3907);
			2227: out = 16'(-9818);
			2228: out = 16'(1656);
			2229: out = 16'(-5723);
			2230: out = 16'(3193);
			2231: out = 16'(4500);
			2232: out = 16'(11504);
			2233: out = 16'(-1178);
			2234: out = 16'(6066);
			2235: out = 16'(-2616);
			2236: out = 16'(-4743);
			2237: out = 16'(-3285);
			2238: out = 16'(5127);
			2239: out = 16'(-8131);
			2240: out = 16'(13626);
			2241: out = 16'(-6144);
			2242: out = 16'(-12957);
			2243: out = 16'(16457);
			2244: out = 16'(-4495);
			2245: out = 16'(-3192);
			2246: out = 16'(-9580);
			2247: out = 16'(-8707);
			2248: out = 16'(-2319);
			2249: out = 16'(-10215);
			2250: out = 16'(2402);
			2251: out = 16'(4534);
			2252: out = 16'(8386);
			2253: out = 16'(6022);
			2254: out = 16'(1536);
			2255: out = 16'(-7371);
			2256: out = 16'(-12518);
			2257: out = 16'(1010);
			2258: out = 16'(-8548);
			2259: out = 16'(11517);
			2260: out = 16'(2307);
			2261: out = 16'(10420);
			2262: out = 16'(-1093);
			2263: out = 16'(-10525);
			2264: out = 16'(11600);
			2265: out = 16'(-7082);
			2266: out = 16'(17129);
			2267: out = 16'(10075);
			2268: out = 16'(10838);
			2269: out = 16'(-5588);
			2270: out = 16'(8071);
			2271: out = 16'(-6387);
			2272: out = 16'(13192);
			2273: out = 16'(-4604);
			2274: out = 16'(441);
			2275: out = 16'(9156);
			2276: out = 16'(-1194);
			2277: out = 16'(5111);
			2278: out = 16'(-16067);
			2279: out = 16'(12036);
			2280: out = 16'(-5770);
			2281: out = 16'(4229);
			2282: out = 16'(359);
			2283: out = 16'(-11362);
			2284: out = 16'(252);
			2285: out = 16'(-1325);
			2286: out = 16'(-5480);
			2287: out = 16'(10023);
			2288: out = 16'(197);
			2289: out = 16'(-4995);
			2290: out = 16'(62);
			2291: out = 16'(2863);
			2292: out = 16'(-10295);
			2293: out = 16'(8147);
			2294: out = 16'(3936);
			2295: out = 16'(11830);
			2296: out = 16'(20777);
			2297: out = 16'(-20242);
			2298: out = 16'(-6158);
			2299: out = 16'(-7530);
			2300: out = 16'(277);
			2301: out = 16'(-5870);
			2302: out = 16'(8006);
			2303: out = 16'(4188);
			2304: out = 16'(12538);
			2305: out = 16'(11913);
			2306: out = 16'(2089);
			2307: out = 16'(-6356);
			2308: out = 16'(-12910);
			2309: out = 16'(1111);
			2310: out = 16'(-7909);
			2311: out = 16'(4941);
			2312: out = 16'(14313);
			2313: out = 16'(-8416);
			2314: out = 16'(4946);
			2315: out = 16'(2120);
			2316: out = 16'(-13799);
			2317: out = 16'(13688);
			2318: out = 16'(-8867);
			2319: out = 16'(-259);
			2320: out = 16'(-8599);
			2321: out = 16'(-1274);
			2322: out = 16'(7779);
			2323: out = 16'(11094);
			2324: out = 16'(-342);
			2325: out = 16'(-1834);
			2326: out = 16'(-5595);
			2327: out = 16'(7793);
			2328: out = 16'(-10795);
			2329: out = 16'(9111);
			2330: out = 16'(-8752);
			2331: out = 16'(10866);
			2332: out = 16'(16);
			2333: out = 16'(-12058);
			2334: out = 16'(5875);
			2335: out = 16'(-11005);
			2336: out = 16'(1487);
			2337: out = 16'(-11005);
			2338: out = 16'(2069);
			2339: out = 16'(7922);
			2340: out = 16'(1784);
			2341: out = 16'(3528);
			2342: out = 16'(85);
			2343: out = 16'(11787);
			2344: out = 16'(-7137);
			2345: out = 16'(-3970);
			2346: out = 16'(5255);
			2347: out = 16'(-3855);
			2348: out = 16'(8288);
			2349: out = 16'(-1733);
			2350: out = 16'(10167);
			2351: out = 16'(3022);
			2352: out = 16'(-4942);
			2353: out = 16'(2173);
			2354: out = 16'(14302);
			2355: out = 16'(-1392);
			2356: out = 16'(9018);
			2357: out = 16'(7322);
			2358: out = 16'(12740);
			2359: out = 16'(14132);
			2360: out = 16'(-4743);
			2361: out = 16'(3755);
			2362: out = 16'(8363);
			2363: out = 16'(5931);
			2364: out = 16'(-311);
			2365: out = 16'(2079);
			2366: out = 16'(2211);
			2367: out = 16'(1810);
			2368: out = 16'(8776);
			2369: out = 16'(-8287);
			2370: out = 16'(16590);
			2371: out = 16'(-1274);
			2372: out = 16'(-17631);
			2373: out = 16'(-1490);
			2374: out = 16'(-4052);
			2375: out = 16'(6717);
			2376: out = 16'(1382);
			2377: out = 16'(-7312);
			2378: out = 16'(-769);
			2379: out = 16'(-6164);
			2380: out = 16'(2942);
			2381: out = 16'(-3800);
			2382: out = 16'(5935);
			2383: out = 16'(-7606);
			2384: out = 16'(7002);
			2385: out = 16'(1237);
			2386: out = 16'(8387);
			2387: out = 16'(2157);
			2388: out = 16'(39);
			2389: out = 16'(-6876);
			2390: out = 16'(-12512);
			2391: out = 16'(7131);
			2392: out = 16'(-3005);
			2393: out = 16'(13883);
			2394: out = 16'(3981);
			2395: out = 16'(1418);
			2396: out = 16'(6875);
			2397: out = 16'(-798);
			2398: out = 16'(7881);
			2399: out = 16'(3494);
			2400: out = 16'(5740);
			2401: out = 16'(-2527);
			2402: out = 16'(423);
			2403: out = 16'(2978);
			2404: out = 16'(-471);
			2405: out = 16'(4);
			2406: out = 16'(852);
			2407: out = 16'(13496);
			2408: out = 16'(8089);
			2409: out = 16'(1213);
			2410: out = 16'(11658);
			2411: out = 16'(-11304);
			2412: out = 16'(6770);
			2413: out = 16'(-8014);
			2414: out = 16'(7252);
			2415: out = 16'(-2545);
			2416: out = 16'(-26);
			2417: out = 16'(-9884);
			2418: out = 16'(3865);
			2419: out = 16'(-1524);
			2420: out = 16'(9194);
			2421: out = 16'(-776);
			2422: out = 16'(13189);
			2423: out = 16'(-1321);
			2424: out = 16'(-15072);
			2425: out = 16'(358);
			2426: out = 16'(5206);
			2427: out = 16'(8376);
			2428: out = 16'(-491);
			2429: out = 16'(7006);
			2430: out = 16'(8248);
			2431: out = 16'(5805);
			2432: out = 16'(501);
			2433: out = 16'(-23318);
			2434: out = 16'(5360);
			2435: out = 16'(6023);
			2436: out = 16'(-2310);
			2437: out = 16'(13400);
			2438: out = 16'(-7182);
			2439: out = 16'(-777);
			2440: out = 16'(697);
			2441: out = 16'(-1636);
			2442: out = 16'(8469);
			2443: out = 16'(-438);
			2444: out = 16'(8210);
			2445: out = 16'(4273);
			2446: out = 16'(5985);
			2447: out = 16'(6805);
			2448: out = 16'(-9354);
			2449: out = 16'(-11391);
			2450: out = 16'(4012);
			2451: out = 16'(-11631);
			2452: out = 16'(-339);
			2453: out = 16'(-62);
			2454: out = 16'(-4779);
			2455: out = 16'(8456);
			2456: out = 16'(-765);
			2457: out = 16'(-3088);
			2458: out = 16'(4575);
			2459: out = 16'(11505);
			2460: out = 16'(-16959);
			2461: out = 16'(5848);
			2462: out = 16'(9820);
			2463: out = 16'(6586);
			2464: out = 16'(21067);
			2465: out = 16'(7324);
			2466: out = 16'(6794);
			2467: out = 16'(-18659);
			2468: out = 16'(7945);
			2469: out = 16'(-3154);
			2470: out = 16'(-5316);
			2471: out = 16'(17163);
			2472: out = 16'(7881);
			2473: out = 16'(9839);
			2474: out = 16'(8553);
			2475: out = 16'(-6623);
			2476: out = 16'(-8565);
			2477: out = 16'(-6997);
			2478: out = 16'(1886);
			2479: out = 16'(7246);
			2480: out = 16'(243);
			2481: out = 16'(8519);
			2482: out = 16'(-7170);
			2483: out = 16'(2565);
			2484: out = 16'(10513);
			2485: out = 16'(-3855);
			2486: out = 16'(3353);
			2487: out = 16'(11039);
			2488: out = 16'(-5154);
			2489: out = 16'(-3859);
			2490: out = 16'(-3082);
			2491: out = 16'(3020);
			2492: out = 16'(-571);
			2493: out = 16'(-14971);
			2494: out = 16'(2012);
			2495: out = 16'(-27479);
			2496: out = 16'(11913);
			2497: out = 16'(8132);
			2498: out = 16'(546);
			2499: out = 16'(16387);
			2500: out = 16'(-405);
			2501: out = 16'(4547);
			2502: out = 16'(1912);
			2503: out = 16'(6668);
			2504: out = 16'(-24024);
			2505: out = 16'(11627);
			2506: out = 16'(-4337);
			2507: out = 16'(-445);
			2508: out = 16'(6772);
			2509: out = 16'(-5427);
			2510: out = 16'(2684);
			2511: out = 16'(2903);
			2512: out = 16'(-8607);
			2513: out = 16'(11937);
			2514: out = 16'(-7361);
			2515: out = 16'(6403);
			2516: out = 16'(7098);
			2517: out = 16'(-10192);
			2518: out = 16'(13407);
			2519: out = 16'(-4462);
			2520: out = 16'(-3787);
			2521: out = 16'(-9506);
			2522: out = 16'(-2496);
			2523: out = 16'(1679);
			2524: out = 16'(-699);
			2525: out = 16'(5572);
			2526: out = 16'(16827);
			2527: out = 16'(-5816);
			2528: out = 16'(3011);
			2529: out = 16'(-1759);
			2530: out = 16'(-5642);
			2531: out = 16'(-5022);
			2532: out = 16'(2443);
			2533: out = 16'(-5320);
			2534: out = 16'(8339);
			2535: out = 16'(-3032);
			2536: out = 16'(1357);
			2537: out = 16'(9508);
			2538: out = 16'(-9743);
			2539: out = 16'(3319);
			2540: out = 16'(-17490);
			2541: out = 16'(1090);
			2542: out = 16'(-2500);
			2543: out = 16'(-643);
			2544: out = 16'(10185);
			2545: out = 16'(-5172);
			2546: out = 16'(-16305);
			2547: out = 16'(5120);
			2548: out = 16'(912);
			2549: out = 16'(-8690);
			2550: out = 16'(12398);
			2551: out = 16'(-10708);
			2552: out = 16'(-577);
			2553: out = 16'(128);
			2554: out = 16'(3446);
			2555: out = 16'(5477);
			2556: out = 16'(-2865);
			2557: out = 16'(7667);
			2558: out = 16'(-14076);
			2559: out = 16'(5000);
			2560: out = 16'(-69);
			2561: out = 16'(-6517);
			2562: out = 16'(5178);
			2563: out = 16'(127);
			2564: out = 16'(8635);
			2565: out = 16'(-1267);
			2566: out = 16'(2085);
			2567: out = 16'(7963);
			2568: out = 16'(10309);
			2569: out = 16'(2398);
			2570: out = 16'(-729);
			2571: out = 16'(3139);
			2572: out = 16'(8346);
			2573: out = 16'(3621);
			2574: out = 16'(-615);
			2575: out = 16'(1050);
			2576: out = 16'(4706);
			2577: out = 16'(-16897);
			2578: out = 16'(5046);
			2579: out = 16'(-8650);
			2580: out = 16'(603);
			2581: out = 16'(4612);
			2582: out = 16'(-591);
			2583: out = 16'(-13014);
			2584: out = 16'(6196);
			2585: out = 16'(1940);
			2586: out = 16'(-2294);
			2587: out = 16'(18268);
			2588: out = 16'(-4535);
			2589: out = 16'(3292);
			2590: out = 16'(135);
			2591: out = 16'(-2795);
			2592: out = 16'(-946);
			2593: out = 16'(719);
			2594: out = 16'(12580);
			2595: out = 16'(-20874);
			2596: out = 16'(4151);
			2597: out = 16'(659);
			2598: out = 16'(-14505);
			2599: out = 16'(5434);
			2600: out = 16'(-1609);
			2601: out = 16'(-7185);
			2602: out = 16'(8123);
			2603: out = 16'(-6495);
			2604: out = 16'(-14183);
			2605: out = 16'(-15987);
			2606: out = 16'(15489);
			2607: out = 16'(-13498);
			2608: out = 16'(150);
			2609: out = 16'(12661);
			2610: out = 16'(-14779);
			2611: out = 16'(2539);
			2612: out = 16'(1227);
			2613: out = 16'(-407);
			2614: out = 16'(-904);
			2615: out = 16'(-1684);
			2616: out = 16'(-12120);
			2617: out = 16'(-10889);
			2618: out = 16'(9044);
			2619: out = 16'(4696);
			2620: out = 16'(-11564);
			2621: out = 16'(17465);
			2622: out = 16'(-14284);
			2623: out = 16'(-3243);
			2624: out = 16'(1292);
			2625: out = 16'(-14530);
			2626: out = 16'(5457);
			2627: out = 16'(-2792);
			2628: out = 16'(6528);
			2629: out = 16'(512);
			2630: out = 16'(1854);
			2631: out = 16'(7363);
			2632: out = 16'(-5939);
			2633: out = 16'(-834);
			2634: out = 16'(6023);
			2635: out = 16'(-6476);
			2636: out = 16'(11012);
			2637: out = 16'(-7745);
			2638: out = 16'(2938);
			2639: out = 16'(3130);
			2640: out = 16'(-4910);
			2641: out = 16'(927);
			2642: out = 16'(-360);
			2643: out = 16'(-987);
			2644: out = 16'(-10895);
			2645: out = 16'(8870);
			2646: out = 16'(8630);
			2647: out = 16'(1889);
			2648: out = 16'(2221);
			2649: out = 16'(-10906);
			2650: out = 16'(-1387);
			2651: out = 16'(-16629);
			2652: out = 16'(-7698);
			2653: out = 16'(4362);
			2654: out = 16'(-242);
			2655: out = 16'(11172);
			2656: out = 16'(-3187);
			2657: out = 16'(1007);
			2658: out = 16'(7533);
			2659: out = 16'(4441);
			2660: out = 16'(-3218);
			2661: out = 16'(-4100);
			2662: out = 16'(-5911);
			2663: out = 16'(-231);
			2664: out = 16'(-1719);
			2665: out = 16'(5232);
			2666: out = 16'(-872);
			2667: out = 16'(16981);
			2668: out = 16'(10474);
			2669: out = 16'(4388);
			2670: out = 16'(18291);
			2671: out = 16'(-1354);
			2672: out = 16'(-5228);
			2673: out = 16'(18643);
			2674: out = 16'(1600);
			2675: out = 16'(8929);
			2676: out = 16'(354);
			2677: out = 16'(1462);
			2678: out = 16'(6949);
			2679: out = 16'(-12222);
			2680: out = 16'(-546);
			2681: out = 16'(-312);
			2682: out = 16'(6719);
			2683: out = 16'(-3172);
			2684: out = 16'(2036);
			2685: out = 16'(434);
			2686: out = 16'(-1286);
			2687: out = 16'(-1057);
			2688: out = 16'(-3559);
			2689: out = 16'(1536);
			2690: out = 16'(1364);
			2691: out = 16'(-4243);
			2692: out = 16'(-2976);
			2693: out = 16'(1382);
			2694: out = 16'(2255);
			2695: out = 16'(5014);
			2696: out = 16'(3617);
			2697: out = 16'(7566);
			2698: out = 16'(1251);
			2699: out = 16'(-6982);
			2700: out = 16'(-201);
			2701: out = 16'(-1036);
			2702: out = 16'(-406);
			2703: out = 16'(-5217);
			2704: out = 16'(1872);
			2705: out = 16'(9547);
			2706: out = 16'(-12569);
			2707: out = 16'(-492);
			2708: out = 16'(-6560);
			2709: out = 16'(8639);
			2710: out = 16'(6443);
			2711: out = 16'(-6035);
			2712: out = 16'(-10809);
			2713: out = 16'(-19226);
			2714: out = 16'(5226);
			2715: out = 16'(3006);
			2716: out = 16'(2593);
			2717: out = 16'(6932);
			2718: out = 16'(-1080);
			2719: out = 16'(-4385);
			2720: out = 16'(1078);
			2721: out = 16'(3140);
			2722: out = 16'(1589);
			2723: out = 16'(678);
			2724: out = 16'(489);
			2725: out = 16'(-1556);
			2726: out = 16'(-385);
			2727: out = 16'(3295);
			2728: out = 16'(1734);
			2729: out = 16'(1806);
			2730: out = 16'(-7535);
			2731: out = 16'(455);
			2732: out = 16'(2305);
			2733: out = 16'(-801);
			2734: out = 16'(-5424);
			2735: out = 16'(3002);
			2736: out = 16'(12801);
			2737: out = 16'(1483);
			2738: out = 16'(-1525);
			2739: out = 16'(8960);
			2740: out = 16'(-4524);
			2741: out = 16'(12179);
			2742: out = 16'(1741);
			2743: out = 16'(4372);
			2744: out = 16'(5114);
			2745: out = 16'(-9958);
			2746: out = 16'(-104);
			2747: out = 16'(-2290);
			2748: out = 16'(7319);
			2749: out = 16'(9296);
			2750: out = 16'(356);
			2751: out = 16'(3176);
			2752: out = 16'(1667);
			2753: out = 16'(2278);
			2754: out = 16'(12772);
			2755: out = 16'(-4300);
			2756: out = 16'(402);
			2757: out = 16'(-5613);
			2758: out = 16'(-645);
			2759: out = 16'(13955);
			2760: out = 16'(1571);
			2761: out = 16'(8395);
			2762: out = 16'(14268);
			2763: out = 16'(-700);
			2764: out = 16'(783);
			2765: out = 16'(-1157);
			2766: out = 16'(-4871);
			2767: out = 16'(8825);
			2768: out = 16'(9072);
			2769: out = 16'(10042);
			2770: out = 16'(-8609);
			2771: out = 16'(9755);
			2772: out = 16'(-4930);
			2773: out = 16'(-3471);
			2774: out = 16'(-910);
			2775: out = 16'(691);
			2776: out = 16'(2563);
			2777: out = 16'(2912);
			2778: out = 16'(3878);
			2779: out = 16'(2246);
			2780: out = 16'(1995);
			2781: out = 16'(-4714);
			2782: out = 16'(-10851);
			2783: out = 16'(6183);
			2784: out = 16'(-6068);
			2785: out = 16'(-303);
			2786: out = 16'(-937);
			2787: out = 16'(-5740);
			2788: out = 16'(11673);
			2789: out = 16'(-624);
			2790: out = 16'(8264);
			2791: out = 16'(12337);
			2792: out = 16'(6123);
			2793: out = 16'(10762);
			2794: out = 16'(-386);
			2795: out = 16'(-519);
			2796: out = 16'(9470);
			2797: out = 16'(5122);
			2798: out = 16'(8937);
			2799: out = 16'(-93);
			2800: out = 16'(-5544);
			2801: out = 16'(6587);
			2802: out = 16'(-3438);
			2803: out = 16'(6972);
			2804: out = 16'(-6516);
			2805: out = 16'(-2042);
			2806: out = 16'(4535);
			2807: out = 16'(-4147);
			2808: out = 16'(-5586);
			2809: out = 16'(-11939);
			2810: out = 16'(1488);
			2811: out = 16'(6146);
			2812: out = 16'(-4410);
			2813: out = 16'(-173);
			2814: out = 16'(-6065);
			2815: out = 16'(2214);
			2816: out = 16'(-14355);
			2817: out = 16'(962);
			2818: out = 16'(1880);
			2819: out = 16'(6238);
			2820: out = 16'(152);
			2821: out = 16'(408);
			2822: out = 16'(2098);
			2823: out = 16'(-4336);
			2824: out = 16'(-7210);
			2825: out = 16'(1993);
			2826: out = 16'(-3766);
			2827: out = 16'(7195);
			2828: out = 16'(643);
			2829: out = 16'(-12454);
			2830: out = 16'(4425);
			2831: out = 16'(-5582);
			2832: out = 16'(-11715);
			2833: out = 16'(12890);
			2834: out = 16'(-16428);
			2835: out = 16'(480);
			2836: out = 16'(17857);
			2837: out = 16'(9667);
			2838: out = 16'(12123);
			2839: out = 16'(-17933);
			2840: out = 16'(7537);
			2841: out = 16'(-11810);
			2842: out = 16'(-12987);
			2843: out = 16'(7099);
			2844: out = 16'(-7860);
			2845: out = 16'(7160);
			2846: out = 16'(9150);
			2847: out = 16'(-27978);
			2848: out = 16'(7579);
			2849: out = 16'(12744);
			2850: out = 16'(-8403);
			2851: out = 16'(-8651);
			2852: out = 16'(-5498);
			2853: out = 16'(-869);
			2854: out = 16'(-4901);
			2855: out = 16'(8385);
			2856: out = 16'(11671);
			2857: out = 16'(-7221);
			2858: out = 16'(12972);
			2859: out = 16'(-5434);
			2860: out = 16'(-7249);
			2861: out = 16'(11747);
			2862: out = 16'(13476);
			2863: out = 16'(-966);
			2864: out = 16'(11447);
			2865: out = 16'(-3572);
			2866: out = 16'(-21030);
			2867: out = 16'(18904);
			2868: out = 16'(-11685);
			2869: out = 16'(4001);
			2870: out = 16'(11855);
			2871: out = 16'(-3337);
			2872: out = 16'(3903);
			2873: out = 16'(-13626);
			2874: out = 16'(10023);
			2875: out = 16'(-7025);
			2876: out = 16'(-5008);
			2877: out = 16'(12782);
			2878: out = 16'(-13298);
			2879: out = 16'(371);
			2880: out = 16'(-157);
			2881: out = 16'(-6249);
			2882: out = 16'(-3228);
			2883: out = 16'(4261);
			2884: out = 16'(4660);
			2885: out = 16'(6854);
			2886: out = 16'(7719);
			2887: out = 16'(13077);
			2888: out = 16'(13197);
			2889: out = 16'(12500);
			2890: out = 16'(-1165);
			2891: out = 16'(-5080);
			2892: out = 16'(13183);
			2893: out = 16'(-3858);
			2894: out = 16'(16678);
			2895: out = 16'(-6423);
			2896: out = 16'(9765);
			2897: out = 16'(-4671);
			2898: out = 16'(9969);
			2899: out = 16'(4104);
			2900: out = 16'(-2759);
			2901: out = 16'(11398);
			2902: out = 16'(-11539);
			2903: out = 16'(7578);
			2904: out = 16'(-2656);
			2905: out = 16'(-1712);
			2906: out = 16'(7383);
			2907: out = 16'(7797);
			2908: out = 16'(1579);
			2909: out = 16'(-2898);
			2910: out = 16'(-4827);
			2911: out = 16'(-1243);
			2912: out = 16'(3859);
			2913: out = 16'(-10247);
			2914: out = 16'(8463);
			2915: out = 16'(5946);
			2916: out = 16'(-14307);
			2917: out = 16'(-8877);
			2918: out = 16'(-15492);
			2919: out = 16'(9845);
			2920: out = 16'(-13361);
			2921: out = 16'(1817);
			2922: out = 16'(-3302);
			2923: out = 16'(-7715);
			2924: out = 16'(13405);
			2925: out = 16'(-13844);
			2926: out = 16'(6315);
			2927: out = 16'(-11585);
			2928: out = 16'(4794);
			2929: out = 16'(-7408);
			2930: out = 16'(10293);
			2931: out = 16'(-4286);
			2932: out = 16'(-5825);
			2933: out = 16'(6205);
			2934: out = 16'(-6258);
			2935: out = 16'(2895);
			2936: out = 16'(-508);
			2937: out = 16'(1528);
			2938: out = 16'(3987);
			2939: out = 16'(-231);
			2940: out = 16'(-493);
			2941: out = 16'(-4784);
			2942: out = 16'(1315);
			2943: out = 16'(1350);
			2944: out = 16'(9809);
			2945: out = 16'(8466);
			2946: out = 16'(6671);
			2947: out = 16'(-11473);
			2948: out = 16'(-9089);
			2949: out = 16'(11212);
			2950: out = 16'(-13199);
			2951: out = 16'(18204);
			2952: out = 16'(-20590);
			2953: out = 16'(6141);
			2954: out = 16'(-13067);
			2955: out = 16'(-10668);
			2956: out = 16'(14147);
			2957: out = 16'(-12070);
			2958: out = 16'(9738);
			2959: out = 16'(-27670);
			2960: out = 16'(-12428);
			2961: out = 16'(-9831);
			2962: out = 16'(-6902);
			2963: out = 16'(7264);
			2964: out = 16'(-5404);
			2965: out = 16'(5272);
			2966: out = 16'(7538);
			2967: out = 16'(-3126);
			2968: out = 16'(-11132);
			2969: out = 16'(1);
			2970: out = 16'(-4466);
			2971: out = 16'(-1258);
			2972: out = 16'(12332);
			2973: out = 16'(-16281);
			2974: out = 16'(13981);
			2975: out = 16'(-1726);
			2976: out = 16'(9931);
			2977: out = 16'(-7420);
			2978: out = 16'(4270);
			2979: out = 16'(-1337);
			2980: out = 16'(-1338);
			2981: out = 16'(-1372);
			2982: out = 16'(8203);
			2983: out = 16'(7252);
			2984: out = 16'(-4777);
			2985: out = 16'(4595);
			2986: out = 16'(1798);
			2987: out = 16'(10607);
			2988: out = 16'(6989);
			2989: out = 16'(-8102);
			2990: out = 16'(1702);
			2991: out = 16'(6086);
			2992: out = 16'(-6786);
			2993: out = 16'(1152);
			2994: out = 16'(4647);
			2995: out = 16'(892);
			2996: out = 16'(-4502);
			2997: out = 16'(-3968);
			2998: out = 16'(-1823);
			2999: out = 16'(3560);
			3000: out = 16'(-253);
			3001: out = 16'(2917);
			3002: out = 16'(5779);
			3003: out = 16'(7961);
			3004: out = 16'(-13400);
			3005: out = 16'(-5755);
			3006: out = 16'(-5970);
			3007: out = 16'(9224);
			3008: out = 16'(2972);
			3009: out = 16'(108);
			3010: out = 16'(10358);
			3011: out = 16'(-19837);
			3012: out = 16'(529);
			3013: out = 16'(-695);
			3014: out = 16'(11333);
			3015: out = 16'(11522);
			3016: out = 16'(13208);
			3017: out = 16'(-10044);
			3018: out = 16'(2405);
			3019: out = 16'(-2481);
			3020: out = 16'(-2150);
			3021: out = 16'(8904);
			3022: out = 16'(-4614);
			3023: out = 16'(1622);
			3024: out = 16'(256);
			3025: out = 16'(3906);
			3026: out = 16'(-1565);
			3027: out = 16'(18518);
			3028: out = 16'(-2475);
			3029: out = 16'(3448);
			3030: out = 16'(5884);
			3031: out = 16'(-3545);
			3032: out = 16'(7228);
			3033: out = 16'(6281);
			3034: out = 16'(7687);
			3035: out = 16'(5615);
			3036: out = 16'(-12005);
			3037: out = 16'(9939);
			3038: out = 16'(-14284);
			3039: out = 16'(10760);
			3040: out = 16'(2900);
			3041: out = 16'(-5456);
			3042: out = 16'(1527);
			3043: out = 16'(3200);
			3044: out = 16'(-2239);
			3045: out = 16'(-2978);
			3046: out = 16'(2590);
			3047: out = 16'(-8366);
			3048: out = 16'(892);
			3049: out = 16'(-1728);
			3050: out = 16'(-6243);
			3051: out = 16'(232);
			3052: out = 16'(4012);
			3053: out = 16'(1444);
			3054: out = 16'(-6698);
			3055: out = 16'(-13971);
			3056: out = 16'(-7587);
			3057: out = 16'(-7139);
			3058: out = 16'(6313);
			3059: out = 16'(-8053);
			3060: out = 16'(-6890);
			3061: out = 16'(8739);
			3062: out = 16'(-597);
			3063: out = 16'(2386);
			3064: out = 16'(398);
			3065: out = 16'(5140);
			3066: out = 16'(-634);
			3067: out = 16'(-5686);
			3068: out = 16'(-10944);
			3069: out = 16'(2931);
			3070: out = 16'(8252);
			3071: out = 16'(16986);
			3072: out = 16'(-3564);
			3073: out = 16'(-823);
			3074: out = 16'(9289);
			3075: out = 16'(-12957);
			3076: out = 16'(-17365);
			3077: out = 16'(14389);
			3078: out = 16'(-5233);
			3079: out = 16'(2964);
			3080: out = 16'(3108);
			3081: out = 16'(-9939);
			3082: out = 16'(-690);
			3083: out = 16'(1061);
			3084: out = 16'(-8899);
			3085: out = 16'(6562);
			3086: out = 16'(476);
			3087: out = 16'(1588);
			3088: out = 16'(9429);
			3089: out = 16'(-2987);
			3090: out = 16'(-792);
			3091: out = 16'(-3836);
			3092: out = 16'(-1986);
			3093: out = 16'(-12361);
			3094: out = 16'(1861);
			3095: out = 16'(-621);
			3096: out = 16'(9130);
			3097: out = 16'(-7668);
			3098: out = 16'(4602);
			3099: out = 16'(-2855);
			3100: out = 16'(-2886);
			3101: out = 16'(6110);
			3102: out = 16'(5139);
			3103: out = 16'(10797);
			3104: out = 16'(471);
			3105: out = 16'(15125);
			3106: out = 16'(464);
			3107: out = 16'(-11197);
			3108: out = 16'(5341);
			3109: out = 16'(-2462);
			3110: out = 16'(13827);
			3111: out = 16'(-1796);
			3112: out = 16'(1534);
			3113: out = 16'(12546);
			3114: out = 16'(-148);
			3115: out = 16'(7754);
			3116: out = 16'(14768);
			3117: out = 16'(5585);
			3118: out = 16'(1723);
			3119: out = 16'(-2702);
			3120: out = 16'(-1883);
			3121: out = 16'(11694);
			3122: out = 16'(-181);
			3123: out = 16'(-711);
			3124: out = 16'(-12525);
			3125: out = 16'(-9879);
			3126: out = 16'(5116);
			3127: out = 16'(-13985);
			3128: out = 16'(-5469);
			3129: out = 16'(8582);
			3130: out = 16'(-12491);
			3131: out = 16'(-5084);
			3132: out = 16'(6260);
			3133: out = 16'(-3955);
			3134: out = 16'(442);
			3135: out = 16'(-1345);
			3136: out = 16'(1707);
			3137: out = 16'(1990);
			3138: out = 16'(-9346);
			3139: out = 16'(2124);
			3140: out = 16'(11152);
			3141: out = 16'(3679);
			3142: out = 16'(3861);
			3143: out = 16'(-537);
			3144: out = 16'(12578);
			3145: out = 16'(10080);
			3146: out = 16'(-3513);
			3147: out = 16'(-393);
			3148: out = 16'(7176);
			3149: out = 16'(7664);
			3150: out = 16'(-2329);
			3151: out = 16'(5552);
			3152: out = 16'(-1944);
			3153: out = 16'(5955);
			3154: out = 16'(8360);
			3155: out = 16'(7320);
			3156: out = 16'(-24);
			3157: out = 16'(13047);
			3158: out = 16'(577);
			3159: out = 16'(-5974);
			3160: out = 16'(2261);
			3161: out = 16'(-1330);
			3162: out = 16'(-1379);
			3163: out = 16'(7599);
			3164: out = 16'(1252);
			3165: out = 16'(1905);
			3166: out = 16'(-6000);
			3167: out = 16'(-294);
			3168: out = 16'(6556);
			3169: out = 16'(-7679);
			3170: out = 16'(-383);
			3171: out = 16'(-5978);
			3172: out = 16'(13845);
			3173: out = 16'(-1781);
			3174: out = 16'(4604);
			3175: out = 16'(-365);
			3176: out = 16'(456);
			3177: out = 16'(338);
			3178: out = 16'(-473);
			3179: out = 16'(11427);
			3180: out = 16'(-1734);
			3181: out = 16'(9090);
			3182: out = 16'(-1757);
			3183: out = 16'(5931);
			3184: out = 16'(11735);
			3185: out = 16'(4112);
			3186: out = 16'(10434);
			3187: out = 16'(-2948);
			3188: out = 16'(19041);
			3189: out = 16'(-3605);
			3190: out = 16'(-3274);
			3191: out = 16'(4297);
			3192: out = 16'(4318);
			3193: out = 16'(15111);
			3194: out = 16'(7886);
			3195: out = 16'(3365);
			3196: out = 16'(8805);
			3197: out = 16'(-4);
			3198: out = 16'(-2311);
			3199: out = 16'(-355);
			3200: out = 16'(3975);
			3201: out = 16'(-2902);
			3202: out = 16'(2633);
			3203: out = 16'(-684);
			3204: out = 16'(-2355);
			3205: out = 16'(-93);
			3206: out = 16'(7816);
			3207: out = 16'(-4075);
			3208: out = 16'(8456);
			3209: out = 16'(-25160);
			3210: out = 16'(6024);
			3211: out = 16'(2344);
			3212: out = 16'(-9575);
			3213: out = 16'(289);
			3214: out = 16'(-11408);
			3215: out = 16'(1935);
			3216: out = 16'(-117);
			3217: out = 16'(-7523);
			3218: out = 16'(9663);
			3219: out = 16'(-5694);
			3220: out = 16'(7334);
			3221: out = 16'(-3797);
			3222: out = 16'(2865);
			3223: out = 16'(1178);
			3224: out = 16'(7903);
			3225: out = 16'(7357);
			3226: out = 16'(4957);
			3227: out = 16'(2958);
			3228: out = 16'(-10533);
			3229: out = 16'(630);
			3230: out = 16'(19);
			3231: out = 16'(6600);
			3232: out = 16'(-5369);
			3233: out = 16'(4950);
			3234: out = 16'(-1595);
			3235: out = 16'(5362);
			3236: out = 16'(-1675);
			3237: out = 16'(10798);
			3238: out = 16'(2954);
			3239: out = 16'(4690);
			3240: out = 16'(3372);
			3241: out = 16'(-1346);
			3242: out = 16'(-708);
			3243: out = 16'(2426);
			3244: out = 16'(6072);
			3245: out = 16'(2514);
			3246: out = 16'(4383);
			3247: out = 16'(-8792);
			3248: out = 16'(4354);
			3249: out = 16'(365);
			3250: out = 16'(5442);
			3251: out = 16'(-3475);
			3252: out = 16'(-1978);
			3253: out = 16'(691);
			3254: out = 16'(-9783);
			3255: out = 16'(-12387);
			3256: out = 16'(-1950);
			3257: out = 16'(-4054);
			3258: out = 16'(9803);
			3259: out = 16'(9435);
			3260: out = 16'(1155);
			3261: out = 16'(-5588);
			3262: out = 16'(5088);
			3263: out = 16'(-728);
			3264: out = 16'(2333);
			3265: out = 16'(13460);
			3266: out = 16'(1875);
			3267: out = 16'(3711);
			3268: out = 16'(475);
			3269: out = 16'(2889);
			3270: out = 16'(601);
			3271: out = 16'(-621);
			3272: out = 16'(506);
			3273: out = 16'(13107);
			3274: out = 16'(90);
			3275: out = 16'(12018);
			3276: out = 16'(2838);
			3277: out = 16'(17045);
			3278: out = 16'(-8755);
			3279: out = 16'(1070);
			3280: out = 16'(-12811);
			3281: out = 16'(9063);
			3282: out = 16'(-3577);
			3283: out = 16'(7228);
			3284: out = 16'(-4373);
			3285: out = 16'(-2116);
			3286: out = 16'(9534);
			3287: out = 16'(-10302);
			3288: out = 16'(3849);
			3289: out = 16'(7386);
			3290: out = 16'(7240);
			3291: out = 16'(-1018);
			3292: out = 16'(4466);
			3293: out = 16'(-10765);
			3294: out = 16'(6033);
			3295: out = 16'(-4112);
			3296: out = 16'(4774);
			3297: out = 16'(4065);
			3298: out = 16'(2055);
			3299: out = 16'(-1794);
			3300: out = 16'(-12834);
			3301: out = 16'(5691);
			3302: out = 16'(4810);
			3303: out = 16'(-6421);
			3304: out = 16'(4246);
			3305: out = 16'(-6362);
			3306: out = 16'(-2409);
			3307: out = 16'(3430);
			3308: out = 16'(-1170);
			3309: out = 16'(-3854);
			3310: out = 16'(3341);
			3311: out = 16'(8507);
			3312: out = 16'(-18951);
			3313: out = 16'(3799);
			3314: out = 16'(-10416);
			3315: out = 16'(6577);
			3316: out = 16'(-10230);
			3317: out = 16'(10684);
			3318: out = 16'(-6706);
			3319: out = 16'(-5000);
			3320: out = 16'(3813);
			3321: out = 16'(-9093);
			3322: out = 16'(9773);
			3323: out = 16'(-13244);
			3324: out = 16'(7762);
			3325: out = 16'(-8683);
			3326: out = 16'(6716);
			3327: out = 16'(3017);
			3328: out = 16'(-4945);
			3329: out = 16'(4522);
			3330: out = 16'(-9884);
			3331: out = 16'(-1963);
			3332: out = 16'(-8803);
			3333: out = 16'(893);
			3334: out = 16'(-4000);
			3335: out = 16'(-3876);
			3336: out = 16'(-2387);
			3337: out = 16'(-13271);
			3338: out = 16'(11684);
			3339: out = 16'(-10518);
			3340: out = 16'(12909);
			3341: out = 16'(-9181);
			3342: out = 16'(2608);
			3343: out = 16'(2752);
			3344: out = 16'(-10446);
			3345: out = 16'(9971);
			3346: out = 16'(-7673);
			3347: out = 16'(4906);
			3348: out = 16'(1300);
			3349: out = 16'(6785);
			3350: out = 16'(3538);
			3351: out = 16'(-1062);
			3352: out = 16'(-4106);
			3353: out = 16'(3860);
			3354: out = 16'(5299);
			3355: out = 16'(11475);
			3356: out = 16'(40);
			3357: out = 16'(4518);
			3358: out = 16'(-8798);
			3359: out = 16'(11443);
			3360: out = 16'(5606);
			3361: out = 16'(-1359);
			3362: out = 16'(1111);
			3363: out = 16'(249);
			3364: out = 16'(-3303);
			3365: out = 16'(3251);
			3366: out = 16'(2123);
			3367: out = 16'(4315);
			3368: out = 16'(3865);
			3369: out = 16'(-4921);
			3370: out = 16'(2930);
			3371: out = 16'(-11299);
			3372: out = 16'(3601);
			3373: out = 16'(-6388);
			3374: out = 16'(7509);
			3375: out = 16'(-14126);
			3376: out = 16'(10215);
			3377: out = 16'(-8345);
			3378: out = 16'(-4908);
			3379: out = 16'(3259);
			3380: out = 16'(-1716);
			3381: out = 16'(5163);
			3382: out = 16'(1476);
			3383: out = 16'(-7015);
			3384: out = 16'(1905);
			3385: out = 16'(-7159);
			3386: out = 16'(-9430);
			3387: out = 16'(2150);
			3388: out = 16'(1672);
			3389: out = 16'(925);
			3390: out = 16'(-7147);
			3391: out = 16'(3988);
			3392: out = 16'(-12362);
			3393: out = 16'(529);
			3394: out = 16'(-19284);
			3395: out = 16'(11262);
			3396: out = 16'(-9638);
			3397: out = 16'(-4330);
			3398: out = 16'(587);
			3399: out = 16'(-16106);
			3400: out = 16'(14051);
			3401: out = 16'(-4584);
			3402: out = 16'(-6909);
			3403: out = 16'(-16035);
			3404: out = 16'(-486);
			3405: out = 16'(-423);
			3406: out = 16'(-544);
			3407: out = 16'(3347);
			3408: out = 16'(-3216);
			3409: out = 16'(-6532);
			3410: out = 16'(-1739);
			3411: out = 16'(-2870);
			3412: out = 16'(10275);
			3413: out = 16'(-3382);
			3414: out = 16'(1620);
			3415: out = 16'(-15285);
			3416: out = 16'(1268);
			3417: out = 16'(972);
			3418: out = 16'(-1892);
			3419: out = 16'(9075);
			3420: out = 16'(2796);
			3421: out = 16'(-1675);
			3422: out = 16'(3239);
			3423: out = 16'(-13079);
			3424: out = 16'(5653);
			3425: out = 16'(-18);
			3426: out = 16'(-5245);
			3427: out = 16'(9143);
			3428: out = 16'(-9393);
			3429: out = 16'(18932);
			3430: out = 16'(-14179);
			3431: out = 16'(9438);
			3432: out = 16'(-7104);
			3433: out = 16'(9285);
			3434: out = 16'(-4245);
			3435: out = 16'(-97);
			3436: out = 16'(3308);
			3437: out = 16'(-3671);
			3438: out = 16'(-2837);
			3439: out = 16'(-2775);
			3440: out = 16'(-7775);
			3441: out = 16'(6239);
			3442: out = 16'(-9332);
			3443: out = 16'(10717);
			3444: out = 16'(3136);
			3445: out = 16'(5);
			3446: out = 16'(4867);
			3447: out = 16'(-12192);
			3448: out = 16'(1164);
			3449: out = 16'(-6671);
			3450: out = 16'(4983);
			3451: out = 16'(-516);
			3452: out = 16'(-1281);
			3453: out = 16'(-4561);
			3454: out = 16'(-42);
			3455: out = 16'(-9033);
			3456: out = 16'(5889);
			3457: out = 16'(6948);
			3458: out = 16'(52);
			3459: out = 16'(1620);
			3460: out = 16'(-894);
			3461: out = 16'(-154);
			3462: out = 16'(1892);
			3463: out = 16'(5205);
			3464: out = 16'(-6451);
			3465: out = 16'(13171);
			3466: out = 16'(-12255);
			3467: out = 16'(8004);
			3468: out = 16'(450);
			3469: out = 16'(11399);
			3470: out = 16'(9028);
			3471: out = 16'(1188);
			3472: out = 16'(1903);
			3473: out = 16'(1815);
			3474: out = 16'(3958);
			3475: out = 16'(-142);
			3476: out = 16'(2427);
			3477: out = 16'(-47);
			3478: out = 16'(-8728);
			3479: out = 16'(6900);
			3480: out = 16'(-18541);
			3481: out = 16'(12277);
			3482: out = 16'(-42);
			3483: out = 16'(3065);
			3484: out = 16'(4172);
			3485: out = 16'(-10781);
			3486: out = 16'(2731);
			3487: out = 16'(-6431);
			3488: out = 16'(10465);
			3489: out = 16'(-17196);
			3490: out = 16'(-20);
			3491: out = 16'(-9695);
			3492: out = 16'(-13811);
			3493: out = 16'(9705);
			3494: out = 16'(-11386);
			3495: out = 16'(5179);
			3496: out = 16'(-3961);
			3497: out = 16'(-6500);
			3498: out = 16'(10257);
			3499: out = 16'(-3405);
			3500: out = 16'(4706);
			3501: out = 16'(-5975);
			3502: out = 16'(6488);
			3503: out = 16'(2833);
			3504: out = 16'(-8594);
			3505: out = 16'(8687);
			3506: out = 16'(303);
			3507: out = 16'(2229);
			3508: out = 16'(-2555);
			3509: out = 16'(7247);
			3510: out = 16'(5198);
			3511: out = 16'(3721);
			3512: out = 16'(6213);
			3513: out = 16'(4715);
			3514: out = 16'(4563);
			3515: out = 16'(6262);
			3516: out = 16'(-5960);
			3517: out = 16'(2640);
			3518: out = 16'(635);
			3519: out = 16'(-2321);
			3520: out = 16'(4672);
			3521: out = 16'(-3348);
			3522: out = 16'(11602);
			3523: out = 16'(3649);
			3524: out = 16'(-6222);
			3525: out = 16'(8498);
			3526: out = 16'(-1468);
			3527: out = 16'(16693);
			3528: out = 16'(-3118);
			3529: out = 16'(1247);
			3530: out = 16'(-921);
			3531: out = 16'(-7670);
			3532: out = 16'(-936);
			3533: out = 16'(-11771);
			3534: out = 16'(4440);
			3535: out = 16'(-4773);
			3536: out = 16'(9309);
			3537: out = 16'(-5655);
			3538: out = 16'(3828);
			3539: out = 16'(-10110);
			3540: out = 16'(-3903);
			3541: out = 16'(4510);
			3542: out = 16'(801);
			3543: out = 16'(11269);
			3544: out = 16'(-3638);
			3545: out = 16'(4131);
			3546: out = 16'(-18294);
			3547: out = 16'(10730);
			3548: out = 16'(-9158);
			3549: out = 16'(1898);
			3550: out = 16'(12078);
			3551: out = 16'(6637);
			3552: out = 16'(11416);
			3553: out = 16'(-2756);
			3554: out = 16'(8470);
			3555: out = 16'(8182);
			3556: out = 16'(-2581);
			3557: out = 16'(6818);
			3558: out = 16'(-6744);
			3559: out = 16'(5999);
			3560: out = 16'(-8346);
			3561: out = 16'(9392);
			3562: out = 16'(-3408);
			3563: out = 16'(6664);
			3564: out = 16'(122);
			3565: out = 16'(-3156);
			3566: out = 16'(11775);
			3567: out = 16'(510);
			3568: out = 16'(4167);
			3569: out = 16'(-2904);
			3570: out = 16'(-2790);
			3571: out = 16'(-4692);
			3572: out = 16'(2208);
			3573: out = 16'(-16287);
			3574: out = 16'(5525);
			3575: out = 16'(-12673);
			3576: out = 16'(2039);
			3577: out = 16'(-9236);
			3578: out = 16'(-1940);
			3579: out = 16'(11538);
			3580: out = 16'(-17319);
			3581: out = 16'(5139);
			3582: out = 16'(-15628);
			3583: out = 16'(-4547);
			3584: out = 16'(3099);
			3585: out = 16'(-700);
			3586: out = 16'(770);
			3587: out = 16'(-1142);
			3588: out = 16'(164);
			3589: out = 16'(4838);
			3590: out = 16'(280);
			3591: out = 16'(3168);
			3592: out = 16'(-2665);
			3593: out = 16'(4711);
			3594: out = 16'(-5432);
			3595: out = 16'(-197);
			3596: out = 16'(1513);
			3597: out = 16'(-2711);
			3598: out = 16'(3106);
			3599: out = 16'(7018);
			3600: out = 16'(9255);
			3601: out = 16'(1823);
			3602: out = 16'(-408);
			3603: out = 16'(-1429);
			3604: out = 16'(3888);
			3605: out = 16'(644);
			3606: out = 16'(7931);
			3607: out = 16'(1575);
			3608: out = 16'(1818);
			3609: out = 16'(3100);
			3610: out = 16'(-5725);
			3611: out = 16'(-1639);
			3612: out = 16'(253);
			3613: out = 16'(-2101);
			3614: out = 16'(-2662);
			3615: out = 16'(-737);
			3616: out = 16'(161);
			3617: out = 16'(2677);
			3618: out = 16'(6503);
			3619: out = 16'(-5339);
			3620: out = 16'(-919);
			3621: out = 16'(1276);
			3622: out = 16'(-170);
			3623: out = 16'(3239);
			3624: out = 16'(2506);
			3625: out = 16'(-4307);
			3626: out = 16'(-797);
			3627: out = 16'(-775);
			3628: out = 16'(6707);
			3629: out = 16'(-158);
			3630: out = 16'(-7152);
			3631: out = 16'(8746);
			3632: out = 16'(-6777);
			3633: out = 16'(6118);
			3634: out = 16'(1738);
			3635: out = 16'(-5520);
			3636: out = 16'(-9557);
			3637: out = 16'(4707);
			3638: out = 16'(3089);
			3639: out = 16'(4314);
			3640: out = 16'(10802);
			3641: out = 16'(816);
			3642: out = 16'(-6017);
			3643: out = 16'(1101);
			3644: out = 16'(-15245);
			3645: out = 16'(12920);
			3646: out = 16'(2330);
			3647: out = 16'(2874);
			3648: out = 16'(-2892);
			3649: out = 16'(-6412);
			3650: out = 16'(7022);
			3651: out = 16'(-11871);
			3652: out = 16'(15209);
			3653: out = 16'(-12841);
			3654: out = 16'(3054);
			3655: out = 16'(319);
			3656: out = 16'(-4164);
			3657: out = 16'(14299);
			3658: out = 16'(3234);
			3659: out = 16'(9216);
			3660: out = 16'(-11628);
			3661: out = 16'(8003);
			3662: out = 16'(-10060);
			3663: out = 16'(10644);
			3664: out = 16'(4192);
			3665: out = 16'(3885);
			3666: out = 16'(2402);
			3667: out = 16'(7371);
			3668: out = 16'(-1942);
			3669: out = 16'(7018);
			3670: out = 16'(227);
			3671: out = 16'(11659);
			3672: out = 16'(-2835);
			3673: out = 16'(9274);
			3674: out = 16'(-2823);
			3675: out = 16'(-1833);
			3676: out = 16'(5028);
			3677: out = 16'(4901);
			3678: out = 16'(1556);
			3679: out = 16'(2549);
			3680: out = 16'(4409);
			3681: out = 16'(-1894);
			3682: out = 16'(-10467);
			3683: out = 16'(-5028);
			3684: out = 16'(-4943);
			3685: out = 16'(3642);
			3686: out = 16'(956);
			3687: out = 16'(-12477);
			3688: out = 16'(885);
			3689: out = 16'(-3423);
			3690: out = 16'(-2705);
			3691: out = 16'(661);
			3692: out = 16'(-7338);
			3693: out = 16'(-1221);
			3694: out = 16'(-10860);
			3695: out = 16'(2585);
			3696: out = 16'(-7143);
			3697: out = 16'(6120);
			3698: out = 16'(-1901);
			3699: out = 16'(-32);
			3700: out = 16'(-378);
			3701: out = 16'(-2202);
			3702: out = 16'(2541);
			3703: out = 16'(-1171);
			3704: out = 16'(-2232);
			3705: out = 16'(-4622);
			3706: out = 16'(-5447);
			3707: out = 16'(1321);
			3708: out = 16'(-2767);
			3709: out = 16'(427);
			3710: out = 16'(4319);
			3711: out = 16'(3833);
			3712: out = 16'(6384);
			3713: out = 16'(-279);
			3714: out = 16'(-18086);
			3715: out = 16'(5646);
			3716: out = 16'(968);
			3717: out = 16'(2365);
			3718: out = 16'(4582);
			3719: out = 16'(170);
			3720: out = 16'(-535);
			3721: out = 16'(-5048);
			3722: out = 16'(-8965);
			3723: out = 16'(-1455);
			3724: out = 16'(-1824);
			3725: out = 16'(-6906);
			3726: out = 16'(868);
			3727: out = 16'(-4511);
			3728: out = 16'(4411);
			3729: out = 16'(10405);
			3730: out = 16'(-6376);
			3731: out = 16'(-1584);
			3732: out = 16'(-9140);
			3733: out = 16'(-2615);
			3734: out = 16'(2827);
			3735: out = 16'(-3522);
			3736: out = 16'(5229);
			3737: out = 16'(-4397);
			3738: out = 16'(722);
			3739: out = 16'(-195);
			3740: out = 16'(353);
			3741: out = 16'(7015);
			3742: out = 16'(-9158);
			3743: out = 16'(8094);
			3744: out = 16'(-16937);
			3745: out = 16'(-4005);
			3746: out = 16'(2867);
			3747: out = 16'(4464);
			3748: out = 16'(9338);
			3749: out = 16'(2790);
			3750: out = 16'(-5089);
			3751: out = 16'(-1593);
			3752: out = 16'(-1471);
			3753: out = 16'(-339);
			3754: out = 16'(-3683);
			3755: out = 16'(9400);
			3756: out = 16'(-8009);
			3757: out = 16'(97);
			3758: out = 16'(-8782);
			3759: out = 16'(2799);
			3760: out = 16'(1713);
			3761: out = 16'(-11248);
			3762: out = 16'(-2050);
			3763: out = 16'(-8598);
			3764: out = 16'(-1336);
			3765: out = 16'(-6922);
			3766: out = 16'(-2871);
			3767: out = 16'(353);
			3768: out = 16'(-1040);
			3769: out = 16'(515);
			3770: out = 16'(-4721);
			3771: out = 16'(3614);
			3772: out = 16'(679);
			3773: out = 16'(-5610);
			3774: out = 16'(7192);
			3775: out = 16'(-5809);
			3776: out = 16'(5620);
			3777: out = 16'(4373);
			3778: out = 16'(-5829);
			3779: out = 16'(11895);
			3780: out = 16'(-9058);
			3781: out = 16'(4264);
			3782: out = 16'(180);
			3783: out = 16'(6624);
			3784: out = 16'(-4264);
			3785: out = 16'(12569);
			3786: out = 16'(10993);
			3787: out = 16'(8837);
			3788: out = 16'(7022);
			3789: out = 16'(-9339);
			3790: out = 16'(3651);
			3791: out = 16'(5517);
			3792: out = 16'(938);
			3793: out = 16'(5592);
			3794: out = 16'(-271);
			3795: out = 16'(9645);
			3796: out = 16'(-3466);
			3797: out = 16'(1679);
			3798: out = 16'(-5778);
			3799: out = 16'(7759);
			3800: out = 16'(3015);
			3801: out = 16'(-907);
			3802: out = 16'(7928);
			3803: out = 16'(-10481);
			3804: out = 16'(-2851);
			3805: out = 16'(-9428);
			3806: out = 16'(-8535);
			3807: out = 16'(2614);
			3808: out = 16'(-2318);
			3809: out = 16'(-807);
			3810: out = 16'(-8524);
			3811: out = 16'(-860);
			3812: out = 16'(-8922);
			3813: out = 16'(3609);
			3814: out = 16'(-5163);
			3815: out = 16'(14476);
			3816: out = 16'(-12919);
			3817: out = 16'(-4420);
			3818: out = 16'(-10957);
			3819: out = 16'(-83);
			3820: out = 16'(1698);
			3821: out = 16'(-6290);
			3822: out = 16'(-906);
			3823: out = 16'(4955);
			3824: out = 16'(8333);
			3825: out = 16'(4552);
			3826: out = 16'(4925);
			3827: out = 16'(-4487);
			3828: out = 16'(-7281);
			3829: out = 16'(-1200);
			3830: out = 16'(-6593);
			3831: out = 16'(6542);
			3832: out = 16'(2865);
			3833: out = 16'(6868);
			3834: out = 16'(-2343);
			3835: out = 16'(3409);
			3836: out = 16'(-7945);
			3837: out = 16'(1367);
			3838: out = 16'(4774);
			3839: out = 16'(8839);
			3840: out = 16'(2297);
			3841: out = 16'(7463);
			3842: out = 16'(-6234);
			3843: out = 16'(-535);
			3844: out = 16'(-1963);
			3845: out = 16'(2353);
			3846: out = 16'(-8018);
			3847: out = 16'(8636);
			3848: out = 16'(186);
			3849: out = 16'(3056);
			3850: out = 16'(-6241);
			3851: out = 16'(-2245);
			3852: out = 16'(-5167);
			3853: out = 16'(439);
			3854: out = 16'(1621);
			3855: out = 16'(3795);
			3856: out = 16'(951);
			3857: out = 16'(12757);
			3858: out = 16'(-3565);
			3859: out = 16'(201);
			3860: out = 16'(560);
			3861: out = 16'(946);
			3862: out = 16'(-1425);
			3863: out = 16'(7769);
			3864: out = 16'(1099);
			3865: out = 16'(518);
			3866: out = 16'(-2984);
			3867: out = 16'(-2837);
			3868: out = 16'(331);
			3869: out = 16'(3741);
			3870: out = 16'(-10941);
			3871: out = 16'(9517);
			3872: out = 16'(1878);
			3873: out = 16'(5078);
			3874: out = 16'(-1901);
			3875: out = 16'(-5675);
			3876: out = 16'(-417);
			3877: out = 16'(1061);
			3878: out = 16'(2153);
			3879: out = 16'(-697);
			3880: out = 16'(-1341);
			3881: out = 16'(4915);
			3882: out = 16'(-20447);
			3883: out = 16'(3573);
			3884: out = 16'(-9020);
			3885: out = 16'(9356);
			3886: out = 16'(1003);
			3887: out = 16'(-5487);
			3888: out = 16'(-640);
			3889: out = 16'(-8188);
			3890: out = 16'(-1374);
			3891: out = 16'(1100);
			3892: out = 16'(-919);
			3893: out = 16'(13525);
			3894: out = 16'(-5486);
			3895: out = 16'(8954);
			3896: out = 16'(-3028);
			3897: out = 16'(938);
			3898: out = 16'(-1595);
			3899: out = 16'(-4551);
			3900: out = 16'(-797);
			3901: out = 16'(1078);
			3902: out = 16'(8814);
			3903: out = 16'(5486);
			3904: out = 16'(3234);
			3905: out = 16'(7157);
			3906: out = 16'(4600);
			3907: out = 16'(-426);
			3908: out = 16'(145);
			3909: out = 16'(253);
			3910: out = 16'(6650);
			3911: out = 16'(-5631);
			3912: out = 16'(4168);
			3913: out = 16'(-2777);
			3914: out = 16'(1676);
			3915: out = 16'(1477);
			3916: out = 16'(-1450);
			3917: out = 16'(9789);
			3918: out = 16'(-9797);
			3919: out = 16'(4736);
			3920: out = 16'(667);
			3921: out = 16'(1469);
			3922: out = 16'(-3561);
			3923: out = 16'(-9585);
			3924: out = 16'(4731);
			3925: out = 16'(-4655);
			3926: out = 16'(5619);
			3927: out = 16'(5107);
			3928: out = 16'(136);
			3929: out = 16'(7257);
			3930: out = 16'(-11949);
			3931: out = 16'(380);
			3932: out = 16'(-5649);
			3933: out = 16'(11807);
			3934: out = 16'(3033);
			3935: out = 16'(-1883);
			3936: out = 16'(-2561);
			3937: out = 16'(-9479);
			3938: out = 16'(10266);
			3939: out = 16'(-3564);
			3940: out = 16'(9768);
			3941: out = 16'(-1813);
			3942: out = 16'(3045);
			3943: out = 16'(7064);
			3944: out = 16'(5957);
			3945: out = 16'(6242);
			3946: out = 16'(9588);
			3947: out = 16'(861);
			3948: out = 16'(-101);
			3949: out = 16'(-324);
			3950: out = 16'(719);
			3951: out = 16'(1959);
			3952: out = 16'(1959);
			3953: out = 16'(-1706);
			3954: out = 16'(-3249);
			3955: out = 16'(3468);
			3956: out = 16'(-1992);
			3957: out = 16'(-1584);
			3958: out = 16'(6430);
			3959: out = 16'(750);
			3960: out = 16'(-5325);
			3961: out = 16'(-14646);
			3962: out = 16'(4267);
			3963: out = 16'(783);
			3964: out = 16'(3750);
			3965: out = 16'(-386);
			3966: out = 16'(-8245);
			3967: out = 16'(5456);
			3968: out = 16'(-7701);
			3969: out = 16'(2659);
			3970: out = 16'(-2495);
			3971: out = 16'(3370);
			3972: out = 16'(-63);
			3973: out = 16'(-14023);
			3974: out = 16'(2860);
			3975: out = 16'(-18306);
			3976: out = 16'(8949);
			3977: out = 16'(714);
			3978: out = 16'(-6054);
			3979: out = 16'(5056);
			3980: out = 16'(-4750);
			3981: out = 16'(-7054);
			3982: out = 16'(-2849);
			3983: out = 16'(13594);
			3984: out = 16'(-13704);
			3985: out = 16'(4071);
			3986: out = 16'(-24);
			3987: out = 16'(-2047);
			3988: out = 16'(7647);
			3989: out = 16'(-18755);
			3990: out = 16'(5064);
			3991: out = 16'(3237);
			3992: out = 16'(-5140);
			3993: out = 16'(-9487);
			3994: out = 16'(856);
			3995: out = 16'(6655);
			3996: out = 16'(9104);
			3997: out = 16'(4939);
			3998: out = 16'(-637);
			3999: out = 16'(49);
			4000: out = 16'(2183);
			4001: out = 16'(-8444);
			4002: out = 16'(-790);
			4003: out = 16'(2991);
			4004: out = 16'(61);
			4005: out = 16'(-386);
			4006: out = 16'(-1234);
			4007: out = 16'(12207);
			4008: out = 16'(-613);
			4009: out = 16'(5005);
			4010: out = 16'(-4454);
			4011: out = 16'(-2516);
			4012: out = 16'(2614);
			4013: out = 16'(-8201);
			4014: out = 16'(2444);
			4015: out = 16'(2823);
			4016: out = 16'(4976);
			4017: out = 16'(-5084);
			4018: out = 16'(-2807);
			4019: out = 16'(661);
			4020: out = 16'(289);
			4021: out = 16'(2106);
			4022: out = 16'(5049);
			4023: out = 16'(1747);
			4024: out = 16'(2208);
			4025: out = 16'(-5349);
			4026: out = 16'(758);
			4027: out = 16'(-25);
			4028: out = 16'(10977);
			4029: out = 16'(-460);
			4030: out = 16'(7891);
			4031: out = 16'(-1198);
			4032: out = 16'(-6628);
			4033: out = 16'(-3735);
			4034: out = 16'(-7249);
			4035: out = 16'(3790);
			4036: out = 16'(1415);
			4037: out = 16'(-1337);
			4038: out = 16'(1951);
			4039: out = 16'(1717);
			4040: out = 16'(-1602);
			4041: out = 16'(-63);
			4042: out = 16'(532);
			4043: out = 16'(1192);
			4044: out = 16'(-11489);
			4045: out = 16'(-2003);
			4046: out = 16'(-342);
			4047: out = 16'(5583);
			4048: out = 16'(7727);
			4049: out = 16'(-977);
			4050: out = 16'(-3187);
			4051: out = 16'(-9436);
			4052: out = 16'(-6496);
			4053: out = 16'(-408);
			4054: out = 16'(1331);
			4055: out = 16'(-2205);
			4056: out = 16'(1748);
			4057: out = 16'(-178);
			4058: out = 16'(-168);
			4059: out = 16'(1872);
			4060: out = 16'(-101);
			4061: out = 16'(85);
			4062: out = 16'(8405);
			4063: out = 16'(-1406);
			4064: out = 16'(1138);
			4065: out = 16'(-3249);
			4066: out = 16'(4898);
			4067: out = 16'(229);
			4068: out = 16'(-2156);
			4069: out = 16'(8268);
			4070: out = 16'(-4051);
			4071: out = 16'(7140);
			4072: out = 16'(-572);
			4073: out = 16'(-5066);
			4074: out = 16'(1034);
			4075: out = 16'(-3169);
			4076: out = 16'(2415);
			4077: out = 16'(-4078);
			4078: out = 16'(-14);
			4079: out = 16'(-5003);
			4080: out = 16'(5045);
			4081: out = 16'(4646);
			4082: out = 16'(-4207);
			4083: out = 16'(-3172);
			4084: out = 16'(-2468);
			4085: out = 16'(1938);
			4086: out = 16'(8);
			4087: out = 16'(7143);
			4088: out = 16'(5609);
			4089: out = 16'(-1767);
			4090: out = 16'(4073);
			4091: out = 16'(-3140);
			4092: out = 16'(-12250);
			4093: out = 16'(3284);
			4094: out = 16'(-13436);
			4095: out = 16'(3518);
			4096: out = 16'(1386);
			4097: out = 16'(3936);
			4098: out = 16'(-2412);
			4099: out = 16'(3547);
			4100: out = 16'(3099);
			4101: out = 16'(-3615);
			4102: out = 16'(8133);
			4103: out = 16'(-5458);
			4104: out = 16'(-4156);
			4105: out = 16'(2218);
			4106: out = 16'(-10719);
			4107: out = 16'(2512);
			4108: out = 16'(-5593);
			4109: out = 16'(6655);
			4110: out = 16'(-579);
			4111: out = 16'(3666);
			4112: out = 16'(12859);
			4113: out = 16'(-4591);
			4114: out = 16'(10394);
			4115: out = 16'(-2853);
			4116: out = 16'(-431);
			4117: out = 16'(-1529);
			4118: out = 16'(2967);
			4119: out = 16'(7227);
			4120: out = 16'(-1681);
			4121: out = 16'(9417);
			4122: out = 16'(-4043);
			4123: out = 16'(-760);
			4124: out = 16'(6141);
			4125: out = 16'(-8869);
			4126: out = 16'(1441);
			4127: out = 16'(-5657);
			4128: out = 16'(1888);
			4129: out = 16'(1636);
			4130: out = 16'(1184);
			4131: out = 16'(4);
			4132: out = 16'(83);
			4133: out = 16'(-1847);
			4134: out = 16'(1790);
			4135: out = 16'(-4789);
			4136: out = 16'(1728);
			4137: out = 16'(-3424);
			4138: out = 16'(510);
			4139: out = 16'(-576);
			4140: out = 16'(3252);
			4141: out = 16'(-803);
			4142: out = 16'(21);
			4143: out = 16'(65);
			4144: out = 16'(4827);
			4145: out = 16'(1555);
			4146: out = 16'(5257);
			4147: out = 16'(-2641);
			4148: out = 16'(-43);
			4149: out = 16'(-10381);
			4150: out = 16'(-2723);
			4151: out = 16'(1098);
			4152: out = 16'(10004);
			4153: out = 16'(10293);
			4154: out = 16'(4538);
			4155: out = 16'(-3177);
			4156: out = 16'(598);
			4157: out = 16'(-5332);
			4158: out = 16'(1970);
			4159: out = 16'(4104);
			4160: out = 16'(-3407);
			4161: out = 16'(-2391);
			4162: out = 16'(-3436);
			4163: out = 16'(-5271);
			4164: out = 16'(11460);
			4165: out = 16'(-2643);
			4166: out = 16'(1006);
			4167: out = 16'(-7607);
			4168: out = 16'(11366);
			4169: out = 16'(-1936);
			4170: out = 16'(6159);
			4171: out = 16'(1190);
			4172: out = 16'(-2659);
			4173: out = 16'(4577);
			4174: out = 16'(-1340);
			4175: out = 16'(-2336);
			4176: out = 16'(842);
			4177: out = 16'(-3902);
			4178: out = 16'(-2259);
			4179: out = 16'(-11178);
			4180: out = 16'(9474);
			4181: out = 16'(458);
			4182: out = 16'(-613);
			4183: out = 16'(2282);
			4184: out = 16'(-10621);
			4185: out = 16'(3891);
			4186: out = 16'(4223);
			4187: out = 16'(4128);
			4188: out = 16'(4473);
			4189: out = 16'(-4409);
			4190: out = 16'(5235);
			4191: out = 16'(6710);
			4192: out = 16'(10682);
			4193: out = 16'(3666);
			4194: out = 16'(592);
			4195: out = 16'(313);
			4196: out = 16'(-594);
			4197: out = 16'(-898);
			4198: out = 16'(6109);
			4199: out = 16'(-1221);
			4200: out = 16'(-392);
			4201: out = 16'(-6317);
			4202: out = 16'(-6522);
			4203: out = 16'(-5129);
			4204: out = 16'(7833);
			4205: out = 16'(2312);
			4206: out = 16'(-629);
			4207: out = 16'(4584);
			4208: out = 16'(-920);
			4209: out = 16'(-5130);
			4210: out = 16'(1117);
			4211: out = 16'(516);
			4212: out = 16'(-2628);
			4213: out = 16'(-636);
			4214: out = 16'(4299);
			4215: out = 16'(-6864);
			4216: out = 16'(9443);
			4217: out = 16'(-990);
			4218: out = 16'(2494);
			4219: out = 16'(-1097);
			4220: out = 16'(-8346);
			4221: out = 16'(-1850);
			4222: out = 16'(3367);
			4223: out = 16'(9009);
			4224: out = 16'(10294);
			4225: out = 16'(4031);
			4226: out = 16'(6005);
			4227: out = 16'(-1312);
			4228: out = 16'(4837);
			4229: out = 16'(466);
			4230: out = 16'(4713);
			4231: out = 16'(7480);
			4232: out = 16'(1565);
			4233: out = 16'(2742);
			4234: out = 16'(-8301);
			4235: out = 16'(5637);
			4236: out = 16'(-4088);
			4237: out = 16'(2868);
			4238: out = 16'(-7936);
			4239: out = 16'(-2496);
			4240: out = 16'(6109);
			4241: out = 16'(-5883);
			4242: out = 16'(2211);
			4243: out = 16'(2546);
			4244: out = 16'(-1406);
			4245: out = 16'(1776);
			4246: out = 16'(-8155);
			4247: out = 16'(2037);
			4248: out = 16'(-469);
			4249: out = 16'(-629);
			4250: out = 16'(-5095);
			4251: out = 16'(-4959);
			4252: out = 16'(-146);
			4253: out = 16'(-9798);
			4254: out = 16'(911);
			4255: out = 16'(-4607);
			4256: out = 16'(3727);
			4257: out = 16'(1776);
			4258: out = 16'(-1544);
			4259: out = 16'(7077);
			4260: out = 16'(-7198);
			4261: out = 16'(3044);
			4262: out = 16'(-7165);
			4263: out = 16'(4087);
			4264: out = 16'(-2799);
			4265: out = 16'(-1328);
			4266: out = 16'(4303);
			4267: out = 16'(-4651);
			4268: out = 16'(7936);
			4269: out = 16'(-2599);
			4270: out = 16'(-3166);
			4271: out = 16'(405);
			4272: out = 16'(-4940);
			4273: out = 16'(6163);
			4274: out = 16'(-12345);
			4275: out = 16'(10483);
			4276: out = 16'(929);
			4277: out = 16'(4218);
			4278: out = 16'(3744);
			4279: out = 16'(3926);
			4280: out = 16'(1960);
			4281: out = 16'(-1775);
			4282: out = 16'(336);
			4283: out = 16'(-1119);
			4284: out = 16'(-3216);
			4285: out = 16'(607);
			4286: out = 16'(-6071);
			4287: out = 16'(4819);
			4288: out = 16'(967);
			4289: out = 16'(2088);
			4290: out = 16'(1407);
			4291: out = 16'(1888);
			4292: out = 16'(-367);
			4293: out = 16'(-584);
			4294: out = 16'(-4019);
			4295: out = 16'(3195);
			4296: out = 16'(-574);
			4297: out = 16'(3506);
			4298: out = 16'(2472);
			4299: out = 16'(-678);
			4300: out = 16'(3597);
			4301: out = 16'(-10625);
			4302: out = 16'(479);
			4303: out = 16'(-5996);
			4304: out = 16'(1304);
			4305: out = 16'(-1461);
			4306: out = 16'(-894);
			4307: out = 16'(5120);
			4308: out = 16'(-4522);
			4309: out = 16'(4535);
			4310: out = 16'(2149);
			4311: out = 16'(-1986);
			4312: out = 16'(2402);
			4313: out = 16'(-3104);
			4314: out = 16'(3481);
			4315: out = 16'(-4308);
			4316: out = 16'(3571);
			4317: out = 16'(762);
			4318: out = 16'(2862);
			4319: out = 16'(1178);
			4320: out = 16'(1561);
			4321: out = 16'(6870);
			4322: out = 16'(-10448);
			4323: out = 16'(-510);
			4324: out = 16'(-2792);
			4325: out = 16'(-3393);
			4326: out = 16'(-4915);
			4327: out = 16'(4739);
			4328: out = 16'(-1116);
			4329: out = 16'(-13584);
			4330: out = 16'(11641);
			4331: out = 16'(-12909);
			4332: out = 16'(2934);
			4333: out = 16'(640);
			4334: out = 16'(-1536);
			4335: out = 16'(-1347);
			4336: out = 16'(-763);
			4337: out = 16'(-880);
			4338: out = 16'(1002);
			4339: out = 16'(-132);
			4340: out = 16'(4488);
			4341: out = 16'(-4560);
			4342: out = 16'(8622);
			4343: out = 16'(-3635);
			4344: out = 16'(1522);
			4345: out = 16'(-2491);
			4346: out = 16'(-2091);
			4347: out = 16'(181);
			4348: out = 16'(-1156);
			4349: out = 16'(3723);
			4350: out = 16'(-2806);
			4351: out = 16'(8211);
			4352: out = 16'(5891);
			4353: out = 16'(-9229);
			4354: out = 16'(11018);
			4355: out = 16'(-14630);
			4356: out = 16'(2090);
			4357: out = 16'(2044);
			4358: out = 16'(-6767);
			4359: out = 16'(4112);
			4360: out = 16'(1797);
			4361: out = 16'(1584);
			4362: out = 16'(6168);
			4363: out = 16'(1341);
			4364: out = 16'(-1);
			4365: out = 16'(-15112);
			4366: out = 16'(5140);
			4367: out = 16'(-9259);
			4368: out = 16'(101);
			4369: out = 16'(8108);
			4370: out = 16'(-1634);
			4371: out = 16'(2994);
			4372: out = 16'(-8047);
			4373: out = 16'(-332);
			4374: out = 16'(-3346);
			4375: out = 16'(3676);
			4376: out = 16'(-2313);
			4377: out = 16'(-7722);
			4378: out = 16'(841);
			4379: out = 16'(2595);
			4380: out = 16'(-310);
			4381: out = 16'(6078);
			4382: out = 16'(2385);
			4383: out = 16'(-723);
			4384: out = 16'(-2136);
			4385: out = 16'(2246);
			4386: out = 16'(3258);
			4387: out = 16'(5284);
			4388: out = 16'(-5372);
			4389: out = 16'(1040);
			4390: out = 16'(7018);
			4391: out = 16'(57);
			4392: out = 16'(6898);
			4393: out = 16'(516);
			4394: out = 16'(53);
			4395: out = 16'(4950);
			4396: out = 16'(-133);
			4397: out = 16'(-6153);
			4398: out = 16'(-6578);
			4399: out = 16'(1432);
			4400: out = 16'(-8106);
			4401: out = 16'(6094);
			4402: out = 16'(153);
			4403: out = 16'(-7521);
			4404: out = 16'(1042);
			4405: out = 16'(-1843);
			4406: out = 16'(544);
			4407: out = 16'(-3582);
			4408: out = 16'(638);
			4409: out = 16'(679);
			4410: out = 16'(-10643);
			4411: out = 16'(-1204);
			4412: out = 16'(-1871);
			4413: out = 16'(1388);
			4414: out = 16'(5646);
			4415: out = 16'(-1984);
			4416: out = 16'(464);
			4417: out = 16'(-6800);
			4418: out = 16'(-2728);
			4419: out = 16'(733);
			4420: out = 16'(188);
			4421: out = 16'(5912);
			4422: out = 16'(-955);
			4423: out = 16'(5233);
			4424: out = 16'(-4107);
			4425: out = 16'(-1773);
			4426: out = 16'(-973);
			4427: out = 16'(-5434);
			4428: out = 16'(3886);
			4429: out = 16'(-1053);
			4430: out = 16'(-5546);
			4431: out = 16'(1849);
			4432: out = 16'(-6947);
			4433: out = 16'(5879);
			4434: out = 16'(-2354);
			4435: out = 16'(1471);
			4436: out = 16'(-951);
			4437: out = 16'(-6687);
			4438: out = 16'(-1179);
			4439: out = 16'(-10613);
			4440: out = 16'(-6867);
			4441: out = 16'(-334);
			4442: out = 16'(-7184);
			4443: out = 16'(-1535);
			4444: out = 16'(1592);
			4445: out = 16'(-731);
			4446: out = 16'(-3088);
			4447: out = 16'(2002);
			4448: out = 16'(-5295);
			4449: out = 16'(912);
			4450: out = 16'(-3262);
			4451: out = 16'(1811);
			4452: out = 16'(1932);
			4453: out = 16'(4162);
			4454: out = 16'(-5183);
			4455: out = 16'(-864);
			4456: out = 16'(-1260);
			4457: out = 16'(5346);
			4458: out = 16'(2320);
			4459: out = 16'(-603);
			4460: out = 16'(7306);
			4461: out = 16'(5451);
			4462: out = 16'(-10933);
			4463: out = 16'(640);
			4464: out = 16'(-919);
			4465: out = 16'(8498);
			4466: out = 16'(-2085);
			4467: out = 16'(-2397);
			4468: out = 16'(1467);
			4469: out = 16'(-7131);
			4470: out = 16'(2975);
			4471: out = 16'(1610);
			4472: out = 16'(187);
			4473: out = 16'(569);
			4474: out = 16'(-2024);
			4475: out = 16'(-445);
			4476: out = 16'(-821);
			4477: out = 16'(1857);
			4478: out = 16'(-734);
			4479: out = 16'(-4998);
			4480: out = 16'(-10);
			4481: out = 16'(-8870);
			4482: out = 16'(-6011);
			4483: out = 16'(1106);
			4484: out = 16'(6334);
			4485: out = 16'(7946);
			4486: out = 16'(-424);
			4487: out = 16'(233);
			4488: out = 16'(792);
			4489: out = 16'(-3428);
			4490: out = 16'(-3281);
			4491: out = 16'(1891);
			4492: out = 16'(4049);
			4493: out = 16'(1952);
			4494: out = 16'(34);
			4495: out = 16'(-32);
			4496: out = 16'(4852);
			4497: out = 16'(721);
			4498: out = 16'(1409);
			4499: out = 16'(6036);
			4500: out = 16'(-3977);
			4501: out = 16'(5309);
			4502: out = 16'(1610);
			4503: out = 16'(-1433);
			4504: out = 16'(7175);
			4505: out = 16'(-2052);
			4506: out = 16'(-1075);
			4507: out = 16'(-2127);
			4508: out = 16'(-482);
			4509: out = 16'(5882);
			4510: out = 16'(2904);
			4511: out = 16'(-7015);
			4512: out = 16'(23);
			4513: out = 16'(-4149);
			4514: out = 16'(-5664);
			4515: out = 16'(-1784);
			4516: out = 16'(7143);
			4517: out = 16'(3805);
			4518: out = 16'(1404);
			4519: out = 16'(-938);
			4520: out = 16'(340);
			4521: out = 16'(-4592);
			4522: out = 16'(-3137);
			4523: out = 16'(1645);
			4524: out = 16'(-3970);
			4525: out = 16'(-4610);
			4526: out = 16'(3097);
			4527: out = 16'(-3321);
			4528: out = 16'(3706);
			4529: out = 16'(-3718);
			4530: out = 16'(5516);
			4531: out = 16'(-2747);
			4532: out = 16'(6195);
			4533: out = 16'(-1698);
			4534: out = 16'(54);
			4535: out = 16'(-5877);
			4536: out = 16'(3571);
			4537: out = 16'(8351);
			4538: out = 16'(-1291);
			4539: out = 16'(3268);
			4540: out = 16'(3070);
			4541: out = 16'(-3301);
			4542: out = 16'(4269);
			4543: out = 16'(-4948);
			4544: out = 16'(3057);
			4545: out = 16'(-3956);
			4546: out = 16'(6868);
			4547: out = 16'(-117);
			4548: out = 16'(7173);
			4549: out = 16'(1703);
			4550: out = 16'(-622);
			4551: out = 16'(4103);
			4552: out = 16'(-6009);
			4553: out = 16'(-152);
			4554: out = 16'(2426);
			4555: out = 16'(574);
			4556: out = 16'(2522);
			4557: out = 16'(-2020);
			4558: out = 16'(1800);
			4559: out = 16'(-2927);
			4560: out = 16'(2521);
			4561: out = 16'(5691);
			4562: out = 16'(-3878);
			4563: out = 16'(2305);
			4564: out = 16'(-4902);
			4565: out = 16'(2028);
			4566: out = 16'(291);
			4567: out = 16'(-3931);
			4568: out = 16'(-3201);
			4569: out = 16'(509);
			4570: out = 16'(-1702);
			4571: out = 16'(6036);
			4572: out = 16'(2767);
			4573: out = 16'(-4315);
			4574: out = 16'(-3311);
			4575: out = 16'(7559);
			4576: out = 16'(-3048);
			4577: out = 16'(-3969);
			4578: out = 16'(-4567);
			4579: out = 16'(-2301);
			4580: out = 16'(8146);
			4581: out = 16'(1850);
			4582: out = 16'(5343);
			4583: out = 16'(-500);
			4584: out = 16'(-3161);
			4585: out = 16'(65);
			4586: out = 16'(-13429);
			4587: out = 16'(3588);
			4588: out = 16'(-802);
			4589: out = 16'(-782);
			4590: out = 16'(7341);
			4591: out = 16'(-612);
			4592: out = 16'(1685);
			4593: out = 16'(-415);
			4594: out = 16'(3039);
			4595: out = 16'(-5815);
			4596: out = 16'(502);
			4597: out = 16'(-41);
			4598: out = 16'(573);
			4599: out = 16'(10752);
			4600: out = 16'(-5871);
			4601: out = 16'(3301);
			4602: out = 16'(-6195);
			4603: out = 16'(-164);
			4604: out = 16'(-4116);
			4605: out = 16'(1745);
			4606: out = 16'(-464);
			4607: out = 16'(3339);
			4608: out = 16'(-304);
			4609: out = 16'(377);
			4610: out = 16'(-4540);
			4611: out = 16'(151);
			4612: out = 16'(305);
			4613: out = 16'(4801);
			4614: out = 16'(6902);
			4615: out = 16'(6954);
			4616: out = 16'(-59);
			4617: out = 16'(-2654);
			4618: out = 16'(-1939);
			4619: out = 16'(31);
			4620: out = 16'(-7164);
			4621: out = 16'(7036);
			4622: out = 16'(1475);
			4623: out = 16'(7733);
			4624: out = 16'(1484);
			4625: out = 16'(-3496);
			4626: out = 16'(-9710);
			4627: out = 16'(-1395);
			4628: out = 16'(-6036);
			4629: out = 16'(998);
			4630: out = 16'(785);
			4631: out = 16'(2065);
			4632: out = 16'(3450);
			4633: out = 16'(4936);
			4634: out = 16'(-2573);
			4635: out = 16'(-820);
			4636: out = 16'(-880);
			4637: out = 16'(3798);
			4638: out = 16'(-2572);
			4639: out = 16'(1779);
			4640: out = 16'(3309);
			4641: out = 16'(-4033);
			4642: out = 16'(10801);
			4643: out = 16'(-869);
			4644: out = 16'(-615);
			4645: out = 16'(-116);
			4646: out = 16'(-200);
			4647: out = 16'(30);
			4648: out = 16'(2401);
			4649: out = 16'(627);
			4650: out = 16'(-3170);
			4651: out = 16'(9958);
			4652: out = 16'(-4950);
			4653: out = 16'(7002);
			4654: out = 16'(8521);
			4655: out = 16'(-2243);
			4656: out = 16'(3189);
			4657: out = 16'(-4119);
			4658: out = 16'(-173);
			4659: out = 16'(-6172);
			4660: out = 16'(3971);
			4661: out = 16'(569);
			4662: out = 16'(-1393);
			4663: out = 16'(3780);
			4664: out = 16'(4348);
			4665: out = 16'(-3816);
			4666: out = 16'(1956);
			4667: out = 16'(-5387);
			4668: out = 16'(1848);
			4669: out = 16'(-978);
			4670: out = 16'(-1357);
			4671: out = 16'(4258);
			4672: out = 16'(-383);
			4673: out = 16'(5904);
			4674: out = 16'(6491);
			4675: out = 16'(3201);
			4676: out = 16'(1355);
			4677: out = 16'(3543);
			4678: out = 16'(-180);
			4679: out = 16'(-4157);
			4680: out = 16'(-782);
			4681: out = 16'(-4614);
			4682: out = 16'(-1449);
			4683: out = 16'(-4638);
			4684: out = 16'(6953);
			4685: out = 16'(8649);
			4686: out = 16'(-2308);
			4687: out = 16'(4105);
			4688: out = 16'(-1462);
			4689: out = 16'(103);
			4690: out = 16'(-2669);
			4691: out = 16'(1757);
			4692: out = 16'(6935);
			4693: out = 16'(-1545);
			4694: out = 16'(9164);
			4695: out = 16'(-2244);
			4696: out = 16'(6957);
			4697: out = 16'(-1594);
			4698: out = 16'(1546);
			4699: out = 16'(-4003);
			4700: out = 16'(-2019);
			4701: out = 16'(-2622);
			4702: out = 16'(1304);
			4703: out = 16'(6251);
			4704: out = 16'(-2553);
			4705: out = 16'(6047);
			4706: out = 16'(-1446);
			4707: out = 16'(-6962);
			4708: out = 16'(7282);
			4709: out = 16'(-12765);
			4710: out = 16'(5462);
			4711: out = 16'(-11641);
			4712: out = 16'(-2016);
			4713: out = 16'(4032);
			4714: out = 16'(-7777);
			4715: out = 16'(5172);
			4716: out = 16'(7831);
			4717: out = 16'(-4516);
			4718: out = 16'(4708);
			4719: out = 16'(-7522);
			4720: out = 16'(2374);
			4721: out = 16'(-3025);
			4722: out = 16'(-2111);
			4723: out = 16'(681);
			4724: out = 16'(838);
			4725: out = 16'(1487);
			4726: out = 16'(7775);
			4727: out = 16'(-627);
			4728: out = 16'(648);
			4729: out = 16'(1183);
			4730: out = 16'(-2976);
			4731: out = 16'(-9000);
			4732: out = 16'(-1069);
			4733: out = 16'(-1180);
			4734: out = 16'(6667);
			4735: out = 16'(3997);
			4736: out = 16'(1808);
			4737: out = 16'(9585);
			4738: out = 16'(-4782);
			4739: out = 16'(-1114);
			4740: out = 16'(-522);
			4741: out = 16'(-720);
			4742: out = 16'(-2533);
			4743: out = 16'(531);
			4744: out = 16'(-212);
			4745: out = 16'(-349);
			4746: out = 16'(3699);
			4747: out = 16'(-2878);
			4748: out = 16'(-2342);
			4749: out = 16'(-2241);
			4750: out = 16'(-3251);
			4751: out = 16'(-2469);
			4752: out = 16'(-244);
			4753: out = 16'(5632);
			4754: out = 16'(-7939);
			4755: out = 16'(10460);
			4756: out = 16'(-1043);
			4757: out = 16'(-800);
			4758: out = 16'(3951);
			4759: out = 16'(-9030);
			4760: out = 16'(3365);
			4761: out = 16'(-7518);
			4762: out = 16'(-588);
			4763: out = 16'(-3804);
			4764: out = 16'(-2997);
			4765: out = 16'(4053);
			4766: out = 16'(-7351);
			4767: out = 16'(6214);
			4768: out = 16'(3880);
			4769: out = 16'(-7687);
			4770: out = 16'(1049);
			4771: out = 16'(-2139);
			4772: out = 16'(712);
			4773: out = 16'(5009);
			4774: out = 16'(-1400);
			4775: out = 16'(3606);
			4776: out = 16'(1555);
			4777: out = 16'(963);
			4778: out = 16'(2279);
			4779: out = 16'(1068);
			4780: out = 16'(265);
			4781: out = 16'(-5943);
			4782: out = 16'(5779);
			4783: out = 16'(-956);
			4784: out = 16'(-1154);
			4785: out = 16'(-270);
			4786: out = 16'(-3711);
			4787: out = 16'(10056);
			4788: out = 16'(-2550);
			4789: out = 16'(10339);
			4790: out = 16'(-5804);
			4791: out = 16'(3007);
			4792: out = 16'(-4331);
			4793: out = 16'(-7491);
			4794: out = 16'(2575);
			4795: out = 16'(-2715);
			4796: out = 16'(-466);
			4797: out = 16'(6242);
			4798: out = 16'(-3197);
			4799: out = 16'(7470);
			4800: out = 16'(-2017);
			4801: out = 16'(1353);
			4802: out = 16'(-3230);
			4803: out = 16'(-5501);
			4804: out = 16'(-3139);
			4805: out = 16'(-786);
			4806: out = 16'(-798);
			4807: out = 16'(6032);
			4808: out = 16'(4389);
			4809: out = 16'(-741);
			4810: out = 16'(7114);
			4811: out = 16'(-16627);
			4812: out = 16'(-6);
			4813: out = 16'(-3154);
			4814: out = 16'(-182);
			4815: out = 16'(7109);
			4816: out = 16'(-7493);
			4817: out = 16'(4191);
			4818: out = 16'(-142);
			4819: out = 16'(-423);
			4820: out = 16'(3744);
			4821: out = 16'(-1192);
			4822: out = 16'(3822);
			4823: out = 16'(-7830);
			4824: out = 16'(-3651);
			4825: out = 16'(1033);
			4826: out = 16'(-53);
			4827: out = 16'(3033);
			4828: out = 16'(-2568);
			4829: out = 16'(2484);
			4830: out = 16'(448);
			4831: out = 16'(-264);
			4832: out = 16'(3055);
			4833: out = 16'(-4755);
			4834: out = 16'(6709);
			4835: out = 16'(-1430);
			4836: out = 16'(65);
			4837: out = 16'(3366);
			4838: out = 16'(997);
			4839: out = 16'(6296);
			4840: out = 16'(-6376);
			4841: out = 16'(2025);
			4842: out = 16'(-986);
			4843: out = 16'(-5973);
			4844: out = 16'(6793);
			4845: out = 16'(-3259);
			4846: out = 16'(3138);
			4847: out = 16'(-12807);
			4848: out = 16'(-4830);
			4849: out = 16'(8435);
			4850: out = 16'(-6156);
			4851: out = 16'(946);
			4852: out = 16'(1517);
			4853: out = 16'(-5897);
			4854: out = 16'(5515);
			4855: out = 16'(-5642);
			4856: out = 16'(4754);
			4857: out = 16'(9531);
			4858: out = 16'(4948);
			4859: out = 16'(1232);
			4860: out = 16'(3417);
			4861: out = 16'(-3525);
			4862: out = 16'(2759);
			4863: out = 16'(-4242);
			4864: out = 16'(-2783);
			4865: out = 16'(917);
			4866: out = 16'(-7084);
			4867: out = 16'(4205);
			4868: out = 16'(-2216);
			4869: out = 16'(4048);
			4870: out = 16'(-745);
			4871: out = 16'(794);
			4872: out = 16'(6010);
			4873: out = 16'(-5018);
			4874: out = 16'(1871);
			4875: out = 16'(-3527);
			4876: out = 16'(7851);
			4877: out = 16'(-224);
			4878: out = 16'(3145);
			4879: out = 16'(5269);
			4880: out = 16'(106);
			4881: out = 16'(5024);
			4882: out = 16'(-3968);
			4883: out = 16'(-183);
			4884: out = 16'(6806);
			4885: out = 16'(-11989);
			4886: out = 16'(-995);
			4887: out = 16'(-2528);
			4888: out = 16'(8027);
			4889: out = 16'(-738);
			4890: out = 16'(269);
			4891: out = 16'(1939);
			4892: out = 16'(-236);
			4893: out = 16'(-5881);
			4894: out = 16'(5165);
			4895: out = 16'(-13);
			4896: out = 16'(10384);
			4897: out = 16'(-5611);
			4898: out = 16'(-938);
			4899: out = 16'(5359);
			4900: out = 16'(-1398);
			4901: out = 16'(3617);
			4902: out = 16'(-3028);
			4903: out = 16'(1201);
			4904: out = 16'(41);
			4905: out = 16'(-2424);
			4906: out = 16'(298);
			4907: out = 16'(412);
			4908: out = 16'(3179);
			4909: out = 16'(-7809);
			4910: out = 16'(3083);
			4911: out = 16'(6578);
			4912: out = 16'(2787);
			4913: out = 16'(2985);
			4914: out = 16'(-3122);
			4915: out = 16'(910);
			4916: out = 16'(1355);
			4917: out = 16'(1415);
			4918: out = 16'(3643);
			4919: out = 16'(5944);
			4920: out = 16'(5361);
			4921: out = 16'(-6631);
			4922: out = 16'(-4225);
			4923: out = 16'(4153);
			4924: out = 16'(-1051);
			4925: out = 16'(-1764);
			4926: out = 16'(738);
			4927: out = 16'(114);
			4928: out = 16'(871);
			4929: out = 16'(177);
			4930: out = 16'(8400);
			4931: out = 16'(293);
			4932: out = 16'(6167);
			4933: out = 16'(-284);
			4934: out = 16'(31);
			4935: out = 16'(778);
			4936: out = 16'(461);
			4937: out = 16'(-2394);
			4938: out = 16'(8650);
			4939: out = 16'(-4476);
			4940: out = 16'(3019);
			4941: out = 16'(532);
			4942: out = 16'(1828);
			4943: out = 16'(7270);
			4944: out = 16'(2496);
			4945: out = 16'(-2308);
			4946: out = 16'(-2155);
			4947: out = 16'(-4657);
			4948: out = 16'(834);
			4949: out = 16'(919);
			4950: out = 16'(-2622);
			4951: out = 16'(345);
			4952: out = 16'(-8544);
			4953: out = 16'(-309);
			4954: out = 16'(751);
			4955: out = 16'(-3014);
			4956: out = 16'(-4043);
			4957: out = 16'(-4601);
			4958: out = 16'(2019);
			4959: out = 16'(-881);
			4960: out = 16'(239);
			4961: out = 16'(2001);
			4962: out = 16'(7146);
			4963: out = 16'(1230);
			4964: out = 16'(-3838);
			4965: out = 16'(4932);
			4966: out = 16'(-10964);
			4967: out = 16'(6131);
			4968: out = 16'(-4950);
			4969: out = 16'(94);
			4970: out = 16'(763);
			4971: out = 16'(-7170);
			4972: out = 16'(6054);
			4973: out = 16'(-9510);
			4974: out = 16'(4755);
			4975: out = 16'(-1356);
			4976: out = 16'(-4636);
			4977: out = 16'(-19);
			4978: out = 16'(-5076);
			4979: out = 16'(7476);
			4980: out = 16'(-5913);
			4981: out = 16'(4741);
			4982: out = 16'(3320);
			4983: out = 16'(-8134);
			4984: out = 16'(205);
			4985: out = 16'(2950);
			4986: out = 16'(-1372);
			4987: out = 16'(979);
			4988: out = 16'(-1942);
			4989: out = 16'(-6797);
			4990: out = 16'(5520);
			4991: out = 16'(-12491);
			4992: out = 16'(2179);
			4993: out = 16'(-5214);
			4994: out = 16'(2150);
			4995: out = 16'(-1985);
			4996: out = 16'(-3048);
			4997: out = 16'(-550);
			4998: out = 16'(-1014);
			4999: out = 16'(-352);
			5000: out = 16'(93);
			5001: out = 16'(5813);
			5002: out = 16'(-5205);
			5003: out = 16'(-128);
			5004: out = 16'(-2464);
			5005: out = 16'(-5154);
			5006: out = 16'(3922);
			5007: out = 16'(-1342);
			5008: out = 16'(73);
			5009: out = 16'(766);
			5010: out = 16'(559);
			5011: out = 16'(534);
			5012: out = 16'(197);
			5013: out = 16'(5800);
			5014: out = 16'(3597);
			5015: out = 16'(-2230);
			5016: out = 16'(4244);
			5017: out = 16'(1251);
			5018: out = 16'(-3819);
			5019: out = 16'(533);
			5020: out = 16'(-4277);
			5021: out = 16'(-291);
			5022: out = 16'(316);
			5023: out = 16'(-5399);
			5024: out = 16'(2665);
			5025: out = 16'(-5881);
			5026: out = 16'(366);
			5027: out = 16'(-5280);
			5028: out = 16'(-120);
			5029: out = 16'(1269);
			5030: out = 16'(-16090);
			5031: out = 16'(5096);
			5032: out = 16'(2089);
			5033: out = 16'(3087);
			5034: out = 16'(-450);
			5035: out = 16'(-2766);
			5036: out = 16'(849);
			5037: out = 16'(-1027);
			5038: out = 16'(-245);
			5039: out = 16'(-5037);
			5040: out = 16'(6960);
			5041: out = 16'(-565);
			5042: out = 16'(-2116);
			5043: out = 16'(-4092);
			5044: out = 16'(4376);
			5045: out = 16'(-4610);
			5046: out = 16'(2108);
			5047: out = 16'(1716);
			5048: out = 16'(1219);
			5049: out = 16'(6928);
			5050: out = 16'(-635);
			5051: out = 16'(5624);
			5052: out = 16'(979);
			5053: out = 16'(2987);
			5054: out = 16'(-5979);
			5055: out = 16'(-8463);
			5056: out = 16'(8520);
			5057: out = 16'(-15511);
			5058: out = 16'(9151);
			5059: out = 16'(-7271);
			5060: out = 16'(6068);
			5061: out = 16'(-552);
			5062: out = 16'(-6012);
			5063: out = 16'(202);
			5064: out = 16'(-5159);
			5065: out = 16'(-411);
			5066: out = 16'(-417);
			5067: out = 16'(-3463);
			5068: out = 16'(7016);
			5069: out = 16'(-7627);
			5070: out = 16'(1695);
			5071: out = 16'(1192);
			5072: out = 16'(2597);
			5073: out = 16'(3538);
			5074: out = 16'(-4874);
			5075: out = 16'(-3045);
			5076: out = 16'(4809);
			5077: out = 16'(-2743);
			5078: out = 16'(-1995);
			5079: out = 16'(271);
			5080: out = 16'(-284);
			5081: out = 16'(2986);
			5082: out = 16'(-2122);
			5083: out = 16'(617);
			5084: out = 16'(5943);
			5085: out = 16'(6769);
			5086: out = 16'(-952);
			5087: out = 16'(-5319);
			5088: out = 16'(9853);
			5089: out = 16'(-9229);
			5090: out = 16'(4469);
			5091: out = 16'(-160);
			5092: out = 16'(-1431);
			5093: out = 16'(-847);
			5094: out = 16'(77);
			5095: out = 16'(4509);
			5096: out = 16'(-5041);
			5097: out = 16'(5786);
			5098: out = 16'(-1405);
			5099: out = 16'(-7120);
			5100: out = 16'(4842);
			5101: out = 16'(-10197);
			5102: out = 16'(3168);
			5103: out = 16'(-3079);
			5104: out = 16'(4507);
			5105: out = 16'(-5373);
			5106: out = 16'(-3449);
			5107: out = 16'(-7842);
			5108: out = 16'(-3666);
			5109: out = 16'(-5400);
			5110: out = 16'(6399);
			5111: out = 16'(1480);
			5112: out = 16'(5658);
			5113: out = 16'(3396);
			5114: out = 16'(-9186);
			5115: out = 16'(9486);
			5116: out = 16'(-2280);
			5117: out = 16'(-2994);
			5118: out = 16'(4062);
			5119: out = 16'(-2482);
			5120: out = 16'(3124);
			5121: out = 16'(-2515);
			5122: out = 16'(7442);
			5123: out = 16'(2074);
			5124: out = 16'(2769);
			5125: out = 16'(-1602);
			5126: out = 16'(-4336);
			5127: out = 16'(-515);
			5128: out = 16'(-1709);
			5129: out = 16'(-3918);
			5130: out = 16'(3670);
			5131: out = 16'(2029);
			5132: out = 16'(-139);
			5133: out = 16'(7243);
			5134: out = 16'(-1961);
			5135: out = 16'(1207);
			5136: out = 16'(-119);
			5137: out = 16'(-197);
			5138: out = 16'(1174);
			5139: out = 16'(-94);
			5140: out = 16'(2682);
			5141: out = 16'(-5663);
			5142: out = 16'(2271);
			5143: out = 16'(-2964);
			5144: out = 16'(-440);
			5145: out = 16'(-7559);
			5146: out = 16'(1050);
			5147: out = 16'(3534);
			5148: out = 16'(-8168);
			5149: out = 16'(1758);
			5150: out = 16'(-1779);
			5151: out = 16'(2205);
			5152: out = 16'(1130);
			5153: out = 16'(-4176);
			5154: out = 16'(2422);
			5155: out = 16'(4627);
			5156: out = 16'(2373);
			5157: out = 16'(7201);
			5158: out = 16'(-3488);
			5159: out = 16'(3665);
			5160: out = 16'(-2527);
			5161: out = 16'(-1722);
			5162: out = 16'(-1141);
			5163: out = 16'(1390);
			5164: out = 16'(5104);
			5165: out = 16'(1876);
			5166: out = 16'(-692);
			5167: out = 16'(1490);
			5168: out = 16'(-41);
			5169: out = 16'(-419);
			5170: out = 16'(4481);
			5171: out = 16'(-156);
			5172: out = 16'(3619);
			5173: out = 16'(-3968);
			5174: out = 16'(3454);
			5175: out = 16'(3684);
			5176: out = 16'(2090);
			5177: out = 16'(-1558);
			5178: out = 16'(-2191);
			5179: out = 16'(-1317);
			5180: out = 16'(-9227);
			5181: out = 16'(560);
			5182: out = 16'(-8166);
			5183: out = 16'(-3376);
			5184: out = 16'(2090);
			5185: out = 16'(-4891);
			5186: out = 16'(7604);
			5187: out = 16'(-5017);
			5188: out = 16'(7056);
			5189: out = 16'(-3258);
			5190: out = 16'(-343);
			5191: out = 16'(-1606);
			5192: out = 16'(-5076);
			5193: out = 16'(7632);
			5194: out = 16'(870);
			5195: out = 16'(5754);
			5196: out = 16'(4786);
			5197: out = 16'(-2782);
			5198: out = 16'(3377);
			5199: out = 16'(182);
			5200: out = 16'(1979);
			5201: out = 16'(-1356);
			5202: out = 16'(8387);
			5203: out = 16'(-414);
			5204: out = 16'(1394);
			5205: out = 16'(1655);
			5206: out = 16'(2016);
			5207: out = 16'(123);
			5208: out = 16'(1807);
			5209: out = 16'(2262);
			5210: out = 16'(-5227);
			5211: out = 16'(-2194);
			5212: out = 16'(161);
			5213: out = 16'(697);
			5214: out = 16'(4066);
			5215: out = 16'(480);
			5216: out = 16'(1567);
			5217: out = 16'(3736);
			5218: out = 16'(-3557);
			5219: out = 16'(-10262);
			5220: out = 16'(727);
			5221: out = 16'(-2581);
			5222: out = 16'(-1804);
			5223: out = 16'(-782);
			5224: out = 16'(-1904);
			5225: out = 16'(111);
			5226: out = 16'(-6100);
			5227: out = 16'(-891);
			5228: out = 16'(2848);
			5229: out = 16'(-5631);
			5230: out = 16'(-815);
			5231: out = 16'(-177);
			5232: out = 16'(-4532);
			5233: out = 16'(3905);
			5234: out = 16'(478);
			5235: out = 16'(-199);
			5236: out = 16'(-157);
			5237: out = 16'(2533);
			5238: out = 16'(1710);
			5239: out = 16'(-2842);
			5240: out = 16'(6688);
			5241: out = 16'(3387);
			5242: out = 16'(-4469);
			5243: out = 16'(-1102);
			5244: out = 16'(-536);
			5245: out = 16'(-1982);
			5246: out = 16'(5765);
			5247: out = 16'(1479);
			5248: out = 16'(5900);
			5249: out = 16'(-5044);
			5250: out = 16'(2704);
			5251: out = 16'(-6882);
			5252: out = 16'(4200);
			5253: out = 16'(-3752);
			5254: out = 16'(-4625);
			5255: out = 16'(5759);
			5256: out = 16'(1883);
			5257: out = 16'(3368);
			5258: out = 16'(-129);
			5259: out = 16'(4297);
			5260: out = 16'(2930);
			5261: out = 16'(-4495);
			5262: out = 16'(-5315);
			5263: out = 16'(-8337);
			5264: out = 16'(-1820);
			5265: out = 16'(1037);
			5266: out = 16'(-7391);
			5267: out = 16'(1751);
			5268: out = 16'(1810);
			5269: out = 16'(276);
			5270: out = 16'(-4422);
			5271: out = 16'(-3952);
			5272: out = 16'(-474);
			5273: out = 16'(-2124);
			5274: out = 16'(-3534);
			5275: out = 16'(5838);
			5276: out = 16'(-419);
			5277: out = 16'(12354);
			5278: out = 16'(-8298);
			5279: out = 16'(10871);
			5280: out = 16'(3966);
			5281: out = 16'(-9561);
			5282: out = 16'(-377);
			5283: out = 16'(-151);
			5284: out = 16'(-341);
			5285: out = 16'(-3007);
			5286: out = 16'(1909);
			5287: out = 16'(5176);
			5288: out = 16'(-2796);
			5289: out = 16'(2882);
			5290: out = 16'(-7011);
			5291: out = 16'(874);
			5292: out = 16'(2616);
			5293: out = 16'(429);
			5294: out = 16'(356);
			5295: out = 16'(-2768);
			5296: out = 16'(3716);
			5297: out = 16'(-10111);
			5298: out = 16'(5691);
			5299: out = 16'(1011);
			5300: out = 16'(-3134);
			5301: out = 16'(-4977);
			5302: out = 16'(2799);
			5303: out = 16'(-7005);
			5304: out = 16'(4082);
			5305: out = 16'(-346);
			5306: out = 16'(-6348);
			5307: out = 16'(6644);
			5308: out = 16'(3793);
			5309: out = 16'(1988);
			5310: out = 16'(-3327);
			5311: out = 16'(5266);
			5312: out = 16'(5773);
			5313: out = 16'(-69);
			5314: out = 16'(5199);
			5315: out = 16'(-1384);
			5316: out = 16'(4014);
			5317: out = 16'(3475);
			5318: out = 16'(-215);
			5319: out = 16'(6271);
			5320: out = 16'(-6285);
			5321: out = 16'(5776);
			5322: out = 16'(-2811);
			5323: out = 16'(1385);
			5324: out = 16'(202);
			5325: out = 16'(-4515);
			5326: out = 16'(-1409);
			5327: out = 16'(5264);
			5328: out = 16'(-6703);
			5329: out = 16'(8956);
			5330: out = 16'(-953);
			5331: out = 16'(2253);
			5332: out = 16'(-2490);
			5333: out = 16'(-7253);
			5334: out = 16'(721);
			5335: out = 16'(654);
			5336: out = 16'(-1392);
			5337: out = 16'(0);
			5338: out = 16'(3060);
			5339: out = 16'(6371);
			5340: out = 16'(-4398);
			5341: out = 16'(2333);
			5342: out = 16'(-2442);
			5343: out = 16'(299);
			5344: out = 16'(371);
			5345: out = 16'(-4525);
			5346: out = 16'(2163);
			5347: out = 16'(620);
			5348: out = 16'(-381);
			5349: out = 16'(7086);
			5350: out = 16'(2051);
			5351: out = 16'(2333);
			5352: out = 16'(-8160);
			5353: out = 16'(-3085);
			5354: out = 16'(-912);
			5355: out = 16'(1148);
			5356: out = 16'(4470);
			5357: out = 16'(3308);
			5358: out = 16'(4652);
			5359: out = 16'(-16);
			5360: out = 16'(-7376);
			5361: out = 16'(5272);
			5362: out = 16'(-5943);
			5363: out = 16'(5442);
			5364: out = 16'(-4605);
			5365: out = 16'(-4670);
			5366: out = 16'(1057);
			5367: out = 16'(-2436);
			5368: out = 16'(1783);
			5369: out = 16'(-519);
			5370: out = 16'(699);
			5371: out = 16'(6282);
			5372: out = 16'(-16170);
			5373: out = 16'(7808);
			5374: out = 16'(-1641);
			5375: out = 16'(-1612);
			5376: out = 16'(-3204);
			5377: out = 16'(-2103);
			5378: out = 16'(6631);
			5379: out = 16'(-3985);
			5380: out = 16'(208);
			5381: out = 16'(-5788);
			5382: out = 16'(2362);
			5383: out = 16'(282);
			5384: out = 16'(-5685);
			5385: out = 16'(393);
			5386: out = 16'(2108);
			5387: out = 16'(-116);
			5388: out = 16'(-747);
			5389: out = 16'(5371);
			5390: out = 16'(-2238);
			5391: out = 16'(7750);
			5392: out = 16'(-6066);
			5393: out = 16'(5307);
			5394: out = 16'(-1673);
			5395: out = 16'(678);
			5396: out = 16'(-2655);
			5397: out = 16'(-2352);
			5398: out = 16'(4628);
			5399: out = 16'(-696);
			5400: out = 16'(-652);
			5401: out = 16'(1687);
			5402: out = 16'(3530);
			5403: out = 16'(-74);
			5404: out = 16'(-12600);
			5405: out = 16'(6533);
			5406: out = 16'(-8225);
			5407: out = 16'(6027);
			5408: out = 16'(-19);
			5409: out = 16'(4961);
			5410: out = 16'(4422);
			5411: out = 16'(-1641);
			5412: out = 16'(1567);
			5413: out = 16'(2635);
			5414: out = 16'(-874);
			5415: out = 16'(-5534);
			5416: out = 16'(2920);
			5417: out = 16'(-5112);
			5418: out = 16'(1483);
			5419: out = 16'(-4178);
			5420: out = 16'(1129);
			5421: out = 16'(8276);
			5422: out = 16'(-84);
			5423: out = 16'(273);
			5424: out = 16'(-4273);
			5425: out = 16'(-1651);
			5426: out = 16'(3122);
			5427: out = 16'(3696);
			5428: out = 16'(3314);
			5429: out = 16'(1342);
			5430: out = 16'(3525);
			5431: out = 16'(-2148);
			5432: out = 16'(1715);
			5433: out = 16'(1187);
			5434: out = 16'(229);
			5435: out = 16'(3533);
			5436: out = 16'(-1065);
			5437: out = 16'(694);
			5438: out = 16'(-6355);
			5439: out = 16'(-429);
			5440: out = 16'(-3304);
			5441: out = 16'(-5194);
			5442: out = 16'(176);
			5443: out = 16'(946);
			5444: out = 16'(-4429);
			5445: out = 16'(6083);
			5446: out = 16'(-8040);
			5447: out = 16'(3562);
			5448: out = 16'(-3698);
			5449: out = 16'(-3721);
			5450: out = 16'(2782);
			5451: out = 16'(1493);
			5452: out = 16'(4667);
			5453: out = 16'(-2008);
			5454: out = 16'(-1746);
			5455: out = 16'(137);
			5456: out = 16'(-9215);
			5457: out = 16'(6495);
			5458: out = 16'(2769);
			5459: out = 16'(2181);
			5460: out = 16'(96);
			5461: out = 16'(1476);
			5462: out = 16'(45);
			5463: out = 16'(-128);
			5464: out = 16'(1046);
			5465: out = 16'(-3205);
			5466: out = 16'(-1552);
			5467: out = 16'(779);
			5468: out = 16'(-3817);
			5469: out = 16'(-223);
			5470: out = 16'(-4493);
			5471: out = 16'(5896);
			5472: out = 16'(-3594);
			5473: out = 16'(-1902);
			5474: out = 16'(-4967);
			5475: out = 16'(1900);
			5476: out = 16'(-8797);
			5477: out = 16'(7572);
			5478: out = 16'(-2470);
			5479: out = 16'(3662);
			5480: out = 16'(3253);
			5481: out = 16'(1567);
			5482: out = 16'(4489);
			5483: out = 16'(3974);
			5484: out = 16'(622);
			5485: out = 16'(-659);
			5486: out = 16'(-617);
			5487: out = 16'(3592);
			5488: out = 16'(-8679);
			5489: out = 16'(8022);
			5490: out = 16'(-5597);
			5491: out = 16'(5941);
			5492: out = 16'(-6087);
			5493: out = 16'(1604);
			5494: out = 16'(-174);
			5495: out = 16'(-2794);
			5496: out = 16'(6170);
			5497: out = 16'(-8694);
			5498: out = 16'(-689);
			5499: out = 16'(2007);
			5500: out = 16'(-2778);
			5501: out = 16'(-4521);
			5502: out = 16'(-4737);
			5503: out = 16'(1875);
			5504: out = 16'(188);
			5505: out = 16'(2330);
			5506: out = 16'(1087);
			5507: out = 16'(-1169);
			5508: out = 16'(460);
			5509: out = 16'(-4479);
			5510: out = 16'(2058);
			5511: out = 16'(1794);
			5512: out = 16'(-1347);
			5513: out = 16'(5935);
			5514: out = 16'(3432);
			5515: out = 16'(-5380);
			5516: out = 16'(367);
			5517: out = 16'(-491);
			5518: out = 16'(-1469);
			5519: out = 16'(2515);
			5520: out = 16'(-1240);
			5521: out = 16'(353);
			5522: out = 16'(95);
			5523: out = 16'(2968);
			5524: out = 16'(-4829);
			5525: out = 16'(2740);
			5526: out = 16'(23);
			5527: out = 16'(-3800);
			5528: out = 16'(-4638);
			5529: out = 16'(5860);
			5530: out = 16'(-3603);
			5531: out = 16'(9614);
			5532: out = 16'(1687);
			5533: out = 16'(-3853);
			5534: out = 16'(-3407);
			5535: out = 16'(2167);
			5536: out = 16'(-3358);
			5537: out = 16'(-2807);
			5538: out = 16'(3937);
			5539: out = 16'(3065);
			5540: out = 16'(-7234);
			5541: out = 16'(9819);
			5542: out = 16'(-13728);
			5543: out = 16'(7044);
			5544: out = 16'(-1751);
			5545: out = 16'(-23);
			5546: out = 16'(3964);
			5547: out = 16'(1070);
			5548: out = 16'(5141);
			5549: out = 16'(-1769);
			5550: out = 16'(2770);
			5551: out = 16'(-1995);
			5552: out = 16'(-2724);
			5553: out = 16'(1699);
			5554: out = 16'(-4048);
			5555: out = 16'(3494);
			5556: out = 16'(-1075);
			5557: out = 16'(-2266);
			5558: out = 16'(2725);
			5559: out = 16'(13);
			5560: out = 16'(-2587);
			5561: out = 16'(-396);
			5562: out = 16'(2339);
			5563: out = 16'(2744);
			5564: out = 16'(-7125);
			5565: out = 16'(3423);
			5566: out = 16'(-1838);
			5567: out = 16'(-8071);
			5568: out = 16'(-45);
			5569: out = 16'(-7128);
			5570: out = 16'(8595);
			5571: out = 16'(-1131);
			5572: out = 16'(-6211);
			5573: out = 16'(6808);
			5574: out = 16'(362);
			5575: out = 16'(3955);
			5576: out = 16'(-7778);
			5577: out = 16'(-2891);
			5578: out = 16'(697);
			5579: out = 16'(15);
			5580: out = 16'(3109);
			5581: out = 16'(219);
			5582: out = 16'(2967);
			5583: out = 16'(-830);
			5584: out = 16'(-2574);
			5585: out = 16'(4528);
			5586: out = 16'(-11982);
			5587: out = 16'(-152);
			5588: out = 16'(-6644);
			5589: out = 16'(-128);
			5590: out = 16'(718);
			5591: out = 16'(-604);
			5592: out = 16'(-4069);
			5593: out = 16'(4813);
			5594: out = 16'(1539);
			5595: out = 16'(-2633);
			5596: out = 16'(-8962);
			5597: out = 16'(1987);
			5598: out = 16'(2461);
			5599: out = 16'(-4098);
			5600: out = 16'(3886);
			5601: out = 16'(2007);
			5602: out = 16'(22);
			5603: out = 16'(148);
			5604: out = 16'(-2797);
			5605: out = 16'(2124);
			5606: out = 16'(2316);
			5607: out = 16'(3081);
			5608: out = 16'(1404);
			5609: out = 16'(5071);
			5610: out = 16'(8126);
			5611: out = 16'(-4161);
			5612: out = 16'(2841);
			5613: out = 16'(1063);
			5614: out = 16'(709);
			5615: out = 16'(-194);
			5616: out = 16'(-804);
			5617: out = 16'(2);
			5618: out = 16'(-8347);
			5619: out = 16'(990);
			5620: out = 16'(-3679);
			5621: out = 16'(-6257);
			5622: out = 16'(5915);
			5623: out = 16'(-14790);
			5624: out = 16'(836);
			5625: out = 16'(3150);
			5626: out = 16'(-9352);
			5627: out = 16'(5610);
			5628: out = 16'(-3972);
			5629: out = 16'(6733);
			5630: out = 16'(-656);
			5631: out = 16'(-4061);
			5632: out = 16'(10369);
			5633: out = 16'(-202);
			5634: out = 16'(1629);
			5635: out = 16'(2678);
			5636: out = 16'(-2922);
			5637: out = 16'(0);
			5638: out = 16'(-3522);
			5639: out = 16'(30);
			5640: out = 16'(-76);
			5641: out = 16'(1413);
			5642: out = 16'(-1934);
			5643: out = 16'(1122);
			5644: out = 16'(4392);
			5645: out = 16'(3153);
			5646: out = 16'(1397);
			5647: out = 16'(199);
			5648: out = 16'(-6724);
			5649: out = 16'(3531);
			5650: out = 16'(-2515);
			5651: out = 16'(1538);
			5652: out = 16'(2694);
			5653: out = 16'(849);
			5654: out = 16'(1927);
			5655: out = 16'(-1447);
			5656: out = 16'(-7223);
			5657: out = 16'(3719);
			5658: out = 16'(-3229);
			5659: out = 16'(2902);
			5660: out = 16'(-1199);
			5661: out = 16'(5930);
			5662: out = 16'(-831);
			5663: out = 16'(3076);
			5664: out = 16'(4601);
			5665: out = 16'(712);
			5666: out = 16'(-2559);
			5667: out = 16'(-2405);
			5668: out = 16'(-914);
			5669: out = 16'(1878);
			5670: out = 16'(-6791);
			5671: out = 16'(2372);
			5672: out = 16'(35);
			5673: out = 16'(2725);
			5674: out = 16'(1430);
			5675: out = 16'(-3388);
			5676: out = 16'(-105);
			5677: out = 16'(2416);
			5678: out = 16'(54);
			5679: out = 16'(3128);
			5680: out = 16'(-3044);
			5681: out = 16'(599);
			5682: out = 16'(-1976);
			5683: out = 16'(3342);
			5684: out = 16'(6738);
			5685: out = 16'(2810);
			5686: out = 16'(4995);
			5687: out = 16'(-829);
			5688: out = 16'(2332);
			5689: out = 16'(-1769);
			5690: out = 16'(-2778);
			5691: out = 16'(4439);
			5692: out = 16'(-4868);
			5693: out = 16'(33);
			5694: out = 16'(4593);
			5695: out = 16'(-356);
			5696: out = 16'(5486);
			5697: out = 16'(-6800);
			5698: out = 16'(1643);
			5699: out = 16'(-531);
			5700: out = 16'(-382);
			5701: out = 16'(2010);
			5702: out = 16'(401);
			5703: out = 16'(9119);
			5704: out = 16'(1174);
			5705: out = 16'(-4961);
			5706: out = 16'(1226);
			5707: out = 16'(-1563);
			5708: out = 16'(-1054);
			5709: out = 16'(643);
			5710: out = 16'(646);
			5711: out = 16'(1631);
			5712: out = 16'(-3410);
			5713: out = 16'(1459);
			5714: out = 16'(-5002);
			5715: out = 16'(1842);
			5716: out = 16'(622);
			5717: out = 16'(-3474);
			5718: out = 16'(2116);
			5719: out = 16'(-1278);
			5720: out = 16'(-167);
			5721: out = 16'(-982);
			5722: out = 16'(44);
			5723: out = 16'(5070);
			5724: out = 16'(574);
			5725: out = 16'(-451);
			5726: out = 16'(2067);
			5727: out = 16'(7252);
			5728: out = 16'(-4323);
			5729: out = 16'(5289);
			5730: out = 16'(490);
			5731: out = 16'(1356);
			5732: out = 16'(1683);
			5733: out = 16'(254);
			5734: out = 16'(-592);
			5735: out = 16'(5981);
			5736: out = 16'(463);
			5737: out = 16'(-479);
			5738: out = 16'(-1983);
			5739: out = 16'(3900);
			5740: out = 16'(-3206);
			5741: out = 16'(2071);
			5742: out = 16'(2);
			5743: out = 16'(9130);
			5744: out = 16'(-4175);
			5745: out = 16'(3027);
			5746: out = 16'(-1079);
			5747: out = 16'(1374);
			5748: out = 16'(2090);
			5749: out = 16'(-378);
			5750: out = 16'(1509);
			5751: out = 16'(-2156);
			5752: out = 16'(-9537);
			5753: out = 16'(2502);
			5754: out = 16'(-4850);
			5755: out = 16'(2776);
			5756: out = 16'(-6327);
			5757: out = 16'(-1185);
			5758: out = 16'(-1263);
			5759: out = 16'(-8958);
			5760: out = 16'(3852);
			5761: out = 16'(-4920);
			5762: out = 16'(447);
			5763: out = 16'(1755);
			5764: out = 16'(-4283);
			5765: out = 16'(6061);
			5766: out = 16'(-107);
			5767: out = 16'(2525);
			5768: out = 16'(5517);
			5769: out = 16'(-2272);
			5770: out = 16'(-1206);
			5771: out = 16'(-1084);
			5772: out = 16'(5813);
			5773: out = 16'(739);
			5774: out = 16'(2945);
			5775: out = 16'(-173);
			5776: out = 16'(-4639);
			5777: out = 16'(110);
			5778: out = 16'(278);
			5779: out = 16'(-663);
			5780: out = 16'(-240);
			5781: out = 16'(-4681);
			5782: out = 16'(614);
			5783: out = 16'(-58);
			5784: out = 16'(764);
			5785: out = 16'(4136);
			5786: out = 16'(-2874);
			5787: out = 16'(3965);
			5788: out = 16'(-2515);
			5789: out = 16'(-1622);
			5790: out = 16'(-3105);
			5791: out = 16'(-5892);
			5792: out = 16'(-144);
			5793: out = 16'(4489);
			5794: out = 16'(-1905);
			5795: out = 16'(1097);
			5796: out = 16'(-1456);
			5797: out = 16'(4642);
			5798: out = 16'(-5956);
			5799: out = 16'(6552);
			5800: out = 16'(-4432);
			5801: out = 16'(3600);
			5802: out = 16'(-672);
			5803: out = 16'(-7871);
			5804: out = 16'(3089);
			5805: out = 16'(4837);
			5806: out = 16'(2026);
			5807: out = 16'(3635);
			5808: out = 16'(2366);
			5809: out = 16'(105);
			5810: out = 16'(21);
			5811: out = 16'(-127);
			5812: out = 16'(2515);
			5813: out = 16'(1661);
			5814: out = 16'(1446);
			5815: out = 16'(1129);
			5816: out = 16'(-6065);
			5817: out = 16'(6412);
			5818: out = 16'(-5150);
			5819: out = 16'(-4383);
			5820: out = 16'(3485);
			5821: out = 16'(-7192);
			5822: out = 16'(2546);
			5823: out = 16'(5530);
			5824: out = 16'(7459);
			5825: out = 16'(-3097);
			5826: out = 16'(-1916);
			5827: out = 16'(-6905);
			5828: out = 16'(-9586);
			5829: out = 16'(552);
			5830: out = 16'(-3210);
			5831: out = 16'(-1594);
			5832: out = 16'(4285);
			5833: out = 16'(-5560);
			5834: out = 16'(-1381);
			5835: out = 16'(21);
			5836: out = 16'(-277);
			5837: out = 16'(1029);
			5838: out = 16'(-2407);
			5839: out = 16'(2378);
			5840: out = 16'(-11060);
			5841: out = 16'(4657);
			5842: out = 16'(-3911);
			5843: out = 16'(1147);
			5844: out = 16'(4160);
			5845: out = 16'(-1598);
			5846: out = 16'(2151);
			5847: out = 16'(2756);
			5848: out = 16'(-3004);
			5849: out = 16'(9100);
			5850: out = 16'(-6826);
			5851: out = 16'(2548);
			5852: out = 16'(-2220);
			5853: out = 16'(510);
			5854: out = 16'(578);
			5855: out = 16'(3);
			5856: out = 16'(2262);
			5857: out = 16'(1564);
			5858: out = 16'(-1335);
			5859: out = 16'(5366);
			5860: out = 16'(-7535);
			5861: out = 16'(-178);
			5862: out = 16'(-318);
			5863: out = 16'(-666);
			5864: out = 16'(921);
			5865: out = 16'(3336);
			5866: out = 16'(2690);
			5867: out = 16'(-563);
			5868: out = 16'(1538);
			5869: out = 16'(1147);
			5870: out = 16'(-2674);
			5871: out = 16'(213);
			5872: out = 16'(-3874);
			5873: out = 16'(-3451);
			5874: out = 16'(-871);
			5875: out = 16'(-963);
			5876: out = 16'(7063);
			5877: out = 16'(-438);
			5878: out = 16'(321);
			5879: out = 16'(-4313);
			5880: out = 16'(-566);
			5881: out = 16'(1723);
			5882: out = 16'(-6388);
			5883: out = 16'(8654);
			5884: out = 16'(-308);
			5885: out = 16'(3952);
			5886: out = 16'(5172);
			5887: out = 16'(-4813);
			5888: out = 16'(3951);
			5889: out = 16'(4950);
			5890: out = 16'(-4981);
			5891: out = 16'(3102);
			5892: out = 16'(-384);
			5893: out = 16'(4467);
			5894: out = 16'(2388);
			5895: out = 16'(-1662);
			5896: out = 16'(1938);
			5897: out = 16'(-792);
			5898: out = 16'(676);
			5899: out = 16'(-3359);
			5900: out = 16'(-3103);
			5901: out = 16'(6802);
			5902: out = 16'(-5674);
			5903: out = 16'(1089);
			5904: out = 16'(4955);
			5905: out = 16'(-2850);
			5906: out = 16'(-259);
			5907: out = 16'(-119);
			5908: out = 16'(6636);
			5909: out = 16'(-2888);
			5910: out = 16'(885);
			5911: out = 16'(-1479);
			5912: out = 16'(-220);
			5913: out = 16'(1837);
			5914: out = 16'(-3490);
			5915: out = 16'(1793);
			5916: out = 16'(-3093);
			5917: out = 16'(4386);
			5918: out = 16'(293);
			5919: out = 16'(-11338);
			5920: out = 16'(3308);
			5921: out = 16'(-2523);
			5922: out = 16'(4956);
			5923: out = 16'(3044);
			5924: out = 16'(1108);
			5925: out = 16'(4413);
			5926: out = 16'(-1778);
			5927: out = 16'(-1409);
			5928: out = 16'(7001);
			5929: out = 16'(885);
			5930: out = 16'(-2988);
			5931: out = 16'(1923);
			5932: out = 16'(-1569);
			5933: out = 16'(7219);
			5934: out = 16'(-287);
			5935: out = 16'(456);
			5936: out = 16'(1306);
			5937: out = 16'(-3558);
			5938: out = 16'(-7005);
			5939: out = 16'(4195);
			5940: out = 16'(-1477);
			5941: out = 16'(661);
			5942: out = 16'(48);
			5943: out = 16'(661);
			5944: out = 16'(-8389);
			5945: out = 16'(4479);
			5946: out = 16'(4468);
			5947: out = 16'(3169);
			5948: out = 16'(-221);
			5949: out = 16'(2451);
			5950: out = 16'(-4584);
			5951: out = 16'(4740);
			5952: out = 16'(3376);
			5953: out = 16'(4588);
			5954: out = 16'(-3261);
			5955: out = 16'(1078);
			5956: out = 16'(-1883);
			5957: out = 16'(-2136);
			5958: out = 16'(1209);
			5959: out = 16'(472);
			5960: out = 16'(4073);
			5961: out = 16'(-2347);
			5962: out = 16'(-2640);
			5963: out = 16'(498);
			5964: out = 16'(-1142);
			5965: out = 16'(5897);
			5966: out = 16'(-639);
			5967: out = 16'(5694);
			5968: out = 16'(-7604);
			5969: out = 16'(53);
			5970: out = 16'(5873);
			5971: out = 16'(-7400);
			5972: out = 16'(2541);
			5973: out = 16'(-1835);
			5974: out = 16'(-506);
			5975: out = 16'(4602);
			5976: out = 16'(-5365);
			5977: out = 16'(3756);
			5978: out = 16'(3953);
			5979: out = 16'(-59);
			5980: out = 16'(-3003);
			5981: out = 16'(-73);
			5982: out = 16'(-745);
			5983: out = 16'(-3228);
			5984: out = 16'(751);
			5985: out = 16'(1990);
			5986: out = 16'(1706);
			5987: out = 16'(261);
			5988: out = 16'(5109);
			5989: out = 16'(-2333);
			5990: out = 16'(1154);
			5991: out = 16'(3762);
			5992: out = 16'(-5856);
			5993: out = 16'(1094);
			5994: out = 16'(1453);
			5995: out = 16'(-930);
			5996: out = 16'(1088);
			5997: out = 16'(4499);
			5998: out = 16'(-2068);
			5999: out = 16'(-1801);
			6000: out = 16'(-9489);
			6001: out = 16'(-2255);
			6002: out = 16'(-1139);
			6003: out = 16'(-163);
			6004: out = 16'(3692);
			6005: out = 16'(1191);
			6006: out = 16'(2867);
			6007: out = 16'(-6101);
			6008: out = 16'(-5765);
			6009: out = 16'(3402);
			6010: out = 16'(-68);
			6011: out = 16'(1201);
			6012: out = 16'(-4);
			6013: out = 16'(2650);
			6014: out = 16'(-2624);
			6015: out = 16'(3471);
			6016: out = 16'(-6913);
			6017: out = 16'(5420);
			6018: out = 16'(-703);
			6019: out = 16'(-2924);
			6020: out = 16'(-5942);
			6021: out = 16'(-61);
			6022: out = 16'(-1405);
			6023: out = 16'(705);
			6024: out = 16'(249);
			6025: out = 16'(-3524);
			6026: out = 16'(1608);
			6027: out = 16'(1913);
			6028: out = 16'(-7894);
			6029: out = 16'(3562);
			6030: out = 16'(-336);
			6031: out = 16'(-755);
			6032: out = 16'(-530);
			6033: out = 16'(1714);
			6034: out = 16'(-957);
			6035: out = 16'(-5089);
			6036: out = 16'(4927);
			6037: out = 16'(-901);
			6038: out = 16'(4371);
			6039: out = 16'(-3203);
			6040: out = 16'(5388);
			6041: out = 16'(-1308);
			6042: out = 16'(-1601);
			6043: out = 16'(-268);
			6044: out = 16'(-1082);
			6045: out = 16'(-77);
			6046: out = 16'(976);
			6047: out = 16'(-3910);
			6048: out = 16'(4433);
			6049: out = 16'(1821);
			6050: out = 16'(130);
			6051: out = 16'(1684);
			6052: out = 16'(-4254);
			6053: out = 16'(1179);
			6054: out = 16'(3283);
			6055: out = 16'(-206);
			6056: out = 16'(4608);
			6057: out = 16'(5898);
			6058: out = 16'(-1604);
			6059: out = 16'(-5742);
			6060: out = 16'(205);
			6061: out = 16'(-1359);
			6062: out = 16'(-538);
			6063: out = 16'(440);
			6064: out = 16'(-6941);
			6065: out = 16'(4394);
			6066: out = 16'(-3412);
			6067: out = 16'(3109);
			6068: out = 16'(6104);
			6069: out = 16'(712);
			6070: out = 16'(-4451);
			6071: out = 16'(-421);
			6072: out = 16'(284);
			6073: out = 16'(293);
			6074: out = 16'(-508);
			6075: out = 16'(4790);
			6076: out = 16'(1883);
			6077: out = 16'(-4193);
			6078: out = 16'(1659);
			6079: out = 16'(-1491);
			6080: out = 16'(235);
			6081: out = 16'(1311);
			6082: out = 16'(-366);
			6083: out = 16'(3230);
			6084: out = 16'(1368);
			6085: out = 16'(-1610);
			6086: out = 16'(502);
			6087: out = 16'(-4651);
			6088: out = 16'(3637);
			6089: out = 16'(-3746);
			6090: out = 16'(4943);
			6091: out = 16'(-6540);
			6092: out = 16'(2042);
			6093: out = 16'(-3970);
			6094: out = 16'(-2393);
			6095: out = 16'(291);
			6096: out = 16'(684);
			6097: out = 16'(-463);
			6098: out = 16'(-993);
			6099: out = 16'(-154);
			6100: out = 16'(2732);
			6101: out = 16'(-8736);
			6102: out = 16'(-163);
			6103: out = 16'(-1060);
			6104: out = 16'(-5297);
			6105: out = 16'(3097);
			6106: out = 16'(4674);
			6107: out = 16'(1853);
			6108: out = 16'(4174);
			6109: out = 16'(-5644);
			6110: out = 16'(1544);
			6111: out = 16'(-5105);
			6112: out = 16'(-1952);
			6113: out = 16'(3745);
			6114: out = 16'(-1484);
			6115: out = 16'(3484);
			6116: out = 16'(-2191);
			6117: out = 16'(-103);
			6118: out = 16'(-3310);
			6119: out = 16'(-3426);
			6120: out = 16'(446);
			6121: out = 16'(-7114);
			6122: out = 16'(430);
			6123: out = 16'(-4809);
			6124: out = 16'(5148);
			6125: out = 16'(1614);
			6126: out = 16'(4534);
			6127: out = 16'(-162);
			6128: out = 16'(-1128);
			6129: out = 16'(-690);
			6130: out = 16'(-5472);
			6131: out = 16'(122);
			6132: out = 16'(3694);
			6133: out = 16'(1883);
			6134: out = 16'(-401);
			6135: out = 16'(-91);
			6136: out = 16'(-6374);
			6137: out = 16'(1677);
			6138: out = 16'(1566);
			6139: out = 16'(-5093);
			6140: out = 16'(1590);
			6141: out = 16'(5063);
			6142: out = 16'(-4224);
			6143: out = 16'(-5082);
			6144: out = 16'(2321);
			6145: out = 16'(2545);
			6146: out = 16'(-4892);
			6147: out = 16'(4358);
			6148: out = 16'(-2521);
			6149: out = 16'(1393);
			6150: out = 16'(-841);
			6151: out = 16'(-324);
			6152: out = 16'(790);
			6153: out = 16'(2848);
			6154: out = 16'(-5077);
			6155: out = 16'(-5901);
			6156: out = 16'(-675);
			6157: out = 16'(-1118);
			6158: out = 16'(2278);
			6159: out = 16'(553);
			6160: out = 16'(-295);
			6161: out = 16'(-2630);
			6162: out = 16'(-951);
			6163: out = 16'(-3971);
			6164: out = 16'(-5571);
			6165: out = 16'(6525);
			6166: out = 16'(515);
			6167: out = 16'(1497);
			6168: out = 16'(-181);
			6169: out = 16'(1602);
			6170: out = 16'(-2678);
			6171: out = 16'(-4394);
			6172: out = 16'(6093);
			6173: out = 16'(-7875);
			6174: out = 16'(6611);
			6175: out = 16'(-9484);
			6176: out = 16'(8338);
			6177: out = 16'(1804);
			6178: out = 16'(1653);
			6179: out = 16'(-822);
			6180: out = 16'(-4409);
			6181: out = 16'(-708);
			6182: out = 16'(-2227);
			6183: out = 16'(-957);
			6184: out = 16'(1741);
			6185: out = 16'(-5642);
			6186: out = 16'(1652);
			6187: out = 16'(-3160);
			6188: out = 16'(649);
			6189: out = 16'(-382);
			6190: out = 16'(610);
			6191: out = 16'(1102);
			6192: out = 16'(112);
			6193: out = 16'(-4935);
			6194: out = 16'(-1845);
			6195: out = 16'(4984);
			6196: out = 16'(-111);
			6197: out = 16'(1991);
			6198: out = 16'(-1031);
			6199: out = 16'(-3316);
			6200: out = 16'(-382);
			6201: out = 16'(2193);
			6202: out = 16'(-4192);
			6203: out = 16'(380);
			6204: out = 16'(135);
			6205: out = 16'(489);
			6206: out = 16'(-4812);
			6207: out = 16'(-809);
			6208: out = 16'(-3215);
			6209: out = 16'(1870);
			6210: out = 16'(-129);
			6211: out = 16'(-2513);
			6212: out = 16'(-5892);
			6213: out = 16'(-4762);
			6214: out = 16'(-5711);
			6215: out = 16'(2661);
			6216: out = 16'(-1007);
			6217: out = 16'(-2149);
			6218: out = 16'(1030);
			6219: out = 16'(3536);
			6220: out = 16'(-3135);
			6221: out = 16'(2360);
			6222: out = 16'(3619);
			6223: out = 16'(-2990);
			6224: out = 16'(177);
			6225: out = 16'(2055);
			6226: out = 16'(180);
			6227: out = 16'(1443);
			6228: out = 16'(7348);
			6229: out = 16'(210);
			6230: out = 16'(2764);
			6231: out = 16'(1470);
			6232: out = 16'(-7817);
			6233: out = 16'(-1550);
			6234: out = 16'(3802);
			6235: out = 16'(137);
			6236: out = 16'(4927);
			6237: out = 16'(2890);
			6238: out = 16'(-699);
			6239: out = 16'(-5662);
			6240: out = 16'(2499);
			6241: out = 16'(-5456);
			6242: out = 16'(771);
			6243: out = 16'(348);
			6244: out = 16'(-2961);
			6245: out = 16'(-2148);
			6246: out = 16'(3430);
			6247: out = 16'(-2869);
			6248: out = 16'(-661);
			6249: out = 16'(1596);
			6250: out = 16'(2042);
			6251: out = 16'(-2928);
			6252: out = 16'(1337);
			6253: out = 16'(4404);
			6254: out = 16'(2683);
			6255: out = 16'(410);
			6256: out = 16'(-3408);
			6257: out = 16'(1714);
			6258: out = 16'(6580);
			6259: out = 16'(-2226);
			6260: out = 16'(7168);
			6261: out = 16'(-196);
			6262: out = 16'(3926);
			6263: out = 16'(961);
			6264: out = 16'(-7241);
			6265: out = 16'(-603);
			6266: out = 16'(-839);
			6267: out = 16'(4213);
			6268: out = 16'(-3998);
			6269: out = 16'(1920);
			6270: out = 16'(3598);
			6271: out = 16'(-3384);
			6272: out = 16'(-375);
			6273: out = 16'(-4461);
			6274: out = 16'(1650);
			6275: out = 16'(-2634);
			6276: out = 16'(286);
			6277: out = 16'(235);
			6278: out = 16'(-19);
			6279: out = 16'(2661);
			6280: out = 16'(-2732);
			6281: out = 16'(-2280);
			6282: out = 16'(-540);
			6283: out = 16'(-5571);
			6284: out = 16'(-981);
			6285: out = 16'(1176);
			6286: out = 16'(-692);
			6287: out = 16'(-577);
			6288: out = 16'(2624);
			6289: out = 16'(-1629);
			6290: out = 16'(1759);
			6291: out = 16'(-6146);
			6292: out = 16'(1704);
			6293: out = 16'(707);
			6294: out = 16'(-376);
			6295: out = 16'(-2458);
			6296: out = 16'(-3275);
			6297: out = 16'(-2410);
			6298: out = 16'(3255);
			6299: out = 16'(-6147);
			6300: out = 16'(7505);
			6301: out = 16'(-2540);
			6302: out = 16'(272);
			6303: out = 16'(-3968);
			6304: out = 16'(-1357);
			6305: out = 16'(2088);
			6306: out = 16'(1237);
			6307: out = 16'(5155);
			6308: out = 16'(-1949);
			6309: out = 16'(-2050);
			6310: out = 16'(-456);
			6311: out = 16'(-8383);
			6312: out = 16'(5916);
			6313: out = 16'(-5053);
			6314: out = 16'(4164);
			6315: out = 16'(1439);
			6316: out = 16'(-551);
			6317: out = 16'(-391);
			6318: out = 16'(-4857);
			6319: out = 16'(1617);
			6320: out = 16'(1028);
			6321: out = 16'(2119);
			6322: out = 16'(-589);
			6323: out = 16'(-1979);
			6324: out = 16'(6193);
			6325: out = 16'(-5831);
			6326: out = 16'(-3322);
			6327: out = 16'(-4162);
			6328: out = 16'(-2444);
			6329: out = 16'(-477);
			6330: out = 16'(-2628);
			6331: out = 16'(7192);
			6332: out = 16'(-462);
			6333: out = 16'(373);
			6334: out = 16'(-8239);
			6335: out = 16'(-1685);
			6336: out = 16'(-3953);
			6337: out = 16'(3914);
			6338: out = 16'(-1368);
			6339: out = 16'(4564);
			6340: out = 16'(2462);
			6341: out = 16'(-1967);
			6342: out = 16'(845);
			6343: out = 16'(1557);
			6344: out = 16'(1777);
			6345: out = 16'(-1068);
			6346: out = 16'(-224);
			6347: out = 16'(215);
			6348: out = 16'(2255);
			6349: out = 16'(3536);
			6350: out = 16'(804);
			6351: out = 16'(1953);
			6352: out = 16'(1322);
			6353: out = 16'(-6034);
			6354: out = 16'(-1421);
			6355: out = 16'(4566);
			6356: out = 16'(3011);
			6357: out = 16'(-1909);
			6358: out = 16'(1319);
			6359: out = 16'(3120);
			6360: out = 16'(3405);
			6361: out = 16'(-6660);
			6362: out = 16'(1086);
			6363: out = 16'(598);
			6364: out = 16'(6994);
			6365: out = 16'(-1563);
			6366: out = 16'(-310);
			6367: out = 16'(3791);
			6368: out = 16'(-179);
			6369: out = 16'(5372);
			6370: out = 16'(102);
			6371: out = 16'(-36);
			6372: out = 16'(5870);
			6373: out = 16'(-3762);
			6374: out = 16'(-180);
			6375: out = 16'(-4814);
			6376: out = 16'(4246);
			6377: out = 16'(967);
			6378: out = 16'(-4734);
			6379: out = 16'(5121);
			6380: out = 16'(-2442);
			6381: out = 16'(3051);
			6382: out = 16'(897);
			6383: out = 16'(1394);
			6384: out = 16'(4360);
			6385: out = 16'(-375);
			6386: out = 16'(2538);
			6387: out = 16'(-4771);
			6388: out = 16'(1080);
			6389: out = 16'(-1768);
			6390: out = 16'(-113);
			6391: out = 16'(3274);
			6392: out = 16'(-4532);
			6393: out = 16'(5116);
			6394: out = 16'(-2786);
			6395: out = 16'(-2491);
			6396: out = 16'(545);
			6397: out = 16'(-4701);
			6398: out = 16'(6891);
			6399: out = 16'(-337);
			6400: out = 16'(-382);
			6401: out = 16'(5096);
			6402: out = 16'(631);
			6403: out = 16'(1948);
			6404: out = 16'(-3199);
			6405: out = 16'(560);
			6406: out = 16'(-2359);
			6407: out = 16'(1741);
			6408: out = 16'(3898);
			6409: out = 16'(-2363);
			6410: out = 16'(4682);
			6411: out = 16'(-3242);
			6412: out = 16'(752);
			6413: out = 16'(-5620);
			6414: out = 16'(3503);
			6415: out = 16'(2036);
			6416: out = 16'(-1532);
			6417: out = 16'(3133);
			6418: out = 16'(-3708);
			6419: out = 16'(-1926);
			6420: out = 16'(-1175);
			6421: out = 16'(3440);
			6422: out = 16'(1409);
			6423: out = 16'(373);
			6424: out = 16'(-353);
			6425: out = 16'(133);
			6426: out = 16'(1694);
			6427: out = 16'(-5146);
			6428: out = 16'(533);
			6429: out = 16'(3435);
			6430: out = 16'(-1174);
			6431: out = 16'(-3426);
			6432: out = 16'(575);
			6433: out = 16'(-705);
			6434: out = 16'(6421);
			6435: out = 16'(-1423);
			6436: out = 16'(4635);
			6437: out = 16'(-800);
			6438: out = 16'(177);
			6439: out = 16'(334);
			6440: out = 16'(1820);
			6441: out = 16'(2970);
			6442: out = 16'(2747);
			6443: out = 16'(240);
			6444: out = 16'(-1170);
			6445: out = 16'(-2618);
			6446: out = 16'(2720);
			6447: out = 16'(-2041);
			6448: out = 16'(1239);
			6449: out = 16'(-1276);
			6450: out = 16'(527);
			6451: out = 16'(-861);
			6452: out = 16'(1824);
			6453: out = 16'(1119);
			6454: out = 16'(-41);
			6455: out = 16'(3443);
			6456: out = 16'(-5054);
			6457: out = 16'(-4772);
			6458: out = 16'(309);
			6459: out = 16'(-6710);
			6460: out = 16'(1932);
			6461: out = 16'(1893);
			6462: out = 16'(-3769);
			6463: out = 16'(-327);
			6464: out = 16'(332);
			6465: out = 16'(-1008);
			6466: out = 16'(-8093);
			6467: out = 16'(6190);
			6468: out = 16'(1282);
			6469: out = 16'(-3795);
			6470: out = 16'(4484);
			6471: out = 16'(-154);
			6472: out = 16'(327);
			6473: out = 16'(-648);
			6474: out = 16'(702);
			6475: out = 16'(-5203);
			6476: out = 16'(-4336);
			6477: out = 16'(5121);
			6478: out = 16'(-1254);
			6479: out = 16'(1262);
			6480: out = 16'(-1832);
			6481: out = 16'(-2128);
			6482: out = 16'(889);
			6483: out = 16'(-3719);
			6484: out = 16'(187);
			6485: out = 16'(-1991);
			6486: out = 16'(3996);
			6487: out = 16'(-1922);
			6488: out = 16'(-2578);
			6489: out = 16'(93);
			6490: out = 16'(-6023);
			6491: out = 16'(4096);
			6492: out = 16'(4047);
			6493: out = 16'(-3223);
			6494: out = 16'(3294);
			6495: out = 16'(-2123);
			6496: out = 16'(5096);
			6497: out = 16'(-7398);
			6498: out = 16'(6274);
			6499: out = 16'(3731);
			6500: out = 16'(-2407);
			6501: out = 16'(-1449);
			6502: out = 16'(1972);
			6503: out = 16'(4439);
			6504: out = 16'(2258);
			6505: out = 16'(1231);
			6506: out = 16'(6618);
			6507: out = 16'(-803);
			6508: out = 16'(-4061);
			6509: out = 16'(-2252);
			6510: out = 16'(2356);
			6511: out = 16'(-226);
			6512: out = 16'(-115);
			6513: out = 16'(-1769);
			6514: out = 16'(-478);
			6515: out = 16'(-1777);
			6516: out = 16'(1384);
			6517: out = 16'(-1763);
			6518: out = 16'(38);
			6519: out = 16'(2029);
			6520: out = 16'(-252);
			6521: out = 16'(-2070);
			6522: out = 16'(909);
			6523: out = 16'(1703);
			6524: out = 16'(2221);
			6525: out = 16'(-1958);
			6526: out = 16'(2791);
			6527: out = 16'(244);
			6528: out = 16'(-747);
			6529: out = 16'(-1534);
			6530: out = 16'(1364);
			6531: out = 16'(4282);
			6532: out = 16'(-2290);
			6533: out = 16'(920);
			6534: out = 16'(3057);
			6535: out = 16'(-764);
			6536: out = 16'(-1455);
			6537: out = 16'(2817);
			6538: out = 16'(2545);
			6539: out = 16'(-60);
			6540: out = 16'(1363);
			6541: out = 16'(-935);
			6542: out = 16'(-502);
			6543: out = 16'(3801);
			6544: out = 16'(-756);
			6545: out = 16'(1033);
			6546: out = 16'(1223);
			6547: out = 16'(-736);
			6548: out = 16'(2560);
			6549: out = 16'(-1976);
			6550: out = 16'(-983);
			6551: out = 16'(4538);
			6552: out = 16'(1433);
			6553: out = 16'(-6799);
			6554: out = 16'(950);
			6555: out = 16'(3354);
			6556: out = 16'(-223);
			6557: out = 16'(437);
			6558: out = 16'(5742);
			6559: out = 16'(-3514);
			6560: out = 16'(-1248);
			6561: out = 16'(1357);
			6562: out = 16'(-222);
			6563: out = 16'(1252);
			6564: out = 16'(1379);
			6565: out = 16'(2816);
			6566: out = 16'(-4101);
			6567: out = 16'(3763);
			6568: out = 16'(-771);
			6569: out = 16'(-4211);
			6570: out = 16'(3922);
			6571: out = 16'(-4218);
			6572: out = 16'(1735);
			6573: out = 16'(2183);
			6574: out = 16'(-5173);
			6575: out = 16'(-2957);
			6576: out = 16'(2191);
			6577: out = 16'(-6456);
			6578: out = 16'(-4423);
			6579: out = 16'(-3125);
			6580: out = 16'(1537);
			6581: out = 16'(-1143);
			6582: out = 16'(3197);
			6583: out = 16'(3250);
			6584: out = 16'(254);
			6585: out = 16'(83);
			6586: out = 16'(-2821);
			6587: out = 16'(-296);
			6588: out = 16'(-435);
			6589: out = 16'(3179);
			6590: out = 16'(1558);
			6591: out = 16'(1546);
			6592: out = 16'(-1596);
			6593: out = 16'(-668);
			6594: out = 16'(-293);
			6595: out = 16'(203);
			6596: out = 16'(1688);
			6597: out = 16'(-818);
			6598: out = 16'(-2343);
			6599: out = 16'(458);
			6600: out = 16'(7605);
			6601: out = 16'(-5006);
			6602: out = 16'(-787);
			6603: out = 16'(2090);
			6604: out = 16'(-4778);
			6605: out = 16'(-4269);
			6606: out = 16'(-4572);
			6607: out = 16'(-503);
			6608: out = 16'(1131);
			6609: out = 16'(-3152);
			6610: out = 16'(1089);
			6611: out = 16'(-662);
			6612: out = 16'(2048);
			6613: out = 16'(-2225);
			6614: out = 16'(-1145);
			6615: out = 16'(4274);
			6616: out = 16'(-3283);
			6617: out = 16'(343);
			6618: out = 16'(3465);
			6619: out = 16'(-3299);
			6620: out = 16'(3519);
			6621: out = 16'(195);
			6622: out = 16'(96);
			6623: out = 16'(-3669);
			6624: out = 16'(4352);
			6625: out = 16'(4030);
			6626: out = 16'(2782);
			6627: out = 16'(243);
			6628: out = 16'(1026);
			6629: out = 16'(-673);
			6630: out = 16'(-2249);
			6631: out = 16'(-1326);
			6632: out = 16'(5494);
			6633: out = 16'(-1709);
			6634: out = 16'(2747);
			6635: out = 16'(-770);
			6636: out = 16'(-1261);
			6637: out = 16'(-4862);
			6638: out = 16'(-1778);
			6639: out = 16'(3372);
			6640: out = 16'(1839);
			6641: out = 16'(-1650);
			6642: out = 16'(5512);
			6643: out = 16'(-7383);
			6644: out = 16'(717);
			6645: out = 16'(-2198);
			6646: out = 16'(206);
			6647: out = 16'(1803);
			6648: out = 16'(330);
			6649: out = 16'(1732);
			6650: out = 16'(-383);
			6651: out = 16'(-242);
			6652: out = 16'(3237);
			6653: out = 16'(0);
			6654: out = 16'(3679);
			6655: out = 16'(-3079);
			6656: out = 16'(177);
			6657: out = 16'(-4);
			6658: out = 16'(-2306);
			6659: out = 16'(2714);
			6660: out = 16'(1847);
			6661: out = 16'(-3110);
			6662: out = 16'(-843);
			6663: out = 16'(-1241);
			6664: out = 16'(919);
			6665: out = 16'(-652);
			6666: out = 16'(2827);
			6667: out = 16'(-4469);
			6668: out = 16'(-920);
			6669: out = 16'(-3035);
			6670: out = 16'(1734);
			6671: out = 16'(-2901);
			6672: out = 16'(-1105);
			6673: out = 16'(1371);
			6674: out = 16'(3067);
			6675: out = 16'(-4660);
			6676: out = 16'(266);
			6677: out = 16'(1995);
			6678: out = 16'(-428);
			6679: out = 16'(1680);
			6680: out = 16'(-3181);
			6681: out = 16'(1239);
			6682: out = 16'(-1180);
			6683: out = 16'(-787);
			6684: out = 16'(8590);
			6685: out = 16'(-49);
			6686: out = 16'(1187);
			6687: out = 16'(2923);
			6688: out = 16'(-1780);
			6689: out = 16'(-57);
			6690: out = 16'(-5339);
			6691: out = 16'(314);
			6692: out = 16'(512);
			6693: out = 16'(-2001);
			6694: out = 16'(3438);
			6695: out = 16'(-147);
			6696: out = 16'(559);
			6697: out = 16'(385);
			6698: out = 16'(257);
			6699: out = 16'(-2406);
			6700: out = 16'(-1903);
			6701: out = 16'(2840);
			6702: out = 16'(-62);
			6703: out = 16'(-4143);
			6704: out = 16'(3889);
			6705: out = 16'(-912);
			6706: out = 16'(714);
			6707: out = 16'(-5309);
			6708: out = 16'(1427);
			6709: out = 16'(3086);
			6710: out = 16'(-2045);
			6711: out = 16'(1576);
			6712: out = 16'(4482);
			6713: out = 16'(-2821);
			6714: out = 16'(-1969);
			6715: out = 16'(-2602);
			6716: out = 16'(3836);
			6717: out = 16'(-305);
			6718: out = 16'(1258);
			6719: out = 16'(-1154);
			6720: out = 16'(-3151);
			6721: out = 16'(-2127);
			6722: out = 16'(528);
			6723: out = 16'(1004);
			6724: out = 16'(-1505);
			6725: out = 16'(-3532);
			6726: out = 16'(5185);
			6727: out = 16'(-3865);
			6728: out = 16'(287);
			6729: out = 16'(-94);
			6730: out = 16'(-6337);
			6731: out = 16'(-594);
			6732: out = 16'(-5261);
			6733: out = 16'(161);
			6734: out = 16'(-1123);
			6735: out = 16'(1923);
			6736: out = 16'(3623);
			6737: out = 16'(86);
			6738: out = 16'(1082);
			6739: out = 16'(-1166);
			6740: out = 16'(-3064);
			6741: out = 16'(-376);
			6742: out = 16'(-389);
			6743: out = 16'(3968);
			6744: out = 16'(954);
			6745: out = 16'(488);
			6746: out = 16'(-1637);
			6747: out = 16'(382);
			6748: out = 16'(2);
			6749: out = 16'(-3069);
			6750: out = 16'(5001);
			6751: out = 16'(-1310);
			6752: out = 16'(-3151);
			6753: out = 16'(-1055);
			6754: out = 16'(1349);
			6755: out = 16'(-754);
			6756: out = 16'(-3552);
			6757: out = 16'(-2061);
			6758: out = 16'(-4332);
			6759: out = 16'(1187);
			6760: out = 16'(-603);
			6761: out = 16'(696);
			6762: out = 16'(4341);
			6763: out = 16'(-1089);
			6764: out = 16'(-4530);
			6765: out = 16'(278);
			6766: out = 16'(-1440);
			6767: out = 16'(-1647);
			6768: out = 16'(5155);
			6769: out = 16'(-873);
			6770: out = 16'(-1934);
			6771: out = 16'(1100);
			6772: out = 16'(-3273);
			6773: out = 16'(-2265);
			6774: out = 16'(1279);
			6775: out = 16'(4081);
			6776: out = 16'(-557);
			6777: out = 16'(-2036);
			6778: out = 16'(988);
			6779: out = 16'(-2157);
			6780: out = 16'(770);
			6781: out = 16'(1217);
			6782: out = 16'(3172);
			6783: out = 16'(-1156);
			6784: out = 16'(12);
			6785: out = 16'(-3923);
			6786: out = 16'(4045);
			6787: out = 16'(-184);
			6788: out = 16'(3362);
			6789: out = 16'(-3640);
			6790: out = 16'(-732);
			6791: out = 16'(-588);
			6792: out = 16'(-977);
			6793: out = 16'(1064);
			6794: out = 16'(626);
			6795: out = 16'(2239);
			6796: out = 16'(-1447);
			6797: out = 16'(-1510);
			6798: out = 16'(-3028);
			6799: out = 16'(-1286);
			6800: out = 16'(4009);
			6801: out = 16'(-1380);
			6802: out = 16'(-190);
			6803: out = 16'(-141);
			6804: out = 16'(-189);
			6805: out = 16'(647);
			6806: out = 16'(-260);
			6807: out = 16'(4356);
			6808: out = 16'(-2087);
			6809: out = 16'(-282);
			6810: out = 16'(3302);
			6811: out = 16'(56);
			6812: out = 16'(-39);
			6813: out = 16'(330);
			6814: out = 16'(2483);
			6815: out = 16'(-2333);
			6816: out = 16'(-2647);
			6817: out = 16'(2214);
			6818: out = 16'(-2802);
			6819: out = 16'(-274);
			6820: out = 16'(3654);
			6821: out = 16'(-2337);
			6822: out = 16'(-250);
			6823: out = 16'(111);
			6824: out = 16'(183);
			6825: out = 16'(1413);
			6826: out = 16'(64);
			6827: out = 16'(693);
			6828: out = 16'(-214);
			6829: out = 16'(-495);
			6830: out = 16'(-220);
			6831: out = 16'(14);
			6832: out = 16'(869);
			6833: out = 16'(-5127);
			6834: out = 16'(2913);
			6835: out = 16'(-3516);
			6836: out = 16'(153);
			6837: out = 16'(-1381);
			6838: out = 16'(3311);
			6839: out = 16'(1178);
			6840: out = 16'(-1855);
			6841: out = 16'(-789);
			6842: out = 16'(-4275);
			6843: out = 16'(-885);
			6844: out = 16'(-419);
			6845: out = 16'(3459);
			6846: out = 16'(-3357);
			6847: out = 16'(1285);
			6848: out = 16'(-1673);
			6849: out = 16'(-4062);
			6850: out = 16'(-2427);
			6851: out = 16'(-2219);
			6852: out = 16'(6922);
			6853: out = 16'(-1987);
			6854: out = 16'(-287);
			6855: out = 16'(-9);
			6856: out = 16'(-768);
			6857: out = 16'(-836);
			6858: out = 16'(290);
			6859: out = 16'(2589);
			6860: out = 16'(-4604);
			6861: out = 16'(-250);
			6862: out = 16'(912);
			6863: out = 16'(-3025);
			6864: out = 16'(2227);
			6865: out = 16'(-3389);
			6866: out = 16'(2428);
			6867: out = 16'(-3222);
			6868: out = 16'(372);
			6869: out = 16'(2903);
			6870: out = 16'(-1357);
			6871: out = 16'(1763);
			6872: out = 16'(-354);
			6873: out = 16'(-758);
			6874: out = 16'(393);
			6875: out = 16'(-2185);
			6876: out = 16'(1901);
			6877: out = 16'(-568);
			6878: out = 16'(-238);
			6879: out = 16'(77);
			6880: out = 16'(50);
			6881: out = 16'(-2193);
			6882: out = 16'(1349);
			6883: out = 16'(466);
			6884: out = 16'(1804);
			6885: out = 16'(637);
			6886: out = 16'(-1385);
			6887: out = 16'(219);
			6888: out = 16'(1201);
			6889: out = 16'(1993);
			6890: out = 16'(111);
			6891: out = 16'(1224);
			6892: out = 16'(-2715);
			6893: out = 16'(3);
			6894: out = 16'(523);
			6895: out = 16'(921);
			6896: out = 16'(998);
			6897: out = 16'(2481);
			6898: out = 16'(-550);
			6899: out = 16'(-3408);
			6900: out = 16'(2301);
			6901: out = 16'(-2299);
			6902: out = 16'(1336);
			6903: out = 16'(60);
			6904: out = 16'(3193);
			6905: out = 16'(-1155);
			6906: out = 16'(-1283);
			6907: out = 16'(-1467);
			6908: out = 16'(-3572);
			6909: out = 16'(2743);
			6910: out = 16'(364);
			6911: out = 16'(1894);
			6912: out = 16'(-2268);
			6913: out = 16'(-176);
			6914: out = 16'(88);
			6915: out = 16'(-2825);
			6916: out = 16'(-263);
			6917: out = 16'(-1427);
			6918: out = 16'(-1777);
			6919: out = 16'(-1812);
			6920: out = 16'(2193);
			6921: out = 16'(1101);
			6922: out = 16'(3668);
			6923: out = 16'(445);
			6924: out = 16'(-1092);
			6925: out = 16'(-5159);
			6926: out = 16'(1696);
			6927: out = 16'(-2106);
			6928: out = 16'(5298);
			6929: out = 16'(4276);
			6930: out = 16'(-190);
			6931: out = 16'(539);
			6932: out = 16'(-1204);
			6933: out = 16'(1961);
			6934: out = 16'(-1331);
			6935: out = 16'(17);
			6936: out = 16'(5535);
			6937: out = 16'(-1236);
			6938: out = 16'(240);
			6939: out = 16'(-73);
			6940: out = 16'(1901);
			6941: out = 16'(-111);
			6942: out = 16'(-2377);
			6943: out = 16'(1331);
			6944: out = 16'(-4174);
			6945: out = 16'(3121);
			6946: out = 16'(-5897);
			6947: out = 16'(2999);
			6948: out = 16'(1791);
			6949: out = 16'(271);
			6950: out = 16'(1622);
			6951: out = 16'(-343);
			6952: out = 16'(127);
			6953: out = 16'(-889);
			6954: out = 16'(-1431);
			6955: out = 16'(911);
			6956: out = 16'(-1120);
			6957: out = 16'(5130);
			6958: out = 16'(-7598);
			6959: out = 16'(1910);
			6960: out = 16'(-1097);
			6961: out = 16'(1470);
			6962: out = 16'(-1813);
			6963: out = 16'(-685);
			6964: out = 16'(-36);
			6965: out = 16'(416);
			6966: out = 16'(1916);
			6967: out = 16'(2680);
			6968: out = 16'(-145);
			6969: out = 16'(-206);
			6970: out = 16'(-2904);
			6971: out = 16'(-525);
			6972: out = 16'(-1441);
			6973: out = 16'(1057);
			6974: out = 16'(3088);
			6975: out = 16'(-2106);
			6976: out = 16'(-3109);
			6977: out = 16'(-3850);
			6978: out = 16'(-1480);
			6979: out = 16'(-2637);
			6980: out = 16'(470);
			6981: out = 16'(4260);
			6982: out = 16'(-642);
			6983: out = 16'(-121);
			6984: out = 16'(-850);
			6985: out = 16'(-1603);
			6986: out = 16'(462);
			6987: out = 16'(-5934);
			6988: out = 16'(2794);
			6989: out = 16'(2631);
			6990: out = 16'(1384);
			6991: out = 16'(1478);
			6992: out = 16'(1153);
			6993: out = 16'(-297);
			6994: out = 16'(-1976);
			6995: out = 16'(-2087);
			6996: out = 16'(-2403);
			6997: out = 16'(2976);
			6998: out = 16'(3924);
			6999: out = 16'(2014);
			7000: out = 16'(-683);
			7001: out = 16'(-3762);
			7002: out = 16'(191);
			7003: out = 16'(-4090);
			7004: out = 16'(-1436);
			7005: out = 16'(3315);
			7006: out = 16'(-542);
			7007: out = 16'(901);
			7008: out = 16'(-3041);
			7009: out = 16'(-2174);
			7010: out = 16'(-6111);
			7011: out = 16'(-1166);
			7012: out = 16'(-361);
			7013: out = 16'(1264);
			7014: out = 16'(2167);
			7015: out = 16'(88);
			7016: out = 16'(-1581);
			7017: out = 16'(-783);
			7018: out = 16'(12);
			7019: out = 16'(-53);
			7020: out = 16'(-2652);
			7021: out = 16'(2511);
			7022: out = 16'(-3043);
			7023: out = 16'(1851);
			7024: out = 16'(600);
			7025: out = 16'(-609);
			7026: out = 16'(5230);
			7027: out = 16'(-2798);
			7028: out = 16'(-3697);
			7029: out = 16'(9);
			7030: out = 16'(-1562);
			7031: out = 16'(1843);
			7032: out = 16'(-156);
			7033: out = 16'(-646);
			7034: out = 16'(-381);
			7035: out = 16'(-1017);
			7036: out = 16'(210);
			7037: out = 16'(157);
			7038: out = 16'(26);
			7039: out = 16'(-2297);
			7040: out = 16'(227);
			7041: out = 16'(-2048);
			7042: out = 16'(1166);
			7043: out = 16'(-1213);
			7044: out = 16'(513);
			7045: out = 16'(-99);
			7046: out = 16'(361);
			7047: out = 16'(-680);
			7048: out = 16'(1201);
			7049: out = 16'(171);
			7050: out = 16'(3292);
			7051: out = 16'(1833);
			7052: out = 16'(-2965);
			7053: out = 16'(-571);
			7054: out = 16'(-1266);
			7055: out = 16'(-4398);
			7056: out = 16'(446);
			7057: out = 16'(1334);
			7058: out = 16'(-129);
			7059: out = 16'(4430);
			7060: out = 16'(342);
			7061: out = 16'(-1761);
			7062: out = 16'(-281);
			7063: out = 16'(-845);
			7064: out = 16'(-687);
			7065: out = 16'(-62);
			7066: out = 16'(1652);
			7067: out = 16'(1136);
			7068: out = 16'(-1314);
			7069: out = 16'(2373);
			7070: out = 16'(-2553);
			7071: out = 16'(51);
			7072: out = 16'(-1427);
			7073: out = 16'(2045);
			7074: out = 16'(1925);
			7075: out = 16'(-202);
			7076: out = 16'(1462);
			7077: out = 16'(-189);
			7078: out = 16'(813);
			7079: out = 16'(-1471);
			7080: out = 16'(-1487);
			7081: out = 16'(-2017);
			7082: out = 16'(-2524);
			7083: out = 16'(5367);
			7084: out = 16'(-933);
			7085: out = 16'(2311);
			7086: out = 16'(-785);
			7087: out = 16'(-1651);
			7088: out = 16'(950);
			7089: out = 16'(-2230);
			7090: out = 16'(3152);
			7091: out = 16'(-1271);
			7092: out = 16'(4146);
			7093: out = 16'(-2851);
			7094: out = 16'(-3445);
			7095: out = 16'(2917);
			7096: out = 16'(-2711);
			7097: out = 16'(-2024);
			7098: out = 16'(-315);
			7099: out = 16'(-267);
			7100: out = 16'(3775);
			7101: out = 16'(1085);
			7102: out = 16'(1860);
			7103: out = 16'(-1269);
			7104: out = 16'(1003);
			7105: out = 16'(-1478);
			7106: out = 16'(-2132);
			7107: out = 16'(1248);
			7108: out = 16'(1728);
			7109: out = 16'(-1049);
			7110: out = 16'(-511);
			7111: out = 16'(325);
			7112: out = 16'(-93);
			7113: out = 16'(-3630);
			7114: out = 16'(1102);
			7115: out = 16'(-2740);
			7116: out = 16'(76);
			7117: out = 16'(119);
			7118: out = 16'(937);
			7119: out = 16'(-1422);
			7120: out = 16'(61);
			7121: out = 16'(582);
			7122: out = 16'(-2444);
			7123: out = 16'(3584);
			7124: out = 16'(-134);
			7125: out = 16'(4066);
			7126: out = 16'(331);
			7127: out = 16'(3955);
			7128: out = 16'(1236);
			7129: out = 16'(-1312);
			7130: out = 16'(-2616);
			7131: out = 16'(270);
			7132: out = 16'(-878);
			7133: out = 16'(-1602);
			7134: out = 16'(-380);
			7135: out = 16'(4044);
			7136: out = 16'(311);
			7137: out = 16'(2534);
			7138: out = 16'(-2487);
			7139: out = 16'(-2862);
			7140: out = 16'(1629);
			7141: out = 16'(-237);
			7142: out = 16'(2478);
			7143: out = 16'(18);
			7144: out = 16'(-1878);
			7145: out = 16'(-791);
			7146: out = 16'(-7083);
			7147: out = 16'(1858);
			7148: out = 16'(-2886);
			7149: out = 16'(1662);
			7150: out = 16'(461);
			7151: out = 16'(422);
			7152: out = 16'(1649);
			7153: out = 16'(890);
			7154: out = 16'(1873);
			7155: out = 16'(-979);
			7156: out = 16'(-2396);
			7157: out = 16'(271);
			7158: out = 16'(-3640);
			7159: out = 16'(4857);
			7160: out = 16'(683);
			7161: out = 16'(-575);
			7162: out = 16'(122);
			7163: out = 16'(-649);
			7164: out = 16'(-5261);
			7165: out = 16'(-464);
			7166: out = 16'(1036);
			7167: out = 16'(1116);
			7168: out = 16'(968);
			7169: out = 16'(4704);
			7170: out = 16'(-5156);
			7171: out = 16'(4163);
			7172: out = 16'(-4422);
			7173: out = 16'(679);
			7174: out = 16'(-2095);
			7175: out = 16'(-559);
			7176: out = 16'(1843);
			7177: out = 16'(-74);
			7178: out = 16'(2517);
			7179: out = 16'(2112);
			7180: out = 16'(-3953);
			7181: out = 16'(-138);
			7182: out = 16'(-2035);
			7183: out = 16'(-1148);
			7184: out = 16'(1723);
			7185: out = 16'(-317);
			7186: out = 16'(3271);
			7187: out = 16'(628);
			7188: out = 16'(589);
			7189: out = 16'(2092);
			7190: out = 16'(707);
			7191: out = 16'(-1786);
			7192: out = 16'(3414);
			7193: out = 16'(-1335);
			7194: out = 16'(1999);
			7195: out = 16'(933);
			7196: out = 16'(-3546);
			7197: out = 16'(-1097);
			7198: out = 16'(-832);
			7199: out = 16'(2160);
			7200: out = 16'(82);
			7201: out = 16'(3334);
			7202: out = 16'(-86);
			7203: out = 16'(-1545);
			7204: out = 16'(1694);
			7205: out = 16'(-1338);
			7206: out = 16'(-62);
			7207: out = 16'(-2071);
			7208: out = 16'(-2038);
			7209: out = 16'(728);
			7210: out = 16'(1610);
			7211: out = 16'(1601);
			7212: out = 16'(-2025);
			7213: out = 16'(1546);
			7214: out = 16'(-289);
			7215: out = 16'(-3463);
			7216: out = 16'(-1554);
			7217: out = 16'(2226);
			7218: out = 16'(3064);
			7219: out = 16'(1065);
			7220: out = 16'(-6735);
			7221: out = 16'(1799);
			7222: out = 16'(-1477);
			7223: out = 16'(-49);
			7224: out = 16'(2094);
			7225: out = 16'(-2890);
			7226: out = 16'(2754);
			7227: out = 16'(-2827);
			7228: out = 16'(2114);
			7229: out = 16'(-1031);
			7230: out = 16'(-785);
			7231: out = 16'(-224);
			7232: out = 16'(-3543);
			7233: out = 16'(1955);
			7234: out = 16'(2125);
			7235: out = 16'(-997);
			7236: out = 16'(1804);
			7237: out = 16'(1014);
			7238: out = 16'(4469);
			7239: out = 16'(-4716);
			7240: out = 16'(1568);
			7241: out = 16'(-872);
			7242: out = 16'(-363);
			7243: out = 16'(589);
			7244: out = 16'(-3057);
			7245: out = 16'(2461);
			7246: out = 16'(-178);
			7247: out = 16'(2101);
			7248: out = 16'(-838);
			7249: out = 16'(2010);
			7250: out = 16'(176);
			7251: out = 16'(1444);
			7252: out = 16'(854);
			7253: out = 16'(-1467);
			7254: out = 16'(2656);
			7255: out = 16'(-240);
			7256: out = 16'(-255);
			7257: out = 16'(171);
			7258: out = 16'(-1269);
			7259: out = 16'(-1017);
			7260: out = 16'(-1961);
			7261: out = 16'(1413);
			7262: out = 16'(1648);
			7263: out = 16'(2471);
			7264: out = 16'(-1987);
			7265: out = 16'(303);
			7266: out = 16'(-1177);
			7267: out = 16'(-1361);
			7268: out = 16'(-2862);
			7269: out = 16'(3114);
			7270: out = 16'(4064);
			7271: out = 16'(1016);
			7272: out = 16'(-793);
			7273: out = 16'(1766);
			7274: out = 16'(-154);
			7275: out = 16'(564);
			7276: out = 16'(2300);
			7277: out = 16'(-344);
			7278: out = 16'(4494);
			7279: out = 16'(-484);
			7280: out = 16'(1547);
			7281: out = 16'(2236);
			7282: out = 16'(-2915);
			7283: out = 16'(606);
			7284: out = 16'(-5564);
			7285: out = 16'(1330);
			7286: out = 16'(-656);
			7287: out = 16'(457);
			7288: out = 16'(2427);
			7289: out = 16'(-1160);
			7290: out = 16'(-348);
			7291: out = 16'(-3791);
			7292: out = 16'(-2214);
			7293: out = 16'(100);
			7294: out = 16'(-878);
			7295: out = 16'(312);
			7296: out = 16'(485);
			7297: out = 16'(3617);
			7298: out = 16'(-1413);
			7299: out = 16'(-1283);
			7300: out = 16'(2141);
			7301: out = 16'(-2025);
			7302: out = 16'(2852);
			7303: out = 16'(-2422);
			7304: out = 16'(2663);
			7305: out = 16'(-1033);
			7306: out = 16'(584);
			7307: out = 16'(227);
			7308: out = 16'(-1277);
			7309: out = 16'(3284);
			7310: out = 16'(-382);
			7311: out = 16'(77);
			7312: out = 16'(1871);
			7313: out = 16'(870);
			7314: out = 16'(272);
			7315: out = 16'(1341);
			7316: out = 16'(-2587);
			7317: out = 16'(-683);
			7318: out = 16'(-2344);
			7319: out = 16'(1888);
			7320: out = 16'(-1731);
			7321: out = 16'(955);
			7322: out = 16'(1741);
			7323: out = 16'(-730);
			7324: out = 16'(-610);
			7325: out = 16'(16);
			7326: out = 16'(-338);
			7327: out = 16'(-2423);
			7328: out = 16'(3344);
			7329: out = 16'(-25);
			7330: out = 16'(240);
			7331: out = 16'(5391);
			7332: out = 16'(2486);
			7333: out = 16'(1669);
			7334: out = 16'(-1844);
			7335: out = 16'(1675);
			7336: out = 16'(-2990);
			7337: out = 16'(-1923);
			7338: out = 16'(-738);
			7339: out = 16'(997);
			7340: out = 16'(2152);
			7341: out = 16'(1026);
			7342: out = 16'(1006);
			7343: out = 16'(-1882);
			7344: out = 16'(157);
			7345: out = 16'(86);
			7346: out = 16'(107);
			7347: out = 16'(3249);
			7348: out = 16'(-94);
			7349: out = 16'(1130);
			7350: out = 16'(-903);
			7351: out = 16'(-2588);
			7352: out = 16'(289);
			7353: out = 16'(-1984);
			7354: out = 16'(1631);
			7355: out = 16'(1100);
			7356: out = 16'(767);
			7357: out = 16'(1084);
			7358: out = 16'(-1052);
			7359: out = 16'(997);
			7360: out = 16'(-3197);
			7361: out = 16'(537);
			7362: out = 16'(-418);
			7363: out = 16'(1293);
			7364: out = 16'(1452);
			7365: out = 16'(-2944);
			7366: out = 16'(492);
			7367: out = 16'(563);
			7368: out = 16'(-3754);
			7369: out = 16'(-647);
			7370: out = 16'(-3150);
			7371: out = 16'(1182);
			7372: out = 16'(969);
			7373: out = 16'(1976);
			7374: out = 16'(953);
			7375: out = 16'(-3922);
			7376: out = 16'(-87);
			7377: out = 16'(-1625);
			7378: out = 16'(274);
			7379: out = 16'(1735);
			7380: out = 16'(-2543);
			7381: out = 16'(2621);
			7382: out = 16'(-2252);
			7383: out = 16'(4759);
			7384: out = 16'(-466);
			7385: out = 16'(812);
			7386: out = 16'(-1949);
			7387: out = 16'(884);
			7388: out = 16'(-1637);
			7389: out = 16'(-941);
			7390: out = 16'(2235);
			7391: out = 16'(775);
			7392: out = 16'(1122);
			7393: out = 16'(160);
			7394: out = 16'(-4291);
			7395: out = 16'(522);
			7396: out = 16'(-1751);
			7397: out = 16'(2126);
			7398: out = 16'(1715);
			7399: out = 16'(923);
			7400: out = 16'(1590);
			7401: out = 16'(-2920);
			7402: out = 16'(2431);
			7403: out = 16'(-268);
			7404: out = 16'(-1989);
			7405: out = 16'(-892);
			7406: out = 16'(1396);
			7407: out = 16'(-640);
			7408: out = 16'(-107);
			7409: out = 16'(1774);
			7410: out = 16'(-17);
			7411: out = 16'(-961);
			7412: out = 16'(-52);
			7413: out = 16'(-6040);
			7414: out = 16'(3492);
			7415: out = 16'(-1872);
			7416: out = 16'(1707);
			7417: out = 16'(-2424);
			7418: out = 16'(336);
			7419: out = 16'(-714);
			7420: out = 16'(-3074);
			7421: out = 16'(1185);
			7422: out = 16'(51);
			7423: out = 16'(-519);
			7424: out = 16'(1189);
			7425: out = 16'(2733);
			7426: out = 16'(2453);
			7427: out = 16'(-6173);
			7428: out = 16'(-1292);
			7429: out = 16'(848);
			7430: out = 16'(-420);
			7431: out = 16'(2707);
			7432: out = 16'(194);
			7433: out = 16'(2549);
			7434: out = 16'(-1374);
			7435: out = 16'(1723);
			7436: out = 16'(-2949);
			7437: out = 16'(-1022);
			7438: out = 16'(-530);
			7439: out = 16'(-3236);
			7440: out = 16'(2282);
			7441: out = 16'(274);
			7442: out = 16'(3775);
			7443: out = 16'(531);
			7444: out = 16'(179);
			7445: out = 16'(2579);
			7446: out = 16'(-7197);
			7447: out = 16'(2274);
			7448: out = 16'(-365);
			7449: out = 16'(415);
			7450: out = 16'(2511);
			7451: out = 16'(-646);
			7452: out = 16'(-667);
			7453: out = 16'(1740);
			7454: out = 16'(162);
			7455: out = 16'(-3951);
			7456: out = 16'(-629);
			7457: out = 16'(800);
			7458: out = 16'(-208);
			7459: out = 16'(-1014);
			7460: out = 16'(-734);
			7461: out = 16'(2306);
			7462: out = 16'(-901);
			7463: out = 16'(-6);
			7464: out = 16'(-323);
			7465: out = 16'(4030);
			7466: out = 16'(3073);
			7467: out = 16'(2328);
			7468: out = 16'(1064);
			7469: out = 16'(-1443);
			7470: out = 16'(-1132);
			7471: out = 16'(-3506);
			7472: out = 16'(-1239);
			7473: out = 16'(122);
			7474: out = 16'(2254);
			7475: out = 16'(-1856);
			7476: out = 16'(558);
			7477: out = 16'(2001);
			7478: out = 16'(148);
			7479: out = 16'(-924);
			7480: out = 16'(-1980);
			7481: out = 16'(2751);
			7482: out = 16'(290);
			7483: out = 16'(2837);
			7484: out = 16'(88);
			7485: out = 16'(-29);
			7486: out = 16'(1998);
			7487: out = 16'(-5585);
			7488: out = 16'(1782);
			7489: out = 16'(-425);
			7490: out = 16'(1429);
			7491: out = 16'(157);
			7492: out = 16'(2873);
			7493: out = 16'(1446);
			7494: out = 16'(-141);
			7495: out = 16'(3394);
			7496: out = 16'(-2789);
			7497: out = 16'(927);
			7498: out = 16'(-1554);
			7499: out = 16'(-660);
			7500: out = 16'(1010);
			7501: out = 16'(617);
			7502: out = 16'(489);
			7503: out = 16'(-590);
			7504: out = 16'(-1044);
			7505: out = 16'(-2010);
			7506: out = 16'(-555);
			7507: out = 16'(2292);
			7508: out = 16'(937);
			7509: out = 16'(315);
			7510: out = 16'(1472);
			7511: out = 16'(-1740);
			7512: out = 16'(551);
			7513: out = 16'(-540);
			7514: out = 16'(2284);
			7515: out = 16'(-2380);
			7516: out = 16'(2348);
			7517: out = 16'(-1308);
			7518: out = 16'(-46);
			7519: out = 16'(611);
			7520: out = 16'(101);
			7521: out = 16'(-683);
			7522: out = 16'(-255);
			7523: out = 16'(-1590);
			7524: out = 16'(-67);
			7525: out = 16'(-2207);
			7526: out = 16'(4126);
			7527: out = 16'(-958);
			7528: out = 16'(316);
			7529: out = 16'(354);
			7530: out = 16'(-3557);
			7531: out = 16'(1215);
			7532: out = 16'(-625);
			7533: out = 16'(1496);
			7534: out = 16'(1343);
			7535: out = 16'(-3336);
			7536: out = 16'(151);
			7537: out = 16'(-1351);
			7538: out = 16'(-2567);
			7539: out = 16'(-1057);
			7540: out = 16'(212);
			7541: out = 16'(271);
			7542: out = 16'(-741);
			7543: out = 16'(870);
			7544: out = 16'(-136);
			7545: out = 16'(3407);
			7546: out = 16'(-2068);
			7547: out = 16'(2321);
			7548: out = 16'(-676);
			7549: out = 16'(-103);
			7550: out = 16'(-1260);
			7551: out = 16'(2236);
			7552: out = 16'(1315);
			7553: out = 16'(-50);
			7554: out = 16'(465);
			7555: out = 16'(-1017);
			7556: out = 16'(-1187);
			7557: out = 16'(-2632);
			7558: out = 16'(990);
			7559: out = 16'(-471);
			7560: out = 16'(752);
			7561: out = 16'(991);
			7562: out = 16'(-4503);
			7563: out = 16'(273);
			7564: out = 16'(-803);
			7565: out = 16'(1583);
			7566: out = 16'(3470);
			7567: out = 16'(553);
			7568: out = 16'(-1021);
			7569: out = 16'(-64);
			7570: out = 16'(-2666);
			7571: out = 16'(384);
			7572: out = 16'(-1108);
			7573: out = 16'(-788);
			7574: out = 16'(-2379);
			7575: out = 16'(-377);
			7576: out = 16'(1356);
			7577: out = 16'(109);
			7578: out = 16'(135);
			7579: out = 16'(3860);
			7580: out = 16'(-1735);
			7581: out = 16'(-2330);
			7582: out = 16'(-886);
			7583: out = 16'(284);
			7584: out = 16'(-617);
			7585: out = 16'(1487);
			7586: out = 16'(390);
			7587: out = 16'(731);
			7588: out = 16'(2406);
			7589: out = 16'(-2117);
			7590: out = 16'(1141);
			7591: out = 16'(-1762);
			7592: out = 16'(819);
			7593: out = 16'(-1778);
			7594: out = 16'(-1998);
			7595: out = 16'(1872);
			7596: out = 16'(351);
			7597: out = 16'(1368);
			7598: out = 16'(-2330);
			7599: out = 16'(-3470);
			7600: out = 16'(80);
			7601: out = 16'(-3506);
			7602: out = 16'(723);
			7603: out = 16'(4347);
			7604: out = 16'(-726);
			7605: out = 16'(-2553);
			7606: out = 16'(3509);
			7607: out = 16'(-2866);
			7608: out = 16'(1562);
			7609: out = 16'(-1829);
			7610: out = 16'(668);
			7611: out = 16'(1317);
			7612: out = 16'(-974);
			7613: out = 16'(177);
			7614: out = 16'(-602);
			7615: out = 16'(1041);
			7616: out = 16'(2173);
			7617: out = 16'(1768);
			7618: out = 16'(-13);
			7619: out = 16'(-350);
			7620: out = 16'(787);
			7621: out = 16'(-2588);
			7622: out = 16'(63);
			7623: out = 16'(-2337);
			7624: out = 16'(940);
			7625: out = 16'(-2470);
			7626: out = 16'(619);
			7627: out = 16'(662);
			7628: out = 16'(-66);
			7629: out = 16'(-790);
			7630: out = 16'(1269);
			7631: out = 16'(979);
			7632: out = 16'(-774);
			7633: out = 16'(-2434);
			7634: out = 16'(-2205);
			7635: out = 16'(479);
			7636: out = 16'(-401);
			7637: out = 16'(1582);
			7638: out = 16'(825);
			7639: out = 16'(-430);
			7640: out = 16'(1253);
			7641: out = 16'(284);
			7642: out = 16'(351);
			7643: out = 16'(2336);
			7644: out = 16'(-5003);
			7645: out = 16'(3369);
			7646: out = 16'(-2135);
			7647: out = 16'(1667);
			7648: out = 16'(1536);
			7649: out = 16'(1232);
			7650: out = 16'(-88);
			7651: out = 16'(-1664);
			7652: out = 16'(1704);
			7653: out = 16'(-3001);
			7654: out = 16'(2667);
			7655: out = 16'(2081);
			7656: out = 16'(-1362);
			7657: out = 16'(-15);
			7658: out = 16'(517);
			7659: out = 16'(-3299);
			7660: out = 16'(328);
			7661: out = 16'(-286);
			7662: out = 16'(-703);
			7663: out = 16'(-542);
			7664: out = 16'(1108);
			7665: out = 16'(1117);
			7666: out = 16'(-976);
			7667: out = 16'(-2369);
			7668: out = 16'(1897);
			7669: out = 16'(-185);
			7670: out = 16'(2926);
			7671: out = 16'(-476);
			7672: out = 16'(1008);
			7673: out = 16'(-2260);
			7674: out = 16'(785);
			7675: out = 16'(1757);
			7676: out = 16'(-1319);
			7677: out = 16'(-210);
			7678: out = 16'(-197);
			7679: out = 16'(-2547);
			7680: out = 16'(-225);
			7681: out = 16'(1227);
			7682: out = 16'(215);
			7683: out = 16'(-3210);
			7684: out = 16'(33);
			7685: out = 16'(-2535);
			7686: out = 16'(524);
			7687: out = 16'(-1206);
			7688: out = 16'(474);
			7689: out = 16'(-579);
			7690: out = 16'(-326);
			7691: out = 16'(-45);
			7692: out = 16'(15);
			7693: out = 16'(-1049);
			7694: out = 16'(40);
			7695: out = 16'(-1387);
			7696: out = 16'(778);
			7697: out = 16'(1496);
			7698: out = 16'(-1683);
			7699: out = 16'(3654);
			7700: out = 16'(151);
			7701: out = 16'(175);
			7702: out = 16'(982);
			7703: out = 16'(-4119);
			7704: out = 16'(-1314);
			7705: out = 16'(-1517);
			7706: out = 16'(5301);
			7707: out = 16'(-908);
			7708: out = 16'(2702);
			7709: out = 16'(-128);
			7710: out = 16'(-139);
			7711: out = 16'(-1977);
			7712: out = 16'(-436);
			7713: out = 16'(-353);
			7714: out = 16'(-191);
			7715: out = 16'(1579);
			7716: out = 16'(-1925);
			7717: out = 16'(1948);
			7718: out = 16'(705);
			7719: out = 16'(-145);
			7720: out = 16'(589);
			7721: out = 16'(-3341);
			7722: out = 16'(443);
			7723: out = 16'(-915);
			7724: out = 16'(135);
			7725: out = 16'(-205);
			7726: out = 16'(2504);
			7727: out = 16'(143);
			7728: out = 16'(-551);
			7729: out = 16'(1426);
			7730: out = 16'(-92);
			7731: out = 16'(-44);
			7732: out = 16'(-878);
			7733: out = 16'(2093);
			7734: out = 16'(1229);
			7735: out = 16'(-699);
			7736: out = 16'(-1488);
			7737: out = 16'(-1027);
			7738: out = 16'(1940);
			7739: out = 16'(980);
			7740: out = 16'(-344);
			7741: out = 16'(-2900);
			7742: out = 16'(-1388);
			7743: out = 16'(-4020);
			7744: out = 16'(14);
			7745: out = 16'(-3580);
			7746: out = 16'(-321);
			7747: out = 16'(1975);
			7748: out = 16'(-1794);
			7749: out = 16'(3435);
			7750: out = 16'(-1415);
			7751: out = 16'(3963);
			7752: out = 16'(-666);
			7753: out = 16'(-437);
			7754: out = 16'(3092);
			7755: out = 16'(-4587);
			7756: out = 16'(1542);
			7757: out = 16'(870);
			7758: out = 16'(2069);
			7759: out = 16'(2228);
			7760: out = 16'(-3696);
			7761: out = 16'(1666);
			7762: out = 16'(-1169);
			7763: out = 16'(-1512);
			7764: out = 16'(-2447);
			7765: out = 16'(3930);
			7766: out = 16'(9);
			7767: out = 16'(1178);
			7768: out = 16'(422);
			7769: out = 16'(-2172);
			7770: out = 16'(3345);
			7771: out = 16'(-481);
			7772: out = 16'(2584);
			7773: out = 16'(-1926);
			7774: out = 16'(-1779);
			7775: out = 16'(3102);
			7776: out = 16'(-2695);
			7777: out = 16'(5381);
			7778: out = 16'(-2279);
			7779: out = 16'(-497);
			7780: out = 16'(161);
			7781: out = 16'(-4191);
			7782: out = 16'(-1737);
			7783: out = 16'(1611);
			7784: out = 16'(-1556);
			7785: out = 16'(464);
			7786: out = 16'(1075);
			7787: out = 16'(-2452);
			7788: out = 16'(870);
			7789: out = 16'(304);
			7790: out = 16'(724);
			7791: out = 16'(2858);
			7792: out = 16'(1514);
			7793: out = 16'(1829);
			7794: out = 16'(-1464);
			7795: out = 16'(-241);
			7796: out = 16'(-639);
			7797: out = 16'(-822);
			7798: out = 16'(-251);
			7799: out = 16'(-230);
			7800: out = 16'(-2017);
			7801: out = 16'(-259);
			7802: out = 16'(-2321);
			7803: out = 16'(-116);
			7804: out = 16'(2460);
			7805: out = 16'(-5246);
			7806: out = 16'(152);
			7807: out = 16'(-1259);
			7808: out = 16'(-1416);
			7809: out = 16'(4671);
			7810: out = 16'(-1455);
			7811: out = 16'(3123);
			7812: out = 16'(-2246);
			7813: out = 16'(-2145);
			7814: out = 16'(175);
			7815: out = 16'(259);
			7816: out = 16'(-73);
			7817: out = 16'(585);
			7818: out = 16'(-253);
			7819: out = 16'(1764);
			7820: out = 16'(1025);
			7821: out = 16'(-1282);
			7822: out = 16'(1754);
			7823: out = 16'(-259);
			7824: out = 16'(-3523);
			7825: out = 16'(23);
			7826: out = 16'(-6142);
			7827: out = 16'(-82);
			7828: out = 16'(2869);
			7829: out = 16'(-4078);
			7830: out = 16'(1148);
			7831: out = 16'(-1432);
			7832: out = 16'(-943);
			7833: out = 16'(-44);
			7834: out = 16'(-1552);
			7835: out = 16'(4102);
			7836: out = 16'(-857);
			7837: out = 16'(897);
			7838: out = 16'(1776);
			7839: out = 16'(-5441);
			7840: out = 16'(2856);
			7841: out = 16'(-4190);
			7842: out = 16'(562);
			7843: out = 16'(2052);
			7844: out = 16'(-560);
			7845: out = 16'(-432);
			7846: out = 16'(-1337);
			7847: out = 16'(-875);
			7848: out = 16'(-755);
			7849: out = 16'(2329);
			7850: out = 16'(-57);
			7851: out = 16'(1754);
			7852: out = 16'(701);
			7853: out = 16'(-257);
			7854: out = 16'(179);
			7855: out = 16'(-420);
			7856: out = 16'(3194);
			7857: out = 16'(831);
			7858: out = 16'(-1513);
			7859: out = 16'(1704);
			7860: out = 16'(-2030);
			7861: out = 16'(2646);
			7862: out = 16'(-58);
			7863: out = 16'(-1348);
			7864: out = 16'(632);
			7865: out = 16'(-5582);
			7866: out = 16'(1752);
			7867: out = 16'(-1099);
			7868: out = 16'(272);
			7869: out = 16'(988);
			7870: out = 16'(1434);
			7871: out = 16'(-241);
			7872: out = 16'(-248);
			7873: out = 16'(-1005);
			7874: out = 16'(2663);
			7875: out = 16'(112);
			7876: out = 16'(1950);
			7877: out = 16'(1669);
			7878: out = 16'(-3679);
			7879: out = 16'(639);
			7880: out = 16'(2084);
			7881: out = 16'(-1777);
			7882: out = 16'(1008);
			7883: out = 16'(-1854);
			7884: out = 16'(-2544);
			7885: out = 16'(2120);
			7886: out = 16'(-2587);
			7887: out = 16'(242);
			7888: out = 16'(62);
			7889: out = 16'(954);
			7890: out = 16'(108);
			7891: out = 16'(-1765);
			7892: out = 16'(776);
			7893: out = 16'(1934);
			7894: out = 16'(2996);
			7895: out = 16'(2686);
			7896: out = 16'(-1607);
			7897: out = 16'(287);
			7898: out = 16'(-935);
			7899: out = 16'(-627);
			7900: out = 16'(-2463);
			7901: out = 16'(1010);
			7902: out = 16'(1158);
			7903: out = 16'(69);
			7904: out = 16'(36);
			7905: out = 16'(246);
			7906: out = 16'(1676);
			7907: out = 16'(-309);
			7908: out = 16'(1384);
			7909: out = 16'(2317);
			7910: out = 16'(-569);
			7911: out = 16'(-50);
			7912: out = 16'(-1349);
			7913: out = 16'(2365);
			7914: out = 16'(2549);
			7915: out = 16'(272);
			7916: out = 16'(-18);
			7917: out = 16'(-2794);
			7918: out = 16'(4133);
			7919: out = 16'(-792);
			7920: out = 16'(1617);
			7921: out = 16'(2253);
			7922: out = 16'(878);
			7923: out = 16'(-3621);
			7924: out = 16'(-2817);
			7925: out = 16'(67);
			7926: out = 16'(357);
			7927: out = 16'(529);
			7928: out = 16'(-3403);
			7929: out = 16'(2252);
			7930: out = 16'(-3980);
			7931: out = 16'(2437);
			7932: out = 16'(32);
			7933: out = 16'(1958);
			7934: out = 16'(767);
			7935: out = 16'(-4151);
			7936: out = 16'(1028);
			7937: out = 16'(456);
			7938: out = 16'(-92);
			7939: out = 16'(-118);
			7940: out = 16'(1185);
			7941: out = 16'(-142);
			7942: out = 16'(243);
			7943: out = 16'(-634);
			7944: out = 16'(-2283);
			7945: out = 16'(1093);
			7946: out = 16'(-51);
			7947: out = 16'(1338);
			7948: out = 16'(-3269);
			7949: out = 16'(-848);
			7950: out = 16'(767);
			7951: out = 16'(-786);
			7952: out = 16'(-455);
			7953: out = 16'(1811);
			7954: out = 16'(1579);
			7955: out = 16'(855);
			7956: out = 16'(-1608);
			7957: out = 16'(1612);
			7958: out = 16'(-655);
			7959: out = 16'(1441);
			7960: out = 16'(-227);
			7961: out = 16'(-2268);
			7962: out = 16'(-2073);
			7963: out = 16'(-438);
			7964: out = 16'(-2609);
			7965: out = 16'(1185);
			7966: out = 16'(43);
			7967: out = 16'(-1221);
			7968: out = 16'(788);
			7969: out = 16'(-4014);
			7970: out = 16'(-715);
			7971: out = 16'(7);
			7972: out = 16'(243);
			7973: out = 16'(1676);
			7974: out = 16'(249);
			7975: out = 16'(2204);
			7976: out = 16'(-5817);
			7977: out = 16'(627);
			7978: out = 16'(1382);
			7979: out = 16'(-2613);
			7980: out = 16'(405);
			7981: out = 16'(-1726);
			7982: out = 16'(-1148);
			7983: out = 16'(703);
			7984: out = 16'(76);
			7985: out = 16'(215);
			7986: out = 16'(-1196);
			7987: out = 16'(-1721);
			7988: out = 16'(-1768);
			7989: out = 16'(-227);
			7990: out = 16'(-2088);
			7991: out = 16'(2043);
			7992: out = 16'(1185);
			7993: out = 16'(-3194);
			7994: out = 16'(1700);
			7995: out = 16'(-452);
			7996: out = 16'(1377);
			7997: out = 16'(-417);
			7998: out = 16'(1570);
			7999: out = 16'(3871);
			8000: out = 16'(-3062);
			8001: out = 16'(-1999);
			8002: out = 16'(-1830);
			8003: out = 16'(-410);
			8004: out = 16'(424);
			8005: out = 16'(923);
			8006: out = 16'(-2633);
			8007: out = 16'(225);
			8008: out = 16'(-1158);
			8009: out = 16'(-3240);
			8010: out = 16'(-1594);
			8011: out = 16'(-1000);
			8012: out = 16'(1514);
			8013: out = 16'(159);
			8014: out = 16'(-1189);
			8015: out = 16'(99);
			8016: out = 16'(1217);
			8017: out = 16'(-534);
			8018: out = 16'(-470);
			8019: out = 16'(-2045);
			8020: out = 16'(1233);
			8021: out = 16'(-4226);
			8022: out = 16'(592);
			8023: out = 16'(1367);
			8024: out = 16'(14);
			8025: out = 16'(1358);
			8026: out = 16'(-120);
			8027: out = 16'(-674);
			8028: out = 16'(206);
			8029: out = 16'(-2356);
			8030: out = 16'(2566);
			8031: out = 16'(227);
			8032: out = 16'(-1423);
			8033: out = 16'(1814);
			8034: out = 16'(-175);
			8035: out = 16'(1580);
			8036: out = 16'(1884);
			8037: out = 16'(1931);
			8038: out = 16'(-2172);
			8039: out = 16'(2274);
			8040: out = 16'(-2391);
			8041: out = 16'(854);
			8042: out = 16'(222);
			8043: out = 16'(-714);
			8044: out = 16'(1763);
			8045: out = 16'(-4514);
			8046: out = 16'(2214);
			8047: out = 16'(1654);
			8048: out = 16'(-2182);
			8049: out = 16'(2305);
			8050: out = 16'(-1126);
			8051: out = 16'(1054);
			8052: out = 16'(-2290);
			8053: out = 16'(-2757);
			8054: out = 16'(-682);
			8055: out = 16'(-823);
			8056: out = 16'(-209);
			8057: out = 16'(2701);
			8058: out = 16'(-355);
			8059: out = 16'(2222);
			8060: out = 16'(-2437);
			8061: out = 16'(1317);
			8062: out = 16'(76);
			8063: out = 16'(676);
			8064: out = 16'(266);
			8065: out = 16'(-550);
			8066: out = 16'(149);
			8067: out = 16'(-64);
			8068: out = 16'(-687);
			8069: out = 16'(1069);
			8070: out = 16'(432);
			8071: out = 16'(1102);
			8072: out = 16'(-1032);
			8073: out = 16'(743);
			8074: out = 16'(-727);
			8075: out = 16'(-136);
			8076: out = 16'(601);
			8077: out = 16'(636);
			8078: out = 16'(3448);
			8079: out = 16'(-2136);
			8080: out = 16'(-1023);
			8081: out = 16'(1268);
			8082: out = 16'(1573);
			8083: out = 16'(1053);
			8084: out = 16'(-500);
			8085: out = 16'(-28);
			8086: out = 16'(-42);
			8087: out = 16'(-169);
			8088: out = 16'(230);
			8089: out = 16'(2227);
			8090: out = 16'(802);
			8091: out = 16'(-145);
			8092: out = 16'(-3042);
			8093: out = 16'(-1209);
			8094: out = 16'(814);
			8095: out = 16'(1677);
			8096: out = 16'(408);
			8097: out = 16'(1280);
			8098: out = 16'(-895);
			8099: out = 16'(-1308);
			8100: out = 16'(526);
			8101: out = 16'(2617);
			8102: out = 16'(276);
			8103: out = 16'(1103);
			8104: out = 16'(-1581);
			8105: out = 16'(-336);
			8106: out = 16'(138);
			8107: out = 16'(108);
			8108: out = 16'(-1451);
			8109: out = 16'(2095);
			8110: out = 16'(1913);
			8111: out = 16'(932);
			8112: out = 16'(431);
			8113: out = 16'(708);
			8114: out = 16'(1023);
			8115: out = 16'(-2065);
			8116: out = 16'(4379);
			8117: out = 16'(-2120);
			8118: out = 16'(1197);
			8119: out = 16'(1236);
			8120: out = 16'(-1495);
			8121: out = 16'(3796);
			8122: out = 16'(23);
			8123: out = 16'(1092);
			8124: out = 16'(-5404);
			8125: out = 16'(1017);
			8126: out = 16'(1590);
			8127: out = 16'(-279);
			8128: out = 16'(3174);
			8129: out = 16'(-2069);
			8130: out = 16'(1941);
			8131: out = 16'(-3014);
			8132: out = 16'(-1282);
			8133: out = 16'(-1681);
			8134: out = 16'(1401);
			8135: out = 16'(152);
			8136: out = 16'(-2104);
			8137: out = 16'(339);
			8138: out = 16'(-1704);
			8139: out = 16'(2791);
			8140: out = 16'(328);
			8141: out = 16'(-1217);
			8142: out = 16'(1639);
			8143: out = 16'(-445);
			8144: out = 16'(-924);
			8145: out = 16'(2489);
			8146: out = 16'(1071);
			8147: out = 16'(-658);
			8148: out = 16'(1001);
			8149: out = 16'(-32);
			8150: out = 16'(-1224);
			8151: out = 16'(61);
			8152: out = 16'(-1912);
			8153: out = 16'(1652);
			8154: out = 16'(732);
			8155: out = 16'(659);
			8156: out = 16'(-5659);
			8157: out = 16'(-1616);
			8158: out = 16'(-877);
			8159: out = 16'(-404);
			8160: out = 16'(1446);
			8161: out = 16'(865);
			8162: out = 16'(-767);
			8163: out = 16'(-257);
			8164: out = 16'(-933);
			8165: out = 16'(1997);
			8166: out = 16'(-551);
			8167: out = 16'(-1075);
			8168: out = 16'(-672);
			8169: out = 16'(575);
			8170: out = 16'(-1165);
			8171: out = 16'(425);
			8172: out = 16'(-125);
			8173: out = 16'(1506);
			8174: out = 16'(-2640);
			8175: out = 16'(-333);
			8176: out = 16'(-2007);
			8177: out = 16'(-933);
			8178: out = 16'(1679);
			8179: out = 16'(-105);
			8180: out = 16'(718);
			8181: out = 16'(232);
			8182: out = 16'(640);
			8183: out = 16'(-3584);
			8184: out = 16'(514);
			8185: out = 16'(-246);
			8186: out = 16'(-71);
			8187: out = 16'(1749);
			8188: out = 16'(-473);
			8189: out = 16'(-1760);
			8190: out = 16'(1554);
			8191: out = 16'(-742);
			8192: out = 16'(1158);
			8193: out = 16'(301);
			8194: out = 16'(-1829);
			8195: out = 16'(235);
			8196: out = 16'(2071);
			8197: out = 16'(206);
			8198: out = 16'(2386);
			8199: out = 16'(-2429);
			8200: out = 16'(1964);
			8201: out = 16'(-4167);
			8202: out = 16'(924);
			8203: out = 16'(1626);
			8204: out = 16'(-1052);
			8205: out = 16'(1253);
			8206: out = 16'(-278);
			8207: out = 16'(37);
			8208: out = 16'(-3689);
			8209: out = 16'(-609);
			8210: out = 16'(-1700);
			8211: out = 16'(1413);
			8212: out = 16'(10);
			8213: out = 16'(431);
			8214: out = 16'(1530);
			8215: out = 16'(-1955);
			8216: out = 16'(70);
			8217: out = 16'(-690);
			8218: out = 16'(1210);
			8219: out = 16'(-1274);
			8220: out = 16'(-750);
			8221: out = 16'(-115);
			8222: out = 16'(-1360);
			8223: out = 16'(2741);
			8224: out = 16'(-706);
			8225: out = 16'(-804);
			8226: out = 16'(-1289);
			8227: out = 16'(-2031);
			8228: out = 16'(271);
			8229: out = 16'(-386);
			8230: out = 16'(2279);
			8231: out = 16'(1027);
			8232: out = 16'(472);
			8233: out = 16'(-2467);
			8234: out = 16'(-421);
			8235: out = 16'(-32);
			8236: out = 16'(-1180);
			8237: out = 16'(2290);
			8238: out = 16'(-1323);
			8239: out = 16'(3280);
			8240: out = 16'(-2451);
			8241: out = 16'(608);
			8242: out = 16'(-15);
			8243: out = 16'(-1611);
			8244: out = 16'(1772);
			8245: out = 16'(106);
			8246: out = 16'(-918);
			8247: out = 16'(-62);
			8248: out = 16'(-651);
			8249: out = 16'(-243);
			8250: out = 16'(240);
			8251: out = 16'(-36);
			8252: out = 16'(598);
			8253: out = 16'(-2570);
			8254: out = 16'(406);
			8255: out = 16'(758);
			8256: out = 16'(-1809);
			8257: out = 16'(2890);
			8258: out = 16'(-4296);
			8259: out = 16'(1080);
			8260: out = 16'(-2466);
			8261: out = 16'(-539);
			8262: out = 16'(584);
			8263: out = 16'(1291);
			8264: out = 16'(2134);
			8265: out = 16'(-1304);
			8266: out = 16'(1271);
			8267: out = 16'(-1580);
			8268: out = 16'(597);
			8269: out = 16'(1017);
			8270: out = 16'(-158);
			8271: out = 16'(714);
			8272: out = 16'(-1523);
			8273: out = 16'(718);
			8274: out = 16'(-1513);
			8275: out = 16'(791);
			8276: out = 16'(-541);
			8277: out = 16'(-1519);
			8278: out = 16'(81);
			8279: out = 16'(-852);
			8280: out = 16'(3235);
			8281: out = 16'(1392);
			8282: out = 16'(1422);
			8283: out = 16'(-83);
			8284: out = 16'(-522);
			8285: out = 16'(58);
			8286: out = 16'(-900);
			8287: out = 16'(2637);
			8288: out = 16'(-3065);
			8289: out = 16'(375);
			8290: out = 16'(-55);
			8291: out = 16'(-1858);
			8292: out = 16'(716);
			8293: out = 16'(421);
			8294: out = 16'(-1643);
			8295: out = 16'(-209);
			8296: out = 16'(1923);
			8297: out = 16'(-155);
			8298: out = 16'(-202);
			8299: out = 16'(-615);
			8300: out = 16'(-2755);
			8301: out = 16'(2690);
			8302: out = 16'(-79);
			8303: out = 16'(2458);
			8304: out = 16'(-1062);
			8305: out = 16'(92);
			8306: out = 16'(-242);
			8307: out = 16'(411);
			8308: out = 16'(1930);
			8309: out = 16'(-473);
			8310: out = 16'(330);
			8311: out = 16'(-1166);
			8312: out = 16'(-2506);
			8313: out = 16'(982);
			8314: out = 16'(2086);
			8315: out = 16'(-585);
			8316: out = 16'(1766);
			8317: out = 16'(-425);
			8318: out = 16'(-4333);
			8319: out = 16'(-598);
			8320: out = 16'(-1447);
			8321: out = 16'(955);
			8322: out = 16'(-241);
			8323: out = 16'(712);
			8324: out = 16'(-726);
			8325: out = 16'(1170);
			8326: out = 16'(-2002);
			8327: out = 16'(536);
			8328: out = 16'(-1696);
			8329: out = 16'(-1161);
			8330: out = 16'(-973);
			8331: out = 16'(-708);
			8332: out = 16'(-883);
			8333: out = 16'(1422);
			8334: out = 16'(3026);
			8335: out = 16'(1095);
			8336: out = 16'(-1230);
			8337: out = 16'(154);
			8338: out = 16'(-1899);
			8339: out = 16'(-60);
			8340: out = 16'(-128);
			8341: out = 16'(973);
			8342: out = 16'(-807);
			8343: out = 16'(382);
			8344: out = 16'(-472);
			8345: out = 16'(1034);
			8346: out = 16'(849);
			8347: out = 16'(298);
			8348: out = 16'(-1047);
			8349: out = 16'(1032);
			8350: out = 16'(-233);
			8351: out = 16'(359);
			8352: out = 16'(1136);
			8353: out = 16'(-199);
			8354: out = 16'(-1487);
			8355: out = 16'(1245);
			8356: out = 16'(-2151);
			8357: out = 16'(-194);
			8358: out = 16'(-307);
			8359: out = 16'(1229);
			8360: out = 16'(-1652);
			8361: out = 16'(1780);
			8362: out = 16'(-2312);
			8363: out = 16'(-2357);
			8364: out = 16'(646);
			8365: out = 16'(-1406);
			8366: out = 16'(3945);
			8367: out = 16'(-571);
			8368: out = 16'(1638);
			8369: out = 16'(-186);
			8370: out = 16'(1052);
			8371: out = 16'(-331);
			8372: out = 16'(-1038);
			8373: out = 16'(304);
			8374: out = 16'(973);
			8375: out = 16'(367);
			8376: out = 16'(-1210);
			8377: out = 16'(1535);
			8378: out = 16'(9);
			8379: out = 16'(1396);
			8380: out = 16'(252);
			8381: out = 16'(-4371);
			8382: out = 16'(867);
			8383: out = 16'(-982);
			8384: out = 16'(1064);
			8385: out = 16'(744);
			8386: out = 16'(1254);
			8387: out = 16'(210);
			8388: out = 16'(-304);
			8389: out = 16'(-833);
			8390: out = 16'(57);
			8391: out = 16'(-543);
			8392: out = 16'(1118);
			8393: out = 16'(-2669);
			8394: out = 16'(2256);
			8395: out = 16'(-2175);
			8396: out = 16'(33);
			8397: out = 16'(-1450);
			8398: out = 16'(317);
			8399: out = 16'(1335);
			8400: out = 16'(-2646);
			8401: out = 16'(862);
			8402: out = 16'(-1242);
			8403: out = 16'(172);
			8404: out = 16'(1776);
			8405: out = 16'(670);
			8406: out = 16'(323);
			8407: out = 16'(-1032);
			8408: out = 16'(-294);
			8409: out = 16'(1160);
			8410: out = 16'(1008);
			8411: out = 16'(2225);
			8412: out = 16'(50);
			8413: out = 16'(-94);
			8414: out = 16'(319);
			8415: out = 16'(-495);
			8416: out = 16'(1028);
			8417: out = 16'(-1024);
			8418: out = 16'(975);
			8419: out = 16'(-233);
			8420: out = 16'(811);
			8421: out = 16'(-1067);
			8422: out = 16'(662);
			8423: out = 16'(1044);
			8424: out = 16'(-1939);
			8425: out = 16'(2099);
			8426: out = 16'(1126);
			8427: out = 16'(1149);
			8428: out = 16'(126);
			8429: out = 16'(-2123);
			8430: out = 16'(419);
			8431: out = 16'(-936);
			8432: out = 16'(1451);
			8433: out = 16'(475);
			8434: out = 16'(-764);
			8435: out = 16'(1466);
			8436: out = 16'(230);
			8437: out = 16'(3172);
			8438: out = 16'(-1538);
			8439: out = 16'(-45);
			8440: out = 16'(-647);
			8441: out = 16'(-2486);
			8442: out = 16'(322);
			8443: out = 16'(1123);
			8444: out = 16'(-400);
			8445: out = 16'(-1727);
			8446: out = 16'(93);
			8447: out = 16'(-452);
			8448: out = 16'(323);
			8449: out = 16'(1005);
			8450: out = 16'(-808);
			8451: out = 16'(1308);
			8452: out = 16'(-384);
			8453: out = 16'(-34);
			8454: out = 16'(1145);
			8455: out = 16'(-1269);
			8456: out = 16'(931);
			8457: out = 16'(1230);
			8458: out = 16'(588);
			8459: out = 16'(103);
			8460: out = 16'(-1038);
			8461: out = 16'(1568);
			8462: out = 16'(-1237);
			8463: out = 16'(1382);
			8464: out = 16'(-647);
			8465: out = 16'(434);
			8466: out = 16'(-3222);
			8467: out = 16'(664);
			8468: out = 16'(452);
			8469: out = 16'(504);
			8470: out = 16'(667);
			8471: out = 16'(273);
			8472: out = 16'(1359);
			8473: out = 16'(-1889);
			8474: out = 16'(-2105);
			8475: out = 16'(1754);
			8476: out = 16'(-1178);
			8477: out = 16'(941);
			8478: out = 16'(1185);
			8479: out = 16'(-1885);
			8480: out = 16'(-186);
			8481: out = 16'(-703);
			8482: out = 16'(-1996);
			8483: out = 16'(73);
			8484: out = 16'(265);
			8485: out = 16'(2260);
			8486: out = 16'(-2026);
			8487: out = 16'(481);
			8488: out = 16'(112);
			8489: out = 16'(110);
			8490: out = 16'(729);
			8491: out = 16'(550);
			8492: out = 16'(-3130);
			8493: out = 16'(3151);
			8494: out = 16'(-1205);
			8495: out = 16'(1145);
			8496: out = 16'(1528);
			8497: out = 16'(717);
			8498: out = 16'(-3587);
			8499: out = 16'(-398);
			8500: out = 16'(1057);
			8501: out = 16'(19);
			8502: out = 16'(1397);
			8503: out = 16'(554);
			8504: out = 16'(566);
			8505: out = 16'(-705);
			8506: out = 16'(468);
			8507: out = 16'(-2823);
			8508: out = 16'(650);
			8509: out = 16'(2501);
			8510: out = 16'(-3949);
			8511: out = 16'(1699);
			8512: out = 16'(-1927);
			8513: out = 16'(169);
			8514: out = 16'(-231);
			8515: out = 16'(350);
			8516: out = 16'(-674);
			8517: out = 16'(32);
			8518: out = 16'(-1671);
			8519: out = 16'(1282);
			8520: out = 16'(2443);
			8521: out = 16'(1736);
			8522: out = 16'(-1235);
			8523: out = 16'(-65);
			8524: out = 16'(-1131);
			8525: out = 16'(-109);
			8526: out = 16'(-211);
			8527: out = 16'(1369);
			8528: out = 16'(126);
			8529: out = 16'(121);
			8530: out = 16'(947);
			8531: out = 16'(-1317);
			8532: out = 16'(1079);
			8533: out = 16'(1029);
			8534: out = 16'(254);
			8535: out = 16'(-12);
			8536: out = 16'(-1712);
			8537: out = 16'(404);
			8538: out = 16'(-1215);
			8539: out = 16'(942);
			8540: out = 16'(-117);
			8541: out = 16'(-144);
			8542: out = 16'(693);
			8543: out = 16'(-1343);
			8544: out = 16'(32);
			8545: out = 16'(-985);
			8546: out = 16'(1512);
			8547: out = 16'(-196);
			8548: out = 16'(-26);
			8549: out = 16'(-880);
			8550: out = 16'(-2162);
			8551: out = 16'(1485);
			8552: out = 16'(-25);
			8553: out = 16'(1239);
			8554: out = 16'(930);
			8555: out = 16'(-1200);
			8556: out = 16'(-702);
			8557: out = 16'(-1235);
			8558: out = 16'(268);
			8559: out = 16'(-332);
			8560: out = 16'(-1248);
			8561: out = 16'(-908);
			8562: out = 16'(-451);
			8563: out = 16'(611);
			8564: out = 16'(361);
			8565: out = 16'(471);
			8566: out = 16'(-135);
			8567: out = 16'(-436);
			8568: out = 16'(-1429);
			8569: out = 16'(-269);
			8570: out = 16'(1990);
			8571: out = 16'(300);
			8572: out = 16'(-103);
			8573: out = 16'(-1364);
			8574: out = 16'(604);
			8575: out = 16'(-2162);
			8576: out = 16'(531);
			8577: out = 16'(976);
			8578: out = 16'(-688);
			8579: out = 16'(1240);
			8580: out = 16'(-281);
			8581: out = 16'(-133);
			8582: out = 16'(1244);
			8583: out = 16'(-1441);
			8584: out = 16'(-110);
			8585: out = 16'(-1015);
			8586: out = 16'(1284);
			8587: out = 16'(-1272);
			8588: out = 16'(-10);
			8589: out = 16'(-425);
			8590: out = 16'(1831);
			8591: out = 16'(-31);
			8592: out = 16'(-1171);
			8593: out = 16'(591);
			8594: out = 16'(-189);
			8595: out = 16'(992);
			8596: out = 16'(-586);
			8597: out = 16'(1193);
			8598: out = 16'(-379);
			8599: out = 16'(-803);
			8600: out = 16'(597);
			8601: out = 16'(-367);
			8602: out = 16'(1064);
			8603: out = 16'(-137);
			8604: out = 16'(-176);
			8605: out = 16'(-767);
			8606: out = 16'(295);
			8607: out = 16'(-534);
			8608: out = 16'(173);
			8609: out = 16'(-1028);
			8610: out = 16'(-1653);
			8611: out = 16'(1503);
			8612: out = 16'(-3858);
			8613: out = 16'(1058);
			8614: out = 16'(458);
			8615: out = 16'(-1413);
			8616: out = 16'(363);
			8617: out = 16'(-706);
			8618: out = 16'(2537);
			8619: out = 16'(-1780);
			8620: out = 16'(162);
			8621: out = 16'(-1140);
			8622: out = 16'(2134);
			8623: out = 16'(302);
			8624: out = 16'(-512);
			8625: out = 16'(-49);
			8626: out = 16'(257);
			8627: out = 16'(-904);
			8628: out = 16'(-1167);
			8629: out = 16'(1670);
			8630: out = 16'(-1715);
			8631: out = 16'(1969);
			8632: out = 16'(1509);
			8633: out = 16'(-1535);
			8634: out = 16'(2479);
			8635: out = 16'(-239);
			8636: out = 16'(-694);
			8637: out = 16'(211);
			8638: out = 16'(-1092);
			8639: out = 16'(1896);
			8640: out = 16'(-1703);
			8641: out = 16'(2322);
			8642: out = 16'(-1578);
			8643: out = 16'(-141);
			8644: out = 16'(-541);
			8645: out = 16'(-33);
			8646: out = 16'(-446);
			8647: out = 16'(-1758);
			8648: out = 16'(-865);
			8649: out = 16'(-192);
			8650: out = 16'(2982);
			8651: out = 16'(-2930);
			8652: out = 16'(2264);
			8653: out = 16'(852);
			8654: out = 16'(-476);
			8655: out = 16'(958);
			8656: out = 16'(2000);
			8657: out = 16'(1638);
			8658: out = 16'(-95);
			8659: out = 16'(-116);
			8660: out = 16'(-214);
			8661: out = 16'(-43);
			8662: out = 16'(-192);
			8663: out = 16'(1194);
			8664: out = 16'(-2069);
			8665: out = 16'(2261);
			8666: out = 16'(-151);
			8667: out = 16'(-326);
			8668: out = 16'(376);
			8669: out = 16'(-1747);
			8670: out = 16'(699);
			8671: out = 16'(1355);
			8672: out = 16'(-3244);
			8673: out = 16'(2744);
			8674: out = 16'(-2848);
			8675: out = 16'(964);
			8676: out = 16'(-424);
			8677: out = 16'(-1470);
			8678: out = 16'(70);
			8679: out = 16'(-2487);
			8680: out = 16'(308);
			8681: out = 16'(326);
			8682: out = 16'(957);
			8683: out = 16'(196);
			8684: out = 16'(279);
			8685: out = 16'(-1799);
			8686: out = 16'(-584);
			8687: out = 16'(-38);
			8688: out = 16'(204);
			8689: out = 16'(810);
			8690: out = 16'(-792);
			8691: out = 16'(861);
			8692: out = 16'(-1079);
			8693: out = 16'(467);
			8694: out = 16'(2164);
			8695: out = 16'(219);
			8696: out = 16'(-2184);
			8697: out = 16'(2061);
			8698: out = 16'(-1557);
			8699: out = 16'(-43);
			8700: out = 16'(-29);
			8701: out = 16'(-109);
			8702: out = 16'(-418);
			8703: out = 16'(-148);
			8704: out = 16'(-667);
			8705: out = 16'(1112);
			8706: out = 16'(-909);
			8707: out = 16'(-413);
			8708: out = 16'(203);
			8709: out = 16'(1819);
			8710: out = 16'(-561);
			8711: out = 16'(-1253);
			8712: out = 16'(-2320);
			8713: out = 16'(189);
			8714: out = 16'(-948);
			8715: out = 16'(1974);
			8716: out = 16'(-1990);
			8717: out = 16'(542);
			8718: out = 16'(-1314);
			8719: out = 16'(285);
			8720: out = 16'(580);
			8721: out = 16'(830);
			8722: out = 16'(-61);
			8723: out = 16'(1214);
			8724: out = 16'(-519);
			8725: out = 16'(952);
			8726: out = 16'(-985);
			8727: out = 16'(-40);
			8728: out = 16'(-377);
			8729: out = 16'(-2073);
			8730: out = 16'(384);
			8731: out = 16'(-1841);
			8732: out = 16'(156);
			8733: out = 16'(1006);
			8734: out = 16'(1318);
			8735: out = 16'(-2049);
			8736: out = 16'(3103);
			8737: out = 16'(229);
			8738: out = 16'(144);
			8739: out = 16'(973);
			8740: out = 16'(-385);
			8741: out = 16'(-162);
			8742: out = 16'(189);
			8743: out = 16'(422);
			8744: out = 16'(-1198);
			8745: out = 16'(420);
			8746: out = 16'(-1828);
			8747: out = 16'(-440);
			8748: out = 16'(-2177);
			8749: out = 16'(3026);
			8750: out = 16'(-2502);
			8751: out = 16'(1013);
			8752: out = 16'(-76);
			8753: out = 16'(-757);
			8754: out = 16'(-16);
			8755: out = 16'(-1024);
			8756: out = 16'(-1142);
			8757: out = 16'(372);
			8758: out = 16'(559);
			8759: out = 16'(-279);
			8760: out = 16'(-156);
			8761: out = 16'(-5);
			8762: out = 16'(-58);
			8763: out = 16'(-1544);
			8764: out = 16'(26);
			8765: out = 16'(-249);
			8766: out = 16'(-283);
			8767: out = 16'(976);
			8768: out = 16'(2060);
			8769: out = 16'(192);
			8770: out = 16'(845);
			8771: out = 16'(-1575);
			8772: out = 16'(129);
			8773: out = 16'(-269);
			8774: out = 16'(-1916);
			8775: out = 16'(507);
			8776: out = 16'(-138);
			8777: out = 16'(973);
			8778: out = 16'(-1657);
			8779: out = 16'(563);
			8780: out = 16'(11);
			8781: out = 16'(-936);
			8782: out = 16'(589);
			8783: out = 16'(-1296);
			8784: out = 16'(195);
			8785: out = 16'(283);
			8786: out = 16'(1);
			8787: out = 16'(-1389);
			8788: out = 16'(2557);
			8789: out = 16'(-1231);
			8790: out = 16'(-272);
			8791: out = 16'(2053);
			8792: out = 16'(-511);
			8793: out = 16'(1384);
			8794: out = 16'(932);
			8795: out = 16'(-1259);
			8796: out = 16'(837);
			8797: out = 16'(-314);
			8798: out = 16'(-445);
			8799: out = 16'(-185);
			8800: out = 16'(467);
			8801: out = 16'(-111);
			8802: out = 16'(-330);
			8803: out = 16'(21);
			8804: out = 16'(308);
			8805: out = 16'(-550);
			8806: out = 16'(-87);
			8807: out = 16'(825);
			8808: out = 16'(390);
			8809: out = 16'(-180);
			8810: out = 16'(-512);
			8811: out = 16'(-431);
			8812: out = 16'(1565);
			8813: out = 16'(-82);
			8814: out = 16'(901);
			8815: out = 16'(-2645);
			8816: out = 16'(754);
			8817: out = 16'(101);
			8818: out = 16'(192);
			8819: out = 16'(-15);
			8820: out = 16'(1568);
			8821: out = 16'(834);
			8822: out = 16'(4);
			8823: out = 16'(864);
			8824: out = 16'(-1912);
			8825: out = 16'(466);
			8826: out = 16'(381);
			8827: out = 16'(1098);
			8828: out = 16'(-1505);
			8829: out = 16'(-664);
			8830: out = 16'(1527);
			8831: out = 16'(-2692);
			8832: out = 16'(2010);
			8833: out = 16'(-1889);
			8834: out = 16'(-330);
			8835: out = 16'(-988);
			8836: out = 16'(28);
			8837: out = 16'(283);
			8838: out = 16'(94);
			8839: out = 16'(59);
			8840: out = 16'(362);
			8841: out = 16'(23);
			8842: out = 16'(-1373);
			8843: out = 16'(372);
			8844: out = 16'(774);
			8845: out = 16'(1142);
			8846: out = 16'(1562);
			8847: out = 16'(-770);
			8848: out = 16'(362);
			8849: out = 16'(-2329);
			8850: out = 16'(730);
			8851: out = 16'(1136);
			8852: out = 16'(-1216);
			8853: out = 16'(61);
			8854: out = 16'(401);
			8855: out = 16'(-629);
			8856: out = 16'(-523);
			8857: out = 16'(-1914);
			8858: out = 16'(322);
			8859: out = 16'(38);
			8860: out = 16'(-8);
			8861: out = 16'(-143);
			8862: out = 16'(1177);
			8863: out = 16'(184);
			8864: out = 16'(-361);
			8865: out = 16'(407);
			8866: out = 16'(-1241);
			8867: out = 16'(-757);
			8868: out = 16'(-316);
			8869: out = 16'(-94);
			8870: out = 16'(140);
			8871: out = 16'(826);
			8872: out = 16'(-545);
			8873: out = 16'(-1519);
			8874: out = 16'(1033);
			8875: out = 16'(105);
			8876: out = 16'(-1584);
			8877: out = 16'(990);
			8878: out = 16'(-25);
			8879: out = 16'(438);
			8880: out = 16'(-235);
			8881: out = 16'(-1832);
			8882: out = 16'(1635);
			8883: out = 16'(-552);
			8884: out = 16'(752);
			8885: out = 16'(479);
			8886: out = 16'(-1150);
			8887: out = 16'(-402);
			8888: out = 16'(-1239);
			8889: out = 16'(440);
			8890: out = 16'(-546);
			8891: out = 16'(2);
			8892: out = 16'(-465);
			8893: out = 16'(348);
			8894: out = 16'(-1244);
			8895: out = 16'(1676);
			8896: out = 16'(-185);
			8897: out = 16'(-13);
			8898: out = 16'(1004);
			8899: out = 16'(6);
			8900: out = 16'(-384);
			8901: out = 16'(402);
			8902: out = 16'(-165);
			8903: out = 16'(165);
			8904: out = 16'(-452);
			8905: out = 16'(-52);
			8906: out = 16'(267);
			8907: out = 16'(-190);
			8908: out = 16'(497);
			8909: out = 16'(-927);
			8910: out = 16'(370);
			8911: out = 16'(-27);
			8912: out = 16'(-763);
			8913: out = 16'(634);
			8914: out = 16'(39);
			8915: out = 16'(0);
			8916: out = 16'(14);
			8917: out = 16'(-301);
			8918: out = 16'(-491);
			8919: out = 16'(793);
			8920: out = 16'(-1558);
			8921: out = 16'(4);
			8922: out = 16'(-146);
			8923: out = 16'(945);
			8924: out = 16'(190);
			8925: out = 16'(-1375);
			8926: out = 16'(208);
			8927: out = 16'(-341);
			8928: out = 16'(-350);
			8929: out = 16'(934);
			8930: out = 16'(-258);
			8931: out = 16'(-149);
			8932: out = 16'(185);
			8933: out = 16'(-1129);
			8934: out = 16'(2259);
			8935: out = 16'(-961);
			8936: out = 16'(464);
			8937: out = 16'(-75);
			8938: out = 16'(-1116);
			8939: out = 16'(-1415);
			8940: out = 16'(534);
			8941: out = 16'(-197);
			8942: out = 16'(753);
			8943: out = 16'(-659);
			8944: out = 16'(623);
			8945: out = 16'(-1041);
			8946: out = 16'(-486);
			8947: out = 16'(1017);
			8948: out = 16'(-39);
			8949: out = 16'(811);
			8950: out = 16'(28);
			8951: out = 16'(308);
			8952: out = 16'(-731);
			8953: out = 16'(572);
			8954: out = 16'(-492);
			8955: out = 16'(275);
			8956: out = 16'(101);
			8957: out = 16'(257);
			8958: out = 16'(-647);
			8959: out = 16'(-1174);
			8960: out = 16'(560);
			8961: out = 16'(-793);
			8962: out = 16'(753);
			8963: out = 16'(180);
			8964: out = 16'(1197);
			8965: out = 16'(845);
			8966: out = 16'(261);
			8967: out = 16'(-27);
			8968: out = 16'(742);
			8969: out = 16'(-1322);
			8970: out = 16'(104);
			8971: out = 16'(-956);
			8972: out = 16'(323);
			8973: out = 16'(215);
			8974: out = 16'(153);
			8975: out = 16'(113);
			8976: out = 16'(-24);
			8977: out = 16'(-612);
			8978: out = 16'(-780);
			8979: out = 16'(-665);
			8980: out = 16'(-1026);
			8981: out = 16'(-553);
			8982: out = 16'(87);
			8983: out = 16'(148);
			8984: out = 16'(1073);
			8985: out = 16'(-1703);
			8986: out = 16'(1720);
			8987: out = 16'(-1494);
			8988: out = 16'(1327);
			8989: out = 16'(-96);
			8990: out = 16'(-647);
			8991: out = 16'(-298);
			8992: out = 16'(-563);
			8993: out = 16'(127);
			8994: out = 16'(1081);
			8995: out = 16'(1064);
			8996: out = 16'(123);
			8997: out = 16'(-143);
			8998: out = 16'(1272);
			8999: out = 16'(-149);
			9000: out = 16'(-62);
			9001: out = 16'(-51);
			9002: out = 16'(-114);
			9003: out = 16'(370);
			9004: out = 16'(-1015);
			9005: out = 16'(814);
			9006: out = 16'(1153);
			9007: out = 16'(9);
			9008: out = 16'(837);
			9009: out = 16'(-454);
			9010: out = 16'(-16);
			9011: out = 16'(-444);
			9012: out = 16'(1148);
			9013: out = 16'(-1483);
			9014: out = 16'(669);
			9015: out = 16'(87);
			9016: out = 16'(1093);
			9017: out = 16'(-785);
			9018: out = 16'(1647);
			9019: out = 16'(-1522);
			9020: out = 16'(1083);
			9021: out = 16'(-77);
			9022: out = 16'(46);
			9023: out = 16'(-1403);
			9024: out = 16'(204);
			9025: out = 16'(306);
			9026: out = 16'(-732);
			9027: out = 16'(1340);
			9028: out = 16'(-945);
			9029: out = 16'(-490);
			9030: out = 16'(-1221);
			9031: out = 16'(-266);
			9032: out = 16'(-87);
			9033: out = 16'(-303);
			9034: out = 16'(422);
			9035: out = 16'(-479);
			9036: out = 16'(764);
			9037: out = 16'(333);
			9038: out = 16'(-37);
			9039: out = 16'(239);
			9040: out = 16'(-865);
			9041: out = 16'(-1272);
			9042: out = 16'(-115);
			9043: out = 16'(20);
			9044: out = 16'(1053);
			9045: out = 16'(-782);
			9046: out = 16'(2322);
			9047: out = 16'(-3576);
			9048: out = 16'(774);
			9049: out = 16'(-293);
			9050: out = 16'(575);
			9051: out = 16'(1271);
			9052: out = 16'(4);
			9053: out = 16'(1624);
			9054: out = 16'(-2065);
			9055: out = 16'(1458);
			9056: out = 16'(-836);
			9057: out = 16'(-67);
			9058: out = 16'(-884);
			9059: out = 16'(-27);
			9060: out = 16'(1841);
			9061: out = 16'(-1398);
			9062: out = 16'(-209);
			9063: out = 16'(-1217);
			9064: out = 16'(-296);
			9065: out = 16'(155);
			9066: out = 16'(284);
			9067: out = 16'(1501);
			9068: out = 16'(-636);
			9069: out = 16'(1448);
			9070: out = 16'(-540);
			9071: out = 16'(-55);
			9072: out = 16'(-464);
			9073: out = 16'(324);
			9074: out = 16'(924);
			9075: out = 16'(255);
			9076: out = 16'(1541);
			9077: out = 16'(80);
			9078: out = 16'(-87);
			9079: out = 16'(-1132);
			9080: out = 16'(875);
			9081: out = 16'(-2547);
			9082: out = 16'(98);
			9083: out = 16'(387);
			9084: out = 16'(-289);
			9085: out = 16'(-173);
			9086: out = 16'(-256);
			9087: out = 16'(592);
			9088: out = 16'(542);
			9089: out = 16'(-293);
			9090: out = 16'(556);
			9091: out = 16'(-86);
			9092: out = 16'(-159);
			9093: out = 16'(-1503);
			9094: out = 16'(232);
			9095: out = 16'(-599);
			9096: out = 16'(569);
			9097: out = 16'(-516);
			9098: out = 16'(117);
			9099: out = 16'(-707);
			9100: out = 16'(248);
			9101: out = 16'(243);
			9102: out = 16'(181);
			9103: out = 16'(673);
			9104: out = 16'(-257);
			9105: out = 16'(779);
			9106: out = 16'(-29);
			9107: out = 16'(109);
			9108: out = 16'(1262);
			9109: out = 16'(-535);
			9110: out = 16'(478);
			9111: out = 16'(695);
			9112: out = 16'(-566);
			9113: out = 16'(-488);
			9114: out = 16'(122);
			9115: out = 16'(-199);
			9116: out = 16'(-431);
			9117: out = 16'(573);
			9118: out = 16'(0);
			9119: out = 16'(558);
			9120: out = 16'(-998);
			9121: out = 16'(472);
			9122: out = 16'(-362);
			9123: out = 16'(-55);
			9124: out = 16'(1207);
			9125: out = 16'(-1133);
			9126: out = 16'(-216);
			9127: out = 16'(-335);
			9128: out = 16'(-638);
			9129: out = 16'(996);
			9130: out = 16'(655);
			9131: out = 16'(-449);
			9132: out = 16'(602);
			9133: out = 16'(-276);
			9134: out = 16'(606);
			9135: out = 16'(1068);
			9136: out = 16'(-475);
			9137: out = 16'(-520);
			9138: out = 16'(736);
			9139: out = 16'(-286);
			9140: out = 16'(-400);
			9141: out = 16'(4);
			9142: out = 16'(-272);
			9143: out = 16'(-491);
			9144: out = 16'(-462);
			9145: out = 16'(206);
			9146: out = 16'(-866);
			9147: out = 16'(775);
			9148: out = 16'(-30);
			9149: out = 16'(200);
			9150: out = 16'(-1329);
			9151: out = 16'(625);
			9152: out = 16'(-1845);
			9153: out = 16'(-495);
			9154: out = 16'(73);
			9155: out = 16'(-398);
			9156: out = 16'(20);
			9157: out = 16'(798);
			9158: out = 16'(376);
			9159: out = 16'(-155);
			9160: out = 16'(432);
			9161: out = 16'(-389);
			9162: out = 16'(912);
			9163: out = 16'(389);
			9164: out = 16'(-1959);
			9165: out = 16'(141);
			9166: out = 16'(673);
			9167: out = 16'(-316);
			9168: out = 16'(668);
			9169: out = 16'(-103);
			9170: out = 16'(-1497);
			9171: out = 16'(814);
			9172: out = 16'(-8);
			9173: out = 16'(-613);
			9174: out = 16'(270);
			9175: out = 16'(237);
			9176: out = 16'(-376);
			9177: out = 16'(-710);
			9178: out = 16'(-1077);
			9179: out = 16'(325);
			9180: out = 16'(114);
			9181: out = 16'(256);
			9182: out = 16'(41);
			9183: out = 16'(-255);
			9184: out = 16'(1376);
			9185: out = 16'(-768);
			9186: out = 16'(898);
			9187: out = 16'(-110);
			9188: out = 16'(-1071);
			9189: out = 16'(835);
			9190: out = 16'(-241);
			9191: out = 16'(530);
			9192: out = 16'(-706);
			9193: out = 16'(1003);
			9194: out = 16'(-78);
			9195: out = 16'(-460);
			9196: out = 16'(1010);
			9197: out = 16'(-1714);
			9198: out = 16'(815);
			9199: out = 16'(-907);
			9200: out = 16'(1685);
			9201: out = 16'(-1201);
			9202: out = 16'(250);
			9203: out = 16'(58);
			9204: out = 16'(-1388);
			9205: out = 16'(811);
			9206: out = 16'(-627);
			9207: out = 16'(386);
			9208: out = 16'(562);
			9209: out = 16'(-551);
			9210: out = 16'(1439);
			9211: out = 16'(-222);
			9212: out = 16'(1055);
			9213: out = 16'(-1330);
			9214: out = 16'(813);
			9215: out = 16'(-1128);
			9216: out = 16'(616);
			9217: out = 16'(-1945);
			9218: out = 16'(954);
			9219: out = 16'(-697);
			9220: out = 16'(168);
			9221: out = 16'(692);
			9222: out = 16'(-862);
			9223: out = 16'(1838);
			9224: out = 16'(69);
			9225: out = 16'(-1171);
			9226: out = 16'(-244);
			9227: out = 16'(-639);
			9228: out = 16'(850);
			9229: out = 16'(-347);
			9230: out = 16'(1074);
			9231: out = 16'(-592);
			9232: out = 16'(-195);
			9233: out = 16'(-218);
			9234: out = 16'(-8);
			9235: out = 16'(849);
			9236: out = 16'(-1138);
			9237: out = 16'(544);
			9238: out = 16'(-748);
			9239: out = 16'(127);
			9240: out = 16'(-835);
			9241: out = 16'(-891);
			9242: out = 16'(84);
			9243: out = 16'(-165);
			9244: out = 16'(1248);
			9245: out = 16'(-1487);
			9246: out = 16'(694);
			9247: out = 16'(-1031);
			9248: out = 16'(-326);
			9249: out = 16'(-376);
			9250: out = 16'(-324);
			9251: out = 16'(637);
			9252: out = 16'(713);
			9253: out = 16'(-791);
			9254: out = 16'(-255);
			9255: out = 16'(-115);
			9256: out = 16'(-2091);
			9257: out = 16'(-839);
			9258: out = 16'(489);
			9259: out = 16'(-967);
			9260: out = 16'(935);
			9261: out = 16'(-130);
			9262: out = 16'(545);
			9263: out = 16'(408);
			9264: out = 16'(-1116);
			9265: out = 16'(-84);
			9266: out = 16'(-1019);
			9267: out = 16'(793);
			9268: out = 16'(-214);
			9269: out = 16'(642);
			9270: out = 16'(-362);
			9271: out = 16'(652);
			9272: out = 16'(-1105);
			9273: out = 16'(-54);
			9274: out = 16'(-905);
			9275: out = 16'(-81);
			9276: out = 16'(1403);
			9277: out = 16'(-1361);
			9278: out = 16'(555);
			9279: out = 16'(-1057);
			9280: out = 16'(-155);
			9281: out = 16'(-939);
			9282: out = 16'(359);
			9283: out = 16'(-212);
			9284: out = 16'(251);
			9285: out = 16'(404);
			9286: out = 16'(701);
			9287: out = 16'(-246);
			9288: out = 16'(236);
			9289: out = 16'(1738);
			9290: out = 16'(-1397);
			9291: out = 16'(1303);
			9292: out = 16'(814);
			9293: out = 16'(-368);
			9294: out = 16'(995);
			9295: out = 16'(-364);
			9296: out = 16'(186);
			9297: out = 16'(-219);
			9298: out = 16'(533);
			9299: out = 16'(-1048);
			9300: out = 16'(20);
			9301: out = 16'(423);
			9302: out = 16'(-32);
			9303: out = 16'(-344);
			9304: out = 16'(-9);
			9305: out = 16'(-1021);
			9306: out = 16'(103);
			9307: out = 16'(638);
			9308: out = 16'(-168);
			9309: out = 16'(690);
			9310: out = 16'(193);
			9311: out = 16'(-148);
			9312: out = 16'(438);
			9313: out = 16'(-154);
			9314: out = 16'(71);
			9315: out = 16'(-1216);
			9316: out = 16'(1231);
			9317: out = 16'(-133);
			9318: out = 16'(-678);
			9319: out = 16'(-49);
			9320: out = 16'(-493);
			9321: out = 16'(463);
			9322: out = 16'(-424);
			9323: out = 16'(728);
			9324: out = 16'(-312);
			9325: out = 16'(775);
			9326: out = 16'(-363);
			9327: out = 16'(-23);
			9328: out = 16'(29);
			9329: out = 16'(-117);
			9330: out = 16'(-35);
			9331: out = 16'(116);
			9332: out = 16'(136);
			9333: out = 16'(-172);
			9334: out = 16'(408);
			9335: out = 16'(-332);
			9336: out = 16'(553);
			9337: out = 16'(-156);
			9338: out = 16'(92);
			9339: out = 16'(-577);
			9340: out = 16'(122);
			9341: out = 16'(113);
			9342: out = 16'(-1027);
			9343: out = 16'(318);
			9344: out = 16'(-786);
			9345: out = 16'(-48);
			9346: out = 16'(718);
			9347: out = 16'(260);
			9348: out = 16'(-512);
			9349: out = 16'(217);
			9350: out = 16'(-427);
			9351: out = 16'(-142);
			9352: out = 16'(662);
			9353: out = 16'(-329);
			9354: out = 16'(-750);
			9355: out = 16'(586);
			9356: out = 16'(-1728);
			9357: out = 16'(251);
			9358: out = 16'(-333);
			9359: out = 16'(-50);
			9360: out = 16'(-123);
			9361: out = 16'(-781);
			9362: out = 16'(-516);
			9363: out = 16'(-992);
			9364: out = 16'(-15);
			9365: out = 16'(161);
			9366: out = 16'(100);
			9367: out = 16'(-50);
			9368: out = 16'(834);
			9369: out = 16'(53);
			9370: out = 16'(80);
			9371: out = 16'(155);
			9372: out = 16'(534);
			9373: out = 16'(616);
			9374: out = 16'(-350);
			9375: out = 16'(602);
			9376: out = 16'(-132);
			9377: out = 16'(-253);
			9378: out = 16'(-787);
			9379: out = 16'(-43);
			9380: out = 16'(674);
			9381: out = 16'(620);
			9382: out = 16'(-90);
			9383: out = 16'(99);
			9384: out = 16'(-449);
			9385: out = 16'(-267);
			9386: out = 16'(-179);
			9387: out = 16'(-934);
			9388: out = 16'(-79);
			9389: out = 16'(947);
			9390: out = 16'(-466);
			9391: out = 16'(393);
			9392: out = 16'(-388);
			9393: out = 16'(215);
			9394: out = 16'(-59);
			9395: out = 16'(105);
			9396: out = 16'(667);
			9397: out = 16'(94);
			9398: out = 16'(-335);
			9399: out = 16'(-502);
			9400: out = 16'(177);
			9401: out = 16'(22);
			9402: out = 16'(-829);
			9403: out = 16'(1331);
			9404: out = 16'(-221);
			9405: out = 16'(231);
			9406: out = 16'(-590);
			9407: out = 16'(47);
			9408: out = 16'(96);
			9409: out = 16'(417);
			9410: out = 16'(-52);
			9411: out = 16'(-575);
			9412: out = 16'(910);
			9413: out = 16'(-1110);
			9414: out = 16'(1021);
			9415: out = 16'(-944);
			9416: out = 16'(-69);
			9417: out = 16'(-288);
			9418: out = 16'(-389);
			9419: out = 16'(-1354);
			9420: out = 16'(-48);
			9421: out = 16'(122);
			9422: out = 16'(-655);
			9423: out = 16'(-197);
			9424: out = 16'(1222);
			9425: out = 16'(-717);
			9426: out = 16'(-381);
			9427: out = 16'(741);
			9428: out = 16'(769);
			9429: out = 16'(-448);
			9430: out = 16'(-99);
			9431: out = 16'(-164);
			9432: out = 16'(567);
			9433: out = 16'(429);
			9434: out = 16'(432);
			9435: out = 16'(50);
			9436: out = 16'(-106);
			9437: out = 16'(-376);
			9438: out = 16'(-786);
			9439: out = 16'(512);
			9440: out = 16'(-657);
			9441: out = 16'(490);
			9442: out = 16'(-210);
			9443: out = 16'(-127);
			9444: out = 16'(-705);
			9445: out = 16'(-15);
			9446: out = 16'(-406);
			9447: out = 16'(-100);
			9448: out = 16'(113);
			9449: out = 16'(-232);
			9450: out = 16'(-838);
			9451: out = 16'(1114);
			9452: out = 16'(488);
			9453: out = 16'(-1179);
			9454: out = 16'(409);
			9455: out = 16'(573);
			9456: out = 16'(52);
			9457: out = 16'(-609);
			9458: out = 16'(-195);
			9459: out = 16'(-540);
			9460: out = 16'(-101);
			9461: out = 16'(-560);
			9462: out = 16'(-257);
			9463: out = 16'(439);
			9464: out = 16'(-438);
			9465: out = 16'(-177);
			9466: out = 16'(499);
			9467: out = 16'(376);
			9468: out = 16'(-808);
			9469: out = 16'(3);
			9470: out = 16'(162);
			9471: out = 16'(91);
			9472: out = 16'(-604);
			9473: out = 16'(554);
			9474: out = 16'(-712);
			9475: out = 16'(317);
			9476: out = 16'(119);
			9477: out = 16'(-928);
			9478: out = 16'(-333);
			9479: out = 16'(875);
			9480: out = 16'(493);
			9481: out = 16'(-197);
			9482: out = 16'(652);
			9483: out = 16'(-110);
			9484: out = 16'(-443);
			9485: out = 16'(-358);
			9486: out = 16'(483);
			9487: out = 16'(-130);
			9488: out = 16'(163);
			9489: out = 16'(-347);
			9490: out = 16'(-740);
			9491: out = 16'(116);
			9492: out = 16'(-719);
			9493: out = 16'(-466);
			9494: out = 16'(241);
			9495: out = 16'(-71);
			9496: out = 16'(-792);
			9497: out = 16'(323);
			9498: out = 16'(417);
			9499: out = 16'(-196);
			9500: out = 16'(329);
			9501: out = 16'(-179);
			9502: out = 16'(437);
			9503: out = 16'(253);
			9504: out = 16'(-104);
			9505: out = 16'(2);
			9506: out = 16'(-60);
			9507: out = 16'(477);
			9508: out = 16'(-958);
			9509: out = 16'(-78);
			9510: out = 16'(-212);
			9511: out = 16'(286);
			9512: out = 16'(-265);
			9513: out = 16'(-101);
			9514: out = 16'(1232);
			9515: out = 16'(-542);
			9516: out = 16'(-782);
			9517: out = 16'(-522);
			9518: out = 16'(218);
			9519: out = 16'(348);
			9520: out = 16'(-1183);
			9521: out = 16'(-177);
			9522: out = 16'(-243);
			9523: out = 16'(178);
			9524: out = 16'(-1608);
			9525: out = 16'(-226);
			9526: out = 16'(138);
			9527: out = 16'(-154);
			9528: out = 16'(-440);
			9529: out = 16'(-972);
			9530: out = 16'(365);
			9531: out = 16'(-508);
			9532: out = 16'(738);
			9533: out = 16'(-812);
			9534: out = 16'(1121);
			9535: out = 16'(-264);
			9536: out = 16'(-36);
			9537: out = 16'(-157);
			9538: out = 16'(987);
			9539: out = 16'(-176);
			9540: out = 16'(-1134);
			9541: out = 16'(772);
			9542: out = 16'(-279);
			9543: out = 16'(548);
			9544: out = 16'(-57);
			9545: out = 16'(-830);
			9546: out = 16'(166);
			9547: out = 16'(-850);
			9548: out = 16'(-444);
			9549: out = 16'(-740);
			9550: out = 16'(1040);
			9551: out = 16'(-195);
			9552: out = 16'(-291);
			9553: out = 16'(-71);
			9554: out = 16'(-1016);
			9555: out = 16'(450);
			9556: out = 16'(-931);
			9557: out = 16'(1178);
			9558: out = 16'(-846);
			9559: out = 16'(1067);
			9560: out = 16'(-29);
			9561: out = 16'(-739);
			9562: out = 16'(151);
			9563: out = 16'(373);
			9564: out = 16'(-146);
			9565: out = 16'(-210);
			9566: out = 16'(1357);
			9567: out = 16'(-469);
			9568: out = 16'(278);
			9569: out = 16'(266);
			9570: out = 16'(-426);
			9571: out = 16'(659);
			9572: out = 16'(-805);
			9573: out = 16'(108);
			9574: out = 16'(-301);
			9575: out = 16'(-30);
			9576: out = 16'(-94);
			9577: out = 16'(-413);
			9578: out = 16'(121);
			9579: out = 16'(-1336);
			9580: out = 16'(-121);
			9581: out = 16'(-135);
			9582: out = 16'(318);
			9583: out = 16'(939);
			9584: out = 16'(-162);
			9585: out = 16'(36);
			9586: out = 16'(-170);
			9587: out = 16'(-219);
			9588: out = 16'(193);
			9589: out = 16'(-629);
			9590: out = 16'(-6);
			9591: out = 16'(430);
			9592: out = 16'(-1636);
			9593: out = 16'(87);
			9594: out = 16'(13);
			9595: out = 16'(142);
			9596: out = 16'(448);
			9597: out = 16'(465);
			9598: out = 16'(476);
			9599: out = 16'(-265);
			9600: out = 16'(-99);
			9601: out = 16'(72);
			9602: out = 16'(-222);
			9603: out = 16'(587);
			9604: out = 16'(-1418);
			9605: out = 16'(57);
			9606: out = 16'(-330);
			9607: out = 16'(398);
			9608: out = 16'(0);
			9609: out = 16'(245);
			9610: out = 16'(-146);
			9611: out = 16'(-368);
			9612: out = 16'(-169);
			9613: out = 16'(-699);
			9614: out = 16'(-136);
			9615: out = 16'(437);
			9616: out = 16'(404);
			9617: out = 16'(-764);
			9618: out = 16'(-143);
			9619: out = 16'(-518);
			9620: out = 16'(-128);
			9621: out = 16'(-282);
			9622: out = 16'(613);
			9623: out = 16'(-211);
			9624: out = 16'(285);
			9625: out = 16'(714);
			9626: out = 16'(-509);
			9627: out = 16'(-600);
			9628: out = 16'(41);
			9629: out = 16'(-102);
			9630: out = 16'(23);
			9631: out = 16'(-257);
			9632: out = 16'(518);
			9633: out = 16'(-962);
			9634: out = 16'(-43);
			9635: out = 16'(-267);
			9636: out = 16'(-273);
			9637: out = 16'(223);
			9638: out = 16'(-921);
			9639: out = 16'(409);
			9640: out = 16'(-5);
			9641: out = 16'(499);
			9642: out = 16'(-381);
			9643: out = 16'(261);
			9644: out = 16'(-439);
			9645: out = 16'(166);
			9646: out = 16'(449);
			9647: out = 16'(-432);
			9648: out = 16'(9);
			9649: out = 16'(-811);
			9650: out = 16'(85);
			9651: out = 16'(-1014);
			9652: out = 16'(397);
			9653: out = 16'(202);
			9654: out = 16'(-290);
			9655: out = 16'(88);
			9656: out = 16'(-398);
			9657: out = 16'(96);
			9658: out = 16'(-168);
			9659: out = 16'(-52);
			9660: out = 16'(314);
			9661: out = 16'(312);
			9662: out = 16'(-200);
			9663: out = 16'(-628);
			9664: out = 16'(680);
			9665: out = 16'(-680);
			9666: out = 16'(282);
			9667: out = 16'(-125);
			9668: out = 16'(579);
			9669: out = 16'(140);
			9670: out = 16'(-248);
			9671: out = 16'(105);
			9672: out = 16'(-1158);
			9673: out = 16'(-162);
			9674: out = 16'(517);
			9675: out = 16'(21);
			9676: out = 16'(228);
			9677: out = 16'(433);
			9678: out = 16'(-337);
			9679: out = 16'(-296);
			9680: out = 16'(403);
			9681: out = 16'(-509);
			9682: out = 16'(469);
			9683: out = 16'(-482);
			9684: out = 16'(670);
			9685: out = 16'(-466);
			9686: out = 16'(-46);
			9687: out = 16'(140);
			9688: out = 16'(-778);
			9689: out = 16'(-293);
			9690: out = 16'(-825);
			9691: out = 16'(-200);
			9692: out = 16'(59);
			9693: out = 16'(79);
			9694: out = 16'(86);
			9695: out = 16'(106);
			9696: out = 16'(-243);
			9697: out = 16'(-779);
			9698: out = 16'(493);
			9699: out = 16'(658);
			9700: out = 16'(320);
			9701: out = 16'(-327);
			9702: out = 16'(105);
			9703: out = 16'(-58);
			9704: out = 16'(1);
			9705: out = 16'(376);
			9706: out = 16'(96);
			9707: out = 16'(195);
			9708: out = 16'(-478);
			9709: out = 16'(-42);
			9710: out = 16'(446);
			9711: out = 16'(440);
			9712: out = 16'(-289);
			9713: out = 16'(241);
			9714: out = 16'(-141);
			9715: out = 16'(-54);
			9716: out = 16'(522);
			9717: out = 16'(-783);
			9718: out = 16'(376);
			9719: out = 16'(482);
			9720: out = 16'(-220);
			9721: out = 16'(-35);
			9722: out = 16'(-757);
			9723: out = 16'(644);
			9724: out = 16'(-997);
			9725: out = 16'(762);
			9726: out = 16'(320);
			9727: out = 16'(153);
			9728: out = 16'(-116);
			9729: out = 16'(-572);
			9730: out = 16'(224);
			9731: out = 16'(-151);
			9732: out = 16'(220);
			9733: out = 16'(30);
			9734: out = 16'(536);
			9735: out = 16'(-410);
			9736: out = 16'(-143);
			9737: out = 16'(-16);
			9738: out = 16'(738);
			9739: out = 16'(442);
			9740: out = 16'(-102);
			9741: out = 16'(-311);
			9742: out = 16'(379);
			9743: out = 16'(-27);
			9744: out = 16'(-63);
			9745: out = 16'(-285);
			9746: out = 16'(76);
			9747: out = 16'(686);
			9748: out = 16'(-473);
			9749: out = 16'(-13);
			9750: out = 16'(-11);
			9751: out = 16'(109);
			9752: out = 16'(-154);
			9753: out = 16'(251);
			9754: out = 16'(301);
			9755: out = 16'(-120);
			9756: out = 16'(-682);
			9757: out = 16'(240);
			9758: out = 16'(384);
			9759: out = 16'(-75);
			9760: out = 16'(-186);
			9761: out = 16'(417);
			9762: out = 16'(609);
			9763: out = 16'(293);
			9764: out = 16'(269);
			9765: out = 16'(-1);
			9766: out = 16'(192);
			9767: out = 16'(-222);
			9768: out = 16'(-96);
			9769: out = 16'(-277);
			9770: out = 16'(293);
			9771: out = 16'(-231);
			9772: out = 16'(240);
			9773: out = 16'(-51);
			9774: out = 16'(80);
			9775: out = 16'(29);
			9776: out = 16'(-227);
			9777: out = 16'(509);
			9778: out = 16'(402);
			9779: out = 16'(-79);
			9780: out = 16'(-182);
			9781: out = 16'(-260);
			9782: out = 16'(-207);
			9783: out = 16'(389);
			9784: out = 16'(-636);
			9785: out = 16'(-179);
			9786: out = 16'(707);
			9787: out = 16'(-559);
			9788: out = 16'(202);
			9789: out = 16'(-180);
			9790: out = 16'(-46);
			9791: out = 16'(65);
			9792: out = 16'(255);
			9793: out = 16'(-82);
			9794: out = 16'(-71);
			9795: out = 16'(344);
			9796: out = 16'(84);
			9797: out = 16'(13);
			9798: out = 16'(1);
			9799: out = 16'(120);
			9800: out = 16'(-190);
			9801: out = 16'(-464);
			9802: out = 16'(738);
			9803: out = 16'(-741);
			9804: out = 16'(-153);
			9805: out = 16'(-109);
			9806: out = 16'(-597);
			9807: out = 16'(137);
			9808: out = 16'(-953);
			9809: out = 16'(726);
			9810: out = 16'(327);
			9811: out = 16'(16);
			9812: out = 16'(-950);
			9813: out = 16'(-209);
			9814: out = 16'(403);
			9815: out = 16'(-879);
			9816: out = 16'(590);
			9817: out = 16'(-146);
			9818: out = 16'(-36);
			9819: out = 16'(33);
			9820: out = 16'(313);
			9821: out = 16'(-192);
			9822: out = 16'(102);
			9823: out = 16'(-222);
			9824: out = 16'(-357);
			9825: out = 16'(334);
			9826: out = 16'(-2);
			9827: out = 16'(242);
			9828: out = 16'(44);
			9829: out = 16'(388);
			9830: out = 16'(-75);
			9831: out = 16'(-352);
			9832: out = 16'(-73);
			9833: out = 16'(434);
			9834: out = 16'(-492);
			9835: out = 16'(430);
			9836: out = 16'(-549);
			9837: out = 16'(-318);
			9838: out = 16'(837);
			9839: out = 16'(-1121);
			9840: out = 16'(-119);
			9841: out = 16'(561);
			9842: out = 16'(16);
			9843: out = 16'(-242);
			9844: out = 16'(221);
			9845: out = 16'(-218);
			9846: out = 16'(-417);
			9847: out = 16'(-169);
			9848: out = 16'(161);
			9849: out = 16'(401);
			9850: out = 16'(-251);
			9851: out = 16'(216);
			9852: out = 16'(-358);
			9853: out = 16'(-18);
			9854: out = 16'(390);
			9855: out = 16'(-763);
			9856: out = 16'(726);
			9857: out = 16'(229);
			9858: out = 16'(-1001);
			9859: out = 16'(133);
			9860: out = 16'(-13);
			9861: out = 16'(169);
			9862: out = 16'(-19);
			9863: out = 16'(-228);
			9864: out = 16'(-939);
			9865: out = 16'(50);
			9866: out = 16'(-203);
			9867: out = 16'(-217);
			9868: out = 16'(-663);
			9869: out = 16'(529);
			9870: out = 16'(-266);
			9871: out = 16'(-472);
			9872: out = 16'(951);
			9873: out = 16'(-111);
			9874: out = 16'(-122);
			9875: out = 16'(70);
			9876: out = 16'(2);
			9877: out = 16'(585);
			9878: out = 16'(-195);
			9879: out = 16'(71);
			9880: out = 16'(-166);
			9881: out = 16'(314);
			9882: out = 16'(-195);
			9883: out = 16'(-269);
			9884: out = 16'(85);
			9885: out = 16'(373);
			9886: out = 16'(-97);
			9887: out = 16'(108);
			9888: out = 16'(79);
			9889: out = 16'(-777);
			9890: out = 16'(220);
			9891: out = 16'(-316);
			9892: out = 16'(-645);
			9893: out = 16'(150);
			9894: out = 16'(-422);
			9895: out = 16'(134);
			9896: out = 16'(-193);
			9897: out = 16'(-49);
			9898: out = 16'(39);
			9899: out = 16'(-441);
			9900: out = 16'(309);
			9901: out = 16'(221);
			9902: out = 16'(-87);
			9903: out = 16'(-185);
			9904: out = 16'(58);
			9905: out = 16'(-193);
			9906: out = 16'(267);
			9907: out = 16'(-405);
			9908: out = 16'(58);
			9909: out = 16'(520);
			9910: out = 16'(-296);
			9911: out = 16'(313);
			9912: out = 16'(-164);
			9913: out = 16'(156);
			9914: out = 16'(-129);
			9915: out = 16'(-73);
			9916: out = 16'(-32);
			9917: out = 16'(-198);
			9918: out = 16'(216);
			9919: out = 16'(44);
			9920: out = 16'(71);
			9921: out = 16'(-77);
			9922: out = 16'(-12);
			9923: out = 16'(-462);
			9924: out = 16'(-9);
			9925: out = 16'(-80);
			9926: out = 16'(23);
			9927: out = 16'(-124);
			9928: out = 16'(285);
			9929: out = 16'(51);
			9930: out = 16'(-59);
			9931: out = 16'(32);
			9932: out = 16'(-68);
			9933: out = 16'(44);
			9934: out = 16'(-37);
			9935: out = 16'(-334);
			9936: out = 16'(100);
			9937: out = 16'(-74);
			9938: out = 16'(6);
			9939: out = 16'(-204);
			9940: out = 16'(356);
			9941: out = 16'(-400);
			9942: out = 16'(17);
			9943: out = 16'(164);
			9944: out = 16'(-329);
			9945: out = 16'(309);
			9946: out = 16'(-402);
			9947: out = 16'(-88);
			default: out = 0;
		endcase
	end
endmodule
