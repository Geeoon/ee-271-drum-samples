module crash1_lookup(index, out);
	input logic unsigned [15:0] index;
	output logic signed [23:0] out;
	always_comb begin
		case(index)
			0: out = 24'(0);
			1: out = 24'(0);
			2: out = 24'(20);
			3: out = 24'(-340);
			4: out = 24'(8);
			5: out = 24'(-324);
			6: out = 24'(104);
			7: out = 24'(-464);
			8: out = 24'(204);
			9: out = 24'(-620);
			10: out = 24'(432);
			11: out = 24'(-856);
			12: out = 24'(884);
			13: out = 24'(-1420);
			14: out = 24'(-96);
			15: out = 24'(-1576);
			16: out = 24'(29572);
			17: out = 24'(15956);
			18: out = 24'(-8112);
			19: out = 24'(15976);
			20: out = 24'(-31788);
			21: out = 24'(-30000);
			22: out = 24'(-3728);
			23: out = 24'(9280);
			24: out = 24'(-70688);
			25: out = 24'(-65564);
			26: out = 24'(20524);
			27: out = 24'(77024);
			28: out = 24'(4632);
			29: out = 24'(-46852);
			30: out = 24'(-46820);
			31: out = 24'(-8832);
			32: out = 24'(-14244);
			33: out = 24'(-11612);
			34: out = 24'(-8972);
			35: out = 24'(2124);
			36: out = 24'(17348);
			37: out = 24'(2216);
			38: out = 24'(-21480);
			39: out = 24'(-27000);
			40: out = 24'(23056);
			41: out = 24'(-3964);
			42: out = 24'(13220);
			43: out = 24'(4892);
			44: out = 24'(-25720);
			45: out = 24'(-39388);
			46: out = 24'(33832);
			47: out = 24'(58624);
			48: out = 24'(4008);
			49: out = 24'(19672);
			50: out = 24'(4552);
			51: out = 24'(-32368);
			52: out = 24'(-71536);
			53: out = 24'(1304);
			54: out = 24'(43224);
			55: out = 24'(51400);
			56: out = 24'(16892);
			57: out = 24'(-10140);
			58: out = 24'(-34652);
			59: out = 24'(-21328);
			60: out = 24'(5112);
			61: out = 24'(14788);
			62: out = 24'(-3868);
			63: out = 24'(-31252);
			64: out = 24'(-13888);
			65: out = 24'(38340);
			66: out = 24'(9684);
			67: out = 24'(-45872);
			68: out = 24'(-61460);
			69: out = 24'(9000);
			70: out = 24'(-18160);
			71: out = 24'(30652);
			72: out = 24'(28952);
			73: out = 24'(4888);
			74: out = 24'(-50628);
			75: out = 24'(13864);
			76: out = 24'(18344);
			77: out = 24'(-16544);
			78: out = 24'(-8000);
			79: out = 24'(44672);
			80: out = 24'(32640);
			81: out = 24'(-21520);
			82: out = 24'(-29172);
			83: out = 24'(-20276);
			84: out = 24'(10284);
			85: out = 24'(17952);
			86: out = 24'(8840);
			87: out = 24'(-21580);
			88: out = 24'(-17028);
			89: out = 24'(19580);
			90: out = 24'(49664);
			91: out = 24'(19628);
			92: out = 24'(6984);
			93: out = 24'(-216);
			94: out = 24'(-7628);
			95: out = 24'(-1432);
			96: out = 24'(-8628);
			97: out = 24'(26916);
			98: out = 24'(50436);
			99: out = 24'(7260);
			100: out = 24'(-4208);
			101: out = 24'(25476);
			102: out = 24'(47400);
			103: out = 24'(-16776);
			104: out = 24'(4492);
			105: out = 24'(-16156);
			106: out = 24'(-2588);
			107: out = 24'(11856);
			108: out = 24'(20380);
			109: out = 24'(-35624);
			110: out = 24'(-36132);
			111: out = 24'(11764);
			112: out = 24'(-7868);
			113: out = 24'(-31084);
			114: out = 24'(-17288);
			115: out = 24'(15892);
			116: out = 24'(-31980);
			117: out = 24'(-17056);
			118: out = 24'(2328);
			119: out = 24'(3592);
			120: out = 24'(-79544);
			121: out = 24'(5800);
			122: out = 24'(8624);
			123: out = 24'(-7116);
			124: out = 24'(-3096);
			125: out = 24'(17672);
			126: out = 24'(-9228);
			127: out = 24'(-24736);
			128: out = 24'(4008);
			129: out = 24'(14724);
			130: out = 24'(7696);
			131: out = 24'(-7888);
			132: out = 24'(1312);
			133: out = 24'(-6540);
			134: out = 24'(27492);
			135: out = 24'(16552);
			136: out = 24'(-10988);
			137: out = 24'(-35272);
			138: out = 24'(10028);
			139: out = 24'(-5616);
			140: out = 24'(-34988);
			141: out = 24'(4620);
			142: out = 24'(11496);
			143: out = 24'(32328);
			144: out = 24'(20096);
			145: out = 24'(-5360);
			146: out = 24'(-26568);
			147: out = 24'(-11496);
			148: out = 24'(-8528);
			149: out = 24'(-27688);
			150: out = 24'(-1096);
			151: out = 24'(-3472);
			152: out = 24'(-372);
			153: out = 24'(2460);
			154: out = 24'(41484);
			155: out = 24'(-13568);
			156: out = 24'(-19556);
			157: out = 24'(2056);
			158: out = 24'(12496);
			159: out = 24'(-2564);
			160: out = 24'(9296);
			161: out = 24'(20116);
			162: out = 24'(18940);
			163: out = 24'(-4868);
			164: out = 24'(13520);
			165: out = 24'(-9684);
			166: out = 24'(-80020);
			167: out = 24'(-59976);
			168: out = 24'(-25892);
			169: out = 24'(-11024);
			170: out = 24'(-24956);
			171: out = 24'(-8312);
			172: out = 24'(-60);
			173: out = 24'(-9548);
			174: out = 24'(-16640);
			175: out = 24'(23916);
			176: out = 24'(40276);
			177: out = 24'(18724);
			178: out = 24'(-13820);
			179: out = 24'(1236);
			180: out = 24'(-16404);
			181: out = 24'(-12932);
			182: out = 24'(6176);
			183: out = 24'(44860);
			184: out = 24'(21136);
			185: out = 24'(9008);
			186: out = 24'(-9192);
			187: out = 24'(-12356);
			188: out = 24'(-72944);
			189: out = 24'(-11484);
			190: out = 24'(16396);
			191: out = 24'(-1164);
			192: out = 24'(18712);
			193: out = 24'(47560);
			194: out = 24'(71040);
			195: out = 24'(62072);
			196: out = 24'(37960);
			197: out = 24'(-2968);
			198: out = 24'(-16104);
			199: out = 24'(-7404);
			200: out = 24'(7296);
			201: out = 24'(76408);
			202: out = 24'(58392);
			203: out = 24'(-9472);
			204: out = 24'(-76092);
			205: out = 24'(-19332);
			206: out = 24'(-20604);
			207: out = 24'(-33148);
			208: out = 24'(-28512);
			209: out = 24'(17416);
			210: out = 24'(-17620);
			211: out = 24'(-36996);
			212: out = 24'(-14784);
			213: out = 24'(17936);
			214: out = 24'(-1500);
			215: out = 24'(-10420);
			216: out = 24'(15252);
			217: out = 24'(57040);
			218: out = 24'(7672);
			219: out = 24'(15764);
			220: out = 24'(49860);
			221: out = 24'(43616);
			222: out = 24'(37720);
			223: out = 24'(-2288);
			224: out = 24'(1108);
			225: out = 24'(38144);
			226: out = 24'(15008);
			227: out = 24'(-12760);
			228: out = 24'(-47768);
			229: out = 24'(-59748);
			230: out = 24'(-54652);
			231: out = 24'(-39436);
			232: out = 24'(-24756);
			233: out = 24'(-14924);
			234: out = 24'(-59380);
			235: out = 24'(3048);
			236: out = 24'(3808);
			237: out = 24'(-8836);
			238: out = 24'(3280);
			239: out = 24'(68412);
			240: out = 24'(46440);
			241: out = 24'(6560);
			242: out = 24'(-2168);
			243: out = 24'(-1712);
			244: out = 24'(-6704);
			245: out = 24'(26960);
			246: out = 24'(72404);
			247: out = 24'(18380);
			248: out = 24'(-20524);
			249: out = 24'(-39088);
			250: out = 24'(-21744);
			251: out = 24'(-1000);
			252: out = 24'(-72524);
			253: out = 24'(-104400);
			254: out = 24'(-42224);
			255: out = 24'(35880);
			256: out = 24'(-5684);
			257: out = 24'(-49372);
			258: out = 24'(-37668);
			259: out = 24'(7036);
			260: out = 24'(-36884);
			261: out = 24'(-51168);
			262: out = 24'(-31216);
			263: out = 24'(-3876);
			264: out = 24'(-5244);
			265: out = 24'(2512);
			266: out = 24'(-5500);
			267: out = 24'(-27500);
			268: out = 24'(6648);
			269: out = 24'(2936);
			270: out = 24'(7516);
			271: out = 24'(7280);
			272: out = 24'(42656);
			273: out = 24'(-35876);
			274: out = 24'(-12448);
			275: out = 24'(58840);
			276: out = 24'(71720);
			277: out = 24'(64948);
			278: out = 24'(78560);
			279: out = 24'(92940);
			280: out = 24'(58344);
			281: out = 24'(8120);
			282: out = 24'(-5088);
			283: out = 24'(43632);
			284: out = 24'(77828);
			285: out = 24'(14132);
			286: out = 24'(30960);
			287: out = 24'(55084);
			288: out = 24'(28420);
			289: out = 24'(-24780);
			290: out = 24'(-76272);
			291: out = 24'(-51212);
			292: out = 24'(-23528);
			293: out = 24'(-87944);
			294: out = 24'(-88052);
			295: out = 24'(-60500);
			296: out = 24'(-26176);
			297: out = 24'(-26360);
			298: out = 24'(-15924);
			299: out = 24'(-23544);
			300: out = 24'(-43616);
			301: out = 24'(-71680);
			302: out = 24'(-62596);
			303: out = 24'(-39968);
			304: out = 24'(-23560);
			305: out = 24'(-27948);
			306: out = 24'(-24176);
			307: out = 24'(5928);
			308: out = 24'(28316);
			309: out = 24'(13808);
			310: out = 24'(10692);
			311: out = 24'(-35328);
			312: out = 24'(-13708);
			313: out = 24'(33696);
			314: out = 24'(45736);
			315: out = 24'(43052);
			316: out = 24'(31496);
			317: out = 24'(28880);
			318: out = 24'(50896);
			319: out = 24'(66856);
			320: out = 24'(104860);
			321: out = 24'(94072);
			322: out = 24'(57096);
			323: out = 24'(82732);
			324: out = 24'(93240);
			325: out = 24'(52120);
			326: out = 24'(-9112);
			327: out = 24'(55372);
			328: out = 24'(55992);
			329: out = 24'(58020);
			330: out = 24'(34828);
			331: out = 24'(45660);
			332: out = 24'(-33728);
			333: out = 24'(-26352);
			334: out = 24'(-16216);
			335: out = 24'(-60468);
			336: out = 24'(-48280);
			337: out = 24'(-19220);
			338: out = 24'(-27424);
			339: out = 24'(-82000);
			340: out = 24'(-44148);
			341: out = 24'(-11548);
			342: out = 24'(1040);
			343: out = 24'(-30176);
			344: out = 24'(-107012);
			345: out = 24'(-115820);
			346: out = 24'(-91020);
			347: out = 24'(-62368);
			348: out = 24'(-131068);
			349: out = 24'(-32040);
			350: out = 24'(-10004);
			351: out = 24'(-53232);
			352: out = 24'(-72564);
			353: out = 24'(32080);
			354: out = 24'(-7712);
			355: out = 24'(-92312);
			356: out = 24'(-84508);
			357: out = 24'(-46576);
			358: out = 24'(-65240);
			359: out = 24'(-67312);
			360: out = 24'(13144);
			361: out = 24'(-13504);
			362: out = 24'(2056);
			363: out = 24'(940);
			364: out = 24'(-13880);
			365: out = 24'(-5996);
			366: out = 24'(-68036);
			367: out = 24'(-57260);
			368: out = 24'(3196);
			369: out = 24'(16900);
			370: out = 24'(12564);
			371: out = 24'(68720);
			372: out = 24'(100372);
			373: out = 24'(26460);
			374: out = 24'(-22652);
			375: out = 24'(1636);
			376: out = 24'(47156);
			377: out = 24'(11384);
			378: out = 24'(56672);
			379: out = 24'(43640);
			380: out = 24'(54132);
			381: out = 24'(65876);
			382: out = 24'(102624);
			383: out = 24'(69108);
			384: out = 24'(58824);
			385: out = 24'(59916);
			386: out = 24'(36948);
			387: out = 24'(24948);
			388: out = 24'(43840);
			389: out = 24'(80708);
			390: out = 24'(70836);
			391: out = 24'(101860);
			392: out = 24'(58044);
			393: out = 24'(25732);
			394: out = 24'(37084);
			395: out = 24'(62068);
			396: out = 24'(33016);
			397: out = 24'(12556);
			398: out = 24'(37416);
			399: out = 24'(45684);
			400: out = 24'(50124);
			401: out = 24'(50328);
			402: out = 24'(65576);
			403: out = 24'(90964);
			404: out = 24'(44864);
			405: out = 24'(13040);
			406: out = 24'(32164);
			407: out = 24'(73196);
			408: out = 24'(60036);
			409: out = 24'(23352);
			410: out = 24'(-3524);
			411: out = 24'(3260);
			412: out = 24'(15908);
			413: out = 24'(9528);
			414: out = 24'(-23292);
			415: out = 24'(-43048);
			416: out = 24'(-56884);
			417: out = 24'(-23436);
			418: out = 24'(-32012);
			419: out = 24'(-78660);
			420: out = 24'(-90180);
			421: out = 24'(-39016);
			422: out = 24'(-34848);
			423: out = 24'(-97644);
			424: out = 24'(-78472);
			425: out = 24'(-96492);
			426: out = 24'(-75264);
			427: out = 24'(-68792);
			428: out = 24'(-85656);
			429: out = 24'(-102620);
			430: out = 24'(-109720);
			431: out = 24'(-118764);
			432: out = 24'(-110772);
			433: out = 24'(-114008);
			434: out = 24'(-76688);
			435: out = 24'(-77168);
			436: out = 24'(-97704);
			437: out = 24'(-117916);
			438: out = 24'(-49228);
			439: out = 24'(-20284);
			440: out = 24'(-46588);
			441: out = 24'(-92140);
			442: out = 24'(-28572);
			443: out = 24'(-30900);
			444: out = 24'(-80056);
			445: out = 24'(-26576);
			446: out = 24'(12436);
			447: out = 24'(2152);
			448: out = 24'(-38104);
			449: out = 24'(-59312);
			450: out = 24'(-14864);
			451: out = 24'(-45848);
			452: out = 24'(-58396);
			453: out = 24'(21384);
			454: out = 24'(23768);
			455: out = 24'(-13072);
			456: out = 24'(12360);
			457: out = 24'(125360);
			458: out = 24'(91888);
			459: out = 24'(70952);
			460: out = 24'(26996);
			461: out = 24'(17032);
			462: out = 24'(-15232);
			463: out = 24'(56788);
			464: out = 24'(98512);
			465: out = 24'(108064);
			466: out = 24'(89460);
			467: out = 24'(111560);
			468: out = 24'(96896);
			469: out = 24'(63792);
			470: out = 24'(29928);
			471: out = 24'(71128);
			472: out = 24'(69304);
			473: out = 24'(36132);
			474: out = 24'(-8896);
			475: out = 24'(4800);
			476: out = 24'(-884);
			477: out = 24'(26180);
			478: out = 24'(61748);
			479: out = 24'(29464);
			480: out = 24'(-10828);
			481: out = 24'(-44768);
			482: out = 24'(-36828);
			483: out = 24'(-80);
			484: out = 24'(15976);
			485: out = 24'(18200);
			486: out = 24'(42764);
			487: out = 24'(104052);
			488: out = 24'(59724);
			489: out = 24'(43588);
			490: out = 24'(37632);
			491: out = 24'(35516);
			492: out = 24'(-20372);
			493: out = 24'(-21144);
			494: out = 24'(-8320);
			495: out = 24'(3712);
			496: out = 24'(50144);
			497: out = 24'(68616);
			498: out = 24'(40772);
			499: out = 24'(-5288);
			500: out = 24'(548);
			501: out = 24'(-10692);
			502: out = 24'(-23604);
			503: out = 24'(-22968);
			504: out = 24'(8768);
			505: out = 24'(16776);
			506: out = 24'(7268);
			507: out = 24'(13380);
			508: out = 24'(53192);
			509: out = 24'(21848);
			510: out = 24'(-11824);
			511: out = 24'(-42104);
			512: out = 24'(-63084);
			513: out = 24'(-53024);
			514: out = 24'(-47464);
			515: out = 24'(-3032);
			516: out = 24'(50896);
			517: out = 24'(19916);
			518: out = 24'(-5476);
			519: out = 24'(-1692);
			520: out = 24'(5348);
			521: out = 24'(-98308);
			522: out = 24'(-75740);
			523: out = 24'(-31748);
			524: out = 24'(-7972);
			525: out = 24'(-8600);
			526: out = 24'(-28200);
			527: out = 24'(-20356);
			528: out = 24'(-5688);
			529: out = 24'(-7972);
			530: out = 24'(-21352);
			531: out = 24'(-11340);
			532: out = 24'(-25320);
			533: out = 24'(-80240);
			534: out = 24'(-54724);
			535: out = 24'(-20332);
			536: out = 24'(-6348);
			537: out = 24'(-24476);
			538: out = 24'(27712);
			539: out = 24'(13244);
			540: out = 24'(-16020);
			541: out = 24'(-50016);
			542: out = 24'(10348);
			543: out = 24'(-72648);
			544: out = 24'(-55640);
			545: out = 24'(26368);
			546: out = 24'(35192);
			547: out = 24'(-584);
			548: out = 24'(-26460);
			549: out = 24'(-3924);
			550: out = 24'(10288);
			551: out = 24'(31852);
			552: out = 24'(19724);
			553: out = 24'(32800);
			554: out = 24'(49888);
			555: out = 24'(95500);
			556: out = 24'(43488);
			557: out = 24'(27248);
			558: out = 24'(31480);
			559: out = 24'(3828);
			560: out = 24'(-63416);
			561: out = 24'(-40652);
			562: out = 24'(36592);
			563: out = 24'(17880);
			564: out = 24'(10684);
			565: out = 24'(-1876);
			566: out = 24'(-2456);
			567: out = 24'(-22940);
			568: out = 24'(-592);
			569: out = 24'(26140);
			570: out = 24'(52412);
			571: out = 24'(50120);
			572: out = 24'(20036);
			573: out = 24'(16220);
			574: out = 24'(19112);
			575: out = 24'(-208);
			576: out = 24'(-20796);
			577: out = 24'(-18636);
			578: out = 24'(1344);
			579: out = 24'(4508);
			580: out = 24'(2692);
			581: out = 24'(23604);
			582: out = 24'(43604);
			583: out = 24'(31672);
			584: out = 24'(22772);
			585: out = 24'(-3944);
			586: out = 24'(13612);
			587: out = 24'(3088);
			588: out = 24'(-30212);
			589: out = 24'(416);
			590: out = 24'(66344);
			591: out = 24'(66308);
			592: out = 24'(10296);
			593: out = 24'(-12824);
			594: out = 24'(22604);
			595: out = 24'(13132);
			596: out = 24'(-47000);
			597: out = 24'(-49500);
			598: out = 24'(25220);
			599: out = 24'(59500);
			600: out = 24'(20452);
			601: out = 24'(416);
			602: out = 24'(6448);
			603: out = 24'(36036);
			604: out = 24'(49984);
			605: out = 24'(48148);
			606: out = 24'(-3876);
			607: out = 24'(-58476);
			608: out = 24'(-67484);
			609: out = 24'(-10936);
			610: out = 24'(-38480);
			611: out = 24'(-22676);
			612: out = 24'(1084);
			613: out = 24'(21724);
			614: out = 24'(-35832);
			615: out = 24'(-11676);
			616: out = 24'(-14488);
			617: out = 24'(-35916);
			618: out = 24'(-10140);
			619: out = 24'(-6296);
			620: out = 24'(308);
			621: out = 24'(-16928);
			622: out = 24'(-56340);
			623: out = 24'(-41112);
			624: out = 24'(-11932);
			625: out = 24'(-9480);
			626: out = 24'(-54876);
			627: out = 24'(-88776);
			628: out = 24'(-105212);
			629: out = 24'(-77820);
			630: out = 24'(-41364);
			631: out = 24'(-24812);
			632: out = 24'(-37632);
			633: out = 24'(-23592);
			634: out = 24'(23424);
			635: out = 24'(77528);
			636: out = 24'(27628);
			637: out = 24'(11352);
			638: out = 24'(45552);
			639: out = 24'(40420);
			640: out = 24'(48072);
			641: out = 24'(3564);
			642: out = 24'(-12496);
			643: out = 24'(31212);
			644: out = 24'(88288);
			645: out = 24'(70244);
			646: out = 24'(21224);
			647: out = 24'(4112);
			648: out = 24'(16180);
			649: out = 24'(48204);
			650: out = 24'(64256);
			651: out = 24'(68576);
			652: out = 24'(54048);
			653: out = 24'(45604);
			654: out = 24'(2304);
			655: out = 24'(-28572);
			656: out = 24'(55060);
			657: out = 24'(-16140);
			658: out = 24'(-55748);
			659: out = 24'(-52152);
			660: out = 24'(-13632);
			661: out = 24'(-51232);
			662: out = 24'(-39540);
			663: out = 24'(19116);
			664: out = 24'(73032);
			665: out = 24'(4908);
			666: out = 24'(-4420);
			667: out = 24'(-16616);
			668: out = 24'(-55648);
			669: out = 24'(-48668);
			670: out = 24'(-41820);
			671: out = 24'(-21648);
			672: out = 24'(-8044);
			673: out = 24'(296);
			674: out = 24'(-22904);
			675: out = 24'(-34488);
			676: out = 24'(-31912);
			677: out = 24'(-51828);
			678: out = 24'(-104396);
			679: out = 24'(-110632);
			680: out = 24'(-52616);
			681: out = 24'(-11648);
			682: out = 24'(42568);
			683: out = 24'(3076);
			684: out = 24'(-22004);
			685: out = 24'(-576);
			686: out = 24'(1724);
			687: out = 24'(-42580);
			688: out = 24'(-46980);
			689: out = 24'(4532);
			690: out = 24'(-22860);
			691: out = 24'(-26808);
			692: out = 24'(-23812);
			693: out = 24'(-11864);
			694: out = 24'(-12284);
			695: out = 24'(-20280);
			696: out = 24'(1688);
			697: out = 24'(33860);
			698: out = 24'(44344);
			699: out = 24'(15720);
			700: out = 24'(30056);
			701: out = 24'(57880);
			702: out = 24'(56888);
			703: out = 24'(13948);
			704: out = 24'(27512);
			705: out = 24'(66720);
			706: out = 24'(90380);
			707: out = 24'(43972);
			708: out = 24'(86508);
			709: out = 24'(88516);
			710: out = 24'(55088);
			711: out = 24'(73712);
			712: out = 24'(58452);
			713: out = 24'(8124);
			714: out = 24'(-26736);
			715: out = 24'(57352);
			716: out = 24'(52260);
			717: out = 24'(35672);
			718: out = 24'(4900);
			719: out = 24'(3588);
			720: out = 24'(24188);
			721: out = 24'(50216);
			722: out = 24'(21356);
			723: out = 24'(-57360);
			724: out = 24'(8980);
			725: out = 24'(23292);
			726: out = 24'(49336);
			727: out = 24'(65772);
			728: out = 24'(79908);
			729: out = 24'(-28048);
			730: out = 24'(-84292);
			731: out = 24'(-57188);
			732: out = 24'(-44532);
			733: out = 24'(-51020);
			734: out = 24'(-40296);
			735: out = 24'(-10652);
			736: out = 24'(-16996);
			737: out = 24'(-7344);
			738: out = 24'(15904);
			739: out = 24'(30616);
			740: out = 24'(-14288);
			741: out = 24'(-28060);
			742: out = 24'(-88208);
			743: out = 24'(-119432);
			744: out = 24'(-102868);
			745: out = 24'(9964);
			746: out = 24'(65668);
			747: out = 24'(44528);
			748: out = 24'(-8624);
			749: out = 24'(-264);
			750: out = 24'(-70376);
			751: out = 24'(-117600);
			752: out = 24'(-111732);
			753: out = 24'(-98924);
			754: out = 24'(-39156);
			755: out = 24'(-23788);
			756: out = 24'(-9992);
			757: out = 24'(43100);
			758: out = 24'(24928);
			759: out = 24'(-14548);
			760: out = 24'(-65928);
			761: out = 24'(-73932);
			762: out = 24'(-35752);
			763: out = 24'(21292);
			764: out = 24'(36436);
			765: out = 24'(31200);
			766: out = 24'(33144);
			767: out = 24'(43832);
			768: out = 24'(14768);
			769: out = 24'(-33036);
			770: out = 24'(-46424);
			771: out = 24'(-15456);
			772: out = 24'(6888);
			773: out = 24'(8204);
			774: out = 24'(15136);
			775: out = 24'(51248);
			776: out = 24'(56652);
			777: out = 24'(36704);
			778: out = 24'(19252);
			779: out = 24'(24024);
			780: out = 24'(24944);
			781: out = 24'(20716);
			782: out = 24'(3920);
			783: out = 24'(-1568);
			784: out = 24'(-35284);
			785: out = 24'(-28564);
			786: out = 24'(6280);
			787: out = 24'(-4272);
			788: out = 24'(-7892);
			789: out = 24'(25168);
			790: out = 24'(67560);
			791: out = 24'(51212);
			792: out = 24'(15536);
			793: out = 24'(-4236);
			794: out = 24'(4252);
			795: out = 24'(592);
			796: out = 24'(30544);
			797: out = 24'(58572);
			798: out = 24'(79504);
			799: out = 24'(60904);
			800: out = 24'(39208);
			801: out = 24'(4276);
			802: out = 24'(-3440);
			803: out = 24'(-5128);
			804: out = 24'(19976);
			805: out = 24'(-47076);
			806: out = 24'(-61176);
			807: out = 24'(10948);
			808: out = 24'(66176);
			809: out = 24'(22076);
			810: out = 24'(-39832);
			811: out = 24'(-46796);
			812: out = 24'(-5144);
			813: out = 24'(-5844);
			814: out = 24'(-22900);
			815: out = 24'(-13296);
			816: out = 24'(17148);
			817: out = 24'(-15772);
			818: out = 24'(-70112);
			819: out = 24'(-92484);
			820: out = 24'(-38524);
			821: out = 24'(-37220);
			822: out = 24'(10392);
			823: out = 24'(20624);
			824: out = 24'(5548);
			825: out = 24'(-28620);
			826: out = 24'(-4332);
			827: out = 24'(-8848);
			828: out = 24'(-25728);
			829: out = 24'(3876);
			830: out = 24'(15944);
			831: out = 24'(8936);
			832: out = 24'(12552);
			833: out = 24'(55140);
			834: out = 24'(16428);
			835: out = 24'(-12912);
			836: out = 24'(-15176);
			837: out = 24'(5848);
			838: out = 24'(-24180);
			839: out = 24'(-21388);
			840: out = 24'(21768);
			841: out = 24'(62324);
			842: out = 24'(61296);
			843: out = 24'(12368);
			844: out = 24'(-19948);
			845: out = 24'(-18260);
			846: out = 24'(22572);
			847: out = 24'(-4248);
			848: out = 24'(11856);
			849: out = 24'(32464);
			850: out = 24'(15136);
			851: out = 24'(1276);
			852: out = 24'(52820);
			853: out = 24'(68248);
			854: out = 24'(-14564);
			855: out = 24'(31608);
			856: out = 24'(84848);
			857: out = 24'(103852);
			858: out = 24'(53100);
			859: out = 24'(56908);
			860: out = 24'(7708);
			861: out = 24'(-12456);
			862: out = 24'(-15656);
			863: out = 24'(-77452);
			864: out = 24'(-34040);
			865: out = 24'(23408);
			866: out = 24'(50272);
			867: out = 24'(9028);
			868: out = 24'(58376);
			869: out = 24'(6800);
			870: out = 24'(-77716);
			871: out = 24'(-87152);
			872: out = 24'(32452);
			873: out = 24'(88396);
			874: out = 24'(65812);
			875: out = 24'(24784);
			876: out = 24'(-10528);
			877: out = 24'(-76168);
			878: out = 24'(-95816);
			879: out = 24'(-34380);
			880: out = 24'(-80768);
			881: out = 24'(-64492);
			882: out = 24'(-49756);
			883: out = 24'(-21436);
			884: out = 24'(-39580);
			885: out = 24'(-1612);
			886: out = 24'(-51456);
			887: out = 24'(-121296);
			888: out = 24'(-111844);
			889: out = 24'(-117796);
			890: out = 24'(-101096);
			891: out = 24'(-70336);
			892: out = 24'(-32680);
			893: out = 24'(38688);
			894: out = 24'(36840);
			895: out = 24'(-38248);
			896: out = 24'(-119840);
			897: out = 24'(-90332);
			898: out = 24'(-103236);
			899: out = 24'(-113704);
			900: out = 24'(-85532);
			901: out = 24'(11612);
			902: out = 24'(3200);
			903: out = 24'(17820);
			904: out = 24'(56216);
			905: out = 24'(11920);
			906: out = 24'(-11580);
			907: out = 24'(-61736);
			908: out = 24'(-69444);
			909: out = 24'(-26508);
			910: out = 24'(43428);
			911: out = 24'(58852);
			912: out = 24'(76804);
			913: out = 24'(120572);
			914: out = 24'(120912);
			915: out = 24'(70868);
			916: out = 24'(-9660);
			917: out = 24'(-32612);
			918: out = 24'(2556);
			919: out = 24'(88312);
			920: out = 24'(112088);
			921: out = 24'(94252);
			922: out = 24'(64652);
			923: out = 24'(106336);
			924: out = 24'(88628);
			925: out = 24'(49800);
			926: out = 24'(73696);
			927: out = 24'(52672);
			928: out = 24'(44640);
			929: out = 24'(38556);
			930: out = 24'(54132);
			931: out = 24'(87824);
			932: out = 24'(101560);
			933: out = 24'(79792);
			934: out = 24'(38572);
			935: out = 24'(44416);
			936: out = 24'(2264);
			937: out = 24'(-33160);
			938: out = 24'(-36916);
			939: out = 24'(2032);
			940: out = 24'(-11416);
			941: out = 24'(-9108);
			942: out = 24'(18088);
			943: out = 24'(20620);
			944: out = 24'(-5064);
			945: out = 24'(-35304);
			946: out = 24'(-34136);
			947: out = 24'(-13232);
			948: out = 24'(-50816);
			949: out = 24'(-57408);
			950: out = 24'(-24960);
			951: out = 24'(-20728);
			952: out = 24'(-7072);
			953: out = 24'(-60736);
			954: out = 24'(-73468);
			955: out = 24'(-32452);
			956: out = 24'(-32800);
			957: out = 24'(-45956);
			958: out = 24'(-32036);
			959: out = 24'(6136);
			960: out = 24'(39792);
			961: out = 24'(-6284);
			962: out = 24'(-22304);
			963: out = 24'(-6652);
			964: out = 24'(-9180);
			965: out = 24'(-45664);
			966: out = 24'(-23932);
			967: out = 24'(25904);
			968: out = 24'(18304);
			969: out = 24'(24236);
			970: out = 24'(17400);
			971: out = 24'(4672);
			972: out = 24'(-30224);
			973: out = 24'(-93764);
			974: out = 24'(-82060);
			975: out = 24'(-25116);
			976: out = 24'(1476);
			977: out = 24'(-16068);
			978: out = 24'(-35372);
			979: out = 24'(-52664);
			980: out = 24'(-63888);
			981: out = 24'(-40508);
			982: out = 24'(-12016);
			983: out = 24'(7960);
			984: out = 24'(-648);
			985: out = 24'(-37096);
			986: out = 24'(-3848);
			987: out = 24'(14580);
			988: out = 24'(11700);
			989: out = 24'(5948);
			990: out = 24'(-11308);
			991: out = 24'(-33808);
			992: out = 24'(-41332);
			993: out = 24'(-3004);
			994: out = 24'(51592);
			995: out = 24'(90780);
			996: out = 24'(77788);
			997: out = 24'(42432);
			998: out = 24'(46536);
			999: out = 24'(20800);
			1000: out = 24'(3912);
			1001: out = 24'(7736);
			1002: out = 24'(21420);
			1003: out = 24'(4220);
			1004: out = 24'(-23540);
			1005: out = 24'(-6784);
			1006: out = 24'(76840);
			1007: out = 24'(89840);
			1008: out = 24'(74304);
			1009: out = 24'(27060);
			1010: out = 24'(-17768);
			1011: out = 24'(-14120);
			1012: out = 24'(-8516);
			1013: out = 24'(-14156);
			1014: out = 24'(3156);
			1015: out = 24'(82312);
			1016: out = 24'(102452);
			1017: out = 24'(67120);
			1018: out = 24'(24932);
			1019: out = 24'(34220);
			1020: out = 24'(9136);
			1021: out = 24'(-18904);
			1022: out = 24'(-28972);
			1023: out = 24'(-14432);
			1024: out = 24'(39668);
			1025: out = 24'(64792);
			1026: out = 24'(64028);
			1027: out = 24'(36980);
			1028: out = 24'(3264);
			1029: out = 24'(-45024);
			1030: out = 24'(-33332);
			1031: out = 24'(29260);
			1032: out = 24'(26112);
			1033: out = 24'(9396);
			1034: out = 24'(19308);
			1035: out = 24'(34504);
			1036: out = 24'(-36220);
			1037: out = 24'(-92608);
			1038: out = 24'(-73752);
			1039: out = 24'(6244);
			1040: out = 24'(-7640);
			1041: out = 24'(31180);
			1042: out = 24'(32456);
			1043: out = 24'(26876);
			1044: out = 24'(-11932);
			1045: out = 24'(31508);
			1046: out = 24'(-25644);
			1047: out = 24'(-103524);
			1048: out = 24'(-111168);
			1049: out = 24'(-89112);
			1050: out = 24'(-40788);
			1051: out = 24'(-31748);
			1052: out = 24'(-48884);
			1053: out = 24'(-33636);
			1054: out = 24'(-24388);
			1055: out = 24'(-38892);
			1056: out = 24'(-81676);
			1057: out = 24'(-110132);
			1058: out = 24'(-82148);
			1059: out = 24'(-20924);
			1060: out = 24'(11080);
			1061: out = 24'(20680);
			1062: out = 24'(-66580);
			1063: out = 24'(-102492);
			1064: out = 24'(-93864);
			1065: out = 24'(-75176);
			1066: out = 24'(-30756);
			1067: out = 24'(18628);
			1068: out = 24'(28528);
			1069: out = 24'(4992);
			1070: out = 24'(30972);
			1071: out = 24'(25120);
			1072: out = 24'(-25468);
			1073: out = 24'(-79580);
			1074: out = 24'(10260);
			1075: out = 24'(60268);
			1076: out = 24'(92684);
			1077: out = 24'(95728);
			1078: out = 24'(91600);
			1079: out = 24'(102828);
			1080: out = 24'(94520);
			1081: out = 24'(50536);
			1082: out = 24'(-4440);
			1083: out = 24'(16236);
			1084: out = 24'(32844);
			1085: out = 24'(39380);
			1086: out = 24'(54828);
			1087: out = 24'(32376);
			1088: out = 24'(40172);
			1089: out = 24'(24172);
			1090: out = 24'(-12480);
			1091: out = 24'(-92760);
			1092: out = 24'(-23880);
			1093: out = 24'(44000);
			1094: out = 24'(21360);
			1095: out = 24'(-40796);
			1096: out = 24'(-72572);
			1097: out = 24'(-52484);
			1098: out = 24'(-27552);
			1099: out = 24'(-28928);
			1100: out = 24'(-22500);
			1101: out = 24'(-7908);
			1102: out = 24'(16392);
			1103: out = 24'(48140);
			1104: out = 24'(68764);
			1105: out = 24'(71420);
			1106: out = 24'(53304);
			1107: out = 24'(30840);
			1108: out = 24'(20932);
			1109: out = 24'(-13876);
			1110: out = 24'(-37744);
			1111: out = 24'(-24960);
			1112: out = 24'(-83988);
			1113: out = 24'(-18152);
			1114: out = 24'(-9852);
			1115: out = 24'(-23216);
			1116: out = 24'(22436);
			1117: out = 24'(60936);
			1118: out = 24'(24620);
			1119: out = 24'(-38540);
			1120: out = 24'(-41660);
			1121: out = 24'(-10804);
			1122: out = 24'(4788);
			1123: out = 24'(5284);
			1124: out = 24'(26520);
			1125: out = 24'(38820);
			1126: out = 24'(41524);
			1127: out = 24'(44588);
			1128: out = 24'(46836);
			1129: out = 24'(15840);
			1130: out = 24'(-17644);
			1131: out = 24'(-5380);
			1132: out = 24'(32716);
			1133: out = 24'(-14148);
			1134: out = 24'(8032);
			1135: out = 24'(5676);
			1136: out = 24'(-4696);
			1137: out = 24'(-2680);
			1138: out = 24'(-28716);
			1139: out = 24'(-32516);
			1140: out = 24'(-18108);
			1141: out = 24'(7784);
			1142: out = 24'(32464);
			1143: out = 24'(30536);
			1144: out = 24'(-23416);
			1145: out = 24'(-93432);
			1146: out = 24'(-117088);
			1147: out = 24'(-71608);
			1148: out = 24'(-42720);
			1149: out = 24'(-51216);
			1150: out = 24'(-42776);
			1151: out = 24'(55528);
			1152: out = 24'(98816);
			1153: out = 24'(46184);
			1154: out = 24'(-37728);
			1155: out = 24'(-43580);
			1156: out = 24'(-37436);
			1157: out = 24'(-67716);
			1158: out = 24'(-105704);
			1159: out = 24'(-79368);
			1160: out = 24'(-23840);
			1161: out = 24'(-1744);
			1162: out = 24'(-19096);
			1163: out = 24'(44476);
			1164: out = 24'(24504);
			1165: out = 24'(-19336);
			1166: out = 24'(-27816);
			1167: out = 24'(43080);
			1168: out = 24'(53644);
			1169: out = 24'(45584);
			1170: out = 24'(53496);
			1171: out = 24'(66768);
			1172: out = 24'(36600);
			1173: out = 24'(-15484);
			1174: out = 24'(-36816);
			1175: out = 24'(4616);
			1176: out = 24'(-1448);
			1177: out = 24'(-1564);
			1178: out = 24'(12524);
			1179: out = 24'(25424);
			1180: out = 24'(49748);
			1181: out = 24'(27988);
			1182: out = 24'(-11700);
			1183: out = 24'(-53564);
			1184: out = 24'(-20792);
			1185: out = 24'(-37740);
			1186: out = 24'(-24048);
			1187: out = 24'(38944);
			1188: out = 24'(117472);
			1189: out = 24'(85812);
			1190: out = 24'(66180);
			1191: out = 24'(59484);
			1192: out = 24'(45732);
			1193: out = 24'(-47552);
			1194: out = 24'(-50284);
			1195: out = 24'(23152);
			1196: out = 24'(53056);
			1197: out = 24'(43432);
			1198: out = 24'(51336);
			1199: out = 24'(67324);
			1200: out = 24'(39436);
			1201: out = 24'(16200);
			1202: out = 24'(-9204);
			1203: out = 24'(-28436);
			1204: out = 24'(-64180);
			1205: out = 24'(-34488);
			1206: out = 24'(-30068);
			1207: out = 24'(-5644);
			1208: out = 24'(-7604);
			1209: out = 24'(-44700);
			1210: out = 24'(-84916);
			1211: out = 24'(-81692);
			1212: out = 24'(-77416);
			1213: out = 24'(-90700);
			1214: out = 24'(-63952);
			1215: out = 24'(33012);
			1216: out = 24'(96236);
			1217: out = 24'(86816);
			1218: out = 24'(46256);
			1219: out = 24'(35120);
			1220: out = 24'(-28148);
			1221: out = 24'(-118056);
			1222: out = 24'(-114076);
			1223: out = 24'(-47096);
			1224: out = 24'(9852);
			1225: out = 24'(8724);
			1226: out = 24'(57808);
			1227: out = 24'(79924);
			1228: out = 24'(54908);
			1229: out = 24'(-13932);
			1230: out = 24'(-23108);
			1231: out = 24'(-70796);
			1232: out = 24'(-65092);
			1233: out = 24'(-25220);
			1234: out = 24'(27788);
			1235: out = 24'(43540);
			1236: out = 24'(34452);
			1237: out = 24'(35220);
			1238: out = 24'(74164);
			1239: out = 24'(-2256);
			1240: out = 24'(-780);
			1241: out = 24'(-10344);
			1242: out = 24'(-46948);
			1243: out = 24'(-108660);
			1244: out = 24'(-30324);
			1245: out = 24'(74876);
			1246: out = 24'(83164);
			1247: out = 24'(8908);
			1248: out = 24'(-9212);
			1249: out = 24'(3492);
			1250: out = 24'(420);
			1251: out = 24'(-17396);
			1252: out = 24'(-3412);
			1253: out = 24'(49132);
			1254: out = 24'(62004);
			1255: out = 24'(11148);
			1256: out = 24'(3264);
			1257: out = 24'(3624);
			1258: out = 24'(5956);
			1259: out = 24'(-420);
			1260: out = 24'(-1876);
			1261: out = 24'(9348);
			1262: out = 24'(12656);
			1263: out = 24'(2528);
			1264: out = 24'(-30416);
			1265: out = 24'(1076);
			1266: out = 24'(14700);
			1267: out = 24'(4180);
			1268: out = 24'(6664);
			1269: out = 24'(-2960);
			1270: out = 24'(-44400);
			1271: out = 24'(-79320);
			1272: out = 24'(-31416);
			1273: out = 24'(10252);
			1274: out = 24'(23456);
			1275: out = 24'(-7468);
			1276: out = 24'(-12040);
			1277: out = 24'(23908);
			1278: out = 24'(79888);
			1279: out = 24'(57380);
			1280: out = 24'(-22940);
			1281: out = 24'(-79560);
			1282: out = 24'(-22844);
			1283: out = 24'(69252);
			1284: out = 24'(77896);
			1285: out = 24'(-18244);
			1286: out = 24'(-13244);
			1287: out = 24'(37736);
			1288: out = 24'(59956);
			1289: out = 24'(-14740);
			1290: out = 24'(17256);
			1291: out = 24'(-6384);
			1292: out = 24'(-57748);
			1293: out = 24'(-113596);
			1294: out = 24'(-12988);
			1295: out = 24'(10176);
			1296: out = 24'(-7248);
			1297: out = 24'(-23952);
			1298: out = 24'(-11896);
			1299: out = 24'(-57304);
			1300: out = 24'(-63088);
			1301: out = 24'(-10500);
			1302: out = 24'(1780);
			1303: out = 24'(-10604);
			1304: out = 24'(-11404);
			1305: out = 24'(7756);
			1306: out = 24'(-5108);
			1307: out = 24'(-4404);
			1308: out = 24'(20728);
			1309: out = 24'(43232);
			1310: out = 24'(348);
			1311: out = 24'(36548);
			1312: out = 24'(30224);
			1313: out = 24'(12860);
			1314: out = 24'(-23132);
			1315: out = 24'(17152);
			1316: out = 24'(-33320);
			1317: out = 24'(-90860);
			1318: out = 24'(-103532);
			1319: out = 24'(-25564);
			1320: out = 24'(15628);
			1321: out = 24'(40884);
			1322: out = 24'(42444);
			1323: out = 24'(29304);
			1324: out = 24'(-32596);
			1325: out = 24'(-34500);
			1326: out = 24'(8064);
			1327: out = 24'(16672);
			1328: out = 24'(-8232);
			1329: out = 24'(-25084);
			1330: out = 24'(-26416);
			1331: out = 24'(-33232);
			1332: out = 24'(-33064);
			1333: out = 24'(-8412);
			1334: out = 24'(12080);
			1335: out = 24'(12200);
			1336: out = 24'(68908);
			1337: out = 24'(32640);
			1338: out = 24'(-25828);
			1339: out = 24'(-46876);
			1340: out = 24'(15196);
			1341: out = 24'(11348);
			1342: out = 24'(-26068);
			1343: out = 24'(-17976);
			1344: out = 24'(75304);
			1345: out = 24'(67384);
			1346: out = 24'(23412);
			1347: out = 24'(-212);
			1348: out = 24'(25572);
			1349: out = 24'(15084);
			1350: out = 24'(-9132);
			1351: out = 24'(27040);
			1352: out = 24'(124364);
			1353: out = 24'(107008);
			1354: out = 24'(104208);
			1355: out = 24'(68892);
			1356: out = 24'(13820);
			1357: out = 24'(-79552);
			1358: out = 24'(-58972);
			1359: out = 24'(37540);
			1360: out = 24'(107040);
			1361: out = 24'(86592);
			1362: out = 24'(78552);
			1363: out = 24'(59020);
			1364: out = 24'(29116);
			1365: out = 24'(-10236);
			1366: out = 24'(-80544);
			1367: out = 24'(-61356);
			1368: out = 24'(27132);
			1369: out = 24'(67268);
			1370: out = 24'(41516);
			1371: out = 24'(27388);
			1372: out = 24'(54996);
			1373: out = 24'(57792);
			1374: out = 24'(-6876);
			1375: out = 24'(-63716);
			1376: out = 24'(-46168);
			1377: out = 24'(-4652);
			1378: out = 24'(-44084);
			1379: out = 24'(-79568);
			1380: out = 24'(-52816);
			1381: out = 24'(7624);
			1382: out = 24'(-11436);
			1383: out = 24'(2928);
			1384: out = 24'(-6448);
			1385: out = 24'(-19948);
			1386: out = 24'(-38112);
			1387: out = 24'(-81216);
			1388: out = 24'(-78808);
			1389: out = 24'(-35004);
			1390: out = 24'(-4228);
			1391: out = 24'(-45976);
			1392: out = 24'(-61916);
			1393: out = 24'(-59808);
			1394: out = 24'(-58912);
			1395: out = 24'(-42864);
			1396: out = 24'(-32892);
			1397: out = 24'(-10556);
			1398: out = 24'(-3664);
			1399: out = 24'(-85316);
			1400: out = 24'(-21756);
			1401: out = 24'(39344);
			1402: out = 24'(37340);
			1403: out = 24'(-46924);
			1404: out = 24'(-8184);
			1405: out = 24'(-27908);
			1406: out = 24'(-80016);
			1407: out = 24'(-104688);
			1408: out = 24'(-50768);
			1409: out = 24'(-10948);
			1410: out = 24'(-6728);
			1411: out = 24'(-17124);
			1412: out = 24'(3668);
			1413: out = 24'(29772);
			1414: out = 24'(60532);
			1415: out = 24'(49360);
			1416: out = 24'(-1776);
			1417: out = 24'(-30560);
			1418: out = 24'(44348);
			1419: out = 24'(105752);
			1420: out = 24'(20900);
			1421: out = 24'(8408);
			1422: out = 24'(31268);
			1423: out = 24'(39504);
			1424: out = 24'(-34852);
			1425: out = 24'(-33140);
			1426: out = 24'(-14700);
			1427: out = 24'(-10580);
			1428: out = 24'(-45056);
			1429: out = 24'(-8464);
			1430: out = 24'(65760);
			1431: out = 24'(101472);
			1432: out = 24'(54088);
			1433: out = 24'(20316);
			1434: out = 24'(-11176);
			1435: out = 24'(-4028);
			1436: out = 24'(9412);
			1437: out = 24'(50964);
			1438: out = 24'(42708);
			1439: out = 24'(41604);
			1440: out = 24'(28220);
			1441: out = 24'(16712);
			1442: out = 24'(-35300);
			1443: out = 24'(-26520);
			1444: out = 24'(22164);
			1445: out = 24'(64636);
			1446: out = 24'(36508);
			1447: out = 24'(54292);
			1448: out = 24'(57308);
			1449: out = 24'(17376);
			1450: out = 24'(74716);
			1451: out = 24'(41068);
			1452: out = 24'(-17204);
			1453: out = 24'(-61096);
			1454: out = 24'(12492);
			1455: out = 24'(4380);
			1456: out = 24'(-9092);
			1457: out = 24'(18736);
			1458: out = 24'(115012);
			1459: out = 24'(41640);
			1460: out = 24'(-26384);
			1461: out = 24'(-41380);
			1462: out = 24'(29272);
			1463: out = 24'(-21740);
			1464: out = 24'(-20528);
			1465: out = 24'(9420);
			1466: out = 24'(45452);
			1467: out = 24'(-11440);
			1468: out = 24'(-4192);
			1469: out = 24'(-22176);
			1470: out = 24'(-81580);
			1471: out = 24'(-76548);
			1472: out = 24'(-44976);
			1473: out = 24'(-18000);
			1474: out = 24'(-4604);
			1475: out = 24'(29128);
			1476: out = 24'(58184);
			1477: out = 24'(22932);
			1478: out = 24'(-27028);
			1479: out = 24'(35172);
			1480: out = 24'(15624);
			1481: out = 24'(7384);
			1482: out = 24'(-3976);
			1483: out = 24'(31084);
			1484: out = 24'(-77652);
			1485: out = 24'(-69520);
			1486: out = 24'(-28544);
			1487: out = 24'(-14608);
			1488: out = 24'(-82436);
			1489: out = 24'(-40800);
			1490: out = 24'(-19576);
			1491: out = 24'(-100764);
			1492: out = 24'(-112244);
			1493: out = 24'(-112780);
			1494: out = 24'(-42736);
			1495: out = 24'(26444);
			1496: out = 24'(57804);
			1497: out = 24'(20680);
			1498: out = 24'(-8644);
			1499: out = 24'(-12744);
			1500: out = 24'(6156);
			1501: out = 24'(-31560);
			1502: out = 24'(-36052);
			1503: out = 24'(-11652);
			1504: out = 24'(3364);
			1505: out = 24'(-50560);
			1506: out = 24'(-56552);
			1507: out = 24'(-2820);
			1508: out = 24'(50656);
			1509: out = 24'(25344);
			1510: out = 24'(11716);
			1511: out = 24'(16844);
			1512: out = 24'(17876);
			1513: out = 24'(-75764);
			1514: out = 24'(-24564);
			1515: out = 24'(21780);
			1516: out = 24'(25552);
			1517: out = 24'(8832);
			1518: out = 24'(18948);
			1519: out = 24'(33828);
			1520: out = 24'(43304);
			1521: out = 24'(37540);
			1522: out = 24'(12808);
			1523: out = 24'(-2096);
			1524: out = 24'(2216);
			1525: out = 24'(14952);
			1526: out = 24'(55132);
			1527: out = 24'(55336);
			1528: out = 24'(61496);
			1529: out = 24'(58404);
			1530: out = 24'(19128);
			1531: out = 24'(-5504);
			1532: out = 24'(3736);
			1533: out = 24'(-432);
			1534: out = 24'(-81216);
			1535: out = 24'(-33500);
			1536: out = 24'(66148);
			1537: out = 24'(118124);
			1538: out = 24'(89104);
			1539: out = 24'(80560);
			1540: out = 24'(71256);
			1541: out = 24'(38388);
			1542: out = 24'(-33760);
			1543: out = 24'(-14360);
			1544: out = 24'(-1780);
			1545: out = 24'(22252);
			1546: out = 24'(47220);
			1547: out = 24'(81628);
			1548: out = 24'(70880);
			1549: out = 24'(30308);
			1550: out = 24'(-15860);
			1551: out = 24'(-6740);
			1552: out = 24'(-12296);
			1553: out = 24'(1244);
			1554: out = 24'(17916);
			1555: out = 24'(44988);
			1556: out = 24'(57488);
			1557: out = 24'(64728);
			1558: out = 24'(9500);
			1559: out = 24'(-106716);
			1560: out = 24'(-68144);
			1561: out = 24'(-24592);
			1562: out = 24'(-22556);
			1563: out = 24'(-76896);
			1564: out = 24'(-65628);
			1565: out = 24'(-76316);
			1566: out = 24'(-78528);
			1567: out = 24'(-90060);
			1568: out = 24'(-37544);
			1569: out = 24'(-50340);
			1570: out = 24'(-22196);
			1571: out = 24'(-7576);
			1572: out = 24'(-32620);
			1573: out = 24'(-88176);
			1574: out = 24'(-30480);
			1575: out = 24'(46540);
			1576: out = 24'(10300);
			1577: out = 24'(-10364);
			1578: out = 24'(-29464);
			1579: out = 24'(-56556);
			1580: out = 24'(-117136);
			1581: out = 24'(-86600);
			1582: out = 24'(-48296);
			1583: out = 24'(-30468);
			1584: out = 24'(-34008);
			1585: out = 24'(68560);
			1586: out = 24'(36412);
			1587: out = 24'(-41360);
			1588: out = 24'(-105220);
			1589: out = 24'(-29036);
			1590: out = 24'(-31580);
			1591: out = 24'(-36012);
			1592: out = 24'(-11708);
			1593: out = 24'(80044);
			1594: out = 24'(49488);
			1595: out = 24'(40180);
			1596: out = 24'(23028);
			1597: out = 24'(8860);
			1598: out = 24'(-74124);
			1599: out = 24'(-40464);
			1600: out = 24'(21452);
			1601: out = 24'(20720);
			1602: out = 24'(16416);
			1603: out = 24'(28140);
			1604: out = 24'(66472);
			1605: out = 24'(75840);
			1606: out = 24'(25360);
			1607: out = 24'(4228);
			1608: out = 24'(-13264);
			1609: out = 24'(-39800);
			1610: out = 24'(-57188);
			1611: out = 24'(-31932);
			1612: out = 24'(49688);
			1613: out = 24'(121396);
			1614: out = 24'(117528);
			1615: out = 24'(108044);
			1616: out = 24'(40736);
			1617: out = 24'(-12016);
			1618: out = 24'(-21172);
			1619: out = 24'(-50132);
			1620: out = 24'(-1748);
			1621: out = 24'(77520);
			1622: out = 24'(119064);
			1623: out = 24'(119424);
			1624: out = 24'(92672);
			1625: out = 24'(38228);
			1626: out = 24'(-30052);
			1627: out = 24'(-68828);
			1628: out = 24'(-110556);
			1629: out = 24'(-81616);
			1630: out = 24'(8288);
			1631: out = 24'(91636);
			1632: out = 24'(116216);
			1633: out = 24'(122368);
			1634: out = 24'(92316);
			1635: out = 24'(-16620);
			1636: out = 24'(-98096);
			1637: out = 24'(-111176);
			1638: out = 24'(-32584);
			1639: out = 24'(26936);
			1640: out = 24'(24368);
			1641: out = 24'(-7036);
			1642: out = 24'(40140);
			1643: out = 24'(89004);
			1644: out = 24'(-18464);
			1645: out = 24'(-101500);
			1646: out = 24'(-96976);
			1647: out = 24'(-26812);
			1648: out = 24'(-47444);
			1649: out = 24'(-102848);
			1650: out = 24'(-99988);
			1651: out = 24'(-14592);
			1652: out = 24'(28248);
			1653: out = 24'(-33772);
			1654: out = 24'(-103916);
			1655: out = 24'(-91960);
			1656: out = 24'(-6056);
			1657: out = 24'(-2432);
			1658: out = 24'(-21412);
			1659: out = 24'(-54916);
			1660: out = 24'(-60908);
			1661: out = 24'(572);
			1662: out = 24'(12948);
			1663: out = 24'(-39380);
			1664: out = 24'(-88628);
			1665: out = 24'(-13148);
			1666: out = 24'(46152);
			1667: out = 24'(58260);
			1668: out = 24'(2344);
			1669: out = 24'(-86684);
			1670: out = 24'(-48540);
			1671: out = 24'(-344);
			1672: out = 24'(-14580);
			1673: out = 24'(-62744);
			1674: out = 24'(-55668);
			1675: out = 24'(11892);
			1676: out = 24'(52208);
			1677: out = 24'(20060);
			1678: out = 24'(5520);
			1679: out = 24'(14988);
			1680: out = 24'(55088);
			1681: out = 24'(52864);
			1682: out = 24'(20088);
			1683: out = 24'(-4964);
			1684: out = 24'(44784);
			1685: out = 24'(77300);
			1686: out = 24'(24572);
			1687: out = 24'(10168);
			1688: out = 24'(52644);
			1689: out = 24'(65104);
			1690: out = 24'(-22024);
			1691: out = 24'(-43208);
			1692: out = 24'(-2968);
			1693: out = 24'(57420);
			1694: out = 24'(52732);
			1695: out = 24'(71628);
			1696: out = 24'(39240);
			1697: out = 24'(6812);
			1698: out = 24'(-17784);
			1699: out = 24'(34792);
			1700: out = 24'(14744);
			1701: out = 24'(-10784);
			1702: out = 24'(-8712);
			1703: out = 24'(65260);
			1704: out = 24'(55672);
			1705: out = 24'(43908);
			1706: out = 24'(28868);
			1707: out = 24'(28664);
			1708: out = 24'(27768);
			1709: out = 24'(32648);
			1710: out = 24'(8016);
			1711: out = 24'(-23420);
			1712: out = 24'(-24656);
			1713: out = 24'(5304);
			1714: out = 24'(-5240);
			1715: out = 24'(-37300);
			1716: out = 24'(-8808);
			1717: out = 24'(50648);
			1718: out = 24'(49308);
			1719: out = 24'(7072);
			1720: out = 24'(16284);
			1721: out = 24'(1688);
			1722: out = 24'(-64608);
			1723: out = 24'(-103960);
			1724: out = 24'(17696);
			1725: out = 24'(44684);
			1726: out = 24'(6696);
			1727: out = 24'(-26496);
			1728: out = 24'(39592);
			1729: out = 24'(49504);
			1730: out = 24'(24360);
			1731: out = 24'(-31500);
			1732: out = 24'(-37320);
			1733: out = 24'(-75124);
			1734: out = 24'(-71388);
			1735: out = 24'(-94640);
			1736: out = 24'(-87532);
			1737: out = 24'(-10812);
			1738: out = 24'(69608);
			1739: out = 24'(34592);
			1740: out = 24'(-44468);
			1741: out = 24'(-33468);
			1742: out = 24'(-34272);
			1743: out = 24'(-46236);
			1744: out = 24'(-45968);
			1745: out = 24'(3416);
			1746: out = 24'(-15072);
			1747: out = 24'(-39856);
			1748: out = 24'(-5408);
			1749: out = 24'(86044);
			1750: out = 24'(82236);
			1751: out = 24'(29740);
			1752: out = 24'(-9884);
			1753: out = 24'(5132);
			1754: out = 24'(-32708);
			1755: out = 24'(-42028);
			1756: out = 24'(-13988);
			1757: out = 24'(49900);
			1758: out = 24'(45280);
			1759: out = 24'(62760);
			1760: out = 24'(49148);
			1761: out = 24'(19400);
			1762: out = 24'(-60504);
			1763: out = 24'(-48400);
			1764: out = 24'(-26984);
			1765: out = 24'(3324);
			1766: out = 24'(-2488);
			1767: out = 24'(28188);
			1768: out = 24'(1852);
			1769: out = 24'(13280);
			1770: out = 24'(45808);
			1771: out = 24'(31568);
			1772: out = 24'(-74640);
			1773: out = 24'(-96988);
			1774: out = 24'(13564);
			1775: out = 24'(49620);
			1776: out = 24'(45764);
			1777: out = 24'(40436);
			1778: out = 24'(34704);
			1779: out = 24'(-67284);
			1780: out = 24'(-107816);
			1781: out = 24'(-100480);
			1782: out = 24'(-63332);
			1783: out = 24'(-99644);
			1784: out = 24'(-29156);
			1785: out = 24'(28844);
			1786: out = 24'(77428);
			1787: out = 24'(76228);
			1788: out = 24'(68140);
			1789: out = 24'(22928);
			1790: out = 24'(24716);
			1791: out = 24'(47460);
			1792: out = 24'(15480);
			1793: out = 24'(-2812);
			1794: out = 24'(37256);
			1795: out = 24'(82428);
			1796: out = 24'(47652);
			1797: out = 24'(332);
			1798: out = 24'(-160);
			1799: out = 24'(52488);
			1800: out = 24'(86008);
			1801: out = 24'(58820);
			1802: out = 24'(36540);
			1803: out = 24'(19532);
			1804: out = 24'(-13472);
			1805: out = 24'(-2636);
			1806: out = 24'(36572);
			1807: out = 24'(51136);
			1808: out = 24'(1404);
			1809: out = 24'(25448);
			1810: out = 24'(-20384);
			1811: out = 24'(-73696);
			1812: out = 24'(-104756);
			1813: out = 24'(37560);
			1814: out = 24'(11304);
			1815: out = 24'(-2072);
			1816: out = 24'(26108);
			1817: out = 24'(93444);
			1818: out = 24'(-39276);
			1819: out = 24'(-122752);
			1820: out = 24'(-111996);
			1821: out = 24'(-113584);
			1822: out = 24'(-11280);
			1823: out = 24'(88180);
			1824: out = 24'(103028);
			1825: out = 24'(52916);
			1826: out = 24'(-33720);
			1827: out = 24'(-46232);
			1828: out = 24'(-58156);
			1829: out = 24'(-117252);
			1830: out = 24'(-115216);
			1831: out = 24'(-75248);
			1832: out = 24'(2388);
			1833: out = 24'(25488);
			1834: out = 24'(36680);
			1835: out = 24'(9464);
			1836: out = 24'(11192);
			1837: out = 24'(24092);
			1838: out = 24'(48952);
			1839: out = 24'(-45600);
			1840: out = 24'(-93520);
			1841: out = 24'(-67940);
			1842: out = 24'(6408);
			1843: out = 24'(-58484);
			1844: out = 24'(-39800);
			1845: out = 24'(32248);
			1846: out = 24'(61428);
			1847: out = 24'(-35556);
			1848: out = 24'(-99844);
			1849: out = 24'(-100908);
			1850: out = 24'(-31348);
			1851: out = 24'(61080);
			1852: out = 24'(118768);
			1853: out = 24'(109536);
			1854: out = 24'(79588);
			1855: out = 24'(49004);
			1856: out = 24'(54968);
			1857: out = 24'(5004);
			1858: out = 24'(-42816);
			1859: out = 24'(8040);
			1860: out = 24'(62364);
			1861: out = 24'(68448);
			1862: out = 24'(38252);
			1863: out = 24'(51608);
			1864: out = 24'(27656);
			1865: out = 24'(39064);
			1866: out = 24'(3232);
			1867: out = 24'(-50160);
			1868: out = 24'(-64984);
			1869: out = 24'(10784);
			1870: out = 24'(76960);
			1871: out = 24'(76352);
			1872: out = 24'(440);
			1873: out = 24'(46976);
			1874: out = 24'(90372);
			1875: out = 24'(71180);
			1876: out = 24'(-29288);
			1877: out = 24'(-11424);
			1878: out = 24'(-19080);
			1879: out = 24'(-49580);
			1880: out = 24'(-81104);
			1881: out = 24'(44);
			1882: out = 24'(10936);
			1883: out = 24'(-7572);
			1884: out = 24'(-2740);
			1885: out = 24'(-3208);
			1886: out = 24'(-51188);
			1887: out = 24'(-75764);
			1888: out = 24'(-21136);
			1889: out = 24'(-7904);
			1890: out = 24'(-24016);
			1891: out = 24'(-64816);
			1892: out = 24'(-64364);
			1893: out = 24'(-82088);
			1894: out = 24'(-13160);
			1895: out = 24'(-10192);
			1896: out = 24'(-45636);
			1897: out = 24'(-87636);
			1898: out = 24'(3428);
			1899: out = 24'(27848);
			1900: out = 24'(4400);
			1901: out = 24'(1040);
			1902: out = 24'(34640);
			1903: out = 24'(-608);
			1904: out = 24'(-70092);
			1905: out = 24'(-98268);
			1906: out = 24'(-9088);
			1907: out = 24'(5096);
			1908: out = 24'(-16752);
			1909: out = 24'(-2736);
			1910: out = 24'(48796);
			1911: out = 24'(21936);
			1912: out = 24'(-29992);
			1913: out = 24'(-59840);
			1914: out = 24'(-95460);
			1915: out = 24'(-488);
			1916: out = 24'(62548);
			1917: out = 24'(67676);
			1918: out = 24'(40868);
			1919: out = 24'(37552);
			1920: out = 24'(18480);
			1921: out = 24'(-3072);
			1922: out = 24'(-13660);
			1923: out = 24'(35124);
			1924: out = 24'(29528);
			1925: out = 24'(22368);
			1926: out = 24'(50012);
			1927: out = 24'(97216);
			1928: out = 24'(81504);
			1929: out = 24'(34408);
			1930: out = 24'(-10884);
			1931: out = 24'(-44156);
			1932: out = 24'(-37120);
			1933: out = 24'(-18272);
			1934: out = 24'(-4496);
			1935: out = 24'(7720);
			1936: out = 24'(94280);
			1937: out = 24'(124784);
			1938: out = 24'(76112);
			1939: out = 24'(-14428);
			1940: out = 24'(-6956);
			1941: out = 24'(-22360);
			1942: out = 24'(-67884);
			1943: out = 24'(-94948);
			1944: out = 24'(17108);
			1945: out = 24'(105056);
			1946: out = 24'(102316);
			1947: out = 24'(47956);
			1948: out = 24'(20232);
			1949: out = 24'(40288);
			1950: out = 24'(47272);
			1951: out = 24'(14516);
			1952: out = 24'(-2428);
			1953: out = 24'(-12292);
			1954: out = 24'(12940);
			1955: out = 24'(25736);
			1956: out = 24'(17216);
			1957: out = 24'(-36580);
			1958: out = 24'(-35140);
			1959: out = 24'(-1228);
			1960: out = 24'(3836);
			1961: out = 24'(-89812);
			1962: out = 24'(-124572);
			1963: out = 24'(-83704);
			1964: out = 24'(-8704);
			1965: out = 24'(-62224);
			1966: out = 24'(-35296);
			1967: out = 24'(-18452);
			1968: out = 24'(-4284);
			1969: out = 24'(44672);
			1970: out = 24'(500);
			1971: out = 24'(-81364);
			1972: out = 24'(-109508);
			1973: out = 24'(-7140);
			1974: out = 24'(-13748);
			1975: out = 24'(-33924);
			1976: out = 24'(-27632);
			1977: out = 24'(20204);
			1978: out = 24'(-33568);
			1979: out = 24'(-48572);
			1980: out = 24'(-27952);
			1981: out = 24'(33768);
			1982: out = 24'(62072);
			1983: out = 24'(50752);
			1984: out = 24'(-17848);
			1985: out = 24'(-53928);
			1986: out = 24'(13852);
			1987: out = 24'(86164);
			1988: out = 24'(86588);
			1989: out = 24'(60896);
			1990: out = 24'(44444);
			1991: out = 24'(15772);
			1992: out = 24'(-38192);
			1993: out = 24'(-50876);
			1994: out = 24'(-18220);
			1995: out = 24'(-5308);
			1996: out = 24'(-76116);
			1997: out = 24'(-73484);
			1998: out = 24'(48112);
			1999: out = 24'(50528);
			2000: out = 24'(-15296);
			2001: out = 24'(-15128);
			2002: out = 24'(95960);
			2003: out = 24'(54736);
			2004: out = 24'(44544);
			2005: out = 24'(452);
			2006: out = 24'(7736);
			2007: out = 24'(-8620);
			2008: out = 24'(11384);
			2009: out = 24'(-53256);
			2010: out = 24'(-79524);
			2011: out = 24'(-5064);
			2012: out = 24'(44688);
			2013: out = 24'(22844);
			2014: out = 24'(5348);
			2015: out = 24'(19436);
			2016: out = 24'(-11476);
			2017: out = 24'(-71436);
			2018: out = 24'(-63752);
			2019: out = 24'(28136);
			2020: out = 24'(26804);
			2021: out = 24'(14024);
			2022: out = 24'(9400);
			2023: out = 24'(32964);
			2024: out = 24'(14136);
			2025: out = 24'(39884);
			2026: out = 24'(56096);
			2027: out = 24'(38636);
			2028: out = 24'(-49912);
			2029: out = 24'(-110392);
			2030: out = 24'(-95040);
			2031: out = 24'(-17584);
			2032: out = 24'(15280);
			2033: out = 24'(21092);
			2034: out = 24'(22864);
			2035: out = 24'(29136);
			2036: out = 24'(2112);
			2037: out = 24'(9996);
			2038: out = 24'(-27356);
			2039: out = 24'(-15568);
			2040: out = 24'(17692);
			2041: out = 24'(4020);
			2042: out = 24'(-26184);
			2043: out = 24'(-13596);
			2044: out = 24'(44992);
			2045: out = 24'(101388);
			2046: out = 24'(36844);
			2047: out = 24'(-9036);
			2048: out = 24'(-22340);
			2049: out = 24'(-13000);
			2050: out = 24'(-24112);
			2051: out = 24'(37940);
			2052: out = 24'(102056);
			2053: out = 24'(91156);
			2054: out = 24'(52472);
			2055: out = 24'(10456);
			2056: out = 24'(-17056);
			2057: out = 24'(-47672);
			2058: out = 24'(-75596);
			2059: out = 24'(-43304);
			2060: out = 24'(-624);
			2061: out = 24'(-5416);
			2062: out = 24'(5088);
			2063: out = 24'(15560);
			2064: out = 24'(76292);
			2065: out = 24'(95672);
			2066: out = 24'(50312);
			2067: out = 24'(-29884);
			2068: out = 24'(-59460);
			2069: out = 24'(-50108);
			2070: out = 24'(-20920);
			2071: out = 24'(-10168);
			2072: out = 24'(57156);
			2073: out = 24'(96808);
			2074: out = 24'(85684);
			2075: out = 24'(23728);
			2076: out = 24'(3016);
			2077: out = 24'(-69740);
			2078: out = 24'(-117124);
			2079: out = 24'(-120360);
			2080: out = 24'(-11576);
			2081: out = 24'(60716);
			2082: out = 24'(38108);
			2083: out = 24'(58648);
			2084: out = 24'(81148);
			2085: out = 24'(38404);
			2086: out = 24'(-42172);
			2087: out = 24'(6692);
			2088: out = 24'(5356);
			2089: out = 24'(29636);
			2090: out = 24'(-36932);
			2091: out = 24'(-104580);
			2092: out = 24'(-121188);
			2093: out = 24'(936);
			2094: out = 24'(51660);
			2095: out = 24'(2148);
			2096: out = 24'(-36404);
			2097: out = 24'(-21844);
			2098: out = 24'(-62320);
			2099: out = 24'(-123808);
			2100: out = 24'(-77096);
			2101: out = 24'(34260);
			2102: out = 24'(89892);
			2103: out = 24'(63384);
			2104: out = 24'(13520);
			2105: out = 24'(-35908);
			2106: out = 24'(-90180);
			2107: out = 24'(-100124);
			2108: out = 24'(-33720);
			2109: out = 24'(-43044);
			2110: out = 24'(-63216);
			2111: out = 24'(-16012);
			2112: out = 24'(104548);
			2113: out = 24'(106264);
			2114: out = 24'(42588);
			2115: out = 24'(-34500);
			2116: out = 24'(-39668);
			2117: out = 24'(-95624);
			2118: out = 24'(-55068);
			2119: out = 24'(-44624);
			2120: out = 24'(-10704);
			2121: out = 24'(32624);
			2122: out = 24'(63704);
			2123: out = 24'(-42072);
			2124: out = 24'(-118704);
			2125: out = 24'(-47864);
			2126: out = 24'(66988);
			2127: out = 24'(29692);
			2128: out = 24'(-44860);
			2129: out = 24'(-14044);
			2130: out = 24'(50888);
			2131: out = 24'(40624);
			2132: out = 24'(-18992);
			2133: out = 24'(-12668);
			2134: out = 24'(52336);
			2135: out = 24'(86160);
			2136: out = 24'(50184);
			2137: out = 24'(24312);
			2138: out = 24'(57660);
			2139: out = 24'(42668);
			2140: out = 24'(-12808);
			2141: out = 24'(-71856);
			2142: out = 24'(-94772);
			2143: out = 24'(-9228);
			2144: out = 24'(61064);
			2145: out = 24'(68512);
			2146: out = 24'(25320);
			2147: out = 24'(21360);
			2148: out = 24'(24492);
			2149: out = 24'(70112);
			2150: out = 24'(103568);
			2151: out = 24'(87524);
			2152: out = 24'(0);
			2153: out = 24'(-58352);
			2154: out = 24'(-60628);
			2155: out = 24'(-38816);
			2156: out = 24'(-43988);
			2157: out = 24'(17608);
			2158: out = 24'(92004);
			2159: out = 24'(53788);
			2160: out = 24'(3628);
			2161: out = 24'(-21052);
			2162: out = 24'(5156);
			2163: out = 24'(-8152);
			2164: out = 24'(4144);
			2165: out = 24'(-12120);
			2166: out = 24'(-1844);
			2167: out = 24'(-1360);
			2168: out = 24'(4356);
			2169: out = 24'(-33528);
			2170: out = 24'(-6364);
			2171: out = 24'(64532);
			2172: out = 24'(79548);
			2173: out = 24'(53384);
			2174: out = 24'(29540);
			2175: out = 24'(860);
			2176: out = 24'(-51960);
			2177: out = 24'(-73008);
			2178: out = 24'(-4320);
			2179: out = 24'(69504);
			2180: out = 24'(53000);
			2181: out = 24'(10612);
			2182: out = 24'(27380);
			2183: out = 24'(43284);
			2184: out = 24'(-68008);
			2185: out = 24'(-110488);
			2186: out = 24'(-109180);
			2187: out = 24'(-9440);
			2188: out = 24'(68892);
			2189: out = 24'(72564);
			2190: out = 24'(44840);
			2191: out = 24'(25484);
			2192: out = 24'(-2612);
			2193: out = 24'(-36668);
			2194: out = 24'(-89064);
			2195: out = 24'(-63468);
			2196: out = 24'(22636);
			2197: out = 24'(78900);
			2198: out = 24'(74152);
			2199: out = 24'(53108);
			2200: out = 24'(35176);
			2201: out = 24'(27256);
			2202: out = 24'(-90008);
			2203: out = 24'(-118612);
			2204: out = 24'(-116692);
			2205: out = 24'(-103156);
			2206: out = 24'(-17448);
			2207: out = 24'(39036);
			2208: out = 24'(1540);
			2209: out = 24'(-67392);
			2210: out = 24'(-26120);
			2211: out = 24'(29568);
			2212: out = 24'(5992);
			2213: out = 24'(-73272);
			2214: out = 24'(-86944);
			2215: out = 24'(-37808);
			2216: out = 24'(-49236);
			2217: out = 24'(-126360);
			2218: out = 24'(-102988);
			2219: out = 24'(2772);
			2220: out = 24'(117628);
			2221: out = 24'(83232);
			2222: out = 24'(6928);
			2223: out = 24'(-97828);
			2224: out = 24'(-41104);
			2225: out = 24'(-10088);
			2226: out = 24'(-67216);
			2227: out = 24'(-102904);
			2228: out = 24'(6740);
			2229: out = 24'(99668);
			2230: out = 24'(78076);
			2231: out = 24'(29616);
			2232: out = 24'(24048);
			2233: out = 24'(23748);
			2234: out = 24'(-2496);
			2235: out = 24'(-25972);
			2236: out = 24'(20100);
			2237: out = 24'(43056);
			2238: out = 24'(43452);
			2239: out = 24'(66560);
			2240: out = 24'(74612);
			2241: out = 24'(62928);
			2242: out = 24'(42400);
			2243: out = 24'(51144);
			2244: out = 24'(53256);
			2245: out = 24'(33192);
			2246: out = 24'(-7688);
			2247: out = 24'(-20992);
			2248: out = 24'(-27168);
			2249: out = 24'(40544);
			2250: out = 24'(62220);
			2251: out = 24'(13512);
			2252: out = 24'(-112604);
			2253: out = 24'(-53456);
			2254: out = 24'(9472);
			2255: out = 24'(27528);
			2256: out = 24'(12844);
			2257: out = 24'(53688);
			2258: out = 24'(31144);
			2259: out = 24'(14220);
			2260: out = 24'(32656);
			2261: out = 24'(43036);
			2262: out = 24'(15996);
			2263: out = 24'(2976);
			2264: out = 24'(7368);
			2265: out = 24'(940);
			2266: out = 24'(-56016);
			2267: out = 24'(-28112);
			2268: out = 24'(69924);
			2269: out = 24'(56144);
			2270: out = 24'(-6164);
			2271: out = 24'(-72416);
			2272: out = 24'(-71488);
			2273: out = 24'(-59880);
			2274: out = 24'(-68124);
			2275: out = 24'(-52948);
			2276: out = 24'(31868);
			2277: out = 24'(77656);
			2278: out = 24'(95316);
			2279: out = 24'(-25280);
			2280: out = 24'(-121660);
			2281: out = 24'(-106624);
			2282: out = 24'(55368);
			2283: out = 24'(53060);
			2284: out = 24'(-18072);
			2285: out = 24'(-13252);
			2286: out = 24'(97376);
			2287: out = 24'(86852);
			2288: out = 24'(18444);
			2289: out = 24'(-61304);
			2290: out = 24'(-115844);
			2291: out = 24'(-112112);
			2292: out = 24'(-93376);
			2293: out = 24'(-44564);
			2294: out = 24'(6448);
			2295: out = 24'(65532);
			2296: out = 24'(41560);
			2297: out = 24'(-21888);
			2298: out = 24'(-61752);
			2299: out = 24'(-83072);
			2300: out = 24'(-13012);
			2301: out = 24'(55276);
			2302: out = 24'(57148);
			2303: out = 24'(54848);
			2304: out = 24'(44508);
			2305: out = 24'(56856);
			2306: out = 24'(50696);
			2307: out = 24'(31816);
			2308: out = 24'(-44116);
			2309: out = 24'(-61900);
			2310: out = 24'(-22204);
			2311: out = 24'(12984);
			2312: out = 24'(-57808);
			2313: out = 24'(-72332);
			2314: out = 24'(2552);
			2315: out = 24'(65860);
			2316: out = 24'(844);
			2317: out = 24'(-53068);
			2318: out = 24'(-55760);
			2319: out = 24'(-33856);
			2320: out = 24'(-43104);
			2321: out = 24'(-48192);
			2322: out = 24'(-36404);
			2323: out = 24'(-12652);
			2324: out = 24'(51280);
			2325: out = 24'(46896);
			2326: out = 24'(19980);
			2327: out = 24'(-24424);
			2328: out = 24'(-15188);
			2329: out = 24'(-27076);
			2330: out = 24'(46876);
			2331: out = 24'(100444);
			2332: out = 24'(68396);
			2333: out = 24'(-7656);
			2334: out = 24'(-15624);
			2335: out = 24'(9472);
			2336: out = 24'(-556);
			2337: out = 24'(-61400);
			2338: out = 24'(-18368);
			2339: out = 24'(60004);
			2340: out = 24'(61440);
			2341: out = 24'(12400);
			2342: out = 24'(5784);
			2343: out = 24'(27560);
			2344: out = 24'(26164);
			2345: out = 24'(32544);
			2346: out = 24'(37376);
			2347: out = 24'(61620);
			2348: out = 24'(56296);
			2349: out = 24'(13176);
			2350: out = 24'(-57820);
			2351: out = 24'(-60204);
			2352: out = 24'(17128);
			2353: out = 24'(72984);
			2354: out = 24'(60012);
			2355: out = 24'(5012);
			2356: out = 24'(-9468);
			2357: out = 24'(24500);
			2358: out = 24'(14184);
			2359: out = 24'(-53744);
			2360: out = 24'(-99064);
			2361: out = 24'(-29884);
			2362: out = 24'(52468);
			2363: out = 24'(83624);
			2364: out = 24'(33164);
			2365: out = 24'(2052);
			2366: out = 24'(31436);
			2367: out = 24'(69916);
			2368: out = 24'(6060);
			2369: out = 24'(-97332);
			2370: out = 24'(-113776);
			2371: out = 24'(-62796);
			2372: out = 24'(-35456);
			2373: out = 24'(-69644);
			2374: out = 24'(-86544);
			2375: out = 24'(-69652);
			2376: out = 24'(392);
			2377: out = 24'(34620);
			2378: out = 24'(12516);
			2379: out = 24'(640);
			2380: out = 24'(25928);
			2381: out = 24'(64956);
			2382: out = 24'(37216);
			2383: out = 24'(-36732);
			2384: out = 24'(-107852);
			2385: out = 24'(-35328);
			2386: out = 24'(72424);
			2387: out = 24'(36620);
			2388: out = 24'(440);
			2389: out = 24'(16808);
			2390: out = 24'(70044);
			2391: out = 24'(33392);
			2392: out = 24'(-1036);
			2393: out = 24'(-61476);
			2394: out = 24'(-41168);
			2395: out = 24'(15900);
			2396: out = 24'(26704);
			2397: out = 24'(-18720);
			2398: out = 24'(-13536);
			2399: out = 24'(57576);
			2400: out = 24'(96548);
			2401: out = 24'(63120);
			2402: out = 24'(-8144);
			2403: out = 24'(-74708);
			2404: out = 24'(-99144);
			2405: out = 24'(-61212);
			2406: out = 24'(7872);
			2407: out = 24'(27496);
			2408: out = 24'(-13116);
			2409: out = 24'(-22800);
			2410: out = 24'(8884);
			2411: out = 24'(25608);
			2412: out = 24'(-1320);
			2413: out = 24'(-6732);
			2414: out = 24'(40956);
			2415: out = 24'(71276);
			2416: out = 24'(32520);
			2417: out = 24'(-6648);
			2418: out = 24'(-45432);
			2419: out = 24'(-58796);
			2420: out = 24'(-75296);
			2421: out = 24'(-96212);
			2422: out = 24'(-21524);
			2423: out = 24'(69304);
			2424: out = 24'(78196);
			2425: out = 24'(15948);
			2426: out = 24'(-37928);
			2427: out = 24'(-47564);
			2428: out = 24'(-25532);
			2429: out = 24'(-5584);
			2430: out = 24'(-30200);
			2431: out = 24'(-5408);
			2432: out = 24'(26320);
			2433: out = 24'(9520);
			2434: out = 24'(-23772);
			2435: out = 24'(-41228);
			2436: out = 24'(-9324);
			2437: out = 24'(17624);
			2438: out = 24'(7032);
			2439: out = 24'(-46684);
			2440: out = 24'(-41520);
			2441: out = 24'(23756);
			2442: out = 24'(39616);
			2443: out = 24'(60320);
			2444: out = 24'(19272);
			2445: out = 24'(-37708);
			2446: out = 24'(-76500);
			2447: out = 24'(-7616);
			2448: out = 24'(40928);
			2449: out = 24'(53200);
			2450: out = 24'(58884);
			2451: out = 24'(78068);
			2452: out = 24'(88020);
			2453: out = 24'(58500);
			2454: out = 24'(-4076);
			2455: out = 24'(-3020);
			2456: out = 24'(-43088);
			2457: out = 24'(-40720);
			2458: out = 24'(-2752);
			2459: out = 24'(46016);
			2460: out = 24'(29648);
			2461: out = 24'(55268);
			2462: out = 24'(90240);
			2463: out = 24'(45600);
			2464: out = 24'(-76752);
			2465: out = 24'(-130716);
			2466: out = 24'(-63504);
			2467: out = 24'(57600);
			2468: out = 24'(44752);
			2469: out = 24'(11688);
			2470: out = 24'(1060);
			2471: out = 24'(10032);
			2472: out = 24'(-25612);
			2473: out = 24'(-49904);
			2474: out = 24'(-25524);
			2475: out = 24'(34116);
			2476: out = 24'(9244);
			2477: out = 24'(9076);
			2478: out = 24'(-14620);
			2479: out = 24'(-20896);
			2480: out = 24'(-33328);
			2481: out = 24'(32664);
			2482: out = 24'(-14568);
			2483: out = 24'(-102196);
			2484: out = 24'(-89752);
			2485: out = 24'(-16304);
			2486: out = 24'(41560);
			2487: out = 24'(36084);
			2488: out = 24'(33080);
			2489: out = 24'(-60);
			2490: out = 24'(27652);
			2491: out = 24'(23096);
			2492: out = 24'(-16788);
			2493: out = 24'(-101376);
			2494: out = 24'(-28284);
			2495: out = 24'(38560);
			2496: out = 24'(17428);
			2497: out = 24'(-10184);
			2498: out = 24'(42132);
			2499: out = 24'(93524);
			2500: out = 24'(34180);
			2501: out = 24'(-101944);
			2502: out = 24'(-102104);
			2503: out = 24'(-5916);
			2504: out = 24'(48528);
			2505: out = 24'(-3524);
			2506: out = 24'(-32248);
			2507: out = 24'(-21336);
			2508: out = 24'(10444);
			2509: out = 24'(-10648);
			2510: out = 24'(9828);
			2511: out = 24'(16464);
			2512: out = 24'(76796);
			2513: out = 24'(100408);
			2514: out = 24'(69956);
			2515: out = 24'(-12348);
			2516: out = 24'(2492);
			2517: out = 24'(50692);
			2518: out = 24'(9580);
			2519: out = 24'(-75124);
			2520: out = 24'(-91160);
			2521: out = 24'(-35504);
			2522: out = 24'(-23984);
			2523: out = 24'(2060);
			2524: out = 24'(10696);
			2525: out = 24'(10920);
			2526: out = 24'(-14368);
			2527: out = 24'(6956);
			2528: out = 24'(-6220);
			2529: out = 24'(-41212);
			2530: out = 24'(-68424);
			2531: out = 24'(-16816);
			2532: out = 24'(34936);
			2533: out = 24'(53428);
			2534: out = 24'(49884);
			2535: out = 24'(58180);
			2536: out = 24'(38092);
			2537: out = 24'(7196);
			2538: out = 24'(-6272);
			2539: out = 24'(-3084);
			2540: out = 24'(-17676);
			2541: out = 24'(-73936);
			2542: out = 24'(-80960);
			2543: out = 24'(4860);
			2544: out = 24'(3624);
			2545: out = 24'(-21164);
			2546: out = 24'(-16300);
			2547: out = 24'(36252);
			2548: out = 24'(29708);
			2549: out = 24'(-10200);
			2550: out = 24'(-30472);
			2551: out = 24'(27988);
			2552: out = 24'(101372);
			2553: out = 24'(103160);
			2554: out = 24'(32792);
			2555: out = 24'(-63936);
			2556: out = 24'(-108804);
			2557: out = 24'(-90436);
			2558: out = 24'(4084);
			2559: out = 24'(72732);
			2560: out = 24'(72608);
			2561: out = 24'(50820);
			2562: out = 24'(23164);
			2563: out = 24'(-34048);
			2564: out = 24'(-93220);
			2565: out = 24'(7036);
			2566: out = 24'(80368);
			2567: out = 24'(22176);
			2568: out = 24'(-117672);
			2569: out = 24'(-116560);
			2570: out = 24'(-56972);
			2571: out = 24'(45840);
			2572: out = 24'(31344);
			2573: out = 24'(456);
			2574: out = 24'(-13924);
			2575: out = 24'(45524);
			2576: out = 24'(51392);
			2577: out = 24'(20944);
			2578: out = 24'(-81896);
			2579: out = 24'(9448);
			2580: out = 24'(119548);
			2581: out = 24'(65080);
			2582: out = 24'(-88736);
			2583: out = 24'(-76256);
			2584: out = 24'(63524);
			2585: out = 24'(98588);
			2586: out = 24'(-5152);
			2587: out = 24'(-97720);
			2588: out = 24'(-97492);
			2589: out = 24'(-20316);
			2590: out = 24'(11008);
			2591: out = 24'(33200);
			2592: out = 24'(6520);
			2593: out = 24'(-25036);
			2594: out = 24'(-43264);
			2595: out = 24'(-3964);
			2596: out = 24'(2532);
			2597: out = 24'(41108);
			2598: out = 24'(114592);
			2599: out = 24'(123244);
			2600: out = 24'(-2976);
			2601: out = 24'(-128316);
			2602: out = 24'(-97700);
			2603: out = 24'(-7500);
			2604: out = 24'(31156);
			2605: out = 24'(-7220);
			2606: out = 24'(-22788);
			2607: out = 24'(-32456);
			2608: out = 24'(62536);
			2609: out = 24'(97048);
			2610: out = 24'(53480);
			2611: out = 24'(-63088);
			2612: out = 24'(-44196);
			2613: out = 24'(-4436);
			2614: out = 24'(16344);
			2615: out = 24'(1100);
			2616: out = 24'(61480);
			2617: out = 24'(48512);
			2618: out = 24'(14848);
			2619: out = 24'(-1088);
			2620: out = 24'(536);
			2621: out = 24'(-9156);
			2622: out = 24'(9108);
			2623: out = 24'(43768);
			2624: out = 24'(14724);
			2625: out = 24'(-15556);
			2626: out = 24'(-4420);
			2627: out = 24'(49340);
			2628: out = 24'(59652);
			2629: out = 24'(29816);
			2630: out = 24'(-30956);
			2631: out = 24'(-85200);
			2632: out = 24'(-111248);
			2633: out = 24'(-103888);
			2634: out = 24'(-64160);
			2635: out = 24'(-29548);
			2636: out = 24'(-23708);
			2637: out = 24'(38544);
			2638: out = 24'(39188);
			2639: out = 24'(-18804);
			2640: out = 24'(-71116);
			2641: out = 24'(37760);
			2642: out = 24'(92040);
			2643: out = 24'(46272);
			2644: out = 24'(-49124);
			2645: out = 24'(-62496);
			2646: out = 24'(-43524);
			2647: out = 24'(-17920);
			2648: out = 24'(-22696);
			2649: out = 24'(-22120);
			2650: out = 24'(5272);
			2651: out = 24'(33340);
			2652: out = 24'(9712);
			2653: out = 24'(-64600);
			2654: out = 24'(-94544);
			2655: out = 24'(-52092);
			2656: out = 24'(29580);
			2657: out = 24'(51660);
			2658: out = 24'(43692);
			2659: out = 24'(-1524);
			2660: out = 24'(14388);
			2661: out = 24'(56612);
			2662: out = 24'(47728);
			2663: out = 24'(-3736);
			2664: out = 24'(6828);
			2665: out = 24'(63032);
			2666: out = 24'(61444);
			2667: out = 24'(-19120);
			2668: out = 24'(-42176);
			2669: out = 24'(25128);
			2670: out = 24'(48792);
			2671: out = 24'(8856);
			2672: out = 24'(-47540);
			2673: out = 24'(-17212);
			2674: out = 24'(72260);
			2675: out = 24'(80264);
			2676: out = 24'(32416);
			2677: out = 24'(-14744);
			2678: out = 24'(-10284);
			2679: out = 24'(5940);
			2680: out = 24'(10916);
			2681: out = 24'(-31328);
			2682: out = 24'(-59188);
			2683: out = 24'(20812);
			2684: out = 24'(66624);
			2685: out = 24'(42392);
			2686: out = 24'(-9900);
			2687: out = 24'(17236);
			2688: out = 24'(17184);
			2689: out = 24'(23932);
			2690: out = 24'(-5308);
			2691: out = 24'(-29140);
			2692: out = 24'(-46656);
			2693: out = 24'(1164);
			2694: out = 24'(20528);
			2695: out = 24'(-4592);
			2696: out = 24'(-38036);
			2697: out = 24'(6124);
			2698: out = 24'(23132);
			2699: out = 24'(-28720);
			2700: out = 24'(-53612);
			2701: out = 24'(-17004);
			2702: out = 24'(45140);
			2703: out = 24'(49280);
			2704: out = 24'(1976);
			2705: out = 24'(-32040);
			2706: out = 24'(-30748);
			2707: out = 24'(-9552);
			2708: out = 24'(-2548);
			2709: out = 24'(-16048);
			2710: out = 24'(-18292);
			2711: out = 24'(29020);
			2712: out = 24'(84412);
			2713: out = 24'(34708);
			2714: out = 24'(-10112);
			2715: out = 24'(-19528);
			2716: out = 24'(-8736);
			2717: out = 24'(-60324);
			2718: out = 24'(-87196);
			2719: out = 24'(-36896);
			2720: out = 24'(51576);
			2721: out = 24'(35248);
			2722: out = 24'(33944);
			2723: out = 24'(19164);
			2724: out = 24'(-432);
			2725: out = 24'(-83420);
			2726: out = 24'(-34436);
			2727: out = 24'(-19464);
			2728: out = 24'(-37236);
			2729: out = 24'(-62128);
			2730: out = 24'(-20484);
			2731: out = 24'(136);
			2732: out = 24'(7980);
			2733: out = 24'(18804);
			2734: out = 24'(5664);
			2735: out = 24'(11940);
			2736: out = 24'(28040);
			2737: out = 24'(38072);
			2738: out = 24'(-9980);
			2739: out = 24'(-3820);
			2740: out = 24'(4572);
			2741: out = 24'(-3724);
			2742: out = 24'(-39816);
			2743: out = 24'(-16164);
			2744: out = 24'(9732);
			2745: out = 24'(13884);
			2746: out = 24'(-5328);
			2747: out = 24'(-10624);
			2748: out = 24'(1592);
			2749: out = 24'(25736);
			2750: out = 24'(24784);
			2751: out = 24'(23124);
			2752: out = 24'(-22308);
			2753: out = 24'(-33456);
			2754: out = 24'(14352);
			2755: out = 24'(90908);
			2756: out = 24'(47772);
			2757: out = 24'(-14388);
			2758: out = 24'(-27436);
			2759: out = 24'(22592);
			2760: out = 24'(-17140);
			2761: out = 24'(-79640);
			2762: out = 24'(-92288);
			2763: out = 24'(6572);
			2764: out = 24'(82240);
			2765: out = 24'(107072);
			2766: out = 24'(40076);
			2767: out = 24'(-72012);
			2768: out = 24'(-123728);
			2769: out = 24'(-46752);
			2770: out = 24'(29796);
			2771: out = 24'(13752);
			2772: out = 24'(4416);
			2773: out = 24'(68924);
			2774: out = 24'(112512);
			2775: out = 24'(56892);
			2776: out = 24'(-63724);
			2777: out = 24'(-62160);
			2778: out = 24'(8296);
			2779: out = 24'(11556);
			2780: out = 24'(-47576);
			2781: out = 24'(-31724);
			2782: out = 24'(54780);
			2783: out = 24'(89432);
			2784: out = 24'(44032);
			2785: out = 24'(25824);
			2786: out = 24'(39304);
			2787: out = 24'(36236);
			2788: out = 24'(-8832);
			2789: out = 24'(-86656);
			2790: out = 24'(-97540);
			2791: out = 24'(-50016);
			2792: out = 24'(10344);
			2793: out = 24'(43672);
			2794: out = 24'(78988);
			2795: out = 24'(53700);
			2796: out = 24'(-2200);
			2797: out = 24'(-1960);
			2798: out = 24'(34440);
			2799: out = 24'(32008);
			2800: out = 24'(-16376);
			2801: out = 24'(-36012);
			2802: out = 24'(-26796);
			2803: out = 24'(-20096);
			2804: out = 24'(-40860);
			2805: out = 24'(-47468);
			2806: out = 24'(9472);
			2807: out = 24'(32380);
			2808: out = 24'(-3344);
			2809: out = 24'(-41468);
			2810: out = 24'(-10032);
			2811: out = 24'(17160);
			2812: out = 24'(16452);
			2813: out = 24'(16844);
			2814: out = 24'(21788);
			2815: out = 24'(13784);
			2816: out = 24'(-35776);
			2817: out = 24'(-71860);
			2818: out = 24'(-25700);
			2819: out = 24'(-22292);
			2820: out = 24'(-47448);
			2821: out = 24'(-37952);
			2822: out = 24'(41216);
			2823: out = 24'(44864);
			2824: out = 24'(9260);
			2825: out = 24'(-7332);
			2826: out = 24'(27076);
			2827: out = 24'(-12472);
			2828: out = 24'(-70968);
			2829: out = 24'(-79424);
			2830: out = 24'(17744);
			2831: out = 24'(31996);
			2832: out = 24'(42856);
			2833: out = 24'(7984);
			2834: out = 24'(-168);
			2835: out = 24'(-4556);
			2836: out = 24'(39936);
			2837: out = 24'(-5876);
			2838: out = 24'(-72432);
			2839: out = 24'(-54712);
			2840: out = 24'(12100);
			2841: out = 24'(22620);
			2842: out = 24'(-2144);
			2843: out = 24'(11576);
			2844: out = 24'(1656);
			2845: out = 24'(-6344);
			2846: out = 24'(-2392);
			2847: out = 24'(33840);
			2848: out = 24'(20640);
			2849: out = 24'(42588);
			2850: out = 24'(54716);
			2851: out = 24'(42244);
			2852: out = 24'(4556);
			2853: out = 24'(-59732);
			2854: out = 24'(-78804);
			2855: out = 24'(-21880);
			2856: out = 24'(35436);
			2857: out = 24'(45444);
			2858: out = 24'(35248);
			2859: out = 24'(48156);
			2860: out = 24'(54888);
			2861: out = 24'(14972);
			2862: out = 24'(-34484);
			2863: out = 24'(-32964);
			2864: out = 24'(-2512);
			2865: out = 24'(5164);
			2866: out = 24'(-54648);
			2867: out = 24'(-65692);
			2868: out = 24'(18680);
			2869: out = 24'(64896);
			2870: out = 24'(78028);
			2871: out = 24'(47628);
			2872: out = 24'(-5880);
			2873: out = 24'(-70804);
			2874: out = 24'(-97652);
			2875: out = 24'(-57808);
			2876: out = 24'(-9552);
			2877: out = 24'(-19028);
			2878: out = 24'(37364);
			2879: out = 24'(61544);
			2880: out = 24'(21348);
			2881: out = 24'(-46800);
			2882: out = 24'(-21168);
			2883: out = 24'(38840);
			2884: out = 24'(14096);
			2885: out = 24'(-73168);
			2886: out = 24'(-3796);
			2887: out = 24'(72284);
			2888: out = 24'(60552);
			2889: out = 24'(-23520);
			2890: out = 24'(-38780);
			2891: out = 24'(10688);
			2892: out = 24'(54420);
			2893: out = 24'(38496);
			2894: out = 24'(14300);
			2895: out = 24'(-380);
			2896: out = 24'(-23884);
			2897: out = 24'(-50608);
			2898: out = 24'(-32196);
			2899: out = 24'(13248);
			2900: out = 24'(45688);
			2901: out = 24'(42524);
			2902: out = 24'(21420);
			2903: out = 24'(3112);
			2904: out = 24'(-31204);
			2905: out = 24'(-41752);
			2906: out = 24'(-2932);
			2907: out = 24'(54276);
			2908: out = 24'(4608);
			2909: out = 24'(-60160);
			2910: out = 24'(-45616);
			2911: out = 24'(41712);
			2912: out = 24'(10552);
			2913: out = 24'(-62620);
			2914: out = 24'(-71544);
			2915: out = 24'(13872);
			2916: out = 24'(30228);
			2917: out = 24'(9700);
			2918: out = 24'(7892);
			2919: out = 24'(21960);
			2920: out = 24'(-15188);
			2921: out = 24'(-89124);
			2922: out = 24'(-87904);
			2923: out = 24'(17944);
			2924: out = 24'(57784);
			2925: out = 24'(45548);
			2926: out = 24'(4492);
			2927: out = 24'(-34968);
			2928: out = 24'(-44976);
			2929: out = 24'(-71784);
			2930: out = 24'(-39532);
			2931: out = 24'(19388);
			2932: out = 24'(55236);
			2933: out = 24'(21952);
			2934: out = 24'(38140);
			2935: out = 24'(37976);
			2936: out = 24'(-23720);
			2937: out = 24'(-104204);
			2938: out = 24'(-36092);
			2939: out = 24'(73984);
			2940: out = 24'(63296);
			2941: out = 24'(28236);
			2942: out = 24'(9008);
			2943: out = 24'(20560);
			2944: out = 24'(9792);
			2945: out = 24'(5412);
			2946: out = 24'(-25448);
			2947: out = 24'(-39276);
			2948: out = 24'(-23792);
			2949: out = 24'(27872);
			2950: out = 24'(69780);
			2951: out = 24'(66880);
			2952: out = 24'(30128);
			2953: out = 24'(-908);
			2954: out = 24'(-468);
			2955: out = 24'(-32644);
			2956: out = 24'(-80308);
			2957: out = 24'(-62916);
			2958: out = 24'(7556);
			2959: out = 24'(72112);
			2960: out = 24'(56180);
			2961: out = 24'(11236);
			2962: out = 24'(-2704);
			2963: out = 24'(12844);
			2964: out = 24'(-16256);
			2965: out = 24'(-70452);
			2966: out = 24'(-43432);
			2967: out = 24'(34128);
			2968: out = 24'(57412);
			2969: out = 24'(-9576);
			2970: out = 24'(-79812);
			2971: out = 24'(-31216);
			2972: out = 24'(50756);
			2973: out = 24'(37848);
			2974: out = 24'(-28056);
			2975: out = 24'(-110608);
			2976: out = 24'(-27412);
			2977: out = 24'(85664);
			2978: out = 24'(73536);
			2979: out = 24'(-62680);
			2980: out = 24'(-72036);
			2981: out = 24'(39616);
			2982: out = 24'(102732);
			2983: out = 24'(27860);
			2984: out = 24'(-23376);
			2985: out = 24'(-20312);
			2986: out = 24'(23704);
			2987: out = 24'(21312);
			2988: out = 24'(22692);
			2989: out = 24'(-15292);
			2990: out = 24'(-31096);
			2991: out = 24'(-1844);
			2992: out = 24'(-18472);
			2993: out = 24'(-75056);
			2994: out = 24'(-92100);
			2995: out = 24'(-3056);
			2996: out = 24'(10832);
			2997: out = 24'(14940);
			2998: out = 24'(-5504);
			2999: out = 24'(-9700);
			3000: out = 24'(-27996);
			3001: out = 24'(-13284);
			3002: out = 24'(-10616);
			3003: out = 24'(6876);
			3004: out = 24'(38100);
			3005: out = 24'(40984);
			3006: out = 24'(-11096);
			3007: out = 24'(-63176);
			3008: out = 24'(-70060);
			3009: out = 24'(920);
			3010: out = 24'(18392);
			3011: out = 24'(2692);
			3012: out = 24'(6896);
			3013: out = 24'(34456);
			3014: out = 24'(22296);
			3015: out = 24'(20220);
			3016: out = 24'(56280);
			3017: out = 24'(29932);
			3018: out = 24'(-13168);
			3019: out = 24'(-61552);
			3020: out = 24'(-69224);
			3021: out = 24'(-66188);
			3022: out = 24'(-5644);
			3023: out = 24'(54808);
			3024: out = 24'(99016);
			3025: out = 24'(117020);
			3026: out = 24'(77932);
			3027: out = 24'(26956);
			3028: out = 24'(-4676);
			3029: out = 24'(-524);
			3030: out = 24'(-44088);
			3031: out = 24'(-44492);
			3032: out = 24'(-16860);
			3033: out = 24'(10168);
			3034: out = 24'(45748);
			3035: out = 24'(72648);
			3036: out = 24'(77616);
			3037: out = 24'(48248);
			3038: out = 24'(2480);
			3039: out = 24'(-18984);
			3040: out = 24'(-12228);
			3041: out = 24'(-4124);
			3042: out = 24'(4080);
			3043: out = 24'(37388);
			3044: out = 24'(54176);
			3045: out = 24'(48);
			3046: out = 24'(-100392);
			3047: out = 24'(-63484);
			3048: out = 24'(46716);
			3049: out = 24'(70092);
			3050: out = 24'(-7392);
			3051: out = 24'(-32176);
			3052: out = 24'(21324);
			3053: out = 24'(45792);
			3054: out = 24'(-33952);
			3055: out = 24'(-39028);
			3056: out = 24'(-83668);
			3057: out = 24'(-97564);
			3058: out = 24'(-84116);
			3059: out = 24'(-3536);
			3060: out = 24'(20968);
			3061: out = 24'(36840);
			3062: out = 24'(35064);
			3063: out = 24'(13120);
			3064: out = 24'(-51180);
			3065: out = 24'(-102284);
			3066: out = 24'(-96760);
			3067: out = 24'(-19992);
			3068: out = 24'(51340);
			3069: out = 24'(65756);
			3070: out = 24'(18556);
			3071: out = 24'(-40164);
			3072: out = 24'(-17964);
			3073: out = 24'(9716);
			3074: out = 24'(15224);
			3075: out = 24'(16580);
			3076: out = 24'(59520);
			3077: out = 24'(27140);
			3078: out = 24'(-49316);
			3079: out = 24'(-101852);
			3080: out = 24'(-29396);
			3081: out = 24'(-2220);
			3082: out = 24'(3620);
			3083: out = 24'(19964);
			3084: out = 24'(77356);
			3085: out = 24'(66700);
			3086: out = 24'(32000);
			3087: out = 24'(-13560);
			3088: out = 24'(-26124);
			3089: out = 24'(-45236);
			3090: out = 24'(-13620);
			3091: out = 24'(25756);
			3092: out = 24'(52736);
			3093: out = 24'(26920);
			3094: out = 24'(21924);
			3095: out = 24'(-9368);
			3096: out = 24'(-50724);
			3097: out = 24'(-72480);
			3098: out = 24'(-16808);
			3099: out = 24'(36756);
			3100: out = 24'(49820);
			3101: out = 24'(26692);
			3102: out = 24'(30432);
			3103: out = 24'(-6448);
			3104: out = 24'(-62908);
			3105: out = 24'(-95228);
			3106: out = 24'(-48796);
			3107: out = 24'(-4124);
			3108: out = 24'(21444);
			3109: out = 24'(41496);
			3110: out = 24'(82564);
			3111: out = 24'(43476);
			3112: out = 24'(-3328);
			3113: out = 24'(-8852);
			3114: out = 24'(11152);
			3115: out = 24'(7492);
			3116: out = 24'(-7300);
			3117: out = 24'(-1748);
			3118: out = 24'(12908);
			3119: out = 24'(25652);
			3120: out = 24'(29304);
			3121: out = 24'(29252);
			3122: out = 24'(676);
			3123: out = 24'(-8768);
			3124: out = 24'(-36272);
			3125: out = 24'(-41724);
			3126: out = 24'(-25536);
			3127: out = 24'(43488);
			3128: out = 24'(60772);
			3129: out = 24'(69056);
			3130: out = 24'(43440);
			3131: out = 24'(-30972);
			3132: out = 24'(-82428);
			3133: out = 24'(-22820);
			3134: out = 24'(63824);
			3135: out = 24'(76440);
			3136: out = 24'(-7796);
			3137: out = 24'(-13096);
			3138: out = 24'(27188);
			3139: out = 24'(8088);
			3140: out = 24'(-68180);
			3141: out = 24'(-44780);
			3142: out = 24'(25476);
			3143: out = 24'(2996);
			3144: out = 24'(-45884);
			3145: out = 24'(-35620);
			3146: out = 24'(21104);
			3147: out = 24'(24820);
			3148: out = 24'(6564);
			3149: out = 24'(-31308);
			3150: out = 24'(-52340);
			3151: out = 24'(-41964);
			3152: out = 24'(8112);
			3153: out = 24'(47728);
			3154: out = 24'(10636);
			3155: out = 24'(-63420);
			3156: out = 24'(-63712);
			3157: out = 24'(-50680);
			3158: out = 24'(-47256);
			3159: out = 24'(-46032);
			3160: out = 24'(19752);
			3161: out = 24'(84248);
			3162: out = 24'(66880);
			3163: out = 24'(-40960);
			3164: out = 24'(-112684);
			3165: out = 24'(-82992);
			3166: out = 24'(17096);
			3167: out = 24'(42816);
			3168: out = 24'(-704);
			3169: out = 24'(-5708);
			3170: out = 24'(-1500);
			3171: out = 24'(12064);
			3172: out = 24'(3496);
			3173: out = 24'(-42512);
			3174: out = 24'(-59668);
			3175: out = 24'(-40940);
			3176: out = 24'(11292);
			3177: out = 24'(49836);
			3178: out = 24'(82284);
			3179: out = 24'(59072);
			3180: out = 24'(26140);
			3181: out = 24'(1772);
			3182: out = 24'(-6472);
			3183: out = 24'(-17960);
			3184: out = 24'(17532);
			3185: out = 24'(67460);
			3186: out = 24'(23596);
			3187: out = 24'(-34492);
			3188: out = 24'(-42432);
			3189: out = 24'(18340);
			3190: out = 24'(64116);
			3191: out = 24'(25984);
			3192: out = 24'(-12776);
			3193: out = 24'(-3836);
			3194: out = 24'(25164);
			3195: out = 24'(-12304);
			3196: out = 24'(-23104);
			3197: out = 24'(22836);
			3198: out = 24'(63064);
			3199: out = 24'(16124);
			3200: out = 24'(-7984);
			3201: out = 24'(16152);
			3202: out = 24'(34360);
			3203: out = 24'(25856);
			3204: out = 24'(4252);
			3205: out = 24'(18328);
			3206: out = 24'(28812);
			3207: out = 24'(-21044);
			3208: out = 24'(-75116);
			3209: out = 24'(-39928);
			3210: out = 24'(65444);
			3211: out = 24'(90992);
			3212: out = 24'(49296);
			3213: out = 24'(-5292);
			3214: out = 24'(-13236);
			3215: out = 24'(-8988);
			3216: out = 24'(-60404);
			3217: out = 24'(-115688);
			3218: out = 24'(-78204);
			3219: out = 24'(37028);
			3220: out = 24'(91532);
			3221: out = 24'(59412);
			3222: out = 24'(19488);
			3223: out = 24'(9988);
			3224: out = 24'(-13500);
			3225: out = 24'(-22380);
			3226: out = 24'(13476);
			3227: out = 24'(65744);
			3228: out = 24'(22652);
			3229: out = 24'(4264);
			3230: out = 24'(-7216);
			3231: out = 24'(-17504);
			3232: out = 24'(-111120);
			3233: out = 24'(-34684);
			3234: out = 24'(17260);
			3235: out = 24'(-8588);
			3236: out = 24'(-78640);
			3237: out = 24'(-34288);
			3238: out = 24'(27240);
			3239: out = 24'(31580);
			3240: out = 24'(-26664);
			3241: out = 24'(-52036);
			3242: out = 24'(-36908);
			3243: out = 24'(2212);
			3244: out = 24'(3716);
			3245: out = 24'(-12352);
			3246: out = 24'(4300);
			3247: out = 24'(61260);
			3248: out = 24'(56624);
			3249: out = 24'(-52316);
			3250: out = 24'(-104396);
			3251: out = 24'(-37832);
			3252: out = 24'(37008);
			3253: out = 24'(-12204);
			3254: out = 24'(7740);
			3255: out = 24'(35480);
			3256: out = 24'(-4892);
			3257: out = 24'(-114084);
			3258: out = 24'(-119704);
			3259: out = 24'(-59932);
			3260: out = 24'(50396);
			3261: out = 24'(66208);
			3262: out = 24'(47572);
			3263: out = 24'(-80);
			3264: out = 24'(-21076);
			3265: out = 24'(-12188);
			3266: out = 24'(8840);
			3267: out = 24'(6668);
			3268: out = 24'(-25212);
			3269: out = 24'(-35628);
			3270: out = 24'(25384);
			3271: out = 24'(95404);
			3272: out = 24'(91572);
			3273: out = 24'(35812);
			3274: out = 24'(-10424);
			3275: out = 24'(-3556);
			3276: out = 24'(23712);
			3277: out = 24'(43776);
			3278: out = 24'(25916);
			3279: out = 24'(17428);
			3280: out = 24'(-65824);
			3281: out = 24'(-106180);
			3282: out = 24'(-50588);
			3283: out = 24'(39840);
			3284: out = 24'(33840);
			3285: out = 24'(29616);
			3286: out = 24'(45648);
			3287: out = 24'(14440);
			3288: out = 24'(-32680);
			3289: out = 24'(-44648);
			3290: out = 24'(-12744);
			3291: out = 24'(-15648);
			3292: out = 24'(12840);
			3293: out = 24'(12240);
			3294: out = 24'(-14864);
			3295: out = 24'(-59324);
			3296: out = 24'(17940);
			3297: out = 24'(91832);
			3298: out = 24'(84228);
			3299: out = 24'(-16104);
			3300: out = 24'(-52860);
			3301: out = 24'(-60212);
			3302: out = 24'(188);
			3303: out = 24'(36596);
			3304: out = 24'(72944);
			3305: out = 24'(3216);
			3306: out = 24'(-10452);
			3307: out = 24'(-7364);
			3308: out = 24'(-24860);
			3309: out = 24'(-72996);
			3310: out = 24'(-3680);
			3311: out = 24'(80892);
			3312: out = 24'(47348);
			3313: out = 24'(-5692);
			3314: out = 24'(-17984);
			3315: out = 24'(6160);
			3316: out = 24'(-8296);
			3317: out = 24'(-77656);
			3318: out = 24'(-45516);
			3319: out = 24'(46132);
			3320: out = 24'(69268);
			3321: out = 24'(22420);
			3322: out = 24'(-39812);
			3323: out = 24'(-54092);
			3324: out = 24'(-10128);
			3325: out = 24'(52464);
			3326: out = 24'(25868);
			3327: out = 24'(-32508);
			3328: out = 24'(-63584);
			3329: out = 24'(-27244);
			3330: out = 24'(-26700);
			3331: out = 24'(-18920);
			3332: out = 24'(21028);
			3333: out = 24'(71224);
			3334: out = 24'(-4732);
			3335: out = 24'(-56252);
			3336: out = 24'(-25268);
			3337: out = 24'(85176);
			3338: out = 24'(80580);
			3339: out = 24'(68584);
			3340: out = 24'(-260);
			3341: out = 24'(-62384);
			3342: out = 24'(-118456);
			3343: out = 24'(-64592);
			3344: out = 24'(-34332);
			3345: out = 24'(-9132);
			3346: out = 24'(48812);
			3347: out = 24'(107060);
			3348: out = 24'(70248);
			3349: out = 24'(9888);
			3350: out = 24'(-15376);
			3351: out = 24'(-17480);
			3352: out = 24'(-67564);
			3353: out = 24'(-85324);
			3354: out = 24'(-7448);
			3355: out = 24'(23420);
			3356: out = 24'(16100);
			3357: out = 24'(7908);
			3358: out = 24'(49052);
			3359: out = 24'(78068);
			3360: out = 24'(49340);
			3361: out = 24'(-1608);
			3362: out = 24'(-23488);
			3363: out = 24'(-38876);
			3364: out = 24'(-12368);
			3365: out = 24'(-10480);
			3366: out = 24'(-11812);
			3367: out = 24'(468);
			3368: out = 24'(-260);
			3369: out = 24'(23156);
			3370: out = 24'(59688);
			3371: out = 24'(60364);
			3372: out = 24'(-18512);
			3373: out = 24'(-75332);
			3374: out = 24'(-56816);
			3375: out = 24'(4248);
			3376: out = 24'(1744);
			3377: out = 24'(8560);
			3378: out = 24'(29672);
			3379: out = 24'(41868);
			3380: out = 24'(27288);
			3381: out = 24'(-54140);
			3382: out = 24'(-68576);
			3383: out = 24'(7204);
			3384: out = 24'(53648);
			3385: out = 24'(13940);
			3386: out = 24'(-37308);
			3387: out = 24'(-20100);
			3388: out = 24'(38268);
			3389: out = 24'(25972);
			3390: out = 24'(4556);
			3391: out = 24'(1024);
			3392: out = 24'(-9216);
			3393: out = 24'(-53168);
			3394: out = 24'(-96696);
			3395: out = 24'(-42544);
			3396: out = 24'(78104);
			3397: out = 24'(97800);
			3398: out = 24'(67720);
			3399: out = 24'(4136);
			3400: out = 24'(-50232);
			3401: out = 24'(-103604);
			3402: out = 24'(-29664);
			3403: out = 24'(29328);
			3404: out = 24'(22904);
			3405: out = 24'(-3480);
			3406: out = 24'(-28524);
			3407: out = 24'(14736);
			3408: out = 24'(52336);
			3409: out = 24'(39824);
			3410: out = 24'(4908);
			3411: out = 24'(-932);
			3412: out = 24'(-10428);
			3413: out = 24'(-35540);
			3414: out = 24'(-864);
			3415: out = 24'(7264);
			3416: out = 24'(-2448);
			3417: out = 24'(-25700);
			3418: out = 24'(-33248);
			3419: out = 24'(-9520);
			3420: out = 24'(24668);
			3421: out = 24'(54360);
			3422: out = 24'(60872);
			3423: out = 24'(18568);
			3424: out = 24'(-67860);
			3425: out = 24'(-101328);
			3426: out = 24'(-4044);
			3427: out = 24'(40336);
			3428: out = 24'(34444);
			3429: out = 24'(-13608);
			3430: out = 24'(-28396);
			3431: out = 24'(-20776);
			3432: out = 24'(55232);
			3433: out = 24'(89608);
			3434: out = 24'(68060);
			3435: out = 24'(628);
			3436: out = 24'(-52268);
			3437: out = 24'(-96360);
			3438: out = 24'(-78976);
			3439: out = 24'(4236);
			3440: out = 24'(75464);
			3441: out = 24'(35860);
			3442: out = 24'(-42444);
			3443: out = 24'(-57236);
			3444: out = 24'(12548);
			3445: out = 24'(64296);
			3446: out = 24'(69976);
			3447: out = 24'(59264);
			3448: out = 24'(-7396);
			3449: out = 24'(-30484);
			3450: out = 24'(-20668);
			3451: out = 24'(-4400);
			3452: out = 24'(-27020);
			3453: out = 24'(-5768);
			3454: out = 24'(51988);
			3455: out = 24'(78288);
			3456: out = 24'(-1556);
			3457: out = 24'(-4908);
			3458: out = 24'(-1328);
			3459: out = 24'(-22944);
			3460: out = 24'(-97868);
			3461: out = 24'(-45128);
			3462: out = 24'(51560);
			3463: out = 24'(99192);
			3464: out = 24'(42008);
			3465: out = 24'(-48184);
			3466: out = 24'(-115248);
			3467: out = 24'(-74564);
			3468: out = 24'(15460);
			3469: out = 24'(43748);
			3470: out = 24'(36132);
			3471: out = 24'(30004);
			3472: out = 24'(3196);
			3473: out = 24'(-73352);
			3474: out = 24'(-121672);
			3475: out = 24'(-57600);
			3476: out = 24'(53156);
			3477: out = 24'(37976);
			3478: out = 24'(-8956);
			3479: out = 24'(-54148);
			3480: out = 24'(-22580);
			3481: out = 24'(35728);
			3482: out = 24'(82708);
			3483: out = 24'(41980);
			3484: out = 24'(-11728);
			3485: out = 24'(-50652);
			3486: out = 24'(-110728);
			3487: out = 24'(-100284);
			3488: out = 24'(-22328);
			3489: out = 24'(59052);
			3490: out = 24'(62880);
			3491: out = 24'(55192);
			3492: out = 24'(40108);
			3493: out = 24'(31108);
			3494: out = 24'(5928);
			3495: out = 24'(-16900);
			3496: out = 24'(-36556);
			3497: out = 24'(-21448);
			3498: out = 24'(15068);
			3499: out = 24'(24384);
			3500: out = 24'(-7332);
			3501: out = 24'(-45568);
			3502: out = 24'(-50364);
			3503: out = 24'(-5856);
			3504: out = 24'(37500);
			3505: out = 24'(58452);
			3506: out = 24'(53076);
			3507: out = 24'(37108);
			3508: out = 24'(8424);
			3509: out = 24'(1504);
			3510: out = 24'(-6828);
			3511: out = 24'(-100480);
			3512: out = 24'(-52276);
			3513: out = 24'(38692);
			3514: out = 24'(82924);
			3515: out = 24'(41780);
			3516: out = 24'(46776);
			3517: out = 24'(30352);
			3518: out = 24'(12396);
			3519: out = 24'(-3524);
			3520: out = 24'(-14360);
			3521: out = 24'(-8224);
			3522: out = 24'(228);
			3523: out = 24'(-13228);
			3524: out = 24'(-25336);
			3525: out = 24'(11780);
			3526: out = 24'(69336);
			3527: out = 24'(59748);
			3528: out = 24'(28632);
			3529: out = 24'(-82652);
			3530: out = 24'(-75512);
			3531: out = 24'(21732);
			3532: out = 24'(61200);
			3533: out = 24'(13980);
			3534: out = 24'(-7208);
			3535: out = 24'(-30120);
			3536: out = 24'(-107332);
			3537: out = 24'(-122044);
			3538: out = 24'(-24108);
			3539: out = 24'(104504);
			3540: out = 24'(107212);
			3541: out = 24'(48940);
			3542: out = 24'(-31328);
			3543: out = 24'(-65580);
			3544: out = 24'(-50984);
			3545: out = 24'(232);
			3546: out = 24'(40124);
			3547: out = 24'(41752);
			3548: out = 24'(11048);
			3549: out = 24'(-6396);
			3550: out = 24'(-79616);
			3551: out = 24'(-121884);
			3552: out = 24'(-82004);
			3553: out = 24'(23268);
			3554: out = 24'(66476);
			3555: out = 24'(42740);
			3556: out = 24'(9448);
			3557: out = 24'(9284);
			3558: out = 24'(-14800);
			3559: out = 24'(-43732);
			3560: out = 24'(-36660);
			3561: out = 24'(35288);
			3562: out = 24'(44344);
			3563: out = 24'(41088);
			3564: out = 24'(-11600);
			3565: out = 24'(-44684);
			3566: out = 24'(-24448);
			3567: out = 24'(12820);
			3568: out = 24'(-2116);
			3569: out = 24'(-27296);
			3570: out = 24'(-28264);
			3571: out = 24'(-24864);
			3572: out = 24'(-73424);
			3573: out = 24'(-89684);
			3574: out = 24'(15716);
			3575: out = 24'(95052);
			3576: out = 24'(92632);
			3577: out = 24'(31876);
			3578: out = 24'(-28732);
			3579: out = 24'(-43648);
			3580: out = 24'(-47120);
			3581: out = 24'(-6636);
			3582: out = 24'(59172);
			3583: out = 24'(76996);
			3584: out = 24'(11140);
			3585: out = 24'(-55824);
			3586: out = 24'(-63524);
			3587: out = 24'(-34232);
			3588: out = 24'(22376);
			3589: out = 24'(50820);
			3590: out = 24'(46660);
			3591: out = 24'(22660);
			3592: out = 24'(-6016);
			3593: out = 24'(-13792);
			3594: out = 24'(-8708);
			3595: out = 24'(3176);
			3596: out = 24'(-19140);
			3597: out = 24'(41280);
			3598: out = 24'(93824);
			3599: out = 24'(73888);
			3600: out = 24'(15300);
			3601: out = 24'(-50444);
			3602: out = 24'(-79368);
			3603: out = 24'(-50200);
			3604: out = 24'(10108);
			3605: out = 24'(56636);
			3606: out = 24'(42432);
			3607: out = 24'(8584);
			3608: out = 24'(10540);
			3609: out = 24'(40636);
			3610: out = 24'(47060);
			3611: out = 24'(28332);
			3612: out = 24'(7356);
			3613: out = 24'(-59956);
			3614: out = 24'(-102880);
			3615: out = 24'(-86420);
			3616: out = 24'(-8848);
			3617: out = 24'(43276);
			3618: out = 24'(70256);
			3619: out = 24'(55712);
			3620: out = 24'(2328);
			3621: out = 24'(-63264);
			3622: out = 24'(-109796);
			3623: out = 24'(-61228);
			3624: out = 24'(40040);
			3625: out = 24'(68168);
			3626: out = 24'(52112);
			3627: out = 24'(22392);
			3628: out = 24'(12936);
			3629: out = 24'(-3228);
			3630: out = 24'(-30876);
			3631: out = 24'(-61596);
			3632: out = 24'(-45968);
			3633: out = 24'(2244);
			3634: out = 24'(-14808);
			3635: out = 24'(-25172);
			3636: out = 24'(-13148);
			3637: out = 24'(11280);
			3638: out = 24'(5064);
			3639: out = 24'(-9808);
			3640: out = 24'(-19740);
			3641: out = 24'(-14300);
			3642: out = 24'(-3968);
			3643: out = 24'(-18336);
			3644: out = 24'(-3808);
			3645: out = 24'(50672);
			3646: out = 24'(72332);
			3647: out = 24'(52860);
			3648: out = 24'(-33804);
			3649: out = 24'(-78004);
			3650: out = 24'(2600);
			3651: out = 24'(11708);
			3652: out = 24'(13828);
			3653: out = 24'(-360);
			3654: out = 24'(5148);
			3655: out = 24'(-39220);
			3656: out = 24'(16196);
			3657: out = 24'(64908);
			3658: out = 24'(55756);
			3659: out = 24'(-20236);
			3660: out = 24'(-16188);
			3661: out = 24'(5560);
			3662: out = 24'(-844);
			3663: out = 24'(-51936);
			3664: out = 24'(592);
			3665: out = 24'(46920);
			3666: out = 24'(30312);
			3667: out = 24'(-48456);
			3668: out = 24'(-56756);
			3669: out = 24'(-736);
			3670: out = 24'(79136);
			3671: out = 24'(72832);
			3672: out = 24'(22404);
			3673: out = 24'(-52400);
			3674: out = 24'(-1392);
			3675: out = 24'(93356);
			3676: out = 24'(45000);
			3677: out = 24'(-62140);
			3678: out = 24'(-87708);
			3679: out = 24'(-7340);
			3680: out = 24'(-3752);
			3681: out = 24'(2344);
			3682: out = 24'(31028);
			3683: out = 24'(72672);
			3684: out = 24'(54636);
			3685: out = 24'(-7856);
			3686: out = 24'(-44460);
			3687: out = 24'(-40708);
			3688: out = 24'(-33640);
			3689: out = 24'(-7828);
			3690: out = 24'(37400);
			3691: out = 24'(45072);
			3692: out = 24'(4684);
			3693: out = 24'(18476);
			3694: out = 24'(33648);
			3695: out = 24'(17724);
			3696: out = 24'(-29076);
			3697: out = 24'(-36128);
			3698: out = 24'(-16616);
			3699: out = 24'(-22504);
			3700: out = 24'(-51976);
			3701: out = 24'(-25716);
			3702: out = 24'(9492);
			3703: out = 24'(16948);
			3704: out = 24'(932);
			3705: out = 24'(24200);
			3706: out = 24'(2664);
			3707: out = 24'(-9044);
			3708: out = 24'(-29084);
			3709: out = 24'(-31020);
			3710: out = 24'(-5672);
			3711: out = 24'(25024);
			3712: out = 24'(31240);
			3713: out = 24'(16928);
			3714: out = 24'(2188);
			3715: out = 24'(-48736);
			3716: out = 24'(-73828);
			3717: out = 24'(-18404);
			3718: out = 24'(52852);
			3719: out = 24'(52672);
			3720: out = 24'(-13268);
			3721: out = 24'(-32560);
			3722: out = 24'(42204);
			3723: out = 24'(48668);
			3724: out = 24'(-31868);
			3725: out = 24'(-102156);
			3726: out = 24'(-48928);
			3727: out = 24'(-9648);
			3728: out = 24'(7964);
			3729: out = 24'(10804);
			3730: out = 24'(38240);
			3731: out = 24'(9668);
			3732: out = 24'(17748);
			3733: out = 24'(33456);
			3734: out = 24'(49936);
			3735: out = 24'(19584);
			3736: out = 24'(-16012);
			3737: out = 24'(-61312);
			3738: out = 24'(-82428);
			3739: out = 24'(-79232);
			3740: out = 24'(7728);
			3741: out = 24'(79748);
			3742: out = 24'(95216);
			3743: out = 24'(47728);
			3744: out = 24'(-15148);
			3745: out = 24'(-67752);
			3746: out = 24'(-51732);
			3747: out = 24'(1412);
			3748: out = 24'(-19808);
			3749: out = 24'(-54504);
			3750: out = 24'(-36564);
			3751: out = 24'(33540);
			3752: out = 24'(32612);
			3753: out = 24'(29768);
			3754: out = 24'(25012);
			3755: out = 24'(35248);
			3756: out = 24'(6472);
			3757: out = 24'(21776);
			3758: out = 24'(14776);
			3759: out = 24'(1424);
			3760: out = 24'(-37164);
			3761: out = 24'(-2788);
			3762: out = 24'(-14628);
			3763: out = 24'(-21956);
			3764: out = 24'(7200);
			3765: out = 24'(70840);
			3766: out = 24'(57276);
			3767: out = 24'(32520);
			3768: out = 24'(44864);
			3769: out = 24'(82984);
			3770: out = 24'(19400);
			3771: out = 24'(-72776);
			3772: out = 24'(-110312);
			3773: out = 24'(-65296);
			3774: out = 24'(-9656);
			3775: out = 24'(33560);
			3776: out = 24'(58088);
			3777: out = 24'(45228);
			3778: out = 24'(5792);
			3779: out = 24'(-26628);
			3780: out = 24'(-24012);
			3781: out = 24'(-8984);
			3782: out = 24'(17656);
			3783: out = 24'(-2404);
			3784: out = 24'(-41228);
			3785: out = 24'(-72744);
			3786: out = 24'(-25836);
			3787: out = 24'(-7416);
			3788: out = 24'(19740);
			3789: out = 24'(45844);
			3790: out = 24'(20900);
			3791: out = 24'(-21528);
			3792: out = 24'(-62908);
			3793: out = 24'(-63116);
			3794: out = 24'(-13208);
			3795: out = 24'(16480);
			3796: out = 24'(26712);
			3797: out = 24'(14328);
			3798: out = 24'(-12700);
			3799: out = 24'(-42748);
			3800: out = 24'(-33844);
			3801: out = 24'(-17356);
			3802: out = 24'(-31556);
			3803: out = 24'(20856);
			3804: out = 24'(29692);
			3805: out = 24'(25536);
			3806: out = 24'(11552);
			3807: out = 24'(70476);
			3808: out = 24'(-27672);
			3809: out = 24'(-116300);
			3810: out = 24'(-107012);
			3811: out = 24'(11488);
			3812: out = 24'(84864);
			3813: out = 24'(50364);
			3814: out = 24'(-11344);
			3815: out = 24'(-25008);
			3816: out = 24'(-3260);
			3817: out = 24'(49448);
			3818: out = 24'(69636);
			3819: out = 24'(54104);
			3820: out = 24'(-3752);
			3821: out = 24'(-17608);
			3822: out = 24'(-31176);
			3823: out = 24'(-52716);
			3824: out = 24'(-23980);
			3825: out = 24'(53676);
			3826: out = 24'(86052);
			3827: out = 24'(50172);
			3828: out = 24'(26224);
			3829: out = 24'(29992);
			3830: out = 24'(28100);
			3831: out = 24'(-16436);
			3832: out = 24'(-36932);
			3833: out = 24'(-69492);
			3834: out = 24'(-15960);
			3835: out = 24'(53332);
			3836: out = 24'(76152);
			3837: out = 24'(-26852);
			3838: out = 24'(-43392);
			3839: out = 24'(18292);
			3840: out = 24'(59068);
			3841: out = 24'(-15716);
			3842: out = 24'(-21644);
			3843: out = 24'(28952);
			3844: out = 24'(47836);
			3845: out = 24'(-40000);
			3846: out = 24'(-75424);
			3847: out = 24'(-42604);
			3848: out = 24'(23660);
			3849: out = 24'(62876);
			3850: out = 24'(29588);
			3851: out = 24'(-8436);
			3852: out = 24'(-17776);
			3853: out = 24'(7652);
			3854: out = 24'(-368);
			3855: out = 24'(2612);
			3856: out = 24'(11916);
			3857: out = 24'(22272);
			3858: out = 24'(-53836);
			3859: out = 24'(-48704);
			3860: out = 24'(11352);
			3861: out = 24'(63564);
			3862: out = 24'(53012);
			3863: out = 24'(33780);
			3864: out = 24'(-5084);
			3865: out = 24'(-30776);
			3866: out = 24'(-32864);
			3867: out = 24'(21392);
			3868: out = 24'(32444);
			3869: out = 24'(14864);
			3870: out = 24'(10276);
			3871: out = 24'(3788);
			3872: out = 24'(-41704);
			3873: out = 24'(-69040);
			3874: out = 24'(-12000);
			3875: out = 24'(-3984);
			3876: out = 24'(-8556);
			3877: out = 24'(-6464);
			3878: out = 24'(22548);
			3879: out = 24'(20004);
			3880: out = 24'(-14612);
			3881: out = 24'(-32324);
			3882: out = 24'(7216);
			3883: out = 24'(1252);
			3884: out = 24'(-23464);
			3885: out = 24'(-87608);
			3886: out = 24'(-99856);
			3887: out = 24'(-11248);
			3888: out = 24'(70968);
			3889: out = 24'(68160);
			3890: out = 24'(24572);
			3891: out = 24'(-12980);
			3892: out = 24'(-30632);
			3893: out = 24'(-38640);
			3894: out = 24'(-19828);
			3895: out = 24'(17592);
			3896: out = 24'(34576);
			3897: out = 24'(9440);
			3898: out = 24'(-972);
			3899: out = 24'(22568);
			3900: out = 24'(-5256);
			3901: out = 24'(-13312);
			3902: out = 24'(5408);
			3903: out = 24'(43288);
			3904: out = 24'(17152);
			3905: out = 24'(14920);
			3906: out = 24'(-11252);
			3907: out = 24'(-29848);
			3908: out = 24'(-27360);
			3909: out = 24'(15552);
			3910: out = 24'(32376);
			3911: out = 24'(12780);
			3912: out = 24'(-28364);
			3913: out = 24'(-10952);
			3914: out = 24'(-836);
			3915: out = 24'(1396);
			3916: out = 24'(2832);
			3917: out = 24'(41264);
			3918: out = 24'(23344);
			3919: out = 24'(-6292);
			3920: out = 24'(-6212);
			3921: out = 24'(49968);
			3922: out = 24'(37044);
			3923: out = 24'(8788);
			3924: out = 24'(5032);
			3925: out = 24'(33988);
			3926: out = 24'(24508);
			3927: out = 24'(-11056);
			3928: out = 24'(-41872);
			3929: out = 24'(-20732);
			3930: out = 24'(-21276);
			3931: out = 24'(-1656);
			3932: out = 24'(5228);
			3933: out = 24'(9140);
			3934: out = 24'(24404);
			3935: out = 24'(36964);
			3936: out = 24'(-5628);
			3937: out = 24'(-80616);
			3938: out = 24'(-61248);
			3939: out = 24'(-27312);
			3940: out = 24'(19960);
			3941: out = 24'(66560);
			3942: out = 24'(86340);
			3943: out = 24'(54104);
			3944: out = 24'(-39416);
			3945: out = 24'(-103772);
			3946: out = 24'(-28832);
			3947: out = 24'(39212);
			3948: out = 24'(19940);
			3949: out = 24'(-57868);
			3950: out = 24'(-83528);
			3951: out = 24'(-71556);
			3952: out = 24'(-7188);
			3953: out = 24'(44924);
			3954: out = 24'(86900);
			3955: out = 24'(67084);
			3956: out = 24'(31232);
			3957: out = 24'(-46484);
			3958: out = 24'(-82256);
			3959: out = 24'(-40816);
			3960: out = 24'(39916);
			3961: out = 24'(5840);
			3962: out = 24'(-57388);
			3963: out = 24'(-4972);
			3964: out = 24'(70968);
			3965: out = 24'(51612);
			3966: out = 24'(-24048);
			3967: out = 24'(-42260);
			3968: out = 24'(25512);
			3969: out = 24'(20648);
			3970: out = 24'(-55816);
			3971: out = 24'(-84584);
			3972: out = 24'(4716);
			3973: out = 24'(51656);
			3974: out = 24'(-7228);
			3975: out = 24'(-88132);
			3976: out = 24'(-47024);
			3977: out = 24'(6224);
			3978: out = 24'(21712);
			3979: out = 24'(-3732);
			3980: out = 24'(-13504);
			3981: out = 24'(-13276);
			3982: out = 24'(33884);
			3983: out = 24'(74012);
			3984: out = 24'(57344);
			3985: out = 24'(14972);
			3986: out = 24'(-26872);
			3987: out = 24'(-52888);
			3988: out = 24'(-81032);
			3989: out = 24'(-46120);
			3990: out = 24'(-15280);
			3991: out = 24'(23548);
			3992: out = 24'(36836);
			3993: out = 24'(10824);
			3994: out = 24'(-32372);
			3995: out = 24'(-6912);
			3996: out = 24'(63824);
			3997: out = 24'(63744);
			3998: out = 24'(5680);
			3999: out = 24'(-55532);
			4000: out = 24'(-43712);
			4001: out = 24'(31520);
			4002: out = 24'(18456);
			4003: out = 24'(1916);
			4004: out = 24'(31696);
			4005: out = 24'(80740);
			4006: out = 24'(57156);
			4007: out = 24'(3436);
			4008: out = 24'(-44604);
			4009: out = 24'(-55832);
			4010: out = 24'(-40368);
			4011: out = 24'(848);
			4012: out = 24'(36432);
			4013: out = 24'(38140);
			4014: out = 24'(-2116);
			4015: out = 24'(-16368);
			4016: out = 24'(1336);
			4017: out = 24'(25208);
			4018: out = 24'(38836);
			4019: out = 24'(49048);
			4020: out = 24'(48728);
			4021: out = 24'(524);
			4022: out = 24'(-88464);
			4023: out = 24'(-106984);
			4024: out = 24'(-35004);
			4025: out = 24'(41660);
			4026: out = 24'(51404);
			4027: out = 24'(13188);
			4028: out = 24'(33892);
			4029: out = 24'(50540);
			4030: out = 24'(7320);
			4031: out = 24'(-8380);
			4032: out = 24'(-32392);
			4033: out = 24'(-15544);
			4034: out = 24'(9860);
			4035: out = 24'(37072);
			4036: out = 24'(8076);
			4037: out = 24'(-11892);
			4038: out = 24'(-14188);
			4039: out = 24'(-544);
			4040: out = 24'(-1188);
			4041: out = 24'(-10304);
			4042: out = 24'(-27028);
			4043: out = 24'(-17620);
			4044: out = 24'(-9160);
			4045: out = 24'(10952);
			4046: out = 24'(-17372);
			4047: out = 24'(-62112);
			4048: out = 24'(-42872);
			4049: out = 24'(30508);
			4050: out = 24'(40276);
			4051: out = 24'(-20436);
			4052: out = 24'(-57644);
			4053: out = 24'(-21560);
			4054: out = 24'(15876);
			4055: out = 24'(18792);
			4056: out = 24'(57784);
			4057: out = 24'(16740);
			4058: out = 24'(-7124);
			4059: out = 24'(-26792);
			4060: out = 24'(-34404);
			4061: out = 24'(-52904);
			4062: out = 24'(-57088);
			4063: out = 24'(-45448);
			4064: out = 24'(-11612);
			4065: out = 24'(18288);
			4066: out = 24'(38080);
			4067: out = 24'(41556);
			4068: out = 24'(37064);
			4069: out = 24'(2772);
			4070: out = 24'(2228);
			4071: out = 24'(1684);
			4072: out = 24'(2656);
			4073: out = 24'(7072);
			4074: out = 24'(-39792);
			4075: out = 24'(-78404);
			4076: out = 24'(-33064);
			4077: out = 24'(82092);
			4078: out = 24'(88748);
			4079: out = 24'(20368);
			4080: out = 24'(-40896);
			4081: out = 24'(-2688);
			4082: out = 24'(22208);
			4083: out = 24'(44176);
			4084: out = 24'(27772);
			4085: out = 24'(25328);
			4086: out = 24'(30888);
			4087: out = 24'(33280);
			4088: out = 24'(-14240);
			4089: out = 24'(-36828);
			4090: out = 24'(39448);
			4091: out = 24'(83004);
			4092: out = 24'(35544);
			4093: out = 24'(-32032);
			4094: out = 24'(-21864);
			4095: out = 24'(8880);
			4096: out = 24'(8728);
			4097: out = 24'(5416);
			4098: out = 24'(38104);
			4099: out = 24'(-15324);
			4100: out = 24'(-72892);
			4101: out = 24'(-60208);
			4102: out = 24'(45152);
			4103: out = 24'(53500);
			4104: out = 24'(26396);
			4105: out = 24'(2720);
			4106: out = 24'(23628);
			4107: out = 24'(-25828);
			4108: out = 24'(-27652);
			4109: out = 24'(-34372);
			4110: out = 24'(-30052);
			4111: out = 24'(-46876);
			4112: out = 24'(-36748);
			4113: out = 24'(-27156);
			4114: out = 24'(8688);
			4115: out = 24'(40636);
			4116: out = 24'(78116);
			4117: out = 24'(39912);
			4118: out = 24'(-16072);
			4119: out = 24'(-48664);
			4120: out = 24'(14344);
			4121: out = 24'(-12216);
			4122: out = 24'(-78084);
			4123: out = 24'(-102748);
			4124: out = 24'(-38856);
			4125: out = 24'(5388);
			4126: out = 24'(26772);
			4127: out = 24'(36808);
			4128: out = 24'(2284);
			4129: out = 24'(-15152);
			4130: out = 24'(-4564);
			4131: out = 24'(23612);
			4132: out = 24'(-10168);
			4133: out = 24'(15000);
			4134: out = 24'(-11080);
			4135: out = 24'(-57764);
			4136: out = 24'(-98728);
			4137: out = 24'(-11792);
			4138: out = 24'(30124);
			4139: out = 24'(22556);
			4140: out = 24'(13412);
			4141: out = 24'(36104);
			4142: out = 24'(32880);
			4143: out = 24'(5284);
			4144: out = 24'(-17392);
			4145: out = 24'(7052);
			4146: out = 24'(5652);
			4147: out = 24'(-5440);
			4148: out = 24'(-13480);
			4149: out = 24'(-18568);
			4150: out = 24'(-18908);
			4151: out = 24'(-4796);
			4152: out = 24'(33228);
			4153: out = 24'(75168);
			4154: out = 24'(73624);
			4155: out = 24'(37636);
			4156: out = 24'(-27684);
			4157: out = 24'(-106924);
			4158: out = 24'(-26588);
			4159: out = 24'(8964);
			4160: out = 24'(-6216);
			4161: out = 24'(-18724);
			4162: out = 24'(62568);
			4163: out = 24'(75352);
			4164: out = 24'(49472);
			4165: out = 24'(9832);
			4166: out = 24'(-12804);
			4167: out = 24'(-10656);
			4168: out = 24'(4664);
			4169: out = 24'(668);
			4170: out = 24'(-304);
			4171: out = 24'(-50076);
			4172: out = 24'(-46880);
			4173: out = 24'(-27268);
			4174: out = 24'(-24156);
			4175: out = 24'(23480);
			4176: out = 24'(85392);
			4177: out = 24'(92644);
			4178: out = 24'(39168);
			4179: out = 24'(-67352);
			4180: out = 24'(-57096);
			4181: out = 24'(-84);
			4182: out = 24'(17908);
			4183: out = 24'(24564);
			4184: out = 24'(44304);
			4185: out = 24'(34480);
			4186: out = 24'(-24292);
			4187: out = 24'(-83552);
			4188: out = 24'(-45728);
			4189: out = 24'(42076);
			4190: out = 24'(86124);
			4191: out = 24'(59528);
			4192: out = 24'(-7772);
			4193: out = 24'(-82644);
			4194: out = 24'(-92804);
			4195: out = 24'(-17016);
			4196: out = 24'(13868);
			4197: out = 24'(-4872);
			4198: out = 24'(-43280);
			4199: out = 24'(-37884);
			4200: out = 24'(34688);
			4201: out = 24'(46256);
			4202: out = 24'(23464);
			4203: out = 24'(16496);
			4204: out = 24'(26892);
			4205: out = 24'(26128);
			4206: out = 24'(-20900);
			4207: out = 24'(-74812);
			4208: out = 24'(-62832);
			4209: out = 24'(-34164);
			4210: out = 24'(-11012);
			4211: out = 24'(-17524);
			4212: out = 24'(-3588);
			4213: out = 24'(49476);
			4214: out = 24'(90904);
			4215: out = 24'(38020);
			4216: out = 24'(-76632);
			4217: out = 24'(-118812);
			4218: out = 24'(-68308);
			4219: out = 24'(-5972);
			4220: out = 24'(4392);
			4221: out = 24'(16356);
			4222: out = 24'(23800);
			4223: out = 24'(-2648);
			4224: out = 24'(-45176);
			4225: out = 24'(-28052);
			4226: out = 24'(31116);
			4227: out = 24'(65072);
			4228: out = 24'(37540);
			4229: out = 24'(-12736);
			4230: out = 24'(-43596);
			4231: out = 24'(-32056);
			4232: out = 24'(3916);
			4233: out = 24'(19872);
			4234: out = 24'(21756);
			4235: out = 24'(-39372);
			4236: out = 24'(-54016);
			4237: out = 24'(33680);
			4238: out = 24'(92736);
			4239: out = 24'(63328);
			4240: out = 24'(-36604);
			4241: out = 24'(-98816);
			4242: out = 24'(-44944);
			4243: out = 24'(30508);
			4244: out = 24'(37944);
			4245: out = 24'(6760);
			4246: out = 24'(-9384);
			4247: out = 24'(15952);
			4248: out = 24'(14888);
			4249: out = 24'(-1344);
			4250: out = 24'(5980);
			4251: out = 24'(32976);
			4252: out = 24'(43920);
			4253: out = 24'(18908);
			4254: out = 24'(-22372);
			4255: out = 24'(7864);
			4256: out = 24'(-19660);
			4257: out = 24'(-41176);
			4258: out = 24'(-37288);
			4259: out = 24'(-12200);
			4260: out = 24'(15340);
			4261: out = 24'(53860);
			4262: out = 24'(63232);
			4263: out = 24'(19076);
			4264: out = 24'(-34956);
			4265: out = 24'(-37840);
			4266: out = 24'(-1572);
			4267: out = 24'(4808);
			4268: out = 24'(-13180);
			4269: out = 24'(-12520);
			4270: out = 24'(7000);
			4271: out = 24'(-1404);
			4272: out = 24'(12520);
			4273: out = 24'(-652);
			4274: out = 24'(23080);
			4275: out = 24'(59960);
			4276: out = 24'(78524);
			4277: out = 24'(22860);
			4278: out = 24'(-19444);
			4279: out = 24'(-10616);
			4280: out = 24'(45524);
			4281: out = 24'(28684);
			4282: out = 24'(22516);
			4283: out = 24'(13384);
			4284: out = 24'(-25980);
			4285: out = 24'(-42704);
			4286: out = 24'(-28700);
			4287: out = 24'(-6088);
			4288: out = 24'(-16136);
			4289: out = 24'(33372);
			4290: out = 24'(15172);
			4291: out = 24'(-10452);
			4292: out = 24'(-8544);
			4293: out = 24'(40948);
			4294: out = 24'(20044);
			4295: out = 24'(-33916);
			4296: out = 24'(-57544);
			4297: out = 24'(8072);
			4298: out = 24'(45968);
			4299: out = 24'(23928);
			4300: out = 24'(-49980);
			4301: out = 24'(-107188);
			4302: out = 24'(-103204);
			4303: out = 24'(-43960);
			4304: out = 24'(8944);
			4305: out = 24'(27948);
			4306: out = 24'(11504);
			4307: out = 24'(7112);
			4308: out = 24'(6336);
			4309: out = 24'(-836);
			4310: out = 24'(-16916);
			4311: out = 24'(-6888);
			4312: out = 24'(12872);
			4313: out = 24'(19700);
			4314: out = 24'(2456);
			4315: out = 24'(-4940);
			4316: out = 24'(-3016);
			4317: out = 24'(-1976);
			4318: out = 24'(-26312);
			4319: out = 24'(11668);
			4320: out = 24'(16456);
			4321: out = 24'(-7508);
			4322: out = 24'(-15672);
			4323: out = 24'(808);
			4324: out = 24'(19040);
			4325: out = 24'(24996);
			4326: out = 24'(45788);
			4327: out = 24'(77324);
			4328: out = 24'(56700);
			4329: out = 24'(-22432);
			4330: out = 24'(-87392);
			4331: out = 24'(-73784);
			4332: out = 24'(11480);
			4333: out = 24'(28500);
			4334: out = 24'(-20232);
			4335: out = 24'(-66356);
			4336: out = 24'(12236);
			4337: out = 24'(55180);
			4338: out = 24'(23384);
			4339: out = 24'(-112);
			4340: out = 24'(42368);
			4341: out = 24'(73912);
			4342: out = 24'(46944);
			4343: out = 24'(-4232);
			4344: out = 24'(-11228);
			4345: out = 24'(5116);
			4346: out = 24'(22004);
			4347: out = 24'(17972);
			4348: out = 24'(884);
			4349: out = 24'(-30832);
			4350: out = 24'(-25320);
			4351: out = 24'(1748);
			4352: out = 24'(-36484);
			4353: out = 24'(-30316);
			4354: out = 24'(8212);
			4355: out = 24'(55436);
			4356: out = 24'(46188);
			4357: out = 24'(19860);
			4358: out = 24'(-29584);
			4359: out = 24'(-51496);
			4360: out = 24'(-35376);
			4361: out = 24'(25448);
			4362: out = 24'(23748);
			4363: out = 24'(-6352);
			4364: out = 24'(-14516);
			4365: out = 24'(-18684);
			4366: out = 24'(-26040);
			4367: out = 24'(-43392);
			4368: out = 24'(-20028);
			4369: out = 24'(53656);
			4370: out = 24'(78972);
			4371: out = 24'(4040);
			4372: out = 24'(-103348);
			4373: out = 24'(-85296);
			4374: out = 24'(-13192);
			4375: out = 24'(43796);
			4376: out = 24'(20880);
			4377: out = 24'(-8236);
			4378: out = 24'(-45724);
			4379: out = 24'(9884);
			4380: out = 24'(49500);
			4381: out = 24'(8836);
			4382: out = 24'(-91264);
			4383: out = 24'(-85940);
			4384: out = 24'(-4996);
			4385: out = 24'(21480);
			4386: out = 24'(-2408);
			4387: out = 24'(-41564);
			4388: out = 24'(-25452);
			4389: out = 24'(18460);
			4390: out = 24'(40568);
			4391: out = 24'(39312);
			4392: out = 24'(53248);
			4393: out = 24'(63076);
			4394: out = 24'(31748);
			4395: out = 24'(-79972);
			4396: out = 24'(-122016);
			4397: out = 24'(-57400);
			4398: out = 24'(43028);
			4399: out = 24'(71496);
			4400: out = 24'(32752);
			4401: out = 24'(-44356);
			4402: out = 24'(-107280);
			4403: out = 24'(-25784);
			4404: out = 24'(36460);
			4405: out = 24'(56548);
			4406: out = 24'(45468);
			4407: out = 24'(10684);
			4408: out = 24'(-20252);
			4409: out = 24'(-49508);
			4410: out = 24'(-54584);
			4411: out = 24'(-2740);
			4412: out = 24'(67956);
			4413: out = 24'(91432);
			4414: out = 24'(38384);
			4415: out = 24'(-52436);
			4416: out = 24'(-62480);
			4417: out = 24'(-10396);
			4418: out = 24'(24184);
			4419: out = 24'(116);
			4420: out = 24'(10864);
			4421: out = 24'(8452);
			4422: out = 24'(9856);
			4423: out = 24'(12692);
			4424: out = 24'(47996);
			4425: out = 24'(23984);
			4426: out = 24'(-10968);
			4427: out = 24'(-21688);
			4428: out = 24'(18884);
			4429: out = 24'(12464);
			4430: out = 24'(2184);
			4431: out = 24'(3148);
			4432: out = 24'(5588);
			4433: out = 24'(4840);
			4434: out = 24'(-19844);
			4435: out = 24'(-28380);
			4436: out = 24'(14060);
			4437: out = 24'(46132);
			4438: out = 24'(59276);
			4439: out = 24'(35888);
			4440: out = 24'(1116);
			4441: out = 24'(-2248);
			4442: out = 24'(-16032);
			4443: out = 24'(-26008);
			4444: out = 24'(-20880);
			4445: out = 24'(-24604);
			4446: out = 24'(-9600);
			4447: out = 24'(-19764);
			4448: out = 24'(-35252);
			4449: out = 24'(-16944);
			4450: out = 24'(76480);
			4451: out = 24'(94392);
			4452: out = 24'(14508);
			4453: out = 24'(-83864);
			4454: out = 24'(-94548);
			4455: out = 24'(-12096);
			4456: out = 24'(32456);
			4457: out = 24'(-3076);
			4458: out = 24'(2652);
			4459: out = 24'(12748);
			4460: out = 24'(16616);
			4461: out = 24'(-8164);
			4462: out = 24'(-37656);
			4463: out = 24'(-3620);
			4464: out = 24'(36608);
			4465: out = 24'(10312);
			4466: out = 24'(-78624);
			4467: out = 24'(-92424);
			4468: out = 24'(-22276);
			4469: out = 24'(46164);
			4470: out = 24'(35696);
			4471: out = 24'(13288);
			4472: out = 24'(-25300);
			4473: out = 24'(-34304);
			4474: out = 24'(2076);
			4475: out = 24'(47828);
			4476: out = 24'(44564);
			4477: out = 24'(-19248);
			4478: out = 24'(-98624);
			4479: out = 24'(-103816);
			4480: out = 24'(-34676);
			4481: out = 24'(38688);
			4482: out = 24'(58560);
			4483: out = 24'(60416);
			4484: out = 24'(11920);
			4485: out = 24'(-9500);
			4486: out = 24'(768);
			4487: out = 24'(8612);
			4488: out = 24'(11868);
			4489: out = 24'(2228);
			4490: out = 24'(-11660);
			4491: out = 24'(-30116);
			4492: out = 24'(40760);
			4493: out = 24'(33656);
			4494: out = 24'(-15088);
			4495: out = 24'(-50216);
			4496: out = 24'(724);
			4497: out = 24'(42352);
			4498: out = 24'(63356);
			4499: out = 24'(51316);
			4500: out = 24'(12424);
			4501: out = 24'(-59940);
			4502: out = 24'(-95300);
			4503: out = 24'(-61048);
			4504: out = 24'(8152);
			4505: out = 24'(57860);
			4506: out = 24'(65220);
			4507: out = 24'(33536);
			4508: out = 24'(-3132);
			4509: out = 24'(-1348);
			4510: out = 24'(45008);
			4511: out = 24'(48160);
			4512: out = 24'(-21772);
			4513: out = 24'(-25312);
			4514: out = 24'(-14932);
			4515: out = 24'(5904);
			4516: out = 24'(14084);
			4517: out = 24'(89260);
			4518: out = 24'(32704);
			4519: out = 24'(-49104);
			4520: out = 24'(-100560);
			4521: out = 24'(-14988);
			4522: out = 24'(6204);
			4523: out = 24'(29056);
			4524: out = 24'(40580);
			4525: out = 24'(54080);
			4526: out = 24'(-14704);
			4527: out = 24'(-18500);
			4528: out = 24'(5880);
			4529: out = 24'(4272);
			4530: out = 24'(-11620);
			4531: out = 24'(444);
			4532: out = 24'(9164);
			4533: out = 24'(-18776);
			4534: out = 24'(-12260);
			4535: out = 24'(25848);
			4536: out = 24'(67684);
			4537: out = 24'(31968);
			4538: out = 24'(-85380);
			4539: out = 24'(-130020);
			4540: out = 24'(-75664);
			4541: out = 24'(11488);
			4542: out = 24'(29516);
			4543: out = 24'(-16140);
			4544: out = 24'(4348);
			4545: out = 24'(46984);
			4546: out = 24'(35908);
			4547: out = 24'(7196);
			4548: out = 24'(18688);
			4549: out = 24'(39640);
			4550: out = 24'(7144);
			4551: out = 24'(-90008);
			4552: out = 24'(-102784);
			4553: out = 24'(-27700);
			4554: out = 24'(38352);
			4555: out = 24'(40500);
			4556: out = 24'(32624);
			4557: out = 24'(17356);
			4558: out = 24'(-2556);
			4559: out = 24'(-18364);
			4560: out = 24'(-15152);
			4561: out = 24'(-12464);
			4562: out = 24'(-5876);
			4563: out = 24'(20868);
			4564: out = 24'(-2956);
			4565: out = 24'(-36460);
			4566: out = 24'(-50016);
			4567: out = 24'(-12336);
			4568: out = 24'(14424);
			4569: out = 24'(53576);
			4570: out = 24'(59808);
			4571: out = 24'(14412);
			4572: out = 24'(-61280);
			4573: out = 24'(-73840);
			4574: out = 24'(9828);
			4575: out = 24'(83548);
			4576: out = 24'(57216);
			4577: out = 24'(-12256);
			4578: out = 24'(-50336);
			4579: out = 24'(-29072);
			4580: out = 24'(14772);
			4581: out = 24'(38180);
			4582: out = 24'(54524);
			4583: out = 24'(41188);
			4584: out = 24'(-792);
			4585: out = 24'(-49804);
			4586: out = 24'(-24720);
			4587: out = 24'(13972);
			4588: out = 24'(-3660);
			4589: out = 24'(-27528);
			4590: out = 24'(-13116);
			4591: out = 24'(25076);
			4592: out = 24'(38796);
			4593: out = 24'(49076);
			4594: out = 24'(41528);
			4595: out = 24'(19836);
			4596: out = 24'(-17548);
			4597: out = 24'(-41028);
			4598: out = 24'(-40068);
			4599: out = 24'(-37104);
			4600: out = 24'(-38084);
			4601: out = 24'(-3608);
			4602: out = 24'(14780);
			4603: out = 24'(17652);
			4604: out = 24'(7212);
			4605: out = 24'(39380);
			4606: out = 24'(34788);
			4607: out = 24'(57784);
			4608: out = 24'(20396);
			4609: out = 24'(-48764);
			4610: out = 24'(-97732);
			4611: out = 24'(-25564);
			4612: out = 24'(31616);
			4613: out = 24'(11176);
			4614: out = 24'(-10416);
			4615: out = 24'(-16480);
			4616: out = 24'(-10016);
			4617: out = 24'(10496);
			4618: out = 24'(45164);
			4619: out = 24'(58488);
			4620: out = 24'(8264);
			4621: out = 24'(-43888);
			4622: out = 24'(-35944);
			4623: out = 24'(-22216);
			4624: out = 24'(-46332);
			4625: out = 24'(-51268);
			4626: out = 24'(9460);
			4627: out = 24'(45260);
			4628: out = 24'(32700);
			4629: out = 24'(27324);
			4630: out = 24'(45912);
			4631: out = 24'(2040);
			4632: out = 24'(-52652);
			4633: out = 24'(-50928);
			4634: out = 24'(24148);
			4635: out = 24'(29440);
			4636: out = 24'(-1744);
			4637: out = 24'(-66436);
			4638: out = 24'(-75312);
			4639: out = 24'(-18840);
			4640: out = 24'(48984);
			4641: out = 24'(79296);
			4642: out = 24'(76384);
			4643: out = 24'(25372);
			4644: out = 24'(-43716);
			4645: out = 24'(-99280);
			4646: out = 24'(-56424);
			4647: out = 24'(28748);
			4648: out = 24'(7072);
			4649: out = 24'(-43680);
			4650: out = 24'(-42472);
			4651: out = 24'(20932);
			4652: out = 24'(24088);
			4653: out = 24'(30192);
			4654: out = 24'(31920);
			4655: out = 24'(30432);
			4656: out = 24'(-30332);
			4657: out = 24'(-48380);
			4658: out = 24'(-45592);
			4659: out = 24'(3448);
			4660: out = 24'(37536);
			4661: out = 24'(74648);
			4662: out = 24'(3672);
			4663: out = 24'(-60132);
			4664: out = 24'(-30644);
			4665: out = 24'(10380);
			4666: out = 24'(29300);
			4667: out = 24'(6988);
			4668: out = 24'(-5124);
			4669: out = 24'(-22928);
			4670: out = 24'(12992);
			4671: out = 24'(13832);
			4672: out = 24'(2872);
			4673: out = 24'(5052);
			4674: out = 24'(26516);
			4675: out = 24'(320);
			4676: out = 24'(-27680);
			4677: out = 24'(-2132);
			4678: out = 24'(68212);
			4679: out = 24'(48292);
			4680: out = 24'(-24692);
			4681: out = 24'(-65496);
			4682: out = 24'(-6444);
			4683: out = 24'(33540);
			4684: out = 24'(28840);
			4685: out = 24'(-1344);
			4686: out = 24'(-49704);
			4687: out = 24'(-49708);
			4688: out = 24'(348);
			4689: out = 24'(36504);
			4690: out = 24'(-3580);
			4691: out = 24'(30940);
			4692: out = 24'(80336);
			4693: out = 24'(64084);
			4694: out = 24'(-51632);
			4695: out = 24'(-108044);
			4696: out = 24'(-65332);
			4697: out = 24'(21544);
			4698: out = 24'(10416);
			4699: out = 24'(-17744);
			4700: out = 24'(-50376);
			4701: out = 24'(-6344);
			4702: out = 24'(54756);
			4703: out = 24'(72536);
			4704: out = 24'(43844);
			4705: out = 24'(22320);
			4706: out = 24'(988);
			4707: out = 24'(3984);
			4708: out = 24'(-63136);
			4709: out = 24'(-50036);
			4710: out = 24'(24148);
			4711: out = 24'(44284);
			4712: out = 24'(17508);
			4713: out = 24'(12316);
			4714: out = 24'(19776);
			4715: out = 24'(-25328);
			4716: out = 24'(56);
			4717: out = 24'(-1312);
			4718: out = 24'(3800);
			4719: out = 24'(7116);
			4720: out = 24'(30068);
			4721: out = 24'(-19076);
			4722: out = 24'(-89156);
			4723: out = 24'(-103008);
			4724: out = 24'(7624);
			4725: out = 24'(79352);
			4726: out = 24'(55460);
			4727: out = 24'(-10644);
			4728: out = 24'(-14572);
			4729: out = 24'(-7176);
			4730: out = 24'(-1232);
			4731: out = 24'(-33596);
			4732: out = 24'(-46204);
			4733: out = 24'(-23788);
			4734: out = 24'(52908);
			4735: out = 24'(67512);
			4736: out = 24'(14164);
			4737: out = 24'(-59968);
			4738: out = 24'(-21200);
			4739: out = 24'(30008);
			4740: out = 24'(-4692);
			4741: out = 24'(-42468);
			4742: out = 24'(-27420);
			4743: out = 24'(40628);
			4744: out = 24'(53880);
			4745: out = 24'(9304);
			4746: out = 24'(-46088);
			4747: out = 24'(-14096);
			4748: out = 24'(64708);
			4749: out = 24'(82652);
			4750: out = 24'(-16200);
			4751: out = 24'(-100360);
			4752: out = 24'(-65420);
			4753: out = 24'(68356);
			4754: out = 24'(62036);
			4755: out = 24'(15516);
			4756: out = 24'(-36068);
			4757: out = 24'(-34980);
			4758: out = 24'(-27632);
			4759: out = 24'(12664);
			4760: out = 24'(7428);
			4761: out = 24'(-20608);
			4762: out = 24'(-20236);
			4763: out = 24'(34752);
			4764: out = 24'(51092);
			4765: out = 24'(27412);
			4766: out = 24'(39040);
			4767: out = 24'(35028);
			4768: out = 24'(14952);
			4769: out = 24'(-33428);
			4770: out = 24'(-58384);
			4771: out = 24'(-19440);
			4772: out = 24'(23620);
			4773: out = 24'(5016);
			4774: out = 24'(-46916);
			4775: out = 24'(-117616);
			4776: out = 24'(-37344);
			4777: out = 24'(92084);
			4778: out = 24'(108272);
			4779: out = 24'(18712);
			4780: out = 24'(-79712);
			4781: out = 24'(-117332);
			4782: out = 24'(-73444);
			4783: out = 24'(16476);
			4784: out = 24'(64920);
			4785: out = 24'(65576);
			4786: out = 24'(48320);
			4787: out = 24'(22672);
			4788: out = 24'(-33492);
			4789: out = 24'(-73804);
			4790: out = 24'(-18272);
			4791: out = 24'(90752);
			4792: out = 24'(55596);
			4793: out = 24'(-39296);
			4794: out = 24'(-90672);
			4795: out = 24'(-13008);
			4796: out = 24'(5364);
			4797: out = 24'(43076);
			4798: out = 24'(50980);
			4799: out = 24'(44192);
			4800: out = 24'(-45412);
			4801: out = 24'(-21708);
			4802: out = 24'(5424);
			4803: out = 24'(12900);
			4804: out = 24'(68);
			4805: out = 24'(7488);
			4806: out = 24'(-3020);
			4807: out = 24'(-15576);
			4808: out = 24'(-12900);
			4809: out = 24'(-1916);
			4810: out = 24'(-6680);
			4811: out = 24'(-11548);
			4812: out = 24'(2668);
			4813: out = 24'(436);
			4814: out = 24'(23724);
			4815: out = 24'(49980);
			4816: out = 24'(44456);
			4817: out = 24'(-67352);
			4818: out = 24'(-69228);
			4819: out = 24'(-6600);
			4820: out = 24'(35064);
			4821: out = 24'(-12756);
			4822: out = 24'(-61204);
			4823: out = 24'(-58304);
			4824: out = 24'(14192);
			4825: out = 24'(42464);
			4826: out = 24'(59428);
			4827: out = 24'(11144);
			4828: out = 24'(12964);
			4829: out = 24'(59460);
			4830: out = 24'(20472);
			4831: out = 24'(-73864);
			4832: out = 24'(-92840);
			4833: out = 24'(12932);
			4834: out = 24'(27268);
			4835: out = 24'(15788);
			4836: out = 24'(-888);
			4837: out = 24'(12156);
			4838: out = 24'(12168);
			4839: out = 24'(5204);
			4840: out = 24'(14092);
			4841: out = 24'(46120);
			4842: out = 24'(48496);
			4843: out = 24'(42676);
			4844: out = 24'(2792);
			4845: out = 24'(-50332);
			4846: out = 24'(-93040);
			4847: out = 24'(-57676);
			4848: out = 24'(24216);
			4849: out = 24'(71484);
			4850: out = 24'(39312);
			4851: out = 24'(-32868);
			4852: out = 24'(-64920);
			4853: out = 24'(-27992);
			4854: out = 24'(14808);
			4855: out = 24'(2056);
			4856: out = 24'(15364);
			4857: out = 24'(39644);
			4858: out = 24'(22204);
			4859: out = 24'(-79816);
			4860: out = 24'(-35692);
			4861: out = 24'(42888);
			4862: out = 24'(59880);
			4863: out = 24'(19168);
			4864: out = 24'(-11740);
			4865: out = 24'(5028);
			4866: out = 24'(8064);
			4867: out = 24'(-41528);
			4868: out = 24'(-86888);
			4869: out = 24'(-54640);
			4870: out = 24'(25128);
			4871: out = 24'(66576);
			4872: out = 24'(69904);
			4873: out = 24'(15764);
			4874: out = 24'(-43444);
			4875: out = 24'(-52952);
			4876: out = 24'(2124);
			4877: out = 24'(60064);
			4878: out = 24'(43284);
			4879: out = 24'(-9316);
			4880: out = 24'(-33036);
			4881: out = 24'(-7860);
			4882: out = 24'(-1400);
			4883: out = 24'(-5396);
			4884: out = 24'(8352);
			4885: out = 24'(30388);
			4886: out = 24'(-31984);
			4887: out = 24'(-104692);
			4888: out = 24'(-65548);
			4889: out = 24'(34204);
			4890: out = 24'(104544);
			4891: out = 24'(62764);
			4892: out = 24'(-23336);
			4893: out = 24'(-80580);
			4894: out = 24'(-41336);
			4895: out = 24'(11260);
			4896: out = 24'(18756);
			4897: out = 24'(23856);
			4898: out = 24'(1300);
			4899: out = 24'(16540);
			4900: out = 24'(34292);
			4901: out = 24'(30004);
			4902: out = 24'(8684);
			4903: out = 24'(14968);
			4904: out = 24'(22752);
			4905: out = 24'(-6060);
			4906: out = 24'(-90344);
			4907: out = 24'(-99804);
			4908: out = 24'(-25204);
			4909: out = 24'(45392);
			4910: out = 24'(65608);
			4911: out = 24'(25092);
			4912: out = 24'(7148);
			4913: out = 24'(26168);
			4914: out = 24'(32444);
			4915: out = 24'(-708);
			4916: out = 24'(-67644);
			4917: out = 24'(-99668);
			4918: out = 24'(-14064);
			4919: out = 24'(24384);
			4920: out = 24'(64604);
			4921: out = 24'(50876);
			4922: out = 24'(-5968);
			4923: out = 24'(-92352);
			4924: out = 24'(-87524);
			4925: out = 24'(-23076);
			4926: out = 24'(30476);
			4927: out = 24'(71940);
			4928: out = 24'(66764);
			4929: out = 24'(16632);
			4930: out = 24'(-53124);
			4931: out = 24'(-81492);
			4932: out = 24'(-22068);
			4933: out = 24'(27700);
			4934: out = 24'(12288);
			4935: out = 24'(8220);
			4936: out = 24'(-52596);
			4937: out = 24'(-32008);
			4938: out = 24'(23296);
			4939: out = 24'(55508);
			4940: out = 24'(31132);
			4941: out = 24'(33544);
			4942: out = 24'(31368);
			4943: out = 24'(348);
			4944: out = 24'(-47404);
			4945: out = 24'(-43044);
			4946: out = 24'(-11876);
			4947: out = 24'(4516);
			4948: out = 24'(39620);
			4949: out = 24'(29740);
			4950: out = 24'(20104);
			4951: out = 24'(1280);
			4952: out = 24'(-10476);
			4953: out = 24'(-37776);
			4954: out = 24'(-19704);
			4955: out = 24'(29920);
			4956: out = 24'(78692);
			4957: out = 24'(44408);
			4958: out = 24'(5400);
			4959: out = 24'(-33664);
			4960: out = 24'(-28192);
			4961: out = 24'(-24784);
			4962: out = 24'(51600);
			4963: out = 24'(67228);
			4964: out = 24'(19780);
			4965: out = 24'(-32312);
			4966: out = 24'(-13224);
			4967: out = 24'(-18044);
			4968: out = 24'(-48544);
			4969: out = 24'(-8056);
			4970: out = 24'(48492);
			4971: out = 24'(37956);
			4972: out = 24'(-26980);
			4973: out = 24'(-43716);
			4974: out = 24'(-42908);
			4975: out = 24'(-11536);
			4976: out = 24'(28272);
			4977: out = 24'(72628);
			4978: out = 24'(21900);
			4979: out = 24'(-32676);
			4980: out = 24'(-70148);
			4981: out = 24'(-47588);
			4982: out = 24'(-26280);
			4983: out = 24'(3588);
			4984: out = 24'(13540);
			4985: out = 24'(21812);
			4986: out = 24'(712);
			4987: out = 24'(-5200);
			4988: out = 24'(-15184);
			4989: out = 24'(7640);
			4990: out = 24'(32396);
			4991: out = 24'(47424);
			4992: out = 24'(-27476);
			4993: out = 24'(-100576);
			4994: out = 24'(-60532);
			4995: out = 24'(43352);
			4996: out = 24'(44636);
			4997: out = 24'(-32812);
			4998: out = 24'(-64708);
			4999: out = 24'(-21132);
			5000: out = 24'(54916);
			5001: out = 24'(59444);
			5002: out = 24'(15772);
			5003: out = 24'(-74992);
			5004: out = 24'(-22932);
			5005: out = 24'(48164);
			5006: out = 24'(50576);
			5007: out = 24'(6228);
			5008: out = 24'(-44172);
			5009: out = 24'(-75612);
			5010: out = 24'(-78492);
			5011: out = 24'(-47484);
			5012: out = 24'(18084);
			5013: out = 24'(73948);
			5014: out = 24'(82992);
			5015: out = 24'(37052);
			5016: out = 24'(-21272);
			5017: out = 24'(-68848);
			5018: out = 24'(-54392);
			5019: out = 24'(2992);
			5020: out = 24'(22652);
			5021: out = 24'(31116);
			5022: out = 24'(46180);
			5023: out = 24'(49388);
			5024: out = 24'(6400);
			5025: out = 24'(-18100);
			5026: out = 24'(19544);
			5027: out = 24'(77244);
			5028: out = 24'(45536);
			5029: out = 24'(-27204);
			5030: out = 24'(-92560);
			5031: out = 24'(-45728);
			5032: out = 24'(62892);
			5033: out = 24'(67672);
			5034: out = 24'(7908);
			5035: out = 24'(-26112);
			5036: out = 24'(5188);
			5037: out = 24'(32900);
			5038: out = 24'(40688);
			5039: out = 24'(48416);
			5040: out = 24'(53232);
			5041: out = 24'(37708);
			5042: out = 24'(-42336);
			5043: out = 24'(-91340);
			5044: out = 24'(-55876);
			5045: out = 24'(648);
			5046: out = 24'(20880);
			5047: out = 24'(10968);
			5048: out = 24'(-10968);
			5049: out = 24'(-61460);
			5050: out = 24'(-13024);
			5051: out = 24'(17616);
			5052: out = 24'(12096);
			5053: out = 24'(-12152);
			5054: out = 24'(-3060);
			5055: out = 24'(23152);
			5056: out = 24'(44360);
			5057: out = 24'(41668);
			5058: out = 24'(-14236);
			5059: out = 24'(-11972);
			5060: out = 24'(4812);
			5061: out = 24'(8512);
			5062: out = 24'(35472);
			5063: out = 24'(24572);
			5064: out = 24'(-12088);
			5065: out = 24'(-70988);
			5066: out = 24'(-73968);
			5067: out = 24'(-100292);
			5068: out = 24'(-44300);
			5069: out = 24'(22836);
			5070: out = 24'(23728);
			5071: out = 24'(-25572);
			5072: out = 24'(-34744);
			5073: out = 24'(-4284);
			5074: out = 24'(11844);
			5075: out = 24'(48304);
			5076: out = 24'(58212);
			5077: out = 24'(46284);
			5078: out = 24'(-4884);
			5079: out = 24'(-31012);
			5080: out = 24'(-79816);
			5081: out = 24'(-52964);
			5082: out = 24'(16468);
			5083: out = 24'(37220);
			5084: out = 24'(13468);
			5085: out = 24'(-5516);
			5086: out = 24'(-2652);
			5087: out = 24'(636);
			5088: out = 24'(-9508);
			5089: out = 24'(4432);
			5090: out = 24'(28340);
			5091: out = 24'(21272);
			5092: out = 24'(-22000);
			5093: out = 24'(-32512);
			5094: out = 24'(-224);
			5095: out = 24'(21160);
			5096: out = 24'(35760);
			5097: out = 24'(21308);
			5098: out = 24'(29944);
			5099: out = 24'(31012);
			5100: out = 24'(3148);
			5101: out = 24'(-60104);
			5102: out = 24'(-69496);
			5103: out = 24'(-28128);
			5104: out = 24'(1136);
			5105: out = 24'(27508);
			5106: out = 24'(43628);
			5107: out = 24'(33288);
			5108: out = 24'(456);
			5109: out = 24'(-36640);
			5110: out = 24'(-14576);
			5111: out = 24'(20488);
			5112: out = 24'(33912);
			5113: out = 24'(35256);
			5114: out = 24'(20712);
			5115: out = 24'(-44952);
			5116: out = 24'(-107588);
			5117: out = 24'(-41816);
			5118: out = 24'(26072);
			5119: out = 24'(26384);
			5120: out = 24'(7228);
			5121: out = 24'(37732);
			5122: out = 24'(61424);
			5123: out = 24'(7084);
			5124: out = 24'(-46672);
			5125: out = 24'(16192);
			5126: out = 24'(71360);
			5127: out = 24'(45608);
			5128: out = 24'(-33540);
			5129: out = 24'(-69676);
			5130: out = 24'(-109036);
			5131: out = 24'(-47068);
			5132: out = 24'(50368);
			5133: out = 24'(97196);
			5134: out = 24'(42524);
			5135: out = 24'(-660);
			5136: out = 24'(-8420);
			5137: out = 24'(5460);
			5138: out = 24'(-20400);
			5139: out = 24'(-29064);
			5140: out = 24'(7700);
			5141: out = 24'(51640);
			5142: out = 24'(11968);
			5143: out = 24'(-8012);
			5144: out = 24'(-30300);
			5145: out = 24'(-436);
			5146: out = 24'(37784);
			5147: out = 24'(77616);
			5148: out = 24'(34456);
			5149: out = 24'(-13708);
			5150: out = 24'(-37532);
			5151: out = 24'(-22796);
			5152: out = 24'(-24760);
			5153: out = 24'(-5216);
			5154: out = 24'(20904);
			5155: out = 24'(19192);
			5156: out = 24'(20088);
			5157: out = 24'(33388);
			5158: out = 24'(16796);
			5159: out = 24'(-55848);
			5160: out = 24'(-104516);
			5161: out = 24'(-57664);
			5162: out = 24'(35936);
			5163: out = 24'(55348);
			5164: out = 24'(-8040);
			5165: out = 24'(-49080);
			5166: out = 24'(-30124);
			5167: out = 24'(8484);
			5168: out = 24'(8296);
			5169: out = 24'(27120);
			5170: out = 24'(36200);
			5171: out = 24'(10548);
			5172: out = 24'(-14612);
			5173: out = 24'(-35184);
			5174: out = 24'(-18392);
			5175: out = 24'(6560);
			5176: out = 24'(19004);
			5177: out = 24'(-45184);
			5178: out = 24'(-83772);
			5179: out = 24'(-58348);
			5180: out = 24'(-4612);
			5181: out = 24'(12120);
			5182: out = 24'(2928);
			5183: out = 24'(-1700);
			5184: out = 24'(7568);
			5185: out = 24'(61676);
			5186: out = 24'(36384);
			5187: out = 24'(-11404);
			5188: out = 24'(-26908);
			5189: out = 24'(4376);
			5190: out = 24'(25436);
			5191: out = 24'(18676);
			5192: out = 24'(-2204);
			5193: out = 24'(-16788);
			5194: out = 24'(-5472);
			5195: out = 24'(5260);
			5196: out = 24'(624);
			5197: out = 24'(5032);
			5198: out = 24'(27972);
			5199: out = 24'(49452);
			5200: out = 24'(15304);
			5201: out = 24'(-62676);
			5202: out = 24'(-80868);
			5203: out = 24'(-4716);
			5204: out = 24'(68028);
			5205: out = 24'(49992);
			5206: out = 24'(34848);
			5207: out = 24'(15364);
			5208: out = 24'(24916);
			5209: out = 24'(6480);
			5210: out = 24'(-32132);
			5211: out = 24'(-40164);
			5212: out = 24'(41368);
			5213: out = 24'(92796);
			5214: out = 24'(27512);
			5215: out = 24'(-71788);
			5216: out = 24'(-88584);
			5217: out = 24'(-1524);
			5218: out = 24'(46860);
			5219: out = 24'(46304);
			5220: out = 24'(2988);
			5221: out = 24'(-12844);
			5222: out = 24'(928);
			5223: out = 24'(17104);
			5224: out = 24'(-8252);
			5225: out = 24'(-44048);
			5226: out = 24'(-48772);
			5227: out = 24'(6372);
			5228: out = 24'(10252);
			5229: out = 24'(-27784);
			5230: out = 24'(-63040);
			5231: out = 24'(-40080);
			5232: out = 24'(-8428);
			5233: out = 24'(15748);
			5234: out = 24'(22548);
			5235: out = 24'(22384);
			5236: out = 24'(35880);
			5237: out = 24'(23052);
			5238: out = 24'(-15232);
			5239: out = 24'(-43428);
			5240: out = 24'(-21444);
			5241: out = 24'(25568);
			5242: out = 24'(42364);
			5243: out = 24'(7056);
			5244: out = 24'(-88472);
			5245: out = 24'(-110128);
			5246: out = 24'(-52308);
			5247: out = 24'(19176);
			5248: out = 24'(34332);
			5249: out = 24'(56644);
			5250: out = 24'(49524);
			5251: out = 24'(3956);
			5252: out = 24'(-38808);
			5253: out = 24'(-16876);
			5254: out = 24'(56368);
			5255: out = 24'(82152);
			5256: out = 24'(41792);
			5257: out = 24'(-78584);
			5258: out = 24'(-88596);
			5259: out = 24'(-17972);
			5260: out = 24'(14020);
			5261: out = 24'(24768);
			5262: out = 24'(20196);
			5263: out = 24'(15472);
			5264: out = 24'(-9972);
			5265: out = 24'(6716);
			5266: out = 24'(-30496);
			5267: out = 24'(-20944);
			5268: out = 24'(30080);
			5269: out = 24'(60908);
			5270: out = 24'(16840);
			5271: out = 24'(-40628);
			5272: out = 24'(-50948);
			5273: out = 24'(5948);
			5274: out = 24'(55720);
			5275: out = 24'(47976);
			5276: out = 24'(-1832);
			5277: out = 24'(-28252);
			5278: out = 24'(-8300);
			5279: out = 24'(13840);
			5280: out = 24'(-12308);
			5281: out = 24'(-33276);
			5282: out = 24'(-752);
			5283: out = 24'(88428);
			5284: out = 24'(95048);
			5285: out = 24'(34520);
			5286: out = 24'(-25904);
			5287: out = 24'(-33388);
			5288: out = 24'(-63740);
			5289: out = 24'(-87964);
			5290: out = 24'(-16392);
			5291: out = 24'(76196);
			5292: out = 24'(68880);
			5293: out = 24'(-23000);
			5294: out = 24'(-106032);
			5295: out = 24'(-120300);
			5296: out = 24'(-87212);
			5297: out = 24'(31292);
			5298: out = 24'(118880);
			5299: out = 24'(115492);
			5300: out = 24'(22648);
			5301: out = 24'(-70448);
			5302: out = 24'(-81120);
			5303: out = 24'(-5212);
			5304: out = 24'(24292);
			5305: out = 24'(40412);
			5306: out = 24'(49088);
			5307: out = 24'(-10852);
			5308: out = 24'(-90844);
			5309: out = 24'(-110204);
			5310: out = 24'(-17552);
			5311: out = 24'(68260);
			5312: out = 24'(76624);
			5313: out = 24'(12328);
			5314: out = 24'(-30696);
			5315: out = 24'(-20532);
			5316: out = 24'(29040);
			5317: out = 24'(30892);
			5318: out = 24'(30684);
			5319: out = 24'(27236);
			5320: out = 24'(32);
			5321: out = 24'(-39844);
			5322: out = 24'(-27884);
			5323: out = 24'(-464);
			5324: out = 24'(-35964);
			5325: out = 24'(-30696);
			5326: out = 24'(28932);
			5327: out = 24'(55048);
			5328: out = 24'(-20020);
			5329: out = 24'(-73616);
			5330: out = 24'(-44152);
			5331: out = 24'(17700);
			5332: out = 24'(6320);
			5333: out = 24'(6588);
			5334: out = 24'(29180);
			5335: out = 24'(55944);
			5336: out = 24'(29376);
			5337: out = 24'(3528);
			5338: out = 24'(-54072);
			5339: out = 24'(-83964);
			5340: out = 24'(-61280);
			5341: out = 24'(11664);
			5342: out = 24'(53124);
			5343: out = 24'(34268);
			5344: out = 24'(-21016);
			5345: out = 24'(-69460);
			5346: out = 24'(-2244);
			5347: out = 24'(58956);
			5348: out = 24'(70076);
			5349: out = 24'(52692);
			5350: out = 24'(29124);
			5351: out = 24'(-21912);
			5352: out = 24'(-61208);
			5353: out = 24'(-33224);
			5354: out = 24'(51892);
			5355: out = 24'(65984);
			5356: out = 24'(15240);
			5357: out = 24'(-36160);
			5358: out = 24'(-41420);
			5359: out = 24'(-6576);
			5360: out = 24'(9600);
			5361: out = 24'(-3888);
			5362: out = 24'(-14208);
			5363: out = 24'(54840);
			5364: out = 24'(96436);
			5365: out = 24'(59636);
			5366: out = 24'(-7044);
			5367: out = 24'(-84624);
			5368: out = 24'(-48732);
			5369: out = 24'(36880);
			5370: out = 24'(56468);
			5371: out = 24'(12076);
			5372: out = 24'(-14828);
			5373: out = 24'(-9868);
			5374: out = 24'(-8584);
			5375: out = 24'(15568);
			5376: out = 24'(-3816);
			5377: out = 24'(5544);
			5378: out = 24'(27088);
			5379: out = 24'(30240);
			5380: out = 24'(-48000);
			5381: out = 24'(-77056);
			5382: out = 24'(-10624);
			5383: out = 24'(58900);
			5384: out = 24'(85084);
			5385: out = 24'(32252);
			5386: out = 24'(-44176);
			5387: out = 24'(-99764);
			5388: out = 24'(-55288);
			5389: out = 24'(-16156);
			5390: out = 24'(-2632);
			5391: out = 24'(6708);
			5392: out = 24'(33580);
			5393: out = 24'(19456);
			5394: out = 24'(-31480);
			5395: out = 24'(-53468);
			5396: out = 24'(67948);
			5397: out = 24'(60404);
			5398: out = 24'(14968);
			5399: out = 24'(-23612);
			5400: out = 24'(-5324);
			5401: out = 24'(-9828);
			5402: out = 24'(7528);
			5403: out = 24'(13648);
			5404: out = 24'(-23532);
			5405: out = 24'(-12280);
			5406: out = 24'(-32376);
			5407: out = 24'(-48876);
			5408: out = 24'(-33824);
			5409: out = 24'(7620);
			5410: out = 24'(55636);
			5411: out = 24'(77400);
			5412: out = 24'(44592);
			5413: out = 24'(-55976);
			5414: out = 24'(-76588);
			5415: out = 24'(-29560);
			5416: out = 24'(-1080);
			5417: out = 24'(-19484);
			5418: out = 24'(2276);
			5419: out = 24'(64260);
			5420: out = 24'(72460);
			5421: out = 24'(25736);
			5422: out = 24'(-76052);
			5423: out = 24'(-51000);
			5424: out = 24'(8124);
			5425: out = 24'(-16408);
			5426: out = 24'(-29112);
			5427: out = 24'(10228);
			5428: out = 24'(36588);
			5429: out = 24'(-8060);
			5430: out = 24'(-31688);
			5431: out = 24'(6308);
			5432: out = 24'(68972);
			5433: out = 24'(75904);
			5434: out = 24'(21448);
			5435: out = 24'(-7696);
			5436: out = 24'(-50528);
			5437: out = 24'(-86808);
			5438: out = 24'(-65628);
			5439: out = 24'(6432);
			5440: out = 24'(46604);
			5441: out = 24'(47024);
			5442: out = 24'(35216);
			5443: out = 24'(10460);
			5444: out = 24'(-41816);
			5445: out = 24'(-55196);
			5446: out = 24'(10844);
			5447: out = 24'(27088);
			5448: out = 24'(43792);
			5449: out = 24'(32224);
			5450: out = 24'(888);
			5451: out = 24'(-13468);
			5452: out = 24'(-43576);
			5453: out = 24'(-18956);
			5454: out = 24'(25848);
			5455: out = 24'(19808);
			5456: out = 24'(-19380);
			5457: out = 24'(-18768);
			5458: out = 24'(21412);
			5459: out = 24'(35744);
			5460: out = 24'(47536);
			5461: out = 24'(33340);
			5462: out = 24'(9616);
			5463: out = 24'(-688);
			5464: out = 24'(-63784);
			5465: out = 24'(-36920);
			5466: out = 24'(13048);
			5467: out = 24'(37916);
			5468: out = 24'(17500);
			5469: out = 24'(50900);
			5470: out = 24'(47588);
			5471: out = 24'(2100);
			5472: out = 24'(-90120);
			5473: out = 24'(-34384);
			5474: out = 24'(-14400);
			5475: out = 24'(-37672);
			5476: out = 24'(18976);
			5477: out = 24'(81364);
			5478: out = 24'(62992);
			5479: out = 24'(-36264);
			5480: out = 24'(-105136);
			5481: out = 24'(-53700);
			5482: out = 24'(25280);
			5483: out = 24'(32436);
			5484: out = 24'(-2044);
			5485: out = 24'(-28780);
			5486: out = 24'(-35396);
			5487: out = 24'(-18900);
			5488: out = 24'(15480);
			5489: out = 24'(28760);
			5490: out = 24'(20440);
			5491: out = 24'(-14688);
			5492: out = 24'(-36632);
			5493: out = 24'(-6668);
			5494: out = 24'(-8432);
			5495: out = 24'(-13716);
			5496: out = 24'(-4240);
			5497: out = 24'(15204);
			5498: out = 24'(26980);
			5499: out = 24'(14020);
			5500: out = 24'(-4380);
			5501: out = 24'(-13404);
			5502: out = 24'(-34708);
			5503: out = 24'(-24716);
			5504: out = 24'(23804);
			5505: out = 24'(62732);
			5506: out = 24'(36572);
			5507: out = 24'(3596);
			5508: out = 24'(1560);
			5509: out = 24'(19220);
			5510: out = 24'(1192);
			5511: out = 24'(-2184);
			5512: out = 24'(8744);
			5513: out = 24'(16072);
			5514: out = 24'(-1644);
			5515: out = 24'(-34180);
			5516: out = 24'(-35060);
			5517: out = 24'(-10588);
			5518: out = 24'(15440);
			5519: out = 24'(15460);
			5520: out = 24'(55556);
			5521: out = 24'(65956);
			5522: out = 24'(692);
			5523: out = 24'(-90356);
			5524: out = 24'(-112020);
			5525: out = 24'(-32416);
			5526: out = 24'(64380);
			5527: out = 24'(63648);
			5528: out = 24'(68896);
			5529: out = 24'(28700);
			5530: out = 24'(-30076);
			5531: out = 24'(-75048);
			5532: out = 24'(4300);
			5533: out = 24'(53636);
			5534: out = 24'(26796);
			5535: out = 24'(-18716);
			5536: out = 24'(-2776);
			5537: out = 24'(4104);
			5538: out = 24'(-28576);
			5539: out = 24'(-53876);
			5540: out = 24'(52832);
			5541: out = 24'(53856);
			5542: out = 24'(-46340);
			5543: out = 24'(-115232);
			5544: out = 24'(-40864);
			5545: out = 24'(60828);
			5546: out = 24'(52408);
			5547: out = 24'(1204);
			5548: out = 24'(5040);
			5549: out = 24'(26900);
			5550: out = 24'(688);
			5551: out = 24'(-27056);
			5552: out = 24'(51884);
			5553: out = 24'(82788);
			5554: out = 24'(45372);
			5555: out = 24'(-61972);
			5556: out = 24'(-106888);
			5557: out = 24'(-111952);
			5558: out = 24'(-11620);
			5559: out = 24'(46748);
			5560: out = 24'(29620);
			5561: out = 24'(-20796);
			5562: out = 24'(108);
			5563: out = 24'(26016);
			5564: out = 24'(13836);
			5565: out = 24'(9968);
			5566: out = 24'(12000);
			5567: out = 24'(24688);
			5568: out = 24'(15904);
			5569: out = 24'(-5972);
			5570: out = 24'(3248);
			5571: out = 24'(28204);
			5572: out = 24'(20460);
			5573: out = 24'(-35264);
			5574: out = 24'(-106400);
			5575: out = 24'(-72904);
			5576: out = 24'(44256);
			5577: out = 24'(95844);
			5578: out = 24'(61716);
			5579: out = 24'(-32500);
			5580: out = 24'(-99620);
			5581: out = 24'(-91776);
			5582: out = 24'(-13876);
			5583: out = 24'(31888);
			5584: out = 24'(56428);
			5585: out = 24'(60220);
			5586: out = 24'(46116);
			5587: out = 24'(-30456);
			5588: out = 24'(-66564);
			5589: out = 24'(-40404);
			5590: out = 24'(972);
			5591: out = 24'(6760);
			5592: out = 24'(25432);
			5593: out = 24'(18704);
			5594: out = 24'(-59884);
			5595: out = 24'(3344);
			5596: out = 24'(22376);
			5597: out = 24'(46188);
			5598: out = 24'(20060);
			5599: out = 24'(-25140);
			5600: out = 24'(-105016);
			5601: out = 24'(-56384);
			5602: out = 24'(52540);
			5603: out = 24'(62848);
			5604: out = 24'(19780);
			5605: out = 24'(12548);
			5606: out = 24'(8240);
			5607: out = 24'(-31872);
			5608: out = 24'(-95368);
			5609: out = 24'(-41488);
			5610: out = 24'(40032);
			5611: out = 24'(46996);
			5612: out = 24'(9136);
			5613: out = 24'(56044);
			5614: out = 24'(61572);
			5615: out = 24'(-20828);
			5616: out = 24'(-85544);
			5617: out = 24'(-16080);
			5618: out = 24'(28856);
			5619: out = 24'(-28772);
			5620: out = 24'(6352);
			5621: out = 24'(36160);
			5622: out = 24'(37312);
			5623: out = 24'(-22104);
			5624: out = 24'(-9720);
			5625: out = 24'(16108);
			5626: out = 24'(50760);
			5627: out = 24'(5764);
			5628: out = 24'(-56840);
			5629: out = 24'(-84624);
			5630: out = 24'(-28980);
			5631: out = 24'(496);
			5632: out = 24'(-5148);
			5633: out = 24'(38976);
			5634: out = 24'(69372);
			5635: out = 24'(17236);
			5636: out = 24'(-77464);
			5637: out = 24'(-91920);
			5638: out = 24'(-100);
			5639: out = 24'(67280);
			5640: out = 24'(53932);
			5641: out = 24'(22252);
			5642: out = 24'(6444);
			5643: out = 24'(-17464);
			5644: out = 24'(-21800);
			5645: out = 24'(39176);
			5646: out = 24'(46760);
			5647: out = 24'(13588);
			5648: out = 24'(-37372);
			5649: out = 24'(-49860);
			5650: out = 24'(-8608);
			5651: out = 24'(16856);
			5652: out = 24'(16976);
			5653: out = 24'(4748);
			5654: out = 24'(4620);
			5655: out = 24'(-37896);
			5656: out = 24'(-39788);
			5657: out = 24'(11464);
			5658: out = 24'(28628);
			5659: out = 24'(-11996);
			5660: out = 24'(-21176);
			5661: out = 24'(48876);
			5662: out = 24'(88484);
			5663: out = 24'(67672);
			5664: out = 24'(-41036);
			5665: out = 24'(-120064);
			5666: out = 24'(-111476);
			5667: out = 24'(-85680);
			5668: out = 24'(-32932);
			5669: out = 24'(46420);
			5670: out = 24'(112256);
			5671: out = 24'(59980);
			5672: out = 24'(-15240);
			5673: out = 24'(-93256);
			5674: out = 24'(-106972);
			5675: out = 24'(-53564);
			5676: out = 24'(43272);
			5677: out = 24'(89048);
			5678: out = 24'(73732);
			5679: out = 24'(8576);
			5680: out = 24'(-53148);
			5681: out = 24'(-71904);
			5682: out = 24'(3688);
			5683: out = 24'(96376);
			5684: out = 24'(75808);
			5685: out = 24'(-28276);
			5686: out = 24'(-109024);
			5687: out = 24'(-64972);
			5688: out = 24'(-23420);
			5689: out = 24'(51740);
			5690: out = 24'(95236);
			5691: out = 24'(67916);
			5692: out = 24'(-84960);
			5693: out = 24'(-128472);
			5694: out = 24'(-68900);
			5695: out = 24'(53232);
			5696: out = 24'(63480);
			5697: out = 24'(89996);
			5698: out = 24'(72632);
			5699: out = 24'(4392);
			5700: out = 24'(-101848);
			5701: out = 24'(-93852);
			5702: out = 24'(-10060);
			5703: out = 24'(49688);
			5704: out = 24'(37032);
			5705: out = 24'(25888);
			5706: out = 24'(22220);
			5707: out = 24'(12248);
			5708: out = 24'(-14740);
			5709: out = 24'(-37032);
			5710: out = 24'(-788);
			5711: out = 24'(29460);
			5712: out = 24'(12060);
			5713: out = 24'(-33144);
			5714: out = 24'(4480);
			5715: out = 24'(36372);
			5716: out = 24'(160);
			5717: out = 24'(-67048);
			5718: out = 24'(-51612);
			5719: out = 24'(25264);
			5720: out = 24'(71364);
			5721: out = 24'(55324);
			5722: out = 24'(13540);
			5723: out = 24'(-32572);
			5724: out = 24'(-51748);
			5725: out = 24'(-14464);
			5726: out = 24'(32812);
			5727: out = 24'(67400);
			5728: out = 24'(28628);
			5729: out = 24'(-48736);
			5730: out = 24'(-65284);
			5731: out = 24'(-42648);
			5732: out = 24'(-796);
			5733: out = 24'(26052);
			5734: out = 24'(20480);
			5735: out = 24'(11948);
			5736: out = 24'(-13044);
			5737: out = 24'(-21900);
			5738: out = 24'(-16076);
			5739: out = 24'(78308);
			5740: out = 24'(54276);
			5741: out = 24'(-25424);
			5742: out = 24'(-75912);
			5743: out = 24'(25808);
			5744: out = 24'(43520);
			5745: out = 24'(5752);
			5746: out = 24'(-22908);
			5747: out = 24'(12924);
			5748: out = 24'(6276);
			5749: out = 24'(-844);
			5750: out = 24'(-13740);
			5751: out = 24'(-46492);
			5752: out = 24'(-37380);
			5753: out = 24'(38428);
			5754: out = 24'(78988);
			5755: out = 24'(33248);
			5756: out = 24'(-8676);
			5757: out = 24'(21252);
			5758: out = 24'(24948);
			5759: out = 24'(-79488);
			5760: out = 24'(-76096);
			5761: out = 24'(33328);
			5762: out = 24'(110108);
			5763: out = 24'(28700);
			5764: out = 24'(-37268);
			5765: out = 24'(-109448);
			5766: out = 24'(-87848);
			5767: out = 24'(-24196);
			5768: out = 24'(64520);
			5769: out = 24'(70216);
			5770: out = 24'(53760);
			5771: out = 24'(6468);
			5772: out = 24'(2504);
			5773: out = 24'(-47908);
			5774: out = 24'(14384);
			5775: out = 24'(83468);
			5776: out = 24'(63436);
			5777: out = 24'(-53056);
			5778: out = 24'(-109304);
			5779: out = 24'(-77036);
			5780: out = 24'(-4704);
			5781: out = 24'(25824);
			5782: out = 24'(60504);
			5783: out = 24'(39652);
			5784: out = 24'(-16472);
			5785: out = 24'(-13468);
			5786: out = 24'(13588);
			5787: out = 24'(488);
			5788: out = 24'(-20592);
			5789: out = 24'(77516);
			5790: out = 24'(66656);
			5791: out = 24'(3376);
			5792: out = 24'(-77588);
			5793: out = 24'(-64544);
			5794: out = 24'(-81180);
			5795: out = 24'(-36536);
			5796: out = 24'(32400);
			5797: out = 24'(74488);
			5798: out = 24'(-6400);
			5799: out = 24'(-60016);
			5800: out = 24'(-39436);
			5801: out = 24'(32852);
			5802: out = 24'(10480);
			5803: out = 24'(364);
			5804: out = 24'(3812);
			5805: out = 24'(23240);
			5806: out = 24'(1284);
			5807: out = 24'(-32244);
			5808: out = 24'(-73944);
			5809: out = 24'(-65588);
			5810: out = 24'(9872);
			5811: out = 24'(4308);
			5812: out = 24'(5368);
			5813: out = 24'(53288);
			5814: out = 24'(108232);
			5815: out = 24'(25492);
			5816: out = 24'(-72588);
			5817: out = 24'(-110372);
			5818: out = 24'(-34540);
			5819: out = 24'(65992);
			5820: out = 24'(97196);
			5821: out = 24'(54452);
			5822: out = 24'(-3632);
			5823: out = 24'(-16584);
			5824: out = 24'(-2000);
			5825: out = 24'(11568);
			5826: out = 24'(-3164);
			5827: out = 24'(-50392);
			5828: out = 24'(-39824);
			5829: out = 24'(-22052);
			5830: out = 24'(-13372);
			5831: out = 24'(10632);
			5832: out = 24'(65324);
			5833: out = 24'(92216);
			5834: out = 24'(57208);
			5835: out = 24'(-7208);
			5836: out = 24'(-108452);
			5837: out = 24'(-60500);
			5838: out = 24'(43720);
			5839: out = 24'(72084);
			5840: out = 24'(12836);
			5841: out = 24'(104);
			5842: out = 24'(-10688);
			5843: out = 24'(-43952);
			5844: out = 24'(-78840);
			5845: out = 24'(-23900);
			5846: out = 24'(54312);
			5847: out = 24'(70272);
			5848: out = 24'(20068);
			5849: out = 24'(9232);
			5850: out = 24'(29756);
			5851: out = 24'(57548);
			5852: out = 24'(28948);
			5853: out = 24'(-44900);
			5854: out = 24'(-107000);
			5855: out = 24'(-53136);
			5856: out = 24'(45280);
			5857: out = 24'(38488);
			5858: out = 24'(-70776);
			5859: out = 24'(-94240);
			5860: out = 24'(30464);
			5861: out = 24'(91576);
			5862: out = 24'(76932);
			5863: out = 24'(33052);
			5864: out = 24'(2004);
			5865: out = 24'(-57796);
			5866: out = 24'(-107876);
			5867: out = 24'(-92700);
			5868: out = 24'(5368);
			5869: out = 24'(62244);
			5870: out = 24'(72488);
			5871: out = 24'(25672);
			5872: out = 24'(-6116);
			5873: out = 24'(-11640);
			5874: out = 24'(8976);
			5875: out = 24'(-20344);
			5876: out = 24'(-43668);
			5877: out = 24'(-35692);
			5878: out = 24'(-31180);
			5879: out = 24'(-3128);
			5880: out = 24'(36300);
			5881: out = 24'(61988);
			5882: out = 24'(48164);
			5883: out = 24'(412);
			5884: out = 24'(-33716);
			5885: out = 24'(-36612);
			5886: out = 24'(-30416);
			5887: out = 24'(-2768);
			5888: out = 24'(25328);
			5889: out = 24'(39176);
			5890: out = 24'(16712);
			5891: out = 24'(2552);
			5892: out = 24'(-29336);
			5893: out = 24'(-26532);
			5894: out = 24'(12220);
			5895: out = 24'(2348);
			5896: out = 24'(26952);
			5897: out = 24'(51328);
			5898: out = 24'(63124);
			5899: out = 24'(44944);
			5900: out = 24'(22408);
			5901: out = 24'(-45380);
			5902: out = 24'(-119888);
			5903: out = 24'(-106976);
			5904: out = 24'(-38360);
			5905: out = 24'(62108);
			5906: out = 24'(95536);
			5907: out = 24'(77032);
			5908: out = 24'(40576);
			5909: out = 24'(26292);
			5910: out = 24'(-16152);
			5911: out = 24'(-76524);
			5912: out = 24'(-63148);
			5913: out = 24'(27160);
			5914: out = 24'(69872);
			5915: out = 24'(14936);
			5916: out = 24'(-93720);
			5917: out = 24'(-62880);
			5918: out = 24'(27160);
			5919: out = 24'(44472);
			5920: out = 24'(5664);
			5921: out = 24'(-37300);
			5922: out = 24'(-36224);
			5923: out = 24'(-3596);
			5924: out = 24'(40096);
			5925: out = 24'(42008);
			5926: out = 24'(47792);
			5927: out = 24'(37208);
			5928: out = 24'(1752);
			5929: out = 24'(-44336);
			5930: out = 24'(-43072);
			5931: out = 24'(10784);
			5932: out = 24'(50616);
			5933: out = 24'(35592);
			5934: out = 24'(-64404);
			5935: out = 24'(-120816);
			5936: out = 24'(-58704);
			5937: out = 24'(27580);
			5938: out = 24'(72868);
			5939: out = 24'(40172);
			5940: out = 24'(2132);
			5941: out = 24'(-14244);
			5942: out = 24'(-7200);
			5943: out = 24'(-42456);
			5944: out = 24'(-55900);
			5945: out = 24'(9388);
			5946: out = 24'(69376);
			5947: out = 24'(66600);
			5948: out = 24'(35452);
			5949: out = 24'(18280);
			5950: out = 24'(9252);
			5951: out = 24'(-37448);
			5952: out = 24'(-96800);
			5953: out = 24'(-114036);
			5954: out = 24'(-34592);
			5955: out = 24'(29600);
			5956: out = 24'(79384);
			5957: out = 24'(93212);
			5958: out = 24'(53948);
			5959: out = 24'(-38916);
			5960: out = 24'(-65788);
			5961: out = 24'(-18116);
			5962: out = 24'(-4380);
			5963: out = 24'(-11040);
			5964: out = 24'(-13412);
			5965: out = 24'(12844);
			5966: out = 24'(16588);
			5967: out = 24'(-2932);
			5968: out = 24'(-3544);
			5969: out = 24'(41672);
			5970: out = 24'(56064);
			5971: out = 24'(-38308);
			5972: out = 24'(-116900);
			5973: out = 24'(-81028);
			5974: out = 24'(42244);
			5975: out = 24'(84360);
			5976: out = 24'(50604);
			5977: out = 24'(4540);
			5978: out = 24'(-39684);
			5979: out = 24'(-69212);
			5980: out = 24'(-8912);
			5981: out = 24'(89888);
			5982: out = 24'(85364);
			5983: out = 24'(-40508);
			5984: out = 24'(-106492);
			5985: out = 24'(-59452);
			5986: out = 24'(22248);
			5987: out = 24'(13088);
			5988: out = 24'(62208);
			5989: out = 24'(54896);
			5990: out = 24'(40652);
			5991: out = 24'(-2956);
			5992: out = 24'(-13144);
			5993: out = 24'(-27116);
			5994: out = 24'(-3864);
			5995: out = 24'(1516);
			5996: out = 24'(-1304);
			5997: out = 24'(-9024);
			5998: out = 24'(44724);
			5999: out = 24'(74660);
			6000: out = 24'(41676);
			6001: out = 24'(-39708);
			6002: out = 24'(-34416);
			6003: out = 24'(9752);
			6004: out = 24'(-812);
			6005: out = 24'(-45388);
			6006: out = 24'(-10904);
			6007: out = 24'(57924);
			6008: out = 24'(47364);
			6009: out = 24'(11484);
			6010: out = 24'(-73768);
			6011: out = 24'(-64368);
			6012: out = 24'(12876);
			6013: out = 24'(21236);
			6014: out = 24'(-4792);
			6015: out = 24'(-22132);
			6016: out = 24'(8816);
			6017: out = 24'(32760);
			6018: out = 24'(51696);
			6019: out = 24'(7716);
			6020: out = 24'(-16508);
			6021: out = 24'(21424);
			6022: out = 24'(17676);
			6023: out = 24'(-8244);
			6024: out = 24'(-28032);
			6025: out = 24'(7256);
			6026: out = 24'(16300);
			6027: out = 24'(15824);
			6028: out = 24'(-29276);
			6029: out = 24'(-49832);
			6030: out = 24'(-27932);
			6031: out = 24'(25172);
			6032: out = 24'(6732);
			6033: out = 24'(-11920);
			6034: out = 24'(33252);
			6035: out = 24'(14192);
			6036: out = 24'(-55624);
			6037: out = 24'(-69532);
			6038: out = 24'(42196);
			6039: out = 24'(38512);
			6040: out = 24'(9980);
			6041: out = 24'(1040);
			6042: out = 24'(32256);
			6043: out = 24'(27076);
			6044: out = 24'(-44732);
			6045: out = 24'(-89172);
			6046: out = 24'(-40020);
			6047: out = 24'(1788);
			6048: out = 24'(7976);
			6049: out = 24'(13696);
			6050: out = 24'(47044);
			6051: out = 24'(46808);
			6052: out = 24'(-13620);
			6053: out = 24'(-54600);
			6054: out = 24'(-9760);
			6055: out = 24'(56872);
			6056: out = 24'(5620);
			6057: out = 24'(-39992);
			6058: out = 24'(-7992);
			6059: out = 24'(60956);
			6060: out = 24'(7844);
			6061: out = 24'(-7824);
			6062: out = 24'(24528);
			6063: out = 24'(54544);
			6064: out = 24'(-15108);
			6065: out = 24'(-39992);
			6066: out = 24'(-24996);
			6067: out = 24'(544);
			6068: out = 24'(-19604);
			6069: out = 24'(-16944);
			6070: out = 24'(6260);
			6071: out = 24'(22412);
			6072: out = 24'(-8488);
			6073: out = 24'(-16896);
			6074: out = 24'(-1872);
			6075: out = 24'(30236);
			6076: out = 24'(29408);
			6077: out = 24'(-7092);
			6078: out = 24'(-58792);
			6079: out = 24'(-59984);
			6080: out = 24'(6836);
			6081: out = 24'(44472);
			6082: out = 24'(87828);
			6083: out = 24'(81312);
			6084: out = 24'(28464);
			6085: out = 24'(-76424);
			6086: out = 24'(-87896);
			6087: out = 24'(-51188);
			6088: out = 24'(-14252);
			6089: out = 24'(-19220);
			6090: out = 24'(39588);
			6091: out = 24'(52636);
			6092: out = 24'(26124);
			6093: out = 24'(-21176);
			6094: out = 24'(-536);
			6095: out = 24'(-21528);
			6096: out = 24'(-38604);
			6097: out = 24'(-164);
			6098: out = 24'(84432);
			6099: out = 24'(72640);
			6100: out = 24'(928);
			6101: out = 24'(-67952);
			6102: out = 24'(-76532);
			6103: out = 24'(-37468);
			6104: out = 24'(19072);
			6105: out = 24'(48952);
			6106: out = 24'(45888);
			6107: out = 24'(10800);
			6108: out = 24'(-3700);
			6109: out = 24'(-284);
			6110: out = 24'(-188);
			6111: out = 24'(-1052);
			6112: out = 24'(10328);
			6113: out = 24'(14364);
			6114: out = 24'(-3576);
			6115: out = 24'(-14108);
			6116: out = 24'(19896);
			6117: out = 24'(45760);
			6118: out = 24'(-2872);
			6119: out = 24'(-89084);
			6120: out = 24'(-128472);
			6121: out = 24'(-71648);
			6122: out = 24'(13324);
			6123: out = 24'(38680);
			6124: out = 24'(35184);
			6125: out = 24'(58692);
			6126: out = 24'(65568);
			6127: out = 24'(2964);
			6128: out = 24'(-52492);
			6129: out = 24'(-72104);
			6130: out = 24'(-51772);
			6131: out = 24'(-29928);
			6132: out = 24'(-3124);
			6133: out = 24'(40680);
			6134: out = 24'(66856);
			6135: out = 24'(44148);
			6136: out = 24'(7828);
			6137: out = 24'(-39764);
			6138: out = 24'(-74856);
			6139: out = 24'(-70412);
			6140: out = 24'(13776);
			6141: out = 24'(35936);
			6142: out = 24'(15520);
			6143: out = 24'(-2744);
			6144: out = 24'(13748);
			6145: out = 24'(12880);
			6146: out = 24'(180);
			6147: out = 24'(20016);
			6148: out = 24'(72308);
			6149: out = 24'(9228);
			6150: out = 24'(-75352);
			6151: out = 24'(-87680);
			6152: out = 24'(18184);
			6153: out = 24'(38020);
			6154: out = 24'(39084);
			6155: out = 24'(29728);
			6156: out = 24'(28196);
			6157: out = 24'(-3608);
			6158: out = 24'(-26932);
			6159: out = 24'(-23248);
			6160: out = 24'(8256);
			6161: out = 24'(34148);
			6162: out = 24'(-26176);
			6163: out = 24'(-60328);
			6164: out = 24'(-9832);
			6165: out = 24'(73744);
			6166: out = 24'(24740);
			6167: out = 24'(552);
			6168: out = 24'(35360);
			6169: out = 24'(66660);
			6170: out = 24'(-23488);
			6171: out = 24'(-94200);
			6172: out = 24'(-73536);
			6173: out = 24'(24856);
			6174: out = 24'(51496);
			6175: out = 24'(77024);
			6176: out = 24'(78008);
			6177: out = 24'(52240);
			6178: out = 24'(-1516);
			6179: out = 24'(-91752);
			6180: out = 24'(-121560);
			6181: out = 24'(-102000);
			6182: out = 24'(-8892);
			6183: out = 24'(63016);
			6184: out = 24'(84248);
			6185: out = 24'(54616);
			6186: out = 24'(-9196);
			6187: out = 24'(-31208);
			6188: out = 24'(-21428);
			6189: out = 24'(-2092);
			6190: out = 24'(-1760);
			6191: out = 24'(7648);
			6192: out = 24'(1824);
			6193: out = 24'(1232);
			6194: out = 24'(7956);
			6195: out = 24'(5908);
			6196: out = 24'(2968);
			6197: out = 24'(5124);
			6198: out = 24'(24264);
			6199: out = 24'(24200);
			6200: out = 24'(-1352);
			6201: out = 24'(-56624);
			6202: out = 24'(-62140);
			6203: out = 24'(-3960);
			6204: out = 24'(11812);
			6205: out = 24'(-29460);
			6206: out = 24'(-43400);
			6207: out = 24'(-4416);
			6208: out = 24'(23036);
			6209: out = 24'(-14664);
			6210: out = 24'(-7076);
			6211: out = 24'(60868);
			6212: out = 24'(83740);
			6213: out = 24'(-14808);
			6214: out = 24'(-76436);
			6215: out = 24'(-18208);
			6216: out = 24'(39092);
			6217: out = 24'(63004);
			6218: out = 24'(48060);
			6219: out = 24'(12532);
			6220: out = 24'(-39448);
			6221: out = 24'(-106080);
			6222: out = 24'(-67288);
			6223: out = 24'(27208);
			6224: out = 24'(47372);
			6225: out = 24'(16564);
			6226: out = 24'(16608);
			6227: out = 24'(30984);
			6228: out = 24'(3120);
			6229: out = 24'(-44012);
			6230: out = 24'(-56760);
			6231: out = 24'(-27996);
			6232: out = 24'(9344);
			6233: out = 24'(49924);
			6234: out = 24'(80552);
			6235: out = 24'(69512);
			6236: out = 24'(10796);
			6237: out = 24'(-64192);
			6238: out = 24'(-56568);
			6239: out = 24'(180);
			6240: out = 24'(39960);
			6241: out = 24'(17544);
			6242: out = 24'(-1676);
			6243: out = 24'(-66968);
			6244: out = 24'(-108380);
			6245: out = 24'(-73436);
			6246: out = 24'(12044);
			6247: out = 24'(57072);
			6248: out = 24'(61960);
			6249: out = 24'(47060);
			6250: out = 24'(23140);
			6251: out = 24'(-14000);
			6252: out = 24'(-29656);
			6253: out = 24'(-25684);
			6254: out = 24'(-18700);
			6255: out = 24'(-40684);
			6256: out = 24'(-26240);
			6257: out = 24'(15120);
			6258: out = 24'(36892);
			6259: out = 24'(37160);
			6260: out = 24'(45876);
			6261: out = 24'(42208);
			6262: out = 24'(-2848);
			6263: out = 24'(-89608);
			6264: out = 24'(-111624);
			6265: out = 24'(-60816);
			6266: out = 24'(5376);
			6267: out = 24'(59724);
			6268: out = 24'(71128);
			6269: out = 24'(50264);
			6270: out = 24'(13420);
			6271: out = 24'(9260);
			6272: out = 24'(-25848);
			6273: out = 24'(-62060);
			6274: out = 24'(-76712);
			6275: out = 24'(-15032);
			6276: out = 24'(1444);
			6277: out = 24'(36368);
			6278: out = 24'(55312);
			6279: out = 24'(44332);
			6280: out = 24'(-7520);
			6281: out = 24'(-27832);
			6282: out = 24'(-15292);
			6283: out = 24'(10624);
			6284: out = 24'(6820);
			6285: out = 24'(9752);
			6286: out = 24'(-1992);
			6287: out = 24'(-9972);
			6288: out = 24'(-428);
			6289: out = 24'(13680);
			6290: out = 24'(6460);
			6291: out = 24'(7380);
			6292: out = 24'(32512);
			6293: out = 24'(20540);
			6294: out = 24'(-35088);
			6295: out = 24'(-57004);
			6296: out = 24'(10028);
			6297: out = 24'(52624);
			6298: out = 24'(18188);
			6299: out = 24'(-29168);
			6300: out = 24'(-12800);
			6301: out = 24'(23080);
			6302: out = 24'(19780);
			6303: out = 24'(-1292);
			6304: out = 24'(376);
			6305: out = 24'(-7652);
			6306: out = 24'(-24792);
			6307: out = 24'(-24832);
			6308: out = 24'(5820);
			6309: out = 24'(-1000);
			6310: out = 24'(7404);
			6311: out = 24'(27980);
			6312: out = 24'(64568);
			6313: out = 24'(41420);
			6314: out = 24'(13204);
			6315: out = 24'(-72660);
			6316: out = 24'(-106884);
			6317: out = 24'(-48164);
			6318: out = 24'(35960);
			6319: out = 24'(53792);
			6320: out = 24'(51932);
			6321: out = 24'(37152);
			6322: out = 24'(-3064);
			6323: out = 24'(-84428);
			6324: out = 24'(-78728);
			6325: out = 24'(23280);
			6326: out = 24'(19684);
			6327: out = 24'(12208);
			6328: out = 24'(2824);
			6329: out = 24'(23796);
			6330: out = 24'(-4188);
			6331: out = 24'(6312);
			6332: out = 24'(-5128);
			6333: out = 24'(13016);
			6334: out = 24'(18444);
			6335: out = 24'(24120);
			6336: out = 24'(-53684);
			6337: out = 24'(-114388);
			6338: out = 24'(-105368);
			6339: out = 24'(-26504);
			6340: out = 24'(12692);
			6341: out = 24'(59908);
			6342: out = 24'(91384);
			6343: out = 24'(64228);
			6344: out = 24'(-13556);
			6345: out = 24'(-18976);
			6346: out = 24'(29488);
			6347: out = 24'(408);
			6348: out = 24'(-55596);
			6349: out = 24'(-41116);
			6350: out = 24'(44136);
			6351: out = 24'(50188);
			6352: out = 24'(55168);
			6353: out = 24'(30332);
			6354: out = 24'(17396);
			6355: out = 24'(-23356);
			6356: out = 24'(-80716);
			6357: out = 24'(-115120);
			6358: out = 24'(-66940);
			6359: out = 24'(14356);
			6360: out = 24'(76636);
			6361: out = 24'(56376);
			6362: out = 24'(37220);
			6363: out = 24'(28720);
			6364: out = 24'(21676);
			6365: out = 24'(-37476);
			6366: out = 24'(-58240);
			6367: out = 24'(-8684);
			6368: out = 24'(59264);
			6369: out = 24'(50892);
			6370: out = 24'(-3572);
			6371: out = 24'(-77668);
			6372: out = 24'(-106816);
			6373: out = 24'(-39948);
			6374: out = 24'(56292);
			6375: out = 24'(59992);
			6376: out = 24'(9156);
			6377: out = 24'(4172);
			6378: out = 24'(52980);
			6379: out = 24'(37664);
			6380: out = 24'(-44704);
			6381: out = 24'(-85372);
			6382: out = 24'(-7376);
			6383: out = 24'(57640);
			6384: out = 24'(33012);
			6385: out = 24'(-7124);
			6386: out = 24'(-23860);
			6387: out = 24'(-39376);
			6388: out = 24'(-59856);
			6389: out = 24'(-32576);
			6390: out = 24'(18360);
			6391: out = 24'(49184);
			6392: out = 24'(40804);
			6393: out = 24'(19700);
			6394: out = 24'(11416);
			6395: out = 24'(-8508);
			6396: out = 24'(-14040);
			6397: out = 24'(6540);
			6398: out = 24'(29948);
			6399: out = 24'(-19692);
			6400: out = 24'(-57728);
			6401: out = 24'(-11712);
			6402: out = 24'(43452);
			6403: out = 24'(26920);
			6404: out = 24'(-34612);
			6405: out = 24'(-26964);
			6406: out = 24'(61216);
			6407: out = 24'(41488);
			6408: out = 24'(-67308);
			6409: out = 24'(-114820);
			6410: out = 24'(-27544);
			6411: out = 24'(79936);
			6412: out = 24'(46448);
			6413: out = 24'(-13368);
			6414: out = 24'(-8396);
			6415: out = 24'(55252);
			6416: out = 24'(4548);
			6417: out = 24'(-69760);
			6418: out = 24'(-44876);
			6419: out = 24'(49824);
			6420: out = 24'(72780);
			6421: out = 24'(14540);
			6422: out = 24'(-47872);
			6423: out = 24'(-65060);
			6424: out = 24'(-4948);
			6425: out = 24'(67316);
			6426: out = 24'(95948);
			6427: out = 24'(53988);
			6428: out = 24'(612);
			6429: out = 24'(-63936);
			6430: out = 24'(-71540);
			6431: out = 24'(-15568);
			6432: out = 24'(5648);
			6433: out = 24'(5116);
			6434: out = 24'(476);
			6435: out = 24'(7536);
			6436: out = 24'(55408);
			6437: out = 24'(32456);
			6438: out = 24'(19172);
			6439: out = 24'(32256);
			6440: out = 24'(26676);
			6441: out = 24'(-39272);
			6442: out = 24'(-84756);
			6443: out = 24'(-46308);
			6444: out = 24'(13944);
			6445: out = 24'(26996);
			6446: out = 24'(2524);
			6447: out = 24'(18780);
			6448: out = 24'(57440);
			6449: out = 24'(35708);
			6450: out = 24'(-47592);
			6451: out = 24'(-83884);
			6452: out = 24'(-6888);
			6453: out = 24'(27776);
			6454: out = 24'(20464);
			6455: out = 24'(-24388);
			6456: out = 24'(-39880);
			6457: out = 24'(-3736);
			6458: out = 24'(29688);
			6459: out = 24'(42716);
			6460: out = 24'(47540);
			6461: out = 24'(44000);
			6462: out = 24'(34628);
			6463: out = 24'(1108);
			6464: out = 24'(-44936);
			6465: out = 24'(-76328);
			6466: out = 24'(-81284);
			6467: out = 24'(-39424);
			6468: out = 24'(18656);
			6469: out = 24'(52800);
			6470: out = 24'(33548);
			6471: out = 24'(24464);
			6472: out = 24'(-1192);
			6473: out = 24'(-63716);
			6474: out = 24'(-115208);
			6475: out = 24'(-75868);
			6476: out = 24'(32712);
			6477: out = 24'(90280);
			6478: out = 24'(77116);
			6479: out = 24'(42492);
			6480: out = 24'(4256);
			6481: out = 24'(-46944);
			6482: out = 24'(-95604);
			6483: out = 24'(-99952);
			6484: out = 24'(-38052);
			6485: out = 24'(24840);
			6486: out = 24'(49816);
			6487: out = 24'(8336);
			6488: out = 24'(25900);
			6489: out = 24'(36996);
			6490: out = 24'(16392);
			6491: out = 24'(-15368);
			6492: out = 24'(-15688);
			6493: out = 24'(-39356);
			6494: out = 24'(-69316);
			6495: out = 24'(-16940);
			6496: out = 24'(58804);
			6497: out = 24'(77360);
			6498: out = 24'(37284);
			6499: out = 24'(-2508);
			6500: out = 24'(-6328);
			6501: out = 24'(-13624);
			6502: out = 24'(-31492);
			6503: out = 24'(-42592);
			6504: out = 24'(-2964);
			6505: out = 24'(-13788);
			6506: out = 24'(-29260);
			6507: out = 24'(2800);
			6508: out = 24'(67180);
			6509: out = 24'(87208);
			6510: out = 24'(70368);
			6511: out = 24'(26996);
			6512: out = 24'(-32152);
			6513: out = 24'(-62712);
			6514: out = 24'(-32524);
			6515: out = 24'(-1304);
			6516: out = 24'(-29672);
			6517: out = 24'(-68048);
			6518: out = 24'(-9528);
			6519: out = 24'(96376);
			6520: out = 24'(101628);
			6521: out = 24'(32380);
			6522: out = 24'(-37500);
			6523: out = 24'(-46948);
			6524: out = 24'(-31968);
			6525: out = 24'(2696);
			6526: out = 24'(12);
			6527: out = 24'(14816);
			6528: out = 24'(19656);
			6529: out = 24'(-17164);
			6530: out = 24'(-37744);
			6531: out = 24'(14000);
			6532: out = 24'(71004);
			6533: out = 24'(34988);
			6534: out = 24'(9636);
			6535: out = 24'(-2156);
			6536: out = 24'(-7796);
			6537: out = 24'(-45568);
			6538: out = 24'(-20204);
			6539: out = 24'(9732);
			6540: out = 24'(12660);
			6541: out = 24'(-18860);
			6542: out = 24'(-2028);
			6543: out = 24'(15180);
			6544: out = 24'(13420);
			6545: out = 24'(-5724);
			6546: out = 24'(6864);
			6547: out = 24'(28872);
			6548: out = 24'(26792);
			6549: out = 24'(-10384);
			6550: out = 24'(-48108);
			6551: out = 24'(-34624);
			6552: out = 24'(21636);
			6553: out = 24'(72880);
			6554: out = 24'(68040);
			6555: out = 24'(23092);
			6556: out = 24'(-64624);
			6557: out = 24'(-102748);
			6558: out = 24'(-36584);
			6559: out = 24'(3008);
			6560: out = 24'(-12184);
			6561: out = 24'(-25572);
			6562: out = 24'(20152);
			6563: out = 24'(65352);
			6564: out = 24'(15476);
			6565: out = 24'(-72444);
			6566: out = 24'(-86356);
			6567: out = 24'(-3228);
			6568: out = 24'(48800);
			6569: out = 24'(26936);
			6570: out = 24'(756);
			6571: out = 24'(-6744);
			6572: out = 24'(41424);
			6573: out = 24'(16124);
			6574: out = 24'(-36672);
			6575: out = 24'(-38936);
			6576: out = 24'(36300);
			6577: out = 24'(35904);
			6578: out = 24'(-21668);
			6579: out = 24'(-46092);
			6580: out = 24'(-32668);
			6581: out = 24'(-1788);
			6582: out = 24'(9840);
			6583: out = 24'(37140);
			6584: out = 24'(56552);
			6585: out = 24'(71344);
			6586: out = 24'(21688);
			6587: out = 24'(-36476);
			6588: out = 24'(-19484);
			6589: out = 24'(19208);
			6590: out = 24'(22224);
			6591: out = 24'(-12088);
			6592: out = 24'(-43456);
			6593: out = 24'(-22200);
			6594: out = 24'(6808);
			6595: out = 24'(26792);
			6596: out = 24'(36132);
			6597: out = 24'(51836);
			6598: out = 24'(7752);
			6599: out = 24'(-49908);
			6600: out = 24'(-71720);
			6601: out = 24'(-26804);
			6602: out = 24'(-4240);
			6603: out = 24'(13540);
			6604: out = 24'(49608);
			6605: out = 24'(96164);
			6606: out = 24'(33768);
			6607: out = 24'(-52212);
			6608: out = 24'(-96572);
			6609: out = 24'(-33604);
			6610: out = 24'(-48828);
			6611: out = 24'(-30348);
			6612: out = 24'(25516);
			6613: out = 24'(72592);
			6614: out = 24'(56536);
			6615: out = 24'(33824);
			6616: out = 24'(1404);
			6617: out = 24'(-34628);
			6618: out = 24'(-28644);
			6619: out = 24'(-12868);
			6620: out = 24'(-11312);
			6621: out = 24'(-24828);
			6622: out = 24'(1424);
			6623: out = 24'(6732);
			6624: out = 24'(6236);
			6625: out = 24'(-1240);
			6626: out = 24'(-3888);
			6627: out = 24'(37296);
			6628: out = 24'(51632);
			6629: out = 24'(-3712);
			6630: out = 24'(-106984);
			6631: out = 24'(-62860);
			6632: out = 24'(4320);
			6633: out = 24'(6552);
			6634: out = 24'(-39556);
			6635: out = 24'(36296);
			6636: out = 24'(71664);
			6637: out = 24'(53504);
			6638: out = 24'(10308);
			6639: out = 24'(19872);
			6640: out = 24'(-20992);
			6641: out = 24'(-71116);
			6642: out = 24'(-84492);
			6643: out = 24'(-49044);
			6644: out = 24'(28272);
			6645: out = 24'(59976);
			6646: out = 24'(54224);
			6647: out = 24'(30848);
			6648: out = 24'(67616);
			6649: out = 24'(23444);
			6650: out = 24'(-68068);
			6651: out = 24'(-113876);
			6652: out = 24'(-54696);
			6653: out = 24'(7564);
			6654: out = 24'(28240);
			6655: out = 24'(41380);
			6656: out = 24'(51668);
			6657: out = 24'(7788);
			6658: out = 24'(-51140);
			6659: out = 24'(-52376);
			6660: out = 24'(29228);
			6661: out = 24'(49156);
			6662: out = 24'(21876);
			6663: out = 24'(716);
			6664: out = 24'(6812);
			6665: out = 24'(19188);
			6666: out = 24'(9248);
			6667: out = 24'(3132);
			6668: out = 24'(17332);
			6669: out = 24'(-15444);
			6670: out = 24'(-54476);
			6671: out = 24'(-50684);
			6672: out = 24'(11340);
			6673: out = 24'(-27476);
			6674: out = 24'(-19220);
			6675: out = 24'(27188);
			6676: out = 24'(80084);
			6677: out = 24'(35720);
			6678: out = 24'(30788);
			6679: out = 24'(14576);
			6680: out = 24'(3860);
			6681: out = 24'(-22416);
			6682: out = 24'(-17424);
			6683: out = 24'(-32568);
			6684: out = 24'(-31752);
			6685: out = 24'(2828);
			6686: out = 24'(61916);
			6687: out = 24'(60672);
			6688: out = 24'(38044);
			6689: out = 24'(25528);
			6690: out = 24'(5184);
			6691: out = 24'(-70736);
			6692: out = 24'(-122856);
			6693: out = 24'(-92740);
			6694: out = 24'(-18092);
			6695: out = 24'(19376);
			6696: out = 24'(32836);
			6697: out = 24'(71976);
			6698: out = 24'(93696);
			6699: out = 24'(86060);
			6700: out = 24'(6512);
			6701: out = 24'(-96372);
			6702: out = 24'(-119168);
			6703: out = 24'(-90696);
			6704: out = 24'(-25280);
			6705: out = 24'(30916);
			6706: out = 24'(74464);
			6707: out = 24'(73508);
			6708: out = 24'(43436);
			6709: out = 24'(-3536);
			6710: out = 24'(-41176);
			6711: out = 24'(-35504);
			6712: out = 24'(-23716);
			6713: out = 24'(-18348);
			6714: out = 24'(-12972);
			6715: out = 24'(30192);
			6716: out = 24'(43968);
			6717: out = 24'(36304);
			6718: out = 24'(4600);
			6719: out = 24'(4492);
			6720: out = 24'(-16944);
			6721: out = 24'(6192);
			6722: out = 24'(14544);
			6723: out = 24'(7720);
			6724: out = 24'(-88140);
			6725: out = 24'(-45088);
			6726: out = 24'(47024);
			6727: out = 24'(53080);
			6728: out = 24'(9328);
			6729: out = 24'(6560);
			6730: out = 24'(19456);
			6731: out = 24'(-1600);
			6732: out = 24'(-15776);
			6733: out = 24'(-9672);
			6734: out = 24'(-3280);
			6735: out = 24'(-27244);
			6736: out = 24'(-34276);
			6737: out = 24'(-14232);
			6738: out = 24'(29604);
			6739: out = 24'(39292);
			6740: out = 24'(6296);
			6741: out = 24'(-14080);
			6742: out = 24'(-30812);
			6743: out = 24'(-40320);
			6744: out = 24'(-26924);
			6745: out = 24'(10964);
			6746: out = 24'(35108);
			6747: out = 24'(33072);
			6748: out = 24'(31592);
			6749: out = 24'(16360);
			6750: out = 24'(8068);
			6751: out = 24'(-44252);
			6752: out = 24'(-96340);
			6753: out = 24'(-55360);
			6754: out = 24'(19424);
			6755: out = 24'(48820);
			6756: out = 24'(25408);
			6757: out = 24'(-15956);
			6758: out = 24'(12824);
			6759: out = 24'(4224);
			6760: out = 24'(-15624);
			6761: out = 24'(28372);
			6762: out = 24'(70792);
			6763: out = 24'(55804);
			6764: out = 24'(-19452);
			6765: out = 24'(-72672);
			6766: out = 24'(-95224);
			6767: out = 24'(-54712);
			6768: out = 24'(-30408);
			6769: out = 24'(-3256);
			6770: out = 24'(40980);
			6771: out = 24'(92804);
			6772: out = 24'(57280);
			6773: out = 24'(-11952);
			6774: out = 24'(-29212);
			6775: out = 24'(32376);
			6776: out = 24'(30076);
			6777: out = 24'(-34800);
			6778: out = 24'(-58476);
			6779: out = 24'(-1084);
			6780: out = 24'(39600);
			6781: out = 24'(28428);
			6782: out = 24'(28992);
			6783: out = 24'(14744);
			6784: out = 24'(30036);
			6785: out = 24'(12956);
			6786: out = 24'(-31228);
			6787: out = 24'(-111940);
			6788: out = 24'(-75312);
			6789: out = 24'(5048);
			6790: out = 24'(63772);
			6791: out = 24'(77988);
			6792: out = 24'(68748);
			6793: out = 24'(9148);
			6794: out = 24'(-48252);
			6795: out = 24'(-51152);
			6796: out = 24'(-5100);
			6797: out = 24'(7572);
			6798: out = 24'(96);
			6799: out = 24'(9824);
			6800: out = 24'(46636);
			6801: out = 24'(-2132);
			6802: out = 24'(-77032);
			6803: out = 24'(-75156);
			6804: out = 24'(2932);
			6805: out = 24'(61240);
			6806: out = 24'(49688);
			6807: out = 24'(12748);
			6808: out = 24'(-16008);
			6809: out = 24'(-33232);
			6810: out = 24'(-34500);
			6811: out = 24'(-656);
			6812: out = 24'(57060);
			6813: out = 24'(22316);
			6814: out = 24'(-40796);
			6815: out = 24'(-60888);
			6816: out = 24'(10480);
			6817: out = 24'(-1280);
			6818: out = 24'(-22128);
			6819: out = 24'(-35172);
			6820: out = 24'(-1636);
			6821: out = 24'(36740);
			6822: out = 24'(76768);
			6823: out = 24'(69028);
			6824: out = 24'(31208);
			6825: out = 24'(-33768);
			6826: out = 24'(-41276);
			6827: out = 24'(-48776);
			6828: out = 24'(-67100);
			6829: out = 24'(-50396);
			6830: out = 24'(-7752);
			6831: out = 24'(31464);
			6832: out = 24'(59264);
			6833: out = 24'(94704);
			6834: out = 24'(68324);
			6835: out = 24'(21780);
			6836: out = 24'(-28324);
			6837: out = 24'(-39296);
			6838: out = 24'(-91704);
			6839: out = 24'(-66800);
			6840: out = 24'(-3964);
			6841: out = 24'(31676);
			6842: out = 24'(28480);
			6843: out = 24'(20428);
			6844: out = 24'(21468);
			6845: out = 24'(14284);
			6846: out = 24'(-7940);
			6847: out = 24'(-21108);
			6848: out = 24'(1628);
			6849: out = 24'(23256);
			6850: out = 24'(-5592);
			6851: out = 24'(-16012);
			6852: out = 24'(-14888);
			6853: out = 24'(-17644);
			6854: out = 24'(-39516);
			6855: out = 24'(32004);
			6856: out = 24'(86832);
			6857: out = 24'(69864);
			6858: out = 24'(-10064);
			6859: out = 24'(-76060);
			6860: out = 24'(-73884);
			6861: out = 24'(-19364);
			6862: out = 24'(7924);
			6863: out = 24'(22488);
			6864: out = 24'(-14688);
			6865: out = 24'(-34740);
			6866: out = 24'(-10816);
			6867: out = 24'(53928);
			6868: out = 24'(52276);
			6869: out = 24'(27184);
			6870: out = 24'(1940);
			6871: out = 24'(272);
			6872: out = 24'(-22860);
			6873: out = 24'(-9908);
			6874: out = 24'(32368);
			6875: out = 24'(64844);
			6876: out = 24'(584);
			6877: out = 24'(-54384);
			6878: out = 24'(-77344);
			6879: out = 24'(-54464);
			6880: out = 24'(-25312);
			6881: out = 24'(26164);
			6882: out = 24'(64612);
			6883: out = 24'(77684);
			6884: out = 24'(53668);
			6885: out = 24'(13156);
			6886: out = 24'(-36336);
			6887: out = 24'(-44620);
			6888: out = 24'(808);
			6889: out = 24'(12192);
			6890: out = 24'(-28832);
			6891: out = 24'(-54456);
			6892: out = 24'(-2396);
			6893: out = 24'(29580);
			6894: out = 24'(19800);
			6895: out = 24'(-4120);
			6896: out = 24'(13436);
			6897: out = 24'(51236);
			6898: out = 24'(59472);
			6899: out = 24'(21828);
			6900: out = 24'(-33160);
			6901: out = 24'(-93756);
			6902: out = 24'(-96092);
			6903: out = 24'(-56988);
			6904: out = 24'(-1096);
			6905: out = 24'(61364);
			6906: out = 24'(66320);
			6907: out = 24'(61952);
			6908: out = 24'(47276);
			6909: out = 24'(25648);
			6910: out = 24'(-61960);
			6911: out = 24'(-87212);
			6912: out = 24'(-50500);
			6913: out = 24'(-20868);
			6914: out = 24'(-20852);
			6915: out = 24'(-10144);
			6916: out = 24'(42848);
			6917: out = 24'(94792);
			6918: out = 24'(88728);
			6919: out = 24'(35964);
			6920: out = 24'(-45772);
			6921: out = 24'(-114156);
			6922: out = 24'(-90652);
			6923: out = 24'(-76832);
			6924: out = 24'(-41616);
			6925: out = 24'(-6200);
			6926: out = 24'(25176);
			6927: out = 24'(41948);
			6928: out = 24'(54716);
			6929: out = 24'(29740);
			6930: out = 24'(-10296);
			6931: out = 24'(-50612);
			6932: out = 24'(-1644);
			6933: out = 24'(31940);
			6934: out = 24'(-2876);
			6935: out = 24'(-13572);
			6936: out = 24'(-1200);
			6937: out = 24'(4068);
			6938: out = 24'(-20524);
			6939: out = 24'(-8212);
			6940: out = 24'(18796);
			6941: out = 24'(34200);
			6942: out = 24'(8448);
			6943: out = 24'(-20380);
			6944: out = 24'(-43060);
			6945: out = 24'(-23560);
			6946: out = 24'(21336);
			6947: out = 24'(62000);
			6948: out = 24'(42976);
			6949: out = 24'(4308);
			6950: out = 24'(-19264);
			6951: out = 24'(7048);
			6952: out = 24'(3184);
			6953: out = 24'(8140);
			6954: out = 24'(-13564);
			6955: out = 24'(-15784);
			6956: out = 24'(28748);
			6957: out = 24'(29772);
			6958: out = 24'(-24072);
			6959: out = 24'(-40924);
			6960: out = 24'(55668);
			6961: out = 24'(51776);
			6962: out = 24'(-35548);
			6963: out = 24'(-104652);
			6964: out = 24'(-25708);
			6965: out = 24'(34748);
			6966: out = 24'(29232);
			6967: out = 24'(5248);
			6968: out = 24'(55656);
			6969: out = 24'(44032);
			6970: out = 24'(33088);
			6971: out = 24'(-32380);
			6972: out = 24'(-88664);
			6973: out = 24'(-88228);
			6974: out = 24'(760);
			6975: out = 24'(47996);
			6976: out = 24'(28428);
			6977: out = 24'(4888);
			6978: out = 24'(8136);
			6979: out = 24'(18948);
			6980: out = 24'(23464);
			6981: out = 24'(51920);
			6982: out = 24'(7252);
			6983: out = 24'(6012);
			6984: out = 24'(20788);
			6985: out = 24'(10340);
			6986: out = 24'(-80436);
			6987: out = 24'(-99372);
			6988: out = 24'(-23772);
			6989: out = 24'(38636);
			6990: out = 24'(10504);
			6991: out = 24'(-12944);
			6992: out = 24'(36252);
			6993: out = 24'(83748);
			6994: out = 24'(4044);
			6995: out = 24'(-70896);
			6996: out = 24'(-85056);
			6997: out = 24'(-21704);
			6998: out = 24'(-1548);
			6999: out = 24'(45332);
			7000: out = 24'(58584);
			7001: out = 24'(54688);
			7002: out = 24'(20948);
			7003: out = 24'(35408);
			7004: out = 24'(-3348);
			7005: out = 24'(-70304);
			7006: out = 24'(-113568);
			7007: out = 24'(-85400);
			7008: out = 24'(-20736);
			7009: out = 24'(20448);
			7010: out = 24'(19088);
			7011: out = 24'(5744);
			7012: out = 24'(40932);
			7013: out = 24'(76792);
			7014: out = 24'(48764);
			7015: out = 24'(-42812);
			7016: out = 24'(-47800);
			7017: out = 24'(5908);
			7018: out = 24'(14576);
			7019: out = 24'(-64076);
			7020: out = 24'(-89020);
			7021: out = 24'(-42128);
			7022: out = 24'(21596);
			7023: out = 24'(32456);
			7024: out = 24'(39084);
			7025: out = 24'(45052);
			7026: out = 24'(37424);
			7027: out = 24'(3712);
			7028: out = 24'(-8420);
			7029: out = 24'(-5480);
			7030: out = 24'(1092);
			7031: out = 24'(-7196);
			7032: out = 24'(-3484);
			7033: out = 24'(19388);
			7034: out = 24'(38908);
			7035: out = 24'(26668);
			7036: out = 24'(-5208);
			7037: out = 24'(-42472);
			7038: out = 24'(-53864);
			7039: out = 24'(-28256);
			7040: out = 24'(23856);
			7041: out = 24'(55900);
			7042: out = 24'(51696);
			7043: out = 24'(18992);
			7044: out = 24'(-4072);
			7045: out = 24'(13120);
			7046: out = 24'(16572);
			7047: out = 24'(-21164);
			7048: out = 24'(-65924);
			7049: out = 24'(-22736);
			7050: out = 24'(9508);
			7051: out = 24'(27716);
			7052: out = 24'(43372);
			7053: out = 24'(71140);
			7054: out = 24'(22360);
			7055: out = 24'(-45788);
			7056: out = 24'(-81136);
			7057: out = 24'(-37056);
			7058: out = 24'(6780);
			7059: out = 24'(48020);
			7060: out = 24'(68436);
			7061: out = 24'(49652);
			7062: out = 24'(-23104);
			7063: out = 24'(-54784);
			7064: out = 24'(-2980);
			7065: out = 24'(50576);
			7066: out = 24'(19148);
			7067: out = 24'(-51644);
			7068: out = 24'(-64268);
			7069: out = 24'(-18648);
			7070: out = 24'(5280);
			7071: out = 24'(-53304);
			7072: out = 24'(-45124);
			7073: out = 24'(39140);
			7074: out = 24'(69840);
			7075: out = 24'(42096);
			7076: out = 24'(31804);
			7077: out = 24'(41688);
			7078: out = 24'(-5432);
			7079: out = 24'(-49836);
			7080: out = 24'(-104044);
			7081: out = 24'(-90648);
			7082: out = 24'(-19732);
			7083: out = 24'(68672);
			7084: out = 24'(56480);
			7085: out = 24'(12912);
			7086: out = 24'(-5880);
			7087: out = 24'(46900);
			7088: out = 24'(7332);
			7089: out = 24'(-64732);
			7090: out = 24'(-100828);
			7091: out = 24'(-11892);
			7092: out = 24'(196);
			7093: out = 24'(12752);
			7094: out = 24'(27560);
			7095: out = 24'(49240);
			7096: out = 24'(52700);
			7097: out = 24'(53060);
			7098: out = 24'(3616);
			7099: out = 24'(-93808);
			7100: out = 24'(-72496);
			7101: out = 24'(-28920);
			7102: out = 24'(-1496);
			7103: out = 24'(-22008);
			7104: out = 24'(-11936);
			7105: out = 24'(14856);
			7106: out = 24'(64592);
			7107: out = 24'(47200);
			7108: out = 24'(-61860);
			7109: out = 24'(-81812);
			7110: out = 24'(1736);
			7111: out = 24'(66216);
			7112: out = 24'(34012);
			7113: out = 24'(-34248);
			7114: out = 24'(-30988);
			7115: out = 24'(15296);
			7116: out = 24'(18152);
			7117: out = 24'(11448);
			7118: out = 24'(36260);
			7119: out = 24'(56844);
			7120: out = 24'(13620);
			7121: out = 24'(-72208);
			7122: out = 24'(-120924);
			7123: out = 24'(-89344);
			7124: out = 24'(-9244);
			7125: out = 24'(71244);
			7126: out = 24'(66744);
			7127: out = 24'(41008);
			7128: out = 24'(14972);
			7129: out = 24'(1928);
			7130: out = 24'(-23868);
			7131: out = 24'(-28400);
			7132: out = 24'(-860);
			7133: out = 24'(38244);
			7134: out = 24'(38516);
			7135: out = 24'(32376);
			7136: out = 24'(31784);
			7137: out = 24'(24688);
			7138: out = 24'(-5576);
			7139: out = 24'(-73852);
			7140: out = 24'(-117700);
			7141: out = 24'(-83556);
			7142: out = 24'(12824);
			7143: out = 24'(47852);
			7144: out = 24'(47588);
			7145: out = 24'(54572);
			7146: out = 24'(73292);
			7147: out = 24'(22224);
			7148: out = 24'(-27024);
			7149: out = 24'(-26648);
			7150: out = 24'(17088);
			7151: out = 24'(-2252);
			7152: out = 24'(-57372);
			7153: out = 24'(-75192);
			7154: out = 24'(15100);
			7155: out = 24'(35968);
			7156: out = 24'(70336);
			7157: out = 24'(36760);
			7158: out = 24'(-14380);
			7159: out = 24'(-21984);
			7160: out = 24'(16456);
			7161: out = 24'(-4396);
			7162: out = 24'(-66144);
			7163: out = 24'(-49080);
			7164: out = 24'(-13060);
			7165: out = 24'(2080);
			7166: out = 24'(-6512);
			7167: out = 24'(39268);
			7168: out = 24'(49176);
			7169: out = 24'(70836);
			7170: out = 24'(59692);
			7171: out = 24'(28564);
			7172: out = 24'(-71224);
			7173: out = 24'(-106804);
			7174: out = 24'(-84252);
			7175: out = 24'(-27480);
			7176: out = 24'(15080);
			7177: out = 24'(66996);
			7178: out = 24'(77440);
			7179: out = 24'(44180);
			7180: out = 24'(-1656);
			7181: out = 24'(-23060);
			7182: out = 24'(-27508);
			7183: out = 24'(-40740);
			7184: out = 24'(-77916);
			7185: out = 24'(-35220);
			7186: out = 24'(16492);
			7187: out = 24'(25136);
			7188: out = 24'(-17844);
			7189: out = 24'(-15988);
			7190: out = 24'(13408);
			7191: out = 24'(48360);
			7192: out = 24'(28456);
			7193: out = 24'(14496);
			7194: out = 24'(-20556);
			7195: out = 24'(15528);
			7196: out = 24'(48264);
			7197: out = 24'(-15088);
			7198: out = 24'(-104412);
			7199: out = 24'(-68244);
			7200: out = 24'(50608);
			7201: out = 24'(43536);
			7202: out = 24'(-18724);
			7203: out = 24'(-20348);
			7204: out = 24'(43840);
			7205: out = 24'(21900);
			7206: out = 24'(11344);
			7207: out = 24'(-25412);
			7208: out = 24'(-6424);
			7209: out = 24'(22148);
			7210: out = 24'(80792);
			7211: out = 24'(41228);
			7212: out = 24'(9972);
			7213: out = 24'(668);
			7214: out = 24'(31792);
			7215: out = 24'(-57204);
			7216: out = 24'(-113640);
			7217: out = 24'(-63680);
			7218: out = 24'(41800);
			7219: out = 24'(45308);
			7220: out = 24'(27808);
			7221: out = 24'(16404);
			7222: out = 24'(1180);
			7223: out = 24'(-16300);
			7224: out = 24'(1596);
			7225: out = 24'(18636);
			7226: out = 24'(-6488);
			7227: out = 24'(26984);
			7228: out = 24'(28068);
			7229: out = 24'(-8136);
			7230: out = 24'(-61028);
			7231: out = 24'(47284);
			7232: out = 24'(56024);
			7233: out = 24'(8652);
			7234: out = 24'(-59244);
			7235: out = 24'(-29572);
			7236: out = 24'(-12448);
			7237: out = 24'(8912);
			7238: out = 24'(-10492);
			7239: out = 24'(-22552);
			7240: out = 24'(-11000);
			7241: out = 24'(58440);
			7242: out = 24'(65072);
			7243: out = 24'(8632);
			7244: out = 24'(-22212);
			7245: out = 24'(37360);
			7246: out = 24'(47904);
			7247: out = 24'(-45372);
			7248: out = 24'(-108468);
			7249: out = 24'(-57356);
			7250: out = 24'(14036);
			7251: out = 24'(9256);
			7252: out = 24'(58524);
			7253: out = 24'(72528);
			7254: out = 24'(63432);
			7255: out = 24'(10040);
			7256: out = 24'(-51108);
			7257: out = 24'(-111164);
			7258: out = 24'(-116552);
			7259: out = 24'(-68276);
			7260: out = 24'(65016);
			7261: out = 24'(96380);
			7262: out = 24'(98056);
			7263: out = 24'(66476);
			7264: out = 24'(37944);
			7265: out = 24'(-84640);
			7266: out = 24'(-121368);
			7267: out = 24'(-93732);
			7268: out = 24'(-19432);
			7269: out = 24'(3036);
			7270: out = 24'(42344);
			7271: out = 24'(39908);
			7272: out = 24'(32156);
			7273: out = 24'(57456);
			7274: out = 24'(31168);
			7275: out = 24'(-53904);
			7276: out = 24'(-103976);
			7277: out = 24'(996);
			7278: out = 24'(13492);
			7279: out = 24'(-17920);
			7280: out = 24'(-32108);
			7281: out = 24'(27588);
			7282: out = 24'(65516);
			7283: out = 24'(41344);
			7284: out = 24'(-12644);
			7285: out = 24'(-24720);
			7286: out = 24'(6964);
			7287: out = 24'(4236);
			7288: out = 24'(-20168);
			7289: out = 24'(-10264);
			7290: out = 24'(-2900);
			7291: out = 24'(9256);
			7292: out = 24'(-23152);
			7293: out = 24'(-42052);
			7294: out = 24'(7764);
			7295: out = 24'(61540);
			7296: out = 24'(47744);
			7297: out = 24'(-8076);
			7298: out = 24'(-25420);
			7299: out = 24'(-15040);
			7300: out = 24'(11376);
			7301: out = 24'(10792);
			7302: out = 24'(11284);
			7303: out = 24'(14000);
			7304: out = 24'(38996);
			7305: out = 24'(16784);
			7306: out = 24'(-43736);
			7307: out = 24'(-50616);
			7308: out = 24'(-19000);
			7309: out = 24'(13940);
			7310: out = 24'(21680);
			7311: out = 24'(31616);
			7312: out = 24'(56336);
			7313: out = 24'(58928);
			7314: out = 24'(23912);
			7315: out = 24'(-18516);
			7316: out = 24'(-70360);
			7317: out = 24'(-78648);
			7318: out = 24'(-41136);
			7319: out = 24'(3188);
			7320: out = 24'(29088);
			7321: out = 24'(27656);
			7322: out = 24'(28320);
			7323: out = 24'(34036);
			7324: out = 24'(26372);
			7325: out = 24'(-1344);
			7326: out = 24'(-16952);
			7327: out = 24'(-12524);
			7328: out = 24'(456);
			7329: out = 24'(-41304);
			7330: out = 24'(-55124);
			7331: out = 24'(-9716);
			7332: out = 24'(25996);
			7333: out = 24'(26872);
			7334: out = 24'(9132);
			7335: out = 24'(14044);
			7336: out = 24'(26964);
			7337: out = 24'(8852);
			7338: out = 24'(-6900);
			7339: out = 24'(19480);
			7340: out = 24'(53036);
			7341: out = 24'(-36364);
			7342: out = 24'(-116596);
			7343: out = 24'(-87300);
			7344: out = 24'(63272);
			7345: out = 24'(111016);
			7346: out = 24'(44032);
			7347: out = 24'(-10100);
			7348: out = 24'(11740);
			7349: out = 24'(36108);
			7350: out = 24'(-3836);
			7351: out = 24'(-83752);
			7352: out = 24'(-102200);
			7353: out = 24'(-42352);
			7354: out = 24'(28928);
			7355: out = 24'(20056);
			7356: out = 24'(3012);
			7357: out = 24'(16220);
			7358: out = 24'(58660);
			7359: out = 24'(8628);
			7360: out = 24'(-46536);
			7361: out = 24'(-27368);
			7362: out = 24'(40804);
			7363: out = 24'(29876);
			7364: out = 24'(-21924);
			7365: out = 24'(-52756);
			7366: out = 24'(-46288);
			7367: out = 24'(-3276);
			7368: out = 24'(33200);
			7369: out = 24'(35532);
			7370: out = 24'(8672);
			7371: out = 24'(8260);
			7372: out = 24'(29196);
			7373: out = 24'(18476);
			7374: out = 24'(-42336);
			7375: out = 24'(-95052);
			7376: out = 24'(-52508);
			7377: out = 24'(26732);
			7378: out = 24'(29796);
			7379: out = 24'(4972);
			7380: out = 24'(16472);
			7381: out = 24'(68808);
			7382: out = 24'(62508);
			7383: out = 24'(-6740);
			7384: out = 24'(-86768);
			7385: out = 24'(-70008);
			7386: out = 24'(14672);
			7387: out = 24'(58648);
			7388: out = 24'(26952);
			7389: out = 24'(876);
			7390: out = 24'(-10016);
			7391: out = 24'(-18584);
			7392: out = 24'(-48212);
			7393: out = 24'(-14212);
			7394: out = 24'(31652);
			7395: out = 24'(25796);
			7396: out = 24'(600);
			7397: out = 24'(30112);
			7398: out = 24'(76152);
			7399: out = 24'(56004);
			7400: out = 24'(-7900);
			7401: out = 24'(-61824);
			7402: out = 24'(-47616);
			7403: out = 24'(-9236);
			7404: out = 24'(-20);
			7405: out = 24'(-3476);
			7406: out = 24'(26016);
			7407: out = 24'(59132);
			7408: out = 24'(49020);
			7409: out = 24'(4992);
			7410: out = 24'(-13140);
			7411: out = 24'(13156);
			7412: out = 24'(39828);
			7413: out = 24'(31280);
			7414: out = 24'(-28432);
			7415: out = 24'(-88180);
			7416: out = 24'(-77832);
			7417: out = 24'(-8708);
			7418: out = 24'(35820);
			7419: out = 24'(15764);
			7420: out = 24'(12568);
			7421: out = 24'(70984);
			7422: out = 24'(70488);
			7423: out = 24'(-20740);
			7424: out = 24'(-104216);
			7425: out = 24'(-54496);
			7426: out = 24'(-5972);
			7427: out = 24'(-40512);
			7428: out = 24'(-80208);
			7429: out = 24'(16188);
			7430: out = 24'(100592);
			7431: out = 24'(95540);
			7432: out = 24'(17136);
			7433: out = 24'(-44320);
			7434: out = 24'(-26080);
			7435: out = 24'(-46708);
			7436: out = 24'(-104392);
			7437: out = 24'(-106332);
			7438: out = 24'(32000);
			7439: out = 24'(94960);
			7440: out = 24'(50544);
			7441: out = 24'(-3216);
			7442: out = 24'(2352);
			7443: out = 24'(6900);
			7444: out = 24'(-4192);
			7445: out = 24'(-19000);
			7446: out = 24'(-3460);
			7447: out = 24'(-1172);
			7448: out = 24'(4180);
			7449: out = 24'(-13716);
			7450: out = 24'(-49360);
			7451: out = 24'(-5824);
			7452: out = 24'(9384);
			7453: out = 24'(3936);
			7454: out = 24'(-2376);
			7455: out = 24'(18352);
			7456: out = 24'(38608);
			7457: out = 24'(39460);
			7458: out = 24'(6652);
			7459: out = 24'(-25592);
			7460: out = 24'(-61044);
			7461: out = 24'(-44040);
			7462: out = 24'(8496);
			7463: out = 24'(65212);
			7464: out = 24'(28764);
			7465: out = 24'(124);
			7466: out = 24'(-28188);
			7467: out = 24'(-33800);
			7468: out = 24'(-60616);
			7469: out = 24'(4896);
			7470: out = 24'(60128);
			7471: out = 24'(54940);
			7472: out = 24'(5816);
			7473: out = 24'(16304);
			7474: out = 24'(13292);
			7475: out = 24'(-19360);
			7476: out = 24'(-50476);
			7477: out = 24'(-34936);
			7478: out = 24'(-43468);
			7479: out = 24'(-37816);
			7480: out = 24'(55432);
			7481: out = 24'(102712);
			7482: out = 24'(49816);
			7483: out = 24'(-30144);
			7484: out = 24'(-35156);
			7485: out = 24'(-21508);
			7486: out = 24'(-57324);
			7487: out = 24'(-83192);
			7488: out = 24'(9724);
			7489: out = 24'(12080);
			7490: out = 24'(44212);
			7491: out = 24'(46396);
			7492: out = 24'(52436);
			7493: out = 24'(27320);
			7494: out = 24'(10644);
			7495: out = 24'(-31860);
			7496: out = 24'(-38548);
			7497: out = 24'(24556);
			7498: out = 24'(29144);
			7499: out = 24'(-19744);
			7500: out = 24'(-55324);
			7501: out = 24'(-16028);
			7502: out = 24'(9668);
			7503: out = 24'(11264);
			7504: out = 24'(21808);
			7505: out = 24'(69064);
			7506: out = 24'(76800);
			7507: out = 24'(40652);
			7508: out = 24'(-31688);
			7509: out = 24'(-91220);
			7510: out = 24'(-92000);
			7511: out = 24'(-62012);
			7512: out = 24'(-16816);
			7513: out = 24'(29544);
			7514: out = 24'(43992);
			7515: out = 24'(48192);
			7516: out = 24'(44064);
			7517: out = 24'(39084);
			7518: out = 24'(-2488);
			7519: out = 24'(12504);
			7520: out = 24'(-10440);
			7521: out = 24'(-40568);
			7522: out = 24'(-50668);
			7523: out = 24'(-13700);
			7524: out = 24'(3148);
			7525: out = 24'(16840);
			7526: out = 24'(34268);
			7527: out = 24'(15796);
			7528: out = 24'(-1308);
			7529: out = 24'(-5428);
			7530: out = 24'(3488);
			7531: out = 24'(44168);
			7532: out = 24'(-9380);
			7533: out = 24'(-32576);
			7534: out = 24'(-3952);
			7535: out = 24'(15248);
			7536: out = 24'(-48148);
			7537: out = 24'(-53184);
			7538: out = 24'(35460);
			7539: out = 24'(65668);
			7540: out = 24'(41588);
			7541: out = 24'(-56164);
			7542: out = 24'(-90860);
			7543: out = 24'(-33264);
			7544: out = 24'(41092);
			7545: out = 24'(964);
			7546: out = 24'(-26520);
			7547: out = 24'(19024);
			7548: out = 24'(50384);
			7549: out = 24'(22652);
			7550: out = 24'(-23308);
			7551: out = 24'(-42696);
			7552: out = 24'(-17584);
			7553: out = 24'(-19992);
			7554: out = 24'(3484);
			7555: out = 24'(28924);
			7556: out = 24'(32828);
			7557: out = 24'(42352);
			7558: out = 24'(57644);
			7559: out = 24'(-9016);
			7560: out = 24'(-117568);
			7561: out = 24'(-106596);
			7562: out = 24'(-8384);
			7563: out = 24'(47748);
			7564: out = 24'(-1192);
			7565: out = 24'(47252);
			7566: out = 24'(69324);
			7567: out = 24'(66368);
			7568: out = 24'(7952);
			7569: out = 24'(-11400);
			7570: out = 24'(-36472);
			7571: out = 24'(-18372);
			7572: out = 24'(-9656);
			7573: out = 24'(-16808);
			7574: out = 24'(-36080);
			7575: out = 24'(-28284);
			7576: out = 24'(-12512);
			7577: out = 24'(4548);
			7578: out = 24'(37328);
			7579: out = 24'(47564);
			7580: out = 24'(7508);
			7581: out = 24'(-46852);
			7582: out = 24'(7848);
			7583: out = 24'(29508);
			7584: out = 24'(-26624);
			7585: out = 24'(-108708);
			7586: out = 24'(-24076);
			7587: out = 24'(13468);
			7588: out = 24'(31428);
			7589: out = 24'(61904);
			7590: out = 24'(103204);
			7591: out = 24'(63876);
			7592: out = 24'(-39400);
			7593: out = 24'(-117816);
			7594: out = 24'(-86324);
			7595: out = 24'(-32156);
			7596: out = 24'(-3552);
			7597: out = 24'(18484);
			7598: out = 24'(67060);
			7599: out = 24'(83180);
			7600: out = 24'(38820);
			7601: out = 24'(-28004);
			7602: out = 24'(-54100);
			7603: out = 24'(-18644);
			7604: out = 24'(-27920);
			7605: out = 24'(-47584);
			7606: out = 24'(-7920);
			7607: out = 24'(72128);
			7608: out = 24'(73548);
			7609: out = 24'(21680);
			7610: out = 24'(-10280);
			7611: out = 24'(16368);
			7612: out = 24'(-12020);
			7613: out = 24'(-65896);
			7614: out = 24'(-80848);
			7615: out = 24'(8368);
			7616: out = 24'(4396);
			7617: out = 24'(33468);
			7618: out = 24'(51264);
			7619: out = 24'(51860);
			7620: out = 24'(10420);
			7621: out = 24'(-16872);
			7622: out = 24'(-46916);
			7623: out = 24'(-51728);
			7624: out = 24'(-16536);
			7625: out = 24'(44196);
			7626: out = 24'(63164);
			7627: out = 24'(45368);
			7628: out = 24'(3760);
			7629: out = 24'(-16400);
			7630: out = 24'(-40032);
			7631: out = 24'(-15476);
			7632: out = 24'(52404);
			7633: out = 24'(52704);
			7634: out = 24'(-36316);
			7635: out = 24'(-100504);
			7636: out = 24'(-18996);
			7637: out = 24'(-8824);
			7638: out = 24'(9664);
			7639: out = 24'(-8504);
			7640: out = 24'(6652);
			7641: out = 24'(35796);
			7642: out = 24'(80832);
			7643: out = 24'(31108);
			7644: out = 24'(-66552);
			7645: out = 24'(-114500);
			7646: out = 24'(-48688);
			7647: out = 24'(22576);
			7648: out = 24'(23232);
			7649: out = 24'(-288);
			7650: out = 24'(26140);
			7651: out = 24'(49140);
			7652: out = 24'(18080);
			7653: out = 24'(-66228);
			7654: out = 24'(-18484);
			7655: out = 24'(-4832);
			7656: out = 24'(-7540);
			7657: out = 24'(-16872);
			7658: out = 24'(2980);
			7659: out = 24'(192);
			7660: out = 24'(22780);
			7661: out = 24'(39236);
			7662: out = 24'(-26136);
			7663: out = 24'(-13348);
			7664: out = 24'(36560);
			7665: out = 24'(59676);
			7666: out = 24'(17604);
			7667: out = 24'(-27652);
			7668: out = 24'(-23252);
			7669: out = 24'(-280);
			7670: out = 24'(-34772);
			7671: out = 24'(-1680);
			7672: out = 24'(4944);
			7673: out = 24'(9228);
			7674: out = 24'(10084);
			7675: out = 24'(60936);
			7676: out = 24'(38580);
			7677: out = 24'(-11108);
			7678: out = 24'(-51216);
			7679: out = 24'(-7984);
			7680: out = 24'(-23712);
			7681: out = 24'(-18684);
			7682: out = 24'(38592);
			7683: out = 24'(102936);
			7684: out = 24'(97588);
			7685: out = 24'(26768);
			7686: out = 24'(-56340);
			7687: out = 24'(-84652);
			7688: out = 24'(-54216);
			7689: out = 24'(-11800);
			7690: out = 24'(296);
			7691: out = 24'(4552);
			7692: out = 24'(38284);
			7693: out = 24'(34744);
			7694: out = 24'(-10408);
			7695: out = 24'(-44836);
			7696: out = 24'(20912);
			7697: out = 24'(39816);
			7698: out = 24'(-564);
			7699: out = 24'(-56948);
			7700: out = 24'(-36372);
			7701: out = 24'(28236);
			7702: out = 24'(69828);
			7703: out = 24'(45020);
			7704: out = 24'(3000);
			7705: out = 24'(-6972);
			7706: out = 24'(2996);
			7707: out = 24'(-21324);
			7708: out = 24'(-64436);
			7709: out = 24'(-60676);
			7710: out = 24'(-6292);
			7711: out = 24'(17632);
			7712: out = 24'(-1500);
			7713: out = 24'(-13100);
			7714: out = 24'(47708);
			7715: out = 24'(74712);
			7716: out = 24'(25160);
			7717: out = 24'(-30976);
			7718: out = 24'(-33144);
			7719: out = 24'(-12924);
			7720: out = 24'(-28900);
			7721: out = 24'(-38420);
			7722: out = 24'(-41864);
			7723: out = 24'(17328);
			7724: out = 24'(73512);
			7725: out = 24'(81900);
			7726: out = 24'(940);
			7727: out = 24'(-53792);
			7728: out = 24'(-52992);
			7729: out = 24'(1324);
			7730: out = 24'(-61212);
			7731: out = 24'(-11044);
			7732: out = 24'(54984);
			7733: out = 24'(59572);
			7734: out = 24'(6576);
			7735: out = 24'(7652);
			7736: out = 24'(20188);
			7737: out = 24'(396);
			7738: out = 24'(-34788);
			7739: out = 24'(-39740);
			7740: out = 24'(-15376);
			7741: out = 24'(4320);
			7742: out = 24'(25236);
			7743: out = 24'(7888);
			7744: out = 24'(4968);
			7745: out = 24'(-11564);
			7746: out = 24'(-30876);
			7747: out = 24'(-52984);
			7748: out = 24'(-16004);
			7749: out = 24'(10628);
			7750: out = 24'(-3616);
			7751: out = 24'(-39512);
			7752: out = 24'(-5512);
			7753: out = 24'(36428);
			7754: out = 24'(44712);
			7755: out = 24'(44348);
			7756: out = 24'(11252);
			7757: out = 24'(-30372);
			7758: out = 24'(-31600);
			7759: out = 24'(25032);
			7760: out = 24'(36660);
			7761: out = 24'(-24208);
			7762: out = 24'(-88064);
			7763: out = 24'(-66152);
			7764: out = 24'(12384);
			7765: out = 24'(48364);
			7766: out = 24'(58892);
			7767: out = 24'(74688);
			7768: out = 24'(36064);
			7769: out = 24'(-39224);
			7770: out = 24'(-87848);
			7771: out = 24'(-48744);
			7772: out = 24'(-25988);
			7773: out = 24'(-4904);
			7774: out = 24'(1328);
			7775: out = 24'(33132);
			7776: out = 24'(64860);
			7777: out = 24'(80096);
			7778: out = 24'(48020);
			7779: out = 24'(1408);
			7780: out = 24'(-32072);
			7781: out = 24'(4152);
			7782: out = 24'(13828);
			7783: out = 24'(-26216);
			7784: out = 24'(-68444);
			7785: out = 24'(8552);
			7786: out = 24'(48148);
			7787: out = 24'(-4252);
			7788: out = 24'(-86084);
			7789: out = 24'(-12492);
			7790: out = 24'(58964);
			7791: out = 24'(60176);
			7792: out = 24'(328);
			7793: out = 24'(-53524);
			7794: out = 24'(-32936);
			7795: out = 24'(-5256);
			7796: out = 24'(-23988);
			7797: out = 24'(-38864);
			7798: out = 24'(-15388);
			7799: out = 24'(39460);
			7800: out = 24'(55132);
			7801: out = 24'(31796);
			7802: out = 24'(-12868);
			7803: out = 24'(-12700);
			7804: out = 24'(2560);
			7805: out = 24'(-10492);
			7806: out = 24'(-103808);
			7807: out = 24'(-88412);
			7808: out = 24'(-10184);
			7809: out = 24'(42904);
			7810: out = 24'(55544);
			7811: out = 24'(33132);
			7812: out = 24'(-7064);
			7813: out = 24'(-41024);
			7814: out = 24'(-27980);
			7815: out = 24'(22728);
			7816: out = 24'(59592);
			7817: out = 24'(47508);
			7818: out = 24'(12768);
			7819: out = 24'(788);
			7820: out = 24'(-8468);
			7821: out = 24'(-29252);
			7822: out = 24'(-37264);
			7823: out = 24'(-54136);
			7824: out = 24'(-14960);
			7825: out = 24'(19168);
			7826: out = 24'(31192);
			7827: out = 24'(6808);
			7828: out = 24'(59920);
			7829: out = 24'(64620);
			7830: out = 24'(9820);
			7831: out = 24'(-47292);
			7832: out = 24'(-19352);
			7833: out = 24'(6136);
			7834: out = 24'(-5788);
			7835: out = 24'(1392);
			7836: out = 24'(-38988);
			7837: out = 24'(-38092);
			7838: out = 24'(-8928);
			7839: out = 24'(33888);
			7840: out = 24'(41792);
			7841: out = 24'(44388);
			7842: out = 24'(27136);
			7843: out = 24'(296);
			7844: out = 24'(-36648);
			7845: out = 24'(-33664);
			7846: out = 24'(-26132);
			7847: out = 24'(-34872);
			7848: out = 24'(-28916);
			7849: out = 24'(9272);
			7850: out = 24'(62284);
			7851: out = 24'(75132);
			7852: out = 24'(53160);
			7853: out = 24'(6176);
			7854: out = 24'(-4040);
			7855: out = 24'(-13280);
			7856: out = 24'(-50744);
			7857: out = 24'(-105968);
			7858: out = 24'(-67472);
			7859: out = 24'(26488);
			7860: out = 24'(59884);
			7861: out = 24'(26816);
			7862: out = 24'(23076);
			7863: out = 24'(48632);
			7864: out = 24'(40180);
			7865: out = 24'(-25484);
			7866: out = 24'(-41116);
			7867: out = 24'(-17052);
			7868: out = 24'(-14256);
			7869: out = 24'(-26632);
			7870: out = 24'(-39812);
			7871: out = 24'(16884);
			7872: out = 24'(54484);
			7873: out = 24'(27916);
			7874: out = 24'(856);
			7875: out = 24'(31064);
			7876: out = 24'(44912);
			7877: out = 24'(-6116);
			7878: out = 24'(-70792);
			7879: out = 24'(-63364);
			7880: out = 24'(-25956);
			7881: out = 24'(-17324);
			7882: out = 24'(1256);
			7883: out = 24'(49824);
			7884: out = 24'(61256);
			7885: out = 24'(10256);
			7886: out = 24'(-38872);
			7887: out = 24'(-40944);
			7888: out = 24'(-30108);
			7889: out = 24'(-40444);
			7890: out = 24'(-17940);
			7891: out = 24'(-2700);
			7892: out = 24'(40452);
			7893: out = 24'(54032);
			7894: out = 24'(43584);
			7895: out = 24'(3880);
			7896: out = 24'(9116);
			7897: out = 24'(-9660);
			7898: out = 24'(-71028);
			7899: out = 24'(-51080);
			7900: out = 24'(-11788);
			7901: out = 24'(40748);
			7902: out = 24'(59732);
			7903: out = 24'(60860);
			7904: out = 24'(35348);
			7905: out = 24'(12908);
			7906: out = 24'(-18164);
			7907: out = 24'(-29908);
			7908: out = 24'(-69628);
			7909: out = 24'(-46560);
			7910: out = 24'(5968);
			7911: out = 24'(41416);
			7912: out = 24'(29780);
			7913: out = 24'(34076);
			7914: out = 24'(23156);
			7915: out = 24'(-4448);
			7916: out = 24'(-62272);
			7917: out = 24'(-16212);
			7918: out = 24'(23124);
			7919: out = 24'(-14328);
			7920: out = 24'(-76972);
			7921: out = 24'(-9436);
			7922: out = 24'(80180);
			7923: out = 24'(49308);
			7924: out = 24'(-52352);
			7925: out = 24'(-62072);
			7926: out = 24'(31388);
			7927: out = 24'(64132);
			7928: out = 24'(-8380);
			7929: out = 24'(-70368);
			7930: out = 24'(-54380);
			7931: out = 24'(-20684);
			7932: out = 24'(-24008);
			7933: out = 24'(57036);
			7934: out = 24'(88404);
			7935: out = 24'(36792);
			7936: out = 24'(-46256);
			7937: out = 24'(-18348);
			7938: out = 24'(26684);
			7939: out = 24'(-560);
			7940: out = 24'(-70420);
			7941: out = 24'(-43036);
			7942: out = 24'(43428);
			7943: out = 24'(50176);
			7944: out = 24'(-10984);
			7945: out = 24'(10240);
			7946: out = 24'(31368);
			7947: out = 24'(32288);
			7948: out = 24'(-21828);
			7949: out = 24'(-37564);
			7950: out = 24'(-72400);
			7951: out = 24'(9132);
			7952: out = 24'(62092);
			7953: out = 24'(30828);
			7954: out = 24'(2076);
			7955: out = 24'(-24316);
			7956: out = 24'(-14352);
			7957: out = 24'(9284);
			7958: out = 24'(23196);
			7959: out = 24'(11888);
			7960: out = 24'(6524);
			7961: out = 24'(17344);
			7962: out = 24'(31048);
			7963: out = 24'(680);
			7964: out = 24'(-48780);
			7965: out = 24'(-60352);
			7966: out = 24'(24440);
			7967: out = 24'(18984);
			7968: out = 24'(33528);
			7969: out = 24'(31024);
			7970: out = 24'(31568);
			7971: out = 24'(-54512);
			7972: out = 24'(-40052);
			7973: out = 24'(-33568);
			7974: out = 24'(-48668);
			7975: out = 24'(-23668);
			7976: out = 24'(39564);
			7977: out = 24'(31484);
			7978: out = 24'(-32080);
			7979: out = 24'(-60068);
			7980: out = 24'(20600);
			7981: out = 24'(50060);
			7982: out = 24'(-4624);
			7983: out = 24'(-49192);
			7984: out = 24'(8104);
			7985: out = 24'(46124);
			7986: out = 24'(12688);
			7987: out = 24'(-25908);
			7988: out = 24'(3044);
			7989: out = 24'(45740);
			7990: out = 24'(39112);
			7991: out = 24'(-8316);
			7992: out = 24'(-33916);
			7993: out = 24'(-37816);
			7994: out = 24'(-24316);
			7995: out = 24'(-14920);
			7996: out = 24'(15920);
			7997: out = 24'(14912);
			7998: out = 24'(35492);
			7999: out = 24'(31688);
			8000: out = 24'(-30444);
			8001: out = 24'(-45836);
			8002: out = 24'(-4812);
			8003: out = 24'(52948);
			8004: out = 24'(60412);
			8005: out = 24'(-40992);
			8006: out = 24'(-72672);
			8007: out = 24'(-18112);
			8008: out = 24'(38080);
			8009: out = 24'(55772);
			8010: out = 24'(52728);
			8011: out = 24'(49940);
			8012: out = 24'(17936);
			8013: out = 24'(-45700);
			8014: out = 24'(-114764);
			8015: out = 24'(-94332);
			8016: out = 24'(-14840);
			8017: out = 24'(32688);
			8018: out = 24'(36364);
			8019: out = 24'(69648);
			8020: out = 24'(83516);
			8021: out = 24'(51804);
			8022: out = 24'(-72632);
			8023: out = 24'(-97488);
			8024: out = 24'(-46524);
			8025: out = 24'(-21532);
			8026: out = 24'(-45064);
			8027: out = 24'(-2620);
			8028: out = 24'(71116);
			8029: out = 24'(90776);
			8030: out = 24'(48176);
			8031: out = 24'(24420);
			8032: out = 24'(-2128);
			8033: out = 24'(-47388);
			8034: out = 24'(-96556);
			8035: out = 24'(-47448);
			8036: out = 24'(6196);
			8037: out = 24'(-5320);
			8038: out = 24'(-34332);
			8039: out = 24'(42324);
			8040: out = 24'(107120);
			8041: out = 24'(57928);
			8042: out = 24'(-70564);
			8043: out = 24'(-101348);
			8044: out = 24'(-44104);
			8045: out = 24'(13432);
			8046: out = 24'(-1808);
			8047: out = 24'(11632);
			8048: out = 24'(12660);
			8049: out = 24'(28756);
			8050: out = 24'(25476);
			8051: out = 24'(11368);
			8052: out = 24'(11904);
			8053: out = 24'(29100);
			8054: out = 24'(13072);
			8055: out = 24'(-49120);
			8056: out = 24'(-90968);
			8057: out = 24'(-52676);
			8058: out = 24'(32432);
			8059: out = 24'(65312);
			8060: out = 24'(31136);
			8061: out = 24'(12076);
			8062: out = 24'(28012);
			8063: out = 24'(19200);
			8064: out = 24'(-17920);
			8065: out = 24'(-82140);
			8066: out = 24'(-75072);
			8067: out = 24'(-248);
			8068: out = 24'(66340);
			8069: out = 24'(35456);
			8070: out = 24'(15352);
			8071: out = 24'(17292);
			8072: out = 24'(952);
			8073: out = 24'(-43468);
			8074: out = 24'(-50376);
			8075: out = 24'(-20008);
			8076: out = 24'(-3672);
			8077: out = 24'(24520);
			8078: out = 24'(60592);
			8079: out = 24'(70152);
			8080: out = 24'(23752);
			8081: out = 24'(-37768);
			8082: out = 24'(-29252);
			8083: out = 24'(27852);
			8084: out = 24'(28400);
			8085: out = 24'(-56708);
			8086: out = 24'(-75920);
			8087: out = 24'(-11836);
			8088: out = 24'(37076);
			8089: out = 24'(32988);
			8090: out = 24'(-4848);
			8091: out = 24'(-2772);
			8092: out = 24'(2996);
			8093: out = 24'(-1780);
			8094: out = 24'(-17316);
			8095: out = 24'(36760);
			8096: out = 24'(59972);
			8097: out = 24'(12432);
			8098: out = 24'(-43888);
			8099: out = 24'(-15260);
			8100: out = 24'(8196);
			8101: out = 24'(-26884);
			8102: out = 24'(-2196);
			8103: out = 24'(54008);
			8104: out = 24'(58572);
			8105: out = 24'(-14992);
			8106: out = 24'(-70472);
			8107: out = 24'(-62484);
			8108: out = 24'(-28580);
			8109: out = 24'(-18812);
			8110: out = 24'(23420);
			8111: out = 24'(8940);
			8112: out = 24'(6280);
			8113: out = 24'(2780);
			8114: out = 24'(22760);
			8115: out = 24'(11128);
			8116: out = 24'(32692);
			8117: out = 24'(46208);
			8118: out = 24'(36932);
			8119: out = 24'(-24548);
			8120: out = 24'(-29088);
			8121: out = 24'(-9448);
			8122: out = 24'(-3376);
			8123: out = 24'(-16372);
			8124: out = 24'(11968);
			8125: out = 24'(38816);
			8126: out = 24'(22508);
			8127: out = 24'(3848);
			8128: out = 24'(-51504);
			8129: out = 24'(-29076);
			8130: out = 24'(11848);
			8131: out = 24'(-528);
			8132: out = 24'(-696);
			8133: out = 24'(19136);
			8134: out = 24'(33484);
			8135: out = 24'(13852);
			8136: out = 24'(-3320);
			8137: out = 24'(3108);
			8138: out = 24'(11264);
			8139: out = 24'(-3576);
			8140: out = 24'(-10740);
			8141: out = 24'(5232);
			8142: out = 24'(25488);
			8143: out = 24'(25940);
			8144: out = 24'(28208);
			8145: out = 24'(43884);
			8146: out = 24'(33032);
			8147: out = 24'(-29260);
			8148: out = 24'(-93900);
			8149: out = 24'(-101892);
			8150: out = 24'(-34764);
			8151: out = 24'(15252);
			8152: out = 24'(21120);
			8153: out = 24'(37188);
			8154: out = 24'(68752);
			8155: out = 24'(44480);
			8156: out = 24'(-43112);
			8157: out = 24'(-60140);
			8158: out = 24'(-57740);
			8159: out = 24'(-23100);
			8160: out = 24'(14672);
			8161: out = 24'(35856);
			8162: out = 24'(20372);
			8163: out = 24'(-21844);
			8164: out = 24'(-34592);
			8165: out = 24'(9612);
			8166: out = 24'(43208);
			8167: out = 24'(-912);
			8168: out = 24'(-56316);
			8169: out = 24'(-23528);
			8170: out = 24'(42364);
			8171: out = 24'(37816);
			8172: out = 24'(-32684);
			8173: out = 24'(-79136);
			8174: out = 24'(-44324);
			8175: out = 24'(30216);
			8176: out = 24'(49748);
			8177: out = 24'(10032);
			8178: out = 24'(-10224);
			8179: out = 24'(-68);
			8180: out = 24'(48280);
			8181: out = 24'(53824);
			8182: out = 24'(-6564);
			8183: out = 24'(-67604);
			8184: out = 24'(-54720);
			8185: out = 24'(-14084);
			8186: out = 24'(-28764);
			8187: out = 24'(-6616);
			8188: out = 24'(52348);
			8189: out = 24'(90308);
			8190: out = 24'(58276);
			8191: out = 24'(5808);
			8192: out = 24'(-33332);
			8193: out = 24'(-47988);
			8194: out = 24'(-42456);
			8195: out = 24'(-65960);
			8196: out = 24'(16776);
			8197: out = 24'(71000);
			8198: out = 24'(33488);
			8199: out = 24'(-66488);
			8200: out = 24'(-53656);
			8201: out = 24'(-5684);
			8202: out = 24'(5428);
			8203: out = 24'(4424);
			8204: out = 24'(26304);
			8205: out = 24'(36308);
			8206: out = 24'(7716);
			8207: out = 24'(-33076);
			8208: out = 24'(1596);
			8209: out = 24'(29272);
			8210: out = 24'(12784);
			8211: out = 24'(-31096);
			8212: out = 24'(-8828);
			8213: out = 24'(84);
			8214: out = 24'(-5072);
			8215: out = 24'(-15604);
			8216: out = 24'(18496);
			8217: out = 24'(28496);
			8218: out = 24'(41896);
			8219: out = 24'(33472);
			8220: out = 24'(-9968);
			8221: out = 24'(-70360);
			8222: out = 24'(-73600);
			8223: out = 24'(-21776);
			8224: out = 24'(-468);
			8225: out = 24'(14880);
			8226: out = 24'(27376);
			8227: out = 24'(59592);
			8228: out = 24'(71164);
			8229: out = 24'(50768);
			8230: out = 24'(2760);
			8231: out = 24'(-39008);
			8232: out = 24'(-74068);
			8233: out = 24'(-14948);
			8234: out = 24'(-38936);
			8235: out = 24'(-35948);
			8236: out = 24'(20436);
			8237: out = 24'(95860);
			8238: out = 24'(38028);
			8239: out = 24'(-7460);
			8240: out = 24'(-7584);
			8241: out = 24'(15728);
			8242: out = 24'(-21120);
			8243: out = 24'(-41828);
			8244: out = 24'(-43508);
			8245: out = 24'(-26168);
			8246: out = 24'(-4160);
			8247: out = 24'(62252);
			8248: out = 24'(67556);
			8249: out = 24'(-11864);
			8250: out = 24'(-69344);
			8251: out = 24'(-33792);
			8252: out = 24'(25536);
			8253: out = 24'(7124);
			8254: out = 24'(-8992);
			8255: out = 24'(-12876);
			8256: out = 24'(26016);
			8257: out = 24'(30636);
			8258: out = 24'(3928);
			8259: out = 24'(-44872);
			8260: out = 24'(-24700);
			8261: out = 24'(11728);
			8262: out = 24'(-916);
			8263: out = 24'(-14048);
			8264: out = 24'(-8988);
			8265: out = 24'(5060);
			8266: out = 24'(828);
			8267: out = 24'(7536);
			8268: out = 24'(20804);
			8269: out = 24'(27304);
			8270: out = 24'(7300);
			8271: out = 24'(3216);
			8272: out = 24'(-5052);
			8273: out = 24'(13580);
			8274: out = 24'(24168);
			8275: out = 24'(-6388);
			8276: out = 24'(-31868);
			8277: out = 24'(-33220);
			8278: out = 24'(-11672);
			8279: out = 24'(-1484);
			8280: out = 24'(16876);
			8281: out = 24'(18012);
			8282: out = 24'(19056);
			8283: out = 24'(12548);
			8284: out = 24'(-43920);
			8285: out = 24'(-61120);
			8286: out = 24'(-2188);
			8287: out = 24'(71424);
			8288: out = 24'(54924);
			8289: out = 24'(6296);
			8290: out = 24'(-33764);
			8291: out = 24'(-35728);
			8292: out = 24'(-26720);
			8293: out = 24'(-29080);
			8294: out = 24'(-13872);
			8295: out = 24'(22064);
			8296: out = 24'(13900);
			8297: out = 24'(16212);
			8298: out = 24'(-19688);
			8299: out = 24'(-29596);
			8300: out = 24'(4304);
			8301: out = 24'(41192);
			8302: out = 24'(17232);
			8303: out = 24'(-5716);
			8304: out = 24'(22832);
			8305: out = 24'(-1364);
			8306: out = 24'(-340);
			8307: out = 24'(-17100);
			8308: out = 24'(-18084);
			8309: out = 24'(13464);
			8310: out = 24'(34692);
			8311: out = 24'(9288);
			8312: out = 24'(-33340);
			8313: out = 24'(-42392);
			8314: out = 24'(-45504);
			8315: out = 24'(-22112);
			8316: out = 24'(30344);
			8317: out = 24'(72980);
			8318: out = 24'(42360);
			8319: out = 24'(-23432);
			8320: out = 24'(-52680);
			8321: out = 24'(-4256);
			8322: out = 24'(28596);
			8323: out = 24'(24592);
			8324: out = 24'(10096);
			8325: out = 24'(18092);
			8326: out = 24'(-18924);
			8327: out = 24'(-9616);
			8328: out = 24'(-6344);
			8329: out = 24'(-5656);
			8330: out = 24'(-5764);
			8331: out = 24'(38424);
			8332: out = 24'(59788);
			8333: out = 24'(37188);
			8334: out = 24'(-7700);
			8335: out = 24'(-45748);
			8336: out = 24'(-42676);
			8337: out = 24'(-14460);
			8338: out = 24'(6320);
			8339: out = 24'(6888);
			8340: out = 24'(3064);
			8341: out = 24'(4);
			8342: out = 24'(-4512);
			8343: out = 24'(-78256);
			8344: out = 24'(-46512);
			8345: out = 24'(32124);
			8346: out = 24'(78436);
			8347: out = 24'(56336);
			8348: out = 24'(19704);
			8349: out = 24'(-32888);
			8350: out = 24'(-72560);
			8351: out = 24'(-92704);
			8352: out = 24'(-21552);
			8353: out = 24'(36576);
			8354: out = 24'(53576);
			8355: out = 24'(24468);
			8356: out = 24'(14964);
			8357: out = 24'(-20872);
			8358: out = 24'(-19704);
			8359: out = 24'(4240);
			8360: out = 24'(7872);
			8361: out = 24'(-29576);
			8362: out = 24'(-4556);
			8363: out = 24'(57184);
			8364: out = 24'(42232);
			8365: out = 24'(-38836);
			8366: out = 24'(-51960);
			8367: out = 24'(27564);
			8368: out = 24'(51872);
			8369: out = 24'(4864);
			8370: out = 24'(-20496);
			8371: out = 24'(14936);
			8372: out = 24'(22396);
			8373: out = 24'(19332);
			8374: out = 24'(568);
			8375: out = 24'(-7716);
			8376: out = 24'(-42752);
			8377: out = 24'(-6228);
			8378: out = 24'(-23520);
			8379: out = 24'(-22408);
			8380: out = 24'(5928);
			8381: out = 24'(37684);
			8382: out = 24'(57076);
			8383: out = 24'(75900);
			8384: out = 24'(60564);
			8385: out = 24'(-17548);
			8386: out = 24'(-104200);
			8387: out = 24'(-100544);
			8388: out = 24'(-27708);
			8389: out = 24'(4324);
			8390: out = 24'(17156);
			8391: out = 24'(28192);
			8392: out = 24'(29056);
			8393: out = 24'(5564);
			8394: out = 24'(5496);
			8395: out = 24'(14624);
			8396: out = 24'(4340);
			8397: out = 24'(-35328);
			8398: out = 24'(-43148);
			8399: out = 24'(-5560);
			8400: out = 24'(21448);
			8401: out = 24'(-12588);
			8402: out = 24'(-47432);
			8403: out = 24'(-21836);
			8404: out = 24'(51072);
			8405: out = 24'(65384);
			8406: out = 24'(21500);
			8407: out = 24'(-25764);
			8408: out = 24'(-16056);
			8409: out = 24'(-2212);
			8410: out = 24'(-17452);
			8411: out = 24'(-43872);
			8412: out = 24'(5940);
			8413: out = 24'(46864);
			8414: out = 24'(11036);
			8415: out = 24'(-5876);
			8416: out = 24'(-4508);
			8417: out = 24'(14616);
			8418: out = 24'(15356);
			8419: out = 24'(6580);
			8420: out = 24'(-2404);
			8421: out = 24'(-20696);
			8422: out = 24'(-30564);
			8423: out = 24'(26996);
			8424: out = 24'(12392);
			8425: out = 24'(-42976);
			8426: out = 24'(-91832);
			8427: out = 24'(-16552);
			8428: out = 24'(-2732);
			8429: out = 24'(40028);
			8430: out = 24'(55632);
			8431: out = 24'(53080);
			8432: out = 24'(3784);
			8433: out = 24'(-2400);
			8434: out = 24'(-27912);
			8435: out = 24'(-69292);
			8436: out = 24'(-19536);
			8437: out = 24'(30244);
			8438: out = 24'(42352);
			8439: out = 24'(26080);
			8440: out = 24'(17296);
			8441: out = 24'(12240);
			8442: out = 24'(-27264);
			8443: out = 24'(-61068);
			8444: out = 24'(-4828);
			8445: out = 24'(6316);
			8446: out = 24'(-10260);
			8447: out = 24'(-24368);
			8448: out = 24'(25556);
			8449: out = 24'(34204);
			8450: out = 24'(33340);
			8451: out = 24'(3880);
			8452: out = 24'(-9172);
			8453: out = 24'(-11164);
			8454: out = 24'(9908);
			8455: out = 24'(6184);
			8456: out = 24'(3592);
			8457: out = 24'(13528);
			8458: out = 24'(44472);
			8459: out = 24'(22932);
			8460: out = 24'(-18052);
			8461: out = 24'(-6840);
			8462: out = 24'(-2408);
			8463: out = 24'(-10656);
			8464: out = 24'(-17484);
			8465: out = 24'(412);
			8466: out = 24'(35936);
			8467: out = 24'(41280);
			8468: out = 24'(35696);
			8469: out = 24'(24980);
			8470: out = 24'(-16020);
			8471: out = 24'(-82488);
			8472: out = 24'(-93652);
			8473: out = 24'(-22084);
			8474: out = 24'(-3792);
			8475: out = 24'(20620);
			8476: out = 24'(46748);
			8477: out = 24'(59924);
			8478: out = 24'(56);
			8479: out = 24'(-16748);
			8480: out = 24'(-6440);
			8481: out = 24'(25264);
			8482: out = 24'(33724);
			8483: out = 24'(7136);
			8484: out = 24'(-19160);
			8485: out = 24'(-34000);
			8486: out = 24'(-52640);
			8487: out = 24'(-20088);
			8488: out = 24'(5664);
			8489: out = 24'(23196);
			8490: out = 24'(27800);
			8491: out = 24'(42068);
			8492: out = 24'(-15044);
			8493: out = 24'(-82228);
			8494: out = 24'(-85876);
			8495: out = 24'(-9832);
			8496: out = 24'(33976);
			8497: out = 24'(17580);
			8498: out = 24'(9160);
			8499: out = 24'(41772);
			8500: out = 24'(63028);
			8501: out = 24'(29220);
			8502: out = 24'(-13196);
			8503: out = 24'(-33308);
			8504: out = 24'(12344);
			8505: out = 24'(-23512);
			8506: out = 24'(-65788);
			8507: out = 24'(-44180);
			8508: out = 24'(6192);
			8509: out = 24'(-3788);
			8510: out = 24'(-10360);
			8511: out = 24'(29152);
			8512: out = 24'(59220);
			8513: out = 24'(9104);
			8514: out = 24'(-29564);
			8515: out = 24'(-12608);
			8516: out = 24'(-17344);
			8517: out = 24'(-28700);
			8518: out = 24'(-26744);
			8519: out = 24'(16700);
			8520: out = 24'(16032);
			8521: out = 24'(24004);
			8522: out = 24'(-25272);
			8523: out = 24'(-32796);
			8524: out = 24'(2832);
			8525: out = 24'(66100);
			8526: out = 24'(2468);
			8527: out = 24'(-65952);
			8528: out = 24'(-71468);
			8529: out = 24'(-4864);
			8530: out = 24'(13312);
			8531: out = 24'(45420);
			8532: out = 24'(62740);
			8533: out = 24'(-14244);
			8534: out = 24'(-42880);
			8535: out = 24'(-7008);
			8536: out = 24'(34260);
			8537: out = 24'(-7568);
			8538: out = 24'(-37788);
			8539: out = 24'(13208);
			8540: out = 24'(92848);
			8541: out = 24'(71376);
			8542: out = 24'(-7336);
			8543: out = 24'(-65912);
			8544: out = 24'(-46720);
			8545: out = 24'(-12796);
			8546: out = 24'(7768);
			8547: out = 24'(9852);
			8548: out = 24'(36092);
			8549: out = 24'(52104);
			8550: out = 24'(59296);
			8551: out = 24'(-18228);
			8552: out = 24'(-50372);
			8553: out = 24'(-20376);
			8554: out = 24'(14120);
			8555: out = 24'(-19112);
			8556: out = 24'(-35712);
			8557: out = 24'(-13440);
			8558: out = 24'(12420);
			8559: out = 24'(26736);
			8560: out = 24'(36928);
			8561: out = 24'(40640);
			8562: out = 24'(21116);
			8563: out = 24'(-7988);
			8564: out = 24'(-30204);
			8565: out = 24'(-29336);
			8566: out = 24'(-17284);
			8567: out = 24'(-932);
			8568: out = 24'(11904);
			8569: out = 24'(17128);
			8570: out = 24'(9188);
			8571: out = 24'(18744);
			8572: out = 24'(-5140);
			8573: out = 24'(3340);
			8574: out = 24'(14280);
			8575: out = 24'(-5528);
			8576: out = 24'(-54404);
			8577: out = 24'(-59700);
			8578: out = 24'(-24572);
			8579: out = 24'(-4864);
			8580: out = 24'(54548);
			8581: out = 24'(29532);
			8582: out = 24'(-11880);
			8583: out = 24'(-24132);
			8584: out = 24'(37260);
			8585: out = 24'(37696);
			8586: out = 24'(752);
			8587: out = 24'(-46132);
			8588: out = 24'(-47784);
			8589: out = 24'(-37424);
			8590: out = 24'(10320);
			8591: out = 24'(50560);
			8592: out = 24'(50548);
			8593: out = 24'(11848);
			8594: out = 24'(-8276);
			8595: out = 24'(-3112);
			8596: out = 24'(6540);
			8597: out = 24'(24216);
			8598: out = 24'(15108);
			8599: out = 24'(-31872);
			8600: out = 24'(-94304);
			8601: out = 24'(-45752);
			8602: out = 24'(-6084);
			8603: out = 24'(11696);
			8604: out = 24'(3880);
			8605: out = 24'(-14160);
			8606: out = 24'(-2820);
			8607: out = 24'(31120);
			8608: out = 24'(54276);
			8609: out = 24'(31376);
			8610: out = 24'(10860);
			8611: out = 24'(-13668);
			8612: out = 24'(-12504);
			8613: out = 24'(2804);
			8614: out = 24'(-41636);
			8615: out = 24'(-59560);
			8616: out = 24'(3540);
			8617: out = 24'(71104);
			8618: out = 24'(27852);
			8619: out = 24'(-61792);
			8620: out = 24'(-73872);
			8621: out = 24'(18192);
			8622: out = 24'(26488);
			8623: out = 24'(-6636);
			8624: out = 24'(-31512);
			8625: out = 24'(3412);
			8626: out = 24'(40092);
			8627: out = 24'(29892);
			8628: out = 24'(6880);
			8629: out = 24'(-4124);
			8630: out = 24'(-30808);
			8631: out = 24'(-512);
			8632: out = 24'(21880);
			8633: out = 24'(24080);
			8634: out = 24'(-1396);
			8635: out = 24'(6408);
			8636: out = 24'(10392);
			8637: out = 24'(6648);
			8638: out = 24'(-16296);
			8639: out = 24'(-21584);
			8640: out = 24'(-38400);
			8641: out = 24'(-36512);
			8642: out = 24'(-9440);
			8643: out = 24'(16416);
			8644: out = 24'(50064);
			8645: out = 24'(56140);
			8646: out = 24'(30916);
			8647: out = 24'(-17120);
			8648: out = 24'(-21084);
			8649: out = 24'(-10136);
			8650: out = 24'(8920);
			8651: out = 24'(26996);
			8652: out = 24'(21784);
			8653: out = 24'(-16252);
			8654: out = 24'(-48880);
			8655: out = 24'(-21452);
			8656: out = 24'(30620);
			8657: out = 24'(68676);
			8658: out = 24'(57548);
			8659: out = 24'(34084);
			8660: out = 24'(8916);
			8661: out = 24'(-13652);
			8662: out = 24'(-75920);
			8663: out = 24'(-115628);
			8664: out = 24'(-90640);
			8665: out = 24'(27552);
			8666: out = 24'(82668);
			8667: out = 24'(70860);
			8668: out = 24'(51496);
			8669: out = 24'(33232);
			8670: out = 24'(-8456);
			8671: out = 24'(-52888);
			8672: out = 24'(-65128);
			8673: out = 24'(-38412);
			8674: out = 24'(-24828);
			8675: out = 24'(244);
			8676: out = 24'(41732);
			8677: out = 24'(29304);
			8678: out = 24'(11900);
			8679: out = 24'(17404);
			8680: out = 24'(43872);
			8681: out = 24'(25164);
			8682: out = 24'(-23600);
			8683: out = 24'(-51248);
			8684: out = 24'(-21568);
			8685: out = 24'(-7132);
			8686: out = 24'(7448);
			8687: out = 24'(6144);
			8688: out = 24'(24328);
			8689: out = 24'(15016);
			8690: out = 24'(24752);
			8691: out = 24'(-27816);
			8692: out = 24'(-54928);
			8693: out = 24'(-52724);
			8694: out = 24'(-108);
			8695: out = 24'(-32912);
			8696: out = 24'(-12276);
			8697: out = 24'(58884);
			8698: out = 24'(82768);
			8699: out = 24'(-15296);
			8700: out = 24'(-61840);
			8701: out = 24'(-22452);
			8702: out = 24'(-21132);
			8703: out = 24'(-3848);
			8704: out = 24'(30320);
			8705: out = 24'(42188);
			8706: out = 24'(-26984);
			8707: out = 24'(-22384);
			8708: out = 24'(32424);
			8709: out = 24'(74436);
			8710: out = 24'(27916);
			8711: out = 24'(-59068);
			8712: out = 24'(-93772);
			8713: out = 24'(-59468);
			8714: out = 24'(-28316);
			8715: out = 24'(1664);
			8716: out = 24'(5844);
			8717: out = 24'(14800);
			8718: out = 24'(23144);
			8719: out = 24'(40656);
			8720: out = 24'(40440);
			8721: out = 24'(26344);
			8722: out = 24'(-7252);
			8723: out = 24'(-42356);
			8724: out = 24'(-52848);
			8725: out = 24'(-24680);
			8726: out = 24'(18912);
			8727: out = 24'(44532);
			8728: out = 24'(54872);
			8729: out = 24'(22404);
			8730: out = 24'(-16608);
			8731: out = 24'(-30200);
			8732: out = 24'(-21476);
			8733: out = 24'(-1144);
			8734: out = 24'(17012);
			8735: out = 24'(26104);
			8736: out = 24'(-6700);
			8737: out = 24'(-1524);
			8738: out = 24'(-3924);
			8739: out = 24'(-2964);
			8740: out = 24'(12736);
			8741: out = 24'(33176);
			8742: out = 24'(45384);
			8743: out = 24'(54988);
			8744: out = 24'(52152);
			8745: out = 24'(-25948);
			8746: out = 24'(-77340);
			8747: out = 24'(-51876);
			8748: out = 24'(19024);
			8749: out = 24'(2060);
			8750: out = 24'(-14940);
			8751: out = 24'(-3696);
			8752: out = 24'(30272);
			8753: out = 24'(15028);
			8754: out = 24'(-23692);
			8755: out = 24'(-53376);
			8756: out = 24'(-31452);
			8757: out = 24'(1020);
			8758: out = 24'(31888);
			8759: out = 24'(16632);
			8760: out = 24'(-1324);
			8761: out = 24'(7096);
			8762: out = 24'(14624);
			8763: out = 24'(8676);
			8764: out = 24'(-12452);
			8765: out = 24'(-32804);
			8766: out = 24'(-43096);
			8767: out = 24'(-18296);
			8768: out = 24'(20256);
			8769: out = 24'(35048);
			8770: out = 24'(10076);
			8771: out = 24'(-9688);
			8772: out = 24'(1680);
			8773: out = 24'(18832);
			8774: out = 24'(-31556);
			8775: out = 24'(-21912);
			8776: out = 24'(-3912);
			8777: out = 24'(14180);
			8778: out = 24'(-7820);
			8779: out = 24'(50180);
			8780: out = 24'(29952);
			8781: out = 24'(-22988);
			8782: out = 24'(-58468);
			8783: out = 24'(28576);
			8784: out = 24'(37472);
			8785: out = 24'(9968);
			8786: out = 24'(1220);
			8787: out = 24'(-8520);
			8788: out = 24'(-5612);
			8789: out = 24'(-14216);
			8790: out = 24'(-25836);
			8791: out = 24'(-22928);
			8792: out = 24'(18716);
			8793: out = 24'(63032);
			8794: out = 24'(59832);
			8795: out = 24'(5128);
			8796: out = 24'(-41712);
			8797: out = 24'(-30828);
			8798: out = 24'(8884);
			8799: out = 24'(-940);
			8800: out = 24'(3500);
			8801: out = 24'(-12868);
			8802: out = 24'(-3168);
			8803: out = 24'(16988);
			8804: out = 24'(27484);
			8805: out = 24'(-2660);
			8806: out = 24'(-26996);
			8807: out = 24'(-20424);
			8808: out = 24'(8440);
			8809: out = 24'(4792);
			8810: out = 24'(-2080);
			8811: out = 24'(-656);
			8812: out = 24'(-14408);
			8813: out = 24'(-12024);
			8814: out = 24'(-17112);
			8815: out = 24'(-14428);
			8816: out = 24'(1812);
			8817: out = 24'(23716);
			8818: out = 24'(18460);
			8819: out = 24'(-4340);
			8820: out = 24'(-9380);
			8821: out = 24'(-1004);
			8822: out = 24'(21168);
			8823: out = 24'(-2640);
			8824: out = 24'(-58512);
			8825: out = 24'(-14188);
			8826: out = 24'(18640);
			8827: out = 24'(38020);
			8828: out = 24'(15032);
			8829: out = 24'(-24652);
			8830: out = 24'(-47360);
			8831: out = 24'(-2532);
			8832: out = 24'(49044);
			8833: out = 24'(29248);
			8834: out = 24'(34020);
			8835: out = 24'(33052);
			8836: out = 24'(29836);
			8837: out = 24'(-7504);
			8838: out = 24'(-13484);
			8839: out = 24'(-34384);
			8840: out = 24'(-15492);
			8841: out = 24'(13868);
			8842: out = 24'(3596);
			8843: out = 24'(-46968);
			8844: out = 24'(-41888);
			8845: out = 24'(31464);
			8846: out = 24'(49436);
			8847: out = 24'(20756);
			8848: out = 24'(-31120);
			8849: out = 24'(-49700);
			8850: out = 24'(-46092);
			8851: out = 24'(-8244);
			8852: out = 24'(1656);
			8853: out = 24'(4912);
			8854: out = 24'(19916);
			8855: out = 24'(59212);
			8856: out = 24'(37304);
			8857: out = 24'(-23920);
			8858: out = 24'(-68620);
			8859: out = 24'(-46096);
			8860: out = 24'(-9928);
			8861: out = 24'(-916);
			8862: out = 24'(-3780);
			8863: out = 24'(-1768);
			8864: out = 24'(33452);
			8865: out = 24'(29664);
			8866: out = 24'(-7420);
			8867: out = 24'(-2736);
			8868: out = 24'(8552);
			8869: out = 24'(26864);
			8870: out = 24'(21080);
			8871: out = 24'(5356);
			8872: out = 24'(-40452);
			8873: out = 24'(-55020);
			8874: out = 24'(-37540);
			8875: out = 24'(7784);
			8876: out = 24'(56168);
			8877: out = 24'(84556);
			8878: out = 24'(61264);
			8879: out = 24'(3464);
			8880: out = 24'(-70820);
			8881: out = 24'(-56244);
			8882: out = 24'(-17064);
			8883: out = 24'(-17300);
			8884: out = 24'(-13776);
			8885: out = 24'(-9452);
			8886: out = 24'(29036);
			8887: out = 24'(53688);
			8888: out = 24'(50132);
			8889: out = 24'(-15288);
			8890: out = 24'(-35840);
			8891: out = 24'(-17392);
			8892: out = 24'(-4544);
			8893: out = 24'(-53192);
			8894: out = 24'(-36596);
			8895: out = 24'(40172);
			8896: out = 24'(81628);
			8897: out = 24'(14800);
			8898: out = 24'(-8120);
			8899: out = 24'(21820);
			8900: out = 24'(40312);
			8901: out = 24'(-44600);
			8902: out = 24'(-77140);
			8903: out = 24'(-49144);
			8904: out = 24'(15628);
			8905: out = 24'(27976);
			8906: out = 24'(18172);
			8907: out = 24'(-27056);
			8908: out = 24'(-39272);
			8909: out = 24'(14364);
			8910: out = 24'(3252);
			8911: out = 24'(292);
			8912: out = 24'(6624);
			8913: out = 24'(17664);
			8914: out = 24'(8332);
			8915: out = 24'(-8400);
			8916: out = 24'(-22892);
			8917: out = 24'(-22440);
			8918: out = 24'(-18796);
			8919: out = 24'(-5136);
			8920: out = 24'(12772);
			8921: out = 24'(33496);
			8922: out = 24'(31060);
			8923: out = 24'(47660);
			8924: out = 24'(18000);
			8925: out = 24'(-35168);
			8926: out = 24'(-59016);
			8927: out = 24'(-3532);
			8928: out = 24'(46016);
			8929: out = 24'(38356);
			8930: out = 24'(3036);
			8931: out = 24'(-13552);
			8932: out = 24'(-4712);
			8933: out = 24'(-14180);
			8934: out = 24'(-42936);
			8935: out = 24'(-4500);
			8936: out = 24'(24264);
			8937: out = 24'(22132);
			8938: out = 24'(-12980);
			8939: out = 24'(3228);
			8940: out = 24'(-10464);
			8941: out = 24'(11268);
			8942: out = 24'(25976);
			8943: out = 24'(17156);
			8944: out = 24'(-18972);
			8945: out = 24'(-9348);
			8946: out = 24'(16828);
			8947: out = 24'(13464);
			8948: out = 24'(-13140);
			8949: out = 24'(-15872);
			8950: out = 24'(-2312);
			8951: out = 24'(480);
			8952: out = 24'(20508);
			8953: out = 24'(8752);
			8954: out = 24'(-15388);
			8955: out = 24'(-32824);
			8956: out = 24'(-32524);
			8957: out = 24'(-21524);
			8958: out = 24'(-12436);
			8959: out = 24'(13288);
			8960: out = 24'(54504);
			8961: out = 24'(74952);
			8962: out = 24'(36552);
			8963: out = 24'(-15140);
			8964: out = 24'(-24576);
			8965: out = 24'(-17248);
			8966: out = 24'(-27892);
			8967: out = 24'(-52504);
			8968: out = 24'(-51828);
			8969: out = 24'(-8628);
			8970: out = 24'(23880);
			8971: out = 24'(46856);
			8972: out = 24'(65828);
			8973: out = 24'(50624);
			8974: out = 24'(4212);
			8975: out = 24'(-32308);
			8976: out = 24'(-17980);
			8977: out = 24'(-8088);
			8978: out = 24'(-4536);
			8979: out = 24'(-29900);
			8980: out = 24'(-12768);
			8981: out = 24'(42936);
			8982: out = 24'(48776);
			8983: out = 24'(-5336);
			8984: out = 24'(-38320);
			8985: out = 24'(-12976);
			8986: out = 24'(1016);
			8987: out = 24'(-32308);
			8988: out = 24'(-34828);
			8989: out = 24'(26564);
			8990: out = 24'(47828);
			8991: out = 24'(14904);
			8992: out = 24'(-9276);
			8993: out = 24'(20744);
			8994: out = 24'(35292);
			8995: out = 24'(1728);
			8996: out = 24'(-40860);
			8997: out = 24'(-39620);
			8998: out = 24'(-35556);
			8999: out = 24'(10316);
			9000: out = 24'(9608);
			9001: out = 24'(-8984);
			9002: out = 24'(-30436);
			9003: out = 24'(20536);
			9004: out = 24'(18136);
			9005: out = 24'(220);
			9006: out = 24'(4596);
			9007: out = 24'(53972);
			9008: out = 24'(33544);
			9009: out = 24'(-18960);
			9010: out = 24'(-44056);
			9011: out = 24'(26352);
			9012: out = 24'(24088);
			9013: out = 24'(-2180);
			9014: out = 24'(-20228);
			9015: out = 24'(-1908);
			9016: out = 24'(6144);
			9017: out = 24'(6016);
			9018: out = 24'(-32912);
			9019: out = 24'(-105660);
			9020: out = 24'(-29484);
			9021: out = 24'(69188);
			9022: out = 24'(88716);
			9023: out = 24'(29272);
			9024: out = 24'(-50072);
			9025: out = 24'(-55872);
			9026: out = 24'(-13516);
			9027: out = 24'(-2808);
			9028: out = 24'(4040);
			9029: out = 24'(21376);
			9030: out = 24'(47164);
			9031: out = 24'(18008);
			9032: out = 24'(-34192);
			9033: out = 24'(-91316);
			9034: out = 24'(-42972);
			9035: out = 24'(32592);
			9036: out = 24'(46068);
			9037: out = 24'(-7068);
			9038: out = 24'(5444);
			9039: out = 24'(35960);
			9040: out = 24'(9228);
			9041: out = 24'(-62208);
			9042: out = 24'(-43184);
			9043: out = 24'(31580);
			9044: out = 24'(41680);
			9045: out = 24'(-6700);
			9046: out = 24'(-34148);
			9047: out = 24'(-18256);
			9048: out = 24'(-4372);
			9049: out = 24'(19920);
			9050: out = 24'(-24132);
			9051: out = 24'(-56096);
			9052: out = 24'(-42100);
			9053: out = 24'(66512);
			9054: out = 24'(58848);
			9055: out = 24'(68812);
			9056: out = 24'(46400);
			9057: out = 24'(328);
			9058: out = 24'(-42428);
			9059: out = 24'(-20968);
			9060: out = 24'(-28328);
			9061: out = 24'(-96632);
			9062: out = 24'(-58796);
			9063: out = 24'(28964);
			9064: out = 24'(68516);
			9065: out = 24'(25172);
			9066: out = 24'(-33676);
			9067: out = 24'(4468);
			9068: out = 24'(40300);
			9069: out = 24'(-1884);
			9070: out = 24'(-52660);
			9071: out = 24'(-25340);
			9072: out = 24'(43352);
			9073: out = 24'(49288);
			9074: out = 24'(8176);
			9075: out = 24'(-37176);
			9076: out = 24'(-22352);
			9077: out = 24'(4840);
			9078: out = 24'(2332);
			9079: out = 24'(24584);
			9080: out = 24'(32284);
			9081: out = 24'(4872);
			9082: out = 24'(-53864);
			9083: out = 24'(-41148);
			9084: out = 24'(-25548);
			9085: out = 24'(17120);
			9086: out = 24'(60604);
			9087: out = 24'(71528);
			9088: out = 24'(52768);
			9089: out = 24'(21632);
			9090: out = 24'(-548);
			9091: out = 24'(-21344);
			9092: out = 24'(-18416);
			9093: out = 24'(-33092);
			9094: out = 24'(-42936);
			9095: out = 24'(-29776);
			9096: out = 24'(1764);
			9097: out = 24'(3584);
			9098: out = 24'(10460);
			9099: out = 24'(45428);
			9100: out = 24'(36624);
			9101: out = 24'(17660);
			9102: out = 24'(-2832);
			9103: out = 24'(1312);
			9104: out = 24'(-4776);
			9105: out = 24'(212);
			9106: out = 24'(2824);
			9107: out = 24'(21304);
			9108: out = 24'(20444);
			9109: out = 24'(2348);
			9110: out = 24'(-53924);
			9111: out = 24'(-84908);
			9112: out = 24'(-64268);
			9113: out = 24'(5692);
			9114: out = 24'(17540);
			9115: out = 24'(21492);
			9116: out = 24'(48144);
			9117: out = 24'(58492);
			9118: out = 24'(-3044);
			9119: out = 24'(-52180);
			9120: out = 24'(-23080);
			9121: out = 24'(-284);
			9122: out = 24'(9128);
			9123: out = 24'(8248);
			9124: out = 24'(16916);
			9125: out = 24'(-1876);
			9126: out = 24'(-40604);
			9127: out = 24'(-50028);
			9128: out = 24'(1436);
			9129: out = 24'(31976);
			9130: out = 24'(33592);
			9131: out = 24'(-15488);
			9132: out = 24'(-45448);
			9133: out = 24'(-36788);
			9134: out = 24'(-3456);
			9135: out = 24'(-7096);
			9136: out = 24'(1008);
			9137: out = 24'(39640);
			9138: out = 24'(59076);
			9139: out = 24'(31992);
			9140: out = 24'(-5300);
			9141: out = 24'(-18472);
			9142: out = 24'(-14572);
			9143: out = 24'(-16280);
			9144: out = 24'(-21920);
			9145: out = 24'(-25928);
			9146: out = 24'(-28580);
			9147: out = 24'(508);
			9148: out = 24'(40092);
			9149: out = 24'(56224);
			9150: out = 24'(40192);
			9151: out = 24'(11036);
			9152: out = 24'(788);
			9153: out = 24'(-10624);
			9154: out = 24'(-33884);
			9155: out = 24'(-49800);
			9156: out = 24'(-19980);
			9157: out = 24'(7348);
			9158: out = 24'(-3148);
			9159: out = 24'(-14396);
			9160: out = 24'(248);
			9161: out = 24'(24344);
			9162: out = 24'(23688);
			9163: out = 24'(8896);
			9164: out = 24'(11452);
			9165: out = 24'(31868);
			9166: out = 24'(34276);
			9167: out = 24'(-4896);
			9168: out = 24'(-41180);
			9169: out = 24'(-42024);
			9170: out = 24'(-1844);
			9171: out = 24'(13512);
			9172: out = 24'(32588);
			9173: out = 24'(-2296);
			9174: out = 24'(-492);
			9175: out = 24'(25332);
			9176: out = 24'(15744);
			9177: out = 24'(-55800);
			9178: out = 24'(-74644);
			9179: out = 24'(-5900);
			9180: out = 24'(47320);
			9181: out = 24'(-8220);
			9182: out = 24'(-34880);
			9183: out = 24'(31296);
			9184: out = 24'(83108);
			9185: out = 24'(41008);
			9186: out = 24'(-50040);
			9187: out = 24'(-103112);
			9188: out = 24'(-80968);
			9189: out = 24'(2820);
			9190: out = 24'(23856);
			9191: out = 24'(-2132);
			9192: out = 24'(-24632);
			9193: out = 24'(28968);
			9194: out = 24'(18508);
			9195: out = 24'(-20808);
			9196: out = 24'(-30120);
			9197: out = 24'(49144);
			9198: out = 24'(63944);
			9199: out = 24'(40960);
			9200: out = 24'(1108);
			9201: out = 24'(-15864);
			9202: out = 24'(-18420);
			9203: out = 24'(-5444);
			9204: out = 24'(-23480);
			9205: out = 24'(-73532);
			9206: out = 24'(-11908);
			9207: out = 24'(44700);
			9208: out = 24'(32024);
			9209: out = 24'(-23060);
			9210: out = 24'(11960);
			9211: out = 24'(36812);
			9212: out = 24'(16752);
			9213: out = 24'(-25808);
			9214: out = 24'(-2420);
			9215: out = 24'(47696);
			9216: out = 24'(50152);
			9217: out = 24'(-26268);
			9218: out = 24'(-112272);
			9219: out = 24'(-55904);
			9220: out = 24'(47652);
			9221: out = 24'(60620);
			9222: out = 24'(1144);
			9223: out = 24'(-7580);
			9224: out = 24'(8356);
			9225: out = 24'(9408);
			9226: out = 24'(-29256);
			9227: out = 24'(-50408);
			9228: out = 24'(-25424);
			9229: out = 24'(40596);
			9230: out = 24'(61488);
			9231: out = 24'(17528);
			9232: out = 24'(-51640);
			9233: out = 24'(-42880);
			9234: out = 24'(36260);
			9235: out = 24'(75736);
			9236: out = 24'(4444);
			9237: out = 24'(-57016);
			9238: out = 24'(-37444);
			9239: out = 24'(23040);
			9240: out = 24'(-31636);
			9241: out = 24'(-67608);
			9242: out = 24'(-9340);
			9243: out = 24'(70972);
			9244: out = 24'(19764);
			9245: out = 24'(-51284);
			9246: out = 24'(-56700);
			9247: out = 24'(19064);
			9248: out = 24'(57252);
			9249: out = 24'(45764);
			9250: out = 24'(4612);
			9251: out = 24'(-34900);
			9252: out = 24'(-33664);
			9253: out = 24'(-27604);
			9254: out = 24'(12056);
			9255: out = 24'(38680);
			9256: out = 24'(19784);
			9257: out = 24'(-3044);
			9258: out = 24'(16472);
			9259: out = 24'(37120);
			9260: out = 24'(8480);
			9261: out = 24'(-28040);
			9262: out = 24'(-36404);
			9263: out = 24'(-34672);
			9264: out = 24'(-55196);
			9265: out = 24'(-32704);
			9266: out = 24'(17524);
			9267: out = 24'(59752);
			9268: out = 24'(54752);
			9269: out = 24'(5796);
			9270: out = 24'(-17252);
			9271: out = 24'(-32708);
			9272: out = 24'(-35468);
			9273: out = 24'(6748);
			9274: out = 24'(23232);
			9275: out = 24'(11368);
			9276: out = 24'(-1036);
			9277: out = 24'(30844);
			9278: out = 24'(33516);
			9279: out = 24'(6028);
			9280: out = 24'(-34396);
			9281: out = 24'(-24772);
			9282: out = 24'(-24148);
			9283: out = 24'(-1584);
			9284: out = 24'(-5096);
			9285: out = 24'(-4828);
			9286: out = 24'(17616);
			9287: out = 24'(50192);
			9288: out = 24'(31116);
			9289: out = 24'(-12508);
			9290: out = 24'(-29568);
			9291: out = 24'(22428);
			9292: out = 24'(44376);
			9293: out = 24'(11248);
			9294: out = 24'(-40532);
			9295: out = 24'(-27200);
			9296: out = 24'(-1368);
			9297: out = 24'(22056);
			9298: out = 24'(41048);
			9299: out = 24'(32424);
			9300: out = 24'(-7336);
			9301: out = 24'(-35872);
			9302: out = 24'(-24064);
			9303: out = 24'(-31288);
			9304: out = 24'(-22380);
			9305: out = 24'(14400);
			9306: out = 24'(63860);
			9307: out = 24'(71340);
			9308: out = 24'(31172);
			9309: out = 24'(-4356);
			9310: out = 24'(-9320);
			9311: out = 24'(-29080);
			9312: out = 24'(-43180);
			9313: out = 24'(-51388);
			9314: out = 24'(-24520);
			9315: out = 24'(3732);
			9316: out = 24'(36444);
			9317: out = 24'(33968);
			9318: out = 24'(35500);
			9319: out = 24'(28932);
			9320: out = 24'(-35008);
			9321: out = 24'(-72952);
			9322: out = 24'(-19792);
			9323: out = 24'(64872);
			9324: out = 24'(43464);
			9325: out = 24'(-1752);
			9326: out = 24'(-7636);
			9327: out = 24'(30432);
			9328: out = 24'(64);
			9329: out = 24'(-7996);
			9330: out = 24'(-12388);
			9331: out = 24'(-5656);
			9332: out = 24'(-48232);
			9333: out = 24'(-37384);
			9334: out = 24'(-23576);
			9335: out = 24'(15120);
			9336: out = 24'(23500);
			9337: out = 24'(57252);
			9338: out = 24'(-16808);
			9339: out = 24'(-73764);
			9340: out = 24'(-44020);
			9341: out = 24'(51304);
			9342: out = 24'(35132);
			9343: out = 24'(-484);
			9344: out = 24'(5948);
			9345: out = 24'(13124);
			9346: out = 24'(-4220);
			9347: out = 24'(-37856);
			9348: out = 24'(-44020);
			9349: out = 24'(-11628);
			9350: out = 24'(31240);
			9351: out = 24'(48388);
			9352: out = 24'(8276);
			9353: out = 24'(-88716);
			9354: out = 24'(-5628);
			9355: out = 24'(55380);
			9356: out = 24'(31688);
			9357: out = 24'(-54908);
			9358: out = 24'(-43604);
			9359: out = 24'(-17396);
			9360: out = 24'(7136);
			9361: out = 24'(-512);
			9362: out = 24'(10804);
			9363: out = 24'(592);
			9364: out = 24'(14112);
			9365: out = 24'(32452);
			9366: out = 24'(42572);
			9367: out = 24'(23540);
			9368: out = 24'(340);
			9369: out = 24'(-29092);
			9370: out = 24'(-38628);
			9371: out = 24'(-14044);
			9372: out = 24'(47148);
			9373: out = 24'(55268);
			9374: out = 24'(-6588);
			9375: out = 24'(-43684);
			9376: out = 24'(-28548);
			9377: out = 24'(-940);
			9378: out = 24'(-15344);
			9379: out = 24'(4084);
			9380: out = 24'(-15880);
			9381: out = 24'(-31740);
			9382: out = 24'(-34500);
			9383: out = 24'(30228);
			9384: out = 24'(21020);
			9385: out = 24'(27564);
			9386: out = 24'(45576);
			9387: out = 24'(62872);
			9388: out = 24'(-15420);
			9389: out = 24'(-58008);
			9390: out = 24'(-43012);
			9391: out = 24'(2688);
			9392: out = 24'(33152);
			9393: out = 24'(42072);
			9394: out = 24'(18824);
			9395: out = 24'(-28600);
			9396: out = 24'(-6932);
			9397: out = 24'(-22772);
			9398: out = 24'(-36492);
			9399: out = 24'(-27472);
			9400: out = 24'(40668);
			9401: out = 24'(44096);
			9402: out = 24'(36380);
			9403: out = 24'(21528);
			9404: out = 24'(12088);
			9405: out = 24'(-6548);
			9406: out = 24'(-1492);
			9407: out = 24'(-1944);
			9408: out = 24'(-19768);
			9409: out = 24'(-41984);
			9410: out = 24'(-11192);
			9411: out = 24'(24072);
			9412: out = 24'(8692);
			9413: out = 24'(-45316);
			9414: out = 24'(-19792);
			9415: out = 24'(49304);
			9416: out = 24'(57208);
			9417: out = 24'(19180);
			9418: out = 24'(-9904);
			9419: out = 24'(2492);
			9420: out = 24'(-5568);
			9421: out = 24'(-24320);
			9422: out = 24'(-55756);
			9423: out = 24'(-3588);
			9424: out = 24'(36072);
			9425: out = 24'(16780);
			9426: out = 24'(-54056);
			9427: out = 24'(-16364);
			9428: out = 24'(29288);
			9429: out = 24'(-7100);
			9430: out = 24'(-55628);
			9431: out = 24'(-2028);
			9432: out = 24'(50960);
			9433: out = 24'(18204);
			9434: out = 24'(5976);
			9435: out = 24'(37504);
			9436: out = 24'(56528);
			9437: out = 24'(1896);
			9438: out = 24'(-81852);
			9439: out = 24'(-71912);
			9440: out = 24'(-18972);
			9441: out = 24'(6112);
			9442: out = 24'(30680);
			9443: out = 24'(25860);
			9444: out = 24'(15020);
			9445: out = 24'(-31768);
			9446: out = 24'(-85080);
			9447: out = 24'(-17952);
			9448: out = 24'(33452);
			9449: out = 24'(26544);
			9450: out = 24'(2212);
			9451: out = 24'(4732);
			9452: out = 24'(23724);
			9453: out = 24'(18696);
			9454: out = 24'(-1712);
			9455: out = 24'(-6148);
			9456: out = 24'(-1244);
			9457: out = 24'(-6032);
			9458: out = 24'(-9092);
			9459: out = 24'(5764);
			9460: out = 24'(8316);
			9461: out = 24'(540);
			9462: out = 24'(8164);
			9463: out = 24'(29708);
			9464: out = 24'(8844);
			9465: out = 24'(-20452);
			9466: out = 24'(-5580);
			9467: out = 24'(34388);
			9468: out = 24'(7240);
			9469: out = 24'(-62456);
			9470: out = 24'(-65840);
			9471: out = 24'(28168);
			9472: out = 24'(35104);
			9473: out = 24'(23384);
			9474: out = 24'(-8112);
			9475: out = 24'(-11316);
			9476: out = 24'(-33148);
			9477: out = 24'(-4736);
			9478: out = 24'(11280);
			9479: out = 24'(43872);
			9480: out = 24'(66360);
			9481: out = 24'(32916);
			9482: out = 24'(-49504);
			9483: out = 24'(-86988);
			9484: out = 24'(-5096);
			9485: out = 24'(47192);
			9486: out = 24'(47532);
			9487: out = 24'(-17996);
			9488: out = 24'(-70524);
			9489: out = 24'(-15748);
			9490: out = 24'(27320);
			9491: out = 24'(20564);
			9492: out = 24'(-5960);
			9493: out = 24'(-47936);
			9494: out = 24'(8720);
			9495: out = 24'(22856);
			9496: out = 24'(-16208);
			9497: out = 24'(-56864);
			9498: out = 24'(7332);
			9499: out = 24'(43112);
			9500: out = 24'(26868);
			9501: out = 24'(8584);
			9502: out = 24'(13636);
			9503: out = 24'(19884);
			9504: out = 24'(5528);
			9505: out = 24'(-20988);
			9506: out = 24'(-22808);
			9507: out = 24'(-33556);
			9508: out = 24'(-29248);
			9509: out = 24'(-4316);
			9510: out = 24'(26312);
			9511: out = 24'(5924);
			9512: out = 24'(-3076);
			9513: out = 24'(20392);
			9514: out = 24'(23104);
			9515: out = 24'(6580);
			9516: out = 24'(-24656);
			9517: out = 24'(-22084);
			9518: out = 24'(-7416);
			9519: out = 24'(40252);
			9520: out = 24'(11768);
			9521: out = 24'(-11516);
			9522: out = 24'(6688);
			9523: out = 24'(12832);
			9524: out = 24'(-15200);
			9525: out = 24'(-20372);
			9526: out = 24'(20316);
			9527: out = 24'(42828);
			9528: out = 24'(23740);
			9529: out = 24'(8556);
			9530: out = 24'(16664);
			9531: out = 24'(1712);
			9532: out = 24'(-30424);
			9533: out = 24'(-39796);
			9534: out = 24'(-6424);
			9535: out = 24'(7592);
			9536: out = 24'(28008);
			9537: out = 24'(8560);
			9538: out = 24'(-17700);
			9539: out = 24'(-42148);
			9540: out = 24'(4948);
			9541: out = 24'(7248);
			9542: out = 24'(-2148);
			9543: out = 24'(3268);
			9544: out = 24'(33548);
			9545: out = 24'(18520);
			9546: out = 24'(-11612);
			9547: out = 24'(-20468);
			9548: out = 24'(8628);
			9549: out = 24'(23776);
			9550: out = 24'(20380);
			9551: out = 24'(6216);
			9552: out = 24'(156);
			9553: out = 24'(-2684);
			9554: out = 24'(-6188);
			9555: out = 24'(-20388);
			9556: out = 24'(-27504);
			9557: out = 24'(624);
			9558: out = 24'(29920);
			9559: out = 24'(8168);
			9560: out = 24'(-50048);
			9561: out = 24'(-24272);
			9562: out = 24'(41244);
			9563: out = 24'(72528);
			9564: out = 24'(28524);
			9565: out = 24'(-16560);
			9566: out = 24'(-27056);
			9567: out = 24'(-1908);
			9568: out = 24'(-12020);
			9569: out = 24'(-12112);
			9570: out = 24'(-62984);
			9571: out = 24'(-11020);
			9572: out = 24'(55532);
			9573: out = 24'(46048);
			9574: out = 24'(-3668);
			9575: out = 24'(-2028);
			9576: out = 24'(15924);
			9577: out = 24'(1072);
			9578: out = 24'(-18688);
			9579: out = 24'(1388);
			9580: out = 24'(5672);
			9581: out = 24'(-32248);
			9582: out = 24'(-49060);
			9583: out = 24'(-432);
			9584: out = 24'(27500);
			9585: out = 24'(-2780);
			9586: out = 24'(2288);
			9587: out = 24'(4932);
			9588: out = 24'(-3192);
			9589: out = 24'(-38772);
			9590: out = 24'(-11468);
			9591: out = 24'(-11104);
			9592: out = 24'(31524);
			9593: out = 24'(39996);
			9594: out = 24'(27216);
			9595: out = 24'(-2624);
			9596: out = 24'(13976);
			9597: out = 24'(-14932);
			9598: out = 24'(-85012);
			9599: out = 24'(-40124);
			9600: out = 24'(22960);
			9601: out = 24'(23356);
			9602: out = 24'(-32616);
			9603: out = 24'(-27392);
			9604: out = 24'(-10108);
			9605: out = 24'(-3392);
			9606: out = 24'(-17224);
			9607: out = 24'(10012);
			9608: out = 24'(1692);
			9609: out = 24'(1340);
			9610: out = 24'(11380);
			9611: out = 24'(47988);
			9612: out = 24'(11912);
			9613: out = 24'(-5932);
			9614: out = 24'(-9136);
			9615: out = 24'(8056);
			9616: out = 24'(-1884);
			9617: out = 24'(240);
			9618: out = 24'(-5904);
			9619: out = 24'(-11376);
			9620: out = 24'(16);
			9621: out = 24'(4028);
			9622: out = 24'(15060);
			9623: out = 24'(26400);
			9624: out = 24'(3408);
			9625: out = 24'(-2004);
			9626: out = 24'(-8924);
			9627: out = 24'(16776);
			9628: out = 24'(53984);
			9629: out = 24'(9496);
			9630: out = 24'(-54796);
			9631: out = 24'(-54700);
			9632: out = 24'(32356);
			9633: out = 24'(15652);
			9634: out = 24'(6012);
			9635: out = 24'(-2144);
			9636: out = 24'(4852);
			9637: out = 24'(-18824);
			9638: out = 24'(-4360);
			9639: out = 24'(23292);
			9640: out = 24'(46632);
			9641: out = 24'(32948);
			9642: out = 24'(8900);
			9643: out = 24'(-23620);
			9644: out = 24'(-45216);
			9645: out = 24'(-62972);
			9646: out = 24'(-484);
			9647: out = 24'(33736);
			9648: out = 24'(27080);
			9649: out = 24'(-2520);
			9650: out = 24'(-560);
			9651: out = 24'(-19832);
			9652: out = 24'(-32056);
			9653: out = 24'(-12376);
			9654: out = 24'(11348);
			9655: out = 24'(33664);
			9656: out = 24'(29008);
			9657: out = 24'(10492);
			9658: out = 24'(-13020);
			9659: out = 24'(-14800);
			9660: out = 24'(-10180);
			9661: out = 24'(3452);
			9662: out = 24'(13612);
			9663: out = 24'(22316);
			9664: out = 24'(-104);
			9665: out = 24'(-28204);
			9666: out = 24'(-44532);
			9667: out = 24'(-42028);
			9668: out = 24'(-39536);
			9669: out = 24'(-5712);
			9670: out = 24'(47220);
			9671: out = 24'(67200);
			9672: out = 24'(15460);
			9673: out = 24'(-41844);
			9674: out = 24'(-44612);
			9675: out = 24'(31980);
			9676: out = 24'(-6096);
			9677: out = 24'(-29608);
			9678: out = 24'(20528);
			9679: out = 24'(55052);
			9680: out = 24'(36776);
			9681: out = 24'(-36844);
			9682: out = 24'(-73012);
			9683: out = 24'(-36700);
			9684: out = 24'(-3104);
			9685: out = 24'(-8020);
			9686: out = 24'(7844);
			9687: out = 24'(58880);
			9688: out = 24'(52756);
			9689: out = 24'(8132);
			9690: out = 24'(-20476);
			9691: out = 24'(5808);
			9692: out = 24'(-5284);
			9693: out = 24'(-864);
			9694: out = 24'(-22644);
			9695: out = 24'(-46172);
			9696: out = 24'(-60288);
			9697: out = 24'(-5280);
			9698: out = 24'(47692);
			9699: out = 24'(49712);
			9700: out = 24'(1432);
			9701: out = 24'(-2360);
			9702: out = 24'(21968);
			9703: out = 24'(42596);
			9704: out = 24'(20824);
			9705: out = 24'(-5036);
			9706: out = 24'(-9264);
			9707: out = 24'(22284);
			9708: out = 24'(33504);
			9709: out = 24'(6492);
			9710: out = 24'(-31896);
			9711: out = 24'(-25660);
			9712: out = 24'(-1964);
			9713: out = 24'(40);
			9714: out = 24'(-23528);
			9715: out = 24'(-400);
			9716: out = 24'(28024);
			9717: out = 24'(-14260);
			9718: out = 24'(-30028);
			9719: out = 24'(-4240);
			9720: out = 24'(32992);
			9721: out = 24'(22444);
			9722: out = 24'(8868);
			9723: out = 24'(14040);
			9724: out = 24'(23220);
			9725: out = 24'(184);
			9726: out = 24'(10808);
			9727: out = 24'(4104);
			9728: out = 24'(2004);
			9729: out = 24'(-6368);
			9730: out = 24'(-13512);
			9731: out = 24'(-56108);
			9732: out = 24'(-93272);
			9733: out = 24'(-73572);
			9734: out = 24'(6980);
			9735: out = 24'(42208);
			9736: out = 24'(21440);
			9737: out = 24'(1220);
			9738: out = 24'(18360);
			9739: out = 24'(54696);
			9740: out = 24'(24092);
			9741: out = 24'(-29904);
			9742: out = 24'(-38468);
			9743: out = 24'(-9424);
			9744: out = 24'(-9240);
			9745: out = 24'(-36040);
			9746: out = 24'(-31484);
			9747: out = 24'(29036);
			9748: out = 24'(53600);
			9749: out = 24'(30812);
			9750: out = 24'(-8692);
			9751: out = 24'(-40172);
			9752: out = 24'(-28728);
			9753: out = 24'(-3512);
			9754: out = 24'(3868);
			9755: out = 24'(-10816);
			9756: out = 24'(-3108);
			9757: out = 24'(16640);
			9758: out = 24'(27220);
			9759: out = 24'(15216);
			9760: out = 24'(2788);
			9761: out = 24'(2600);
			9762: out = 24'(272);
			9763: out = 24'(-20724);
			9764: out = 24'(-6544);
			9765: out = 24'(3384);
			9766: out = 24'(16608);
			9767: out = 24'(15164);
			9768: out = 24'(33876);
			9769: out = 24'(-6960);
			9770: out = 24'(-15376);
			9771: out = 24'(76);
			9772: out = 24'(-1752);
			9773: out = 24'(-2496);
			9774: out = 24'(24436);
			9775: out = 24'(52744);
			9776: out = 24'(32840);
			9777: out = 24'(-31860);
			9778: out = 24'(-59448);
			9779: out = 24'(-20364);
			9780: out = 24'(17092);
			9781: out = 24'(-4892);
			9782: out = 24'(-41876);
			9783: out = 24'(-29688);
			9784: out = 24'(23940);
			9785: out = 24'(29184);
			9786: out = 24'(29824);
			9787: out = 24'(24352);
			9788: out = 24'(27220);
			9789: out = 24'(27924);
			9790: out = 24'(-26504);
			9791: out = 24'(-69724);
			9792: out = 24'(-37416);
			9793: out = 24'(45416);
			9794: out = 24'(-3796);
			9795: out = 24'(-63992);
			9796: out = 24'(-45564);
			9797: out = 24'(54216);
			9798: out = 24'(21496);
			9799: out = 24'(6748);
			9800: out = 24'(16048);
			9801: out = 24'(33636);
			9802: out = 24'(2300);
			9803: out = 24'(-35920);
			9804: out = 24'(-46524);
			9805: out = 24'(-13248);
			9806: out = 24'(33548);
			9807: out = 24'(16452);
			9808: out = 24'(-1356);
			9809: out = 24'(0);
			9810: out = 24'(-1216);
			9811: out = 24'(-5492);
			9812: out = 24'(-248);
			9813: out = 24'(20336);
			9814: out = 24'(38012);
			9815: out = 24'(4876);
			9816: out = 24'(-19116);
			9817: out = 24'(-22124);
			9818: out = 24'(2668);
			9819: out = 24'(10096);
			9820: out = 24'(33824);
			9821: out = 24'(11736);
			9822: out = 24'(-35180);
			9823: out = 24'(-14640);
			9824: out = 24'(-3060);
			9825: out = 24'(-12300);
			9826: out = 24'(-31996);
			9827: out = 24'(-12108);
			9828: out = 24'(-12352);
			9829: out = 24'(-20436);
			9830: out = 24'(-32256);
			9831: out = 24'(-26692);
			9832: out = 24'(18300);
			9833: out = 24'(32924);
			9834: out = 24'(23800);
			9835: out = 24'(25468);
			9836: out = 24'(46020);
			9837: out = 24'(38992);
			9838: out = 24'(5124);
			9839: out = 24'(-32148);
			9840: out = 24'(-67836);
			9841: out = 24'(-36872);
			9842: out = 24'(13204);
			9843: out = 24'(30172);
			9844: out = 24'(23392);
			9845: out = 24'(-45900);
			9846: out = 24'(-65520);
			9847: out = 24'(-12780);
			9848: out = 24'(39280);
			9849: out = 24'(30632);
			9850: out = 24'(12260);
			9851: out = 24'(19268);
			9852: out = 24'(26344);
			9853: out = 24'(-34740);
			9854: out = 24'(-34148);
			9855: out = 24'(43372);
			9856: out = 24'(84268);
			9857: out = 24'(37548);
			9858: out = 24'(-43040);
			9859: out = 24'(-35292);
			9860: out = 24'(29296);
			9861: out = 24'(-1028);
			9862: out = 24'(-61748);
			9863: out = 24'(-60308);
			9864: out = 24'(27176);
			9865: out = 24'(58544);
			9866: out = 24'(-64);
			9867: out = 24'(-76956);
			9868: out = 24'(-74636);
			9869: out = 24'(4512);
			9870: out = 24'(42936);
			9871: out = 24'(40860);
			9872: out = 24'(31780);
			9873: out = 24'(35908);
			9874: out = 24'(764);
			9875: out = 24'(-9300);
			9876: out = 24'(-12616);
			9877: out = 24'(4328);
			9878: out = 24'(10628);
			9879: out = 24'(22828);
			9880: out = 24'(-21264);
			9881: out = 24'(-80692);
			9882: out = 24'(-108112);
			9883: out = 24'(12180);
			9884: out = 24'(68652);
			9885: out = 24'(26220);
			9886: out = 24'(-36636);
			9887: out = 24'(21508);
			9888: out = 24'(31524);
			9889: out = 24'(-27208);
			9890: out = 24'(-87752);
			9891: out = 24'(-4488);
			9892: out = 24'(39356);
			9893: out = 24'(18672);
			9894: out = 24'(-13620);
			9895: out = 24'(35128);
			9896: out = 24'(34212);
			9897: out = 24'(5048);
			9898: out = 24'(-36460);
			9899: out = 24'(-25528);
			9900: out = 24'(-26492);
			9901: out = 24'(15940);
			9902: out = 24'(39524);
			9903: out = 24'(12176);
			9904: out = 24'(-34260);
			9905: out = 24'(3468);
			9906: out = 24'(62876);
			9907: out = 24'(27944);
			9908: out = 24'(-27988);
			9909: out = 24'(-71552);
			9910: out = 24'(-30968);
			9911: out = 24'(15892);
			9912: out = 24'(7544);
			9913: out = 24'(-26340);
			9914: out = 24'(-312);
			9915: out = 24'(44920);
			9916: out = 24'(28984);
			9917: out = 24'(-36672);
			9918: out = 24'(-62296);
			9919: out = 24'(-28252);
			9920: out = 24'(972);
			9921: out = 24'(-1276);
			9922: out = 24'(6528);
			9923: out = 24'(26052);
			9924: out = 24'(34076);
			9925: out = 24'(27988);
			9926: out = 24'(43616);
			9927: out = 24'(34412);
			9928: out = 24'(-28680);
			9929: out = 24'(-67252);
			9930: out = 24'(-63360);
			9931: out = 24'(-16952);
			9932: out = 24'(10260);
			9933: out = 24'(31068);
			9934: out = 24'(36368);
			9935: out = 24'(50948);
			9936: out = 24'(42052);
			9937: out = 24'(13320);
			9938: out = 24'(-32636);
			9939: out = 24'(-37872);
			9940: out = 24'(-15420);
			9941: out = 24'(7436);
			9942: out = 24'(768);
			9943: out = 24'(11240);
			9944: out = 24'(13412);
			9945: out = 24'(-388);
			9946: out = 24'(-896);
			9947: out = 24'(30192);
			9948: out = 24'(44156);
			9949: out = 24'(20088);
			9950: out = 24'(6856);
			9951: out = 24'(-13608);
			9952: out = 24'(-20616);
			9953: out = 24'(-3292);
			9954: out = 24'(36508);
			9955: out = 24'(30740);
			9956: out = 24'(-15436);
			9957: out = 24'(-48960);
			9958: out = 24'(-12208);
			9959: out = 24'(-1804);
			9960: out = 24'(-12328);
			9961: out = 24'(-22432);
			9962: out = 24'(1484);
			9963: out = 24'(-968);
			9964: out = 24'(12080);
			9965: out = 24'(31944);
			9966: out = 24'(41056);
			9967: out = 24'(4028);
			9968: out = 24'(-2284);
			9969: out = 24'(16168);
			9970: out = 24'(19340);
			9971: out = 24'(2972);
			9972: out = 24'(-59884);
			9973: out = 24'(-62996);
			9974: out = 24'(-11672);
			9975: out = 24'(14764);
			9976: out = 24'(8048);
			9977: out = 24'(12112);
			9978: out = 24'(1968);
			9979: out = 24'(-60000);
			9980: out = 24'(-109916);
			9981: out = 24'(-63960);
			9982: out = 24'(41356);
			9983: out = 24'(70232);
			9984: out = 24'(47652);
			9985: out = 24'(9236);
			9986: out = 24'(172);
			9987: out = 24'(2992);
			9988: out = 24'(32528);
			9989: out = 24'(17572);
			9990: out = 24'(-260);
			9991: out = 24'(-21360);
			9992: out = 24'(2184);
			9993: out = 24'(-86768);
			9994: out = 24'(-88116);
			9995: out = 24'(5120);
			9996: out = 24'(65548);
			9997: out = 24'(41144);
			9998: out = 24'(5156);
			9999: out = 24'(-4160);
			10000: out = 24'(-1620);
			10001: out = 24'(-8472);
			10002: out = 24'(-14228);
			10003: out = 24'(-520);
			10004: out = 24'(18188);
			10005: out = 24'(8344);
			10006: out = 24'(1612);
			10007: out = 24'(2488);
			10008: out = 24'(7648);
			10009: out = 24'(11980);
			10010: out = 24'(-26020);
			10011: out = 24'(-33108);
			10012: out = 24'(26672);
			10013: out = 24'(79840);
			10014: out = 24'(63368);
			10015: out = 24'(-27524);
			10016: out = 24'(-96096);
			10017: out = 24'(-48684);
			10018: out = 24'(-10724);
			10019: out = 24'(30260);
			10020: out = 24'(46508);
			10021: out = 24'(41620);
			10022: out = 24'(-20);
			10023: out = 24'(-26528);
			10024: out = 24'(-17348);
			10025: out = 24'(14920);
			10026: out = 24'(4556);
			10027: out = 24'(2040);
			10028: out = 24'(-1780);
			10029: out = 24'(-2184);
			10030: out = 24'(-24856);
			10031: out = 24'(6880);
			10032: out = 24'(27088);
			10033: out = 24'(28028);
			10034: out = 24'(8616);
			10035: out = 24'(7692);
			10036: out = 24'(-21708);
			10037: out = 24'(-46916);
			10038: out = 24'(-26192);
			10039: out = 24'(-29384);
			10040: out = 24'(10736);
			10041: out = 24'(32868);
			10042: out = 24'(29172);
			10043: out = 24'(-148);
			10044: out = 24'(11612);
			10045: out = 24'(4720);
			10046: out = 24'(-25956);
			10047: out = 24'(-35084);
			10048: out = 24'(-34428);
			10049: out = 24'(-16388);
			10050: out = 24'(18620);
			10051: out = 24'(68424);
			10052: out = 24'(47748);
			10053: out = 24'(11388);
			10054: out = 24'(-27832);
			10055: out = 24'(-48992);
			10056: out = 24'(-29444);
			10057: out = 24'(-16388);
			10058: out = 24'(-2472);
			10059: out = 24'(21528);
			10060: out = 24'(25612);
			10061: out = 24'(28932);
			10062: out = 24'(25428);
			10063: out = 24'(28212);
			10064: out = 24'(28392);
			10065: out = 24'(-5648);
			10066: out = 24'(-66092);
			10067: out = 24'(-99592);
			10068: out = 24'(-40768);
			10069: out = 24'(-14180);
			10070: out = 24'(17828);
			10071: out = 24'(42848);
			10072: out = 24'(53628);
			10073: out = 24'(15096);
			10074: out = 24'(-20856);
			10075: out = 24'(-36640);
			10076: out = 24'(-17848);
			10077: out = 24'(2116);
			10078: out = 24'(8220);
			10079: out = 24'(-10664);
			10080: out = 24'(-15148);
			10081: out = 24'(23616);
			10082: out = 24'(43268);
			10083: out = 24'(11388);
			10084: out = 24'(-38024);
			10085: out = 24'(-38556);
			10086: out = 24'(-19716);
			10087: out = 24'(-7092);
			10088: out = 24'(-9984);
			10089: out = 24'(7188);
			10090: out = 24'(33980);
			10091: out = 24'(41004);
			10092: out = 24'(6716);
			10093: out = 24'(-26736);
			10094: out = 24'(-11544);
			10095: out = 24'(11484);
			10096: out = 24'(-2796);
			10097: out = 24'(-26580);
			10098: out = 24'(-2752);
			10099: out = 24'(30748);
			10100: out = 24'(22288);
			10101: out = 24'(-9420);
			10102: out = 24'(2868);
			10103: out = 24'(50744);
			10104: out = 24'(67308);
			10105: out = 24'(24052);
			10106: out = 24'(-41352);
			10107: out = 24'(-52416);
			10108: out = 24'(-23264);
			10109: out = 24'(6092);
			10110: out = 24'(5184);
			10111: out = 24'(31108);
			10112: out = 24'(12044);
			10113: out = 24'(-4812);
			10114: out = 24'(-7812);
			10115: out = 24'(-11944);
			10116: out = 24'(-7036);
			10117: out = 24'(8624);
			10118: out = 24'(14488);
			10119: out = 24'(13100);
			10120: out = 24'(-22568);
			10121: out = 24'(-16412);
			10122: out = 24'(13468);
			10123: out = 24'(25432);
			10124: out = 24'(-20088);
			10125: out = 24'(-424);
			10126: out = 24'(47944);
			10127: out = 24'(30784);
			10128: out = 24'(9772);
			10129: out = 24'(-42168);
			10130: out = 24'(-69508);
			10131: out = 24'(-72132);
			10132: out = 24'(-21280);
			10133: out = 24'(-4684);
			10134: out = 24'(11696);
			10135: out = 24'(25400);
			10136: out = 24'(33356);
			10137: out = 24'(17036);
			10138: out = 24'(13560);
			10139: out = 24'(12788);
			10140: out = 24'(-12128);
			10141: out = 24'(-30928);
			10142: out = 24'(-26556);
			10143: out = 24'(-2708);
			10144: out = 24'(5428);
			10145: out = 24'(3760);
			10146: out = 24'(-2732);
			10147: out = 24'(12380);
			10148: out = 24'(38032);
			10149: out = 24'(32440);
			10150: out = 24'(-932);
			10151: out = 24'(-39676);
			10152: out = 24'(-38972);
			10153: out = 24'(5316);
			10154: out = 24'(35192);
			10155: out = 24'(25288);
			10156: out = 24'(13276);
			10157: out = 24'(23552);
			10158: out = 24'(-1356);
			10159: out = 24'(-58428);
			10160: out = 24'(-69960);
			10161: out = 24'(30328);
			10162: out = 24'(32904);
			10163: out = 24'(15204);
			10164: out = 24'(4360);
			10165: out = 24'(27680);
			10166: out = 24'(-3236);
			10167: out = 24'(-15212);
			10168: out = 24'(-10000);
			10169: out = 24'(15796);
			10170: out = 24'(23696);
			10171: out = 24'(18440);
			10172: out = 24'(-2572);
			10173: out = 24'(-20700);
			10174: out = 24'(-23140);
			10175: out = 24'(11104);
			10176: out = 24'(40740);
			10177: out = 24'(38240);
			10178: out = 24'(25884);
			10179: out = 24'(-22944);
			10180: out = 24'(-20688);
			10181: out = 24'(8564);
			10182: out = 24'(25888);
			10183: out = 24'(-65616);
			10184: out = 24'(-65220);
			10185: out = 24'(3300);
			10186: out = 24'(48516);
			10187: out = 24'(28860);
			10188: out = 24'(20480);
			10189: out = 24'(21900);
			10190: out = 24'(23656);
			10191: out = 24'(7952);
			10192: out = 24'(3648);
			10193: out = 24'(-33820);
			10194: out = 24'(-85184);
			10195: out = 24'(-86224);
			10196: out = 24'(-34760);
			10197: out = 24'(27144);
			10198: out = 24'(58736);
			10199: out = 24'(69464);
			10200: out = 24'(49592);
			10201: out = 24'(1080);
			10202: out = 24'(-61832);
			10203: out = 24'(-88068);
			10204: out = 24'(-42832);
			10205: out = 24'(4048);
			10206: out = 24'(8628);
			10207: out = 24'(2040);
			10208: out = 24'(-2308);
			10209: out = 24'(29632);
			10210: out = 24'(25968);
			10211: out = 24'(1792);
			10212: out = 24'(512);
			10213: out = 24'(2600);
			10214: out = 24'(-17440);
			10215: out = 24'(-29560);
			10216: out = 24'(13784);
			10217: out = 24'(16588);
			10218: out = 24'(8280);
			10219: out = 24'(4308);
			10220: out = 24'(21908);
			10221: out = 24'(2048);
			10222: out = 24'(-12544);
			10223: out = 24'(-16892);
			10224: out = 24'(-11460);
			10225: out = 24'(472);
			10226: out = 24'(-28696);
			10227: out = 24'(-24508);
			10228: out = 24'(30668);
			10229: out = 24'(43868);
			10230: out = 24'(24028);
			10231: out = 24'(-31636);
			10232: out = 24'(-56304);
			10233: out = 24'(-16488);
			10234: out = 24'(23488);
			10235: out = 24'(33700);
			10236: out = 24'(20000);
			10237: out = 24'(6188);
			10238: out = 24'(348);
			10239: out = 24'(672);
			10240: out = 24'(-276);
			10241: out = 24'(820);
			10242: out = 24'(-428);
			10243: out = 24'(-9488);
			10244: out = 24'(-26068);
			10245: out = 24'(-24476);
			10246: out = 24'(-2464);
			10247: out = 24'(23212);
			10248: out = 24'(20712);
			10249: out = 24'(10748);
			10250: out = 24'(4528);
			10251: out = 24'(33332);
			10252: out = 24'(508);
			10253: out = 24'(-47436);
			10254: out = 24'(-10476);
			10255: out = 24'(5824);
			10256: out = 24'(34540);
			10257: out = 24'(24228);
			10258: out = 24'(-844);
			10259: out = 24'(-13232);
			10260: out = 24'(-5068);
			10261: out = 24'(-1284);
			10262: out = 24'(2812);
			10263: out = 24'(12836);
			10264: out = 24'(8340);
			10265: out = 24'(-22288);
			10266: out = 24'(-36688);
			10267: out = 24'(-3896);
			10268: out = 24'(31852);
			10269: out = 24'(12836);
			10270: out = 24'(-26372);
			10271: out = 24'(-25732);
			10272: out = 24'(41236);
			10273: out = 24'(54144);
			10274: out = 24'(18840);
			10275: out = 24'(728);
			10276: out = 24'(9592);
			10277: out = 24'(9028);
			10278: out = 24'(-18772);
			10279: out = 24'(-33640);
			10280: out = 24'(-2916);
			10281: out = 24'(12496);
			10282: out = 24'(-1288);
			10283: out = 24'(-9584);
			10284: out = 24'(12556);
			10285: out = 24'(6548);
			10286: out = 24'(-20168);
			10287: out = 24'(-18984);
			10288: out = 24'(33384);
			10289: out = 24'(31236);
			10290: out = 24'(-11936);
			10291: out = 24'(-38308);
			10292: out = 24'(14484);
			10293: out = 24'(-2300);
			10294: out = 24'(172);
			10295: out = 24'(-4172);
			10296: out = 24'(-2460);
			10297: out = 24'(-30104);
			10298: out = 24'(-12720);
			10299: out = 24'(4368);
			10300: out = 24'(4200);
			10301: out = 24'(36);
			10302: out = 24'(-21744);
			10303: out = 24'(-23324);
			10304: out = 24'(18824);
			10305: out = 24'(71764);
			10306: out = 24'(39556);
			10307: out = 24'(-29236);
			10308: out = 24'(-67588);
			10309: out = 24'(-27928);
			10310: out = 24'(-2076);
			10311: out = 24'(13232);
			10312: out = 24'(20184);
			10313: out = 24'(22892);
			10314: out = 24'(-11596);
			10315: out = 24'(-37080);
			10316: out = 24'(-34600);
			10317: out = 24'(-18868);
			10318: out = 24'(-37996);
			10319: out = 24'(-32576);
			10320: out = 24'(2412);
			10321: out = 24'(26732);
			10322: out = 24'(2724);
			10323: out = 24'(-11280);
			10324: out = 24'(18448);
			10325: out = 24'(59456);
			10326: out = 24'(59116);
			10327: out = 24'(16692);
			10328: out = 24'(-2364);
			10329: out = 24'(-4820);
			10330: out = 24'(-22880);
			10331: out = 24'(-60824);
			10332: out = 24'(-52056);
			10333: out = 24'(-6412);
			10334: out = 24'(25040);
			10335: out = 24'(37084);
			10336: out = 24'(24784);
			10337: out = 24'(8256);
			10338: out = 24'(1384);
			10339: out = 24'(4228);
			10340: out = 24'(7760);
			10341: out = 24'(-5748);
			10342: out = 24'(-20980);
			10343: out = 24'(-30716);
			10344: out = 24'(-9176);
			10345: out = 24'(-5184);
			10346: out = 24'(19480);
			10347: out = 24'(71724);
			10348: out = 24'(73072);
			10349: out = 24'(7028);
			10350: out = 24'(-65704);
			10351: out = 24'(-67272);
			10352: out = 24'(-18140);
			10353: out = 24'(4572);
			10354: out = 24'(-8304);
			10355: out = 24'(-5260);
			10356: out = 24'(13168);
			10357: out = 24'(38472);
			10358: out = 24'(24500);
			10359: out = 24'(-4280);
			10360: out = 24'(540);
			10361: out = 24'(-24984);
			10362: out = 24'(-23584);
			10363: out = 24'(-8716);
			10364: out = 24'(-11180);
			10365: out = 24'(33796);
			10366: out = 24'(41672);
			10367: out = 24'(24636);
			10368: out = 24'(-3784);
			10369: out = 24'(668);
			10370: out = 24'(-2916);
			10371: out = 24'(1732);
			10372: out = 24'(2876);
			10373: out = 24'(1784);
			10374: out = 24'(-13004);
			10375: out = 24'(9304);
			10376: out = 24'(50320);
			10377: out = 24'(47872);
			10378: out = 24'(-6604);
			10379: out = 24'(-68776);
			10380: out = 24'(-83496);
			10381: out = 24'(-31256);
			10382: out = 24'(-49840);
			10383: out = 24'(-37536);
			10384: out = 24'(16604);
			10385: out = 24'(69096);
			10386: out = 24'(60256);
			10387: out = 24'(36952);
			10388: out = 24'(2636);
			10389: out = 24'(-23144);
			10390: out = 24'(7036);
			10391: out = 24'(-11556);
			10392: out = 24'(-58020);
			10393: out = 24'(-80348);
			10394: out = 24'(-9640);
			10395: out = 24'(23608);
			10396: out = 24'(21736);
			10397: out = 24'(19796);
			10398: out = 24'(58900);
			10399: out = 24'(30412);
			10400: out = 24'(-6436);
			10401: out = 24'(-31476);
			10402: out = 24'(-10060);
			10403: out = 24'(-38924);
			10404: out = 24'(-28740);
			10405: out = 24'(-7484);
			10406: out = 24'(9580);
			10407: out = 24'(15460);
			10408: out = 24'(32492);
			10409: out = 24'(22876);
			10410: out = 24'(-22276);
			10411: out = 24'(-53580);
			10412: out = 24'(-25980);
			10413: out = 24'(28392);
			10414: out = 24'(23056);
			10415: out = 24'(-21060);
			10416: out = 24'(-56732);
			10417: out = 24'(-4180);
			10418: out = 24'(47968);
			10419: out = 24'(33860);
			10420: out = 24'(-63948);
			10421: out = 24'(-62464);
			10422: out = 24'(20096);
			10423: out = 24'(67784);
			10424: out = 24'(61956);
			10425: out = 24'(40164);
			10426: out = 24'(8920);
			10427: out = 24'(-21548);
			10428: out = 24'(-53992);
			10429: out = 24'(-31916);
			10430: out = 24'(-30572);
			10431: out = 24'(-40348);
			10432: out = 24'(600);
			10433: out = 24'(47288);
			10434: out = 24'(40256);
			10435: out = 24'(20724);
			10436: out = 24'(50644);
			10437: out = 24'(72256);
			10438: out = 24'(13228);
			10439: out = 24'(-68432);
			10440: out = 24'(-59116);
			10441: out = 24'(-5204);
			10442: out = 24'(14208);
			10443: out = 24'(-7724);
			10444: out = 24'(10156);
			10445: out = 24'(23052);
			10446: out = 24'(41796);
			10447: out = 24'(21904);
			10448: out = 24'(4908);
			10449: out = 24'(-75432);
			10450: out = 24'(-20776);
			10451: out = 24'(5056);
			10452: out = 24'(-1628);
			10453: out = 24'(-24232);
			10454: out = 24'(34900);
			10455: out = 24'(26132);
			10456: out = 24'(-3616);
			10457: out = 24'(-696);
			10458: out = 24'(17088);
			10459: out = 24'(-9160);
			10460: out = 24'(-6736);
			10461: out = 24'(45048);
			10462: out = 24'(22120);
			10463: out = 24'(-40332);
			10464: out = 24'(-48480);
			10465: out = 24'(22540);
			10466: out = 24'(-12952);
			10467: out = 24'(-40364);
			10468: out = 24'(-43556);
			10469: out = 24'(-4792);
			10470: out = 24'(-19148);
			10471: out = 24'(9736);
			10472: out = 24'(36176);
			10473: out = 24'(43744);
			10474: out = 24'(-900);
			10475: out = 24'(3972);
			10476: out = 24'(18784);
			10477: out = 24'(9824);
			10478: out = 24'(-60372);
			10479: out = 24'(-52900);
			10480: out = 24'(-46256);
			10481: out = 24'(-20204);
			10482: out = 24'(9920);
			10483: out = 24'(60568);
			10484: out = 24'(69860);
			10485: out = 24'(47524);
			10486: out = 24'(-4872);
			10487: out = 24'(-60996);
			10488: out = 24'(-57136);
			10489: out = 24'(-15200);
			10490: out = 24'(-5244);
			10491: out = 24'(-35724);
			10492: out = 24'(-12972);
			10493: out = 24'(43652);
			10494: out = 24'(66756);
			10495: out = 24'(42964);
			10496: out = 24'(5168);
			10497: out = 24'(-6964);
			10498: out = 24'(-31160);
			10499: out = 24'(-75296);
			10500: out = 24'(-58120);
			10501: out = 24'(4480);
			10502: out = 24'(41012);
			10503: out = 24'(23144);
			10504: out = 24'(21828);
			10505: out = 24'(22564);
			10506: out = 24'(31088);
			10507: out = 24'(18720);
			10508: out = 24'(-11168);
			10509: out = 24'(-50056);
			10510: out = 24'(-56024);
			10511: out = 24'(-14720);
			10512: out = 24'(26112);
			10513: out = 24'(41740);
			10514: out = 24'(4884);
			10515: out = 24'(-14960);
			10516: out = 24'(2048);
			10517: out = 24'(4056);
			10518: out = 24'(-33736);
			10519: out = 24'(-43648);
			10520: out = 24'(7416);
			10521: out = 24'(42424);
			10522: out = 24'(36804);
			10523: out = 24'(24188);
			10524: out = 24'(29452);
			10525: out = 24'(29700);
			10526: out = 24'(-13244);
			10527: out = 24'(-37408);
			10528: out = 24'(-23756);
			10529: out = 24'(-19824);
			10530: out = 24'(-296);
			10531: out = 24'(-7108);
			10532: out = 24'(-3336);
			10533: out = 24'(26264);
			10534: out = 24'(33504);
			10535: out = 24'(39564);
			10536: out = 24'(24092);
			10537: out = 24'(1060);
			10538: out = 24'(-13420);
			10539: out = 24'(-11644);
			10540: out = 24'(-25904);
			10541: out = 24'(-34872);
			10542: out = 24'(25220);
			10543: out = 24'(52180);
			10544: out = 24'(44048);
			10545: out = 24'(7956);
			10546: out = 24'(-11600);
			10547: out = 24'(-30492);
			10548: out = 24'(-30980);
			10549: out = 24'(-30528);
			10550: out = 24'(-21908);
			10551: out = 24'(-20592);
			10552: out = 24'(11752);
			10553: out = 24'(47996);
			10554: out = 24'(64636);
			10555: out = 24'(36932);
			10556: out = 24'(12520);
			10557: out = 24'(-22128);
			10558: out = 24'(-53568);
			10559: out = 24'(-62292);
			10560: out = 24'(-19640);
			10561: out = 24'(14680);
			10562: out = 24'(10156);
			10563: out = 24'(-9248);
			10564: out = 24'(3708);
			10565: out = 24'(23412);
			10566: out = 24'(19604);
			10567: out = 24'(-812);
			10568: out = 24'(-1440);
			10569: out = 24'(1420);
			10570: out = 24'(-9252);
			10571: out = 24'(-21784);
			10572: out = 24'(-3948);
			10573: out = 24'(25900);
			10574: out = 24'(32112);
			10575: out = 24'(6760);
			10576: out = 24'(-43580);
			10577: out = 24'(-39736);
			10578: out = 24'(-15972);
			10579: out = 24'(7248);
			10580: out = 24'(35480);
			10581: out = 24'(6520);
			10582: out = 24'(-17820);
			10583: out = 24'(-3828);
			10584: out = 24'(34520);
			10585: out = 24'(23720);
			10586: out = 24'(-9040);
			10587: out = 24'(-17752);
			10588: out = 24'(7556);
			10589: out = 24'(26028);
			10590: out = 24'(-7448);
			10591: out = 24'(-27904);
			10592: out = 24'(8884);
			10593: out = 24'(43624);
			10594: out = 24'(-1360);
			10595: out = 24'(-59912);
			10596: out = 24'(-43624);
			10597: out = 24'(18000);
			10598: out = 24'(36136);
			10599: out = 24'(72);
			10600: out = 24'(-5548);
			10601: out = 24'(36444);
			10602: out = 24'(36340);
			10603: out = 24'(-29868);
			10604: out = 24'(-66516);
			10605: out = 24'(6808);
			10606: out = 24'(22108);
			10607: out = 24'(1580);
			10608: out = 24'(-30792);
			10609: out = 24'(-10844);
			10610: out = 24'(-11836);
			10611: out = 24'(13248);
			10612: out = 24'(17448);
			10613: out = 24'(22256);
			10614: out = 24'(-2188);
			10615: out = 24'(11636);
			10616: out = 24'(-968);
			10617: out = 24'(-10012);
			10618: out = 24'(-2480);
			10619: out = 24'(55604);
			10620: out = 24'(44688);
			10621: out = 24'(1436);
			10622: out = 24'(-17488);
			10623: out = 24'(9520);
			10624: out = 24'(-12748);
			10625: out = 24'(-55100);
			10626: out = 24'(-48780);
			10627: out = 24'(-20716);
			10628: out = 24'(4028);
			10629: out = 24'(11736);
			10630: out = 24'(31104);
			10631: out = 24'(22900);
			10632: out = 24'(30132);
			10633: out = 24'(8296);
			10634: out = 24'(-17744);
			10635: out = 24'(-36424);
			10636: out = 24'(17764);
			10637: out = 24'(36352);
			10638: out = 24'(2956);
			10639: out = 24'(-45548);
			10640: out = 24'(-12872);
			10641: out = 24'(9296);
			10642: out = 24'(-3560);
			10643: out = 24'(-15688);
			10644: out = 24'(-16400);
			10645: out = 24'(4372);
			10646: out = 24'(12624);
			10647: out = 24'(15376);
			10648: out = 24'(-23644);
			10649: out = 24'(9328);
			10650: out = 24'(31836);
			10651: out = 24'(26272);
			10652: out = 24'(-924);
			10653: out = 24'(-7868);
			10654: out = 24'(-22748);
			10655: out = 24'(-18048);
			10656: out = 24'(-6876);
			10657: out = 24'(6456);
			10658: out = 24'(-40916);
			10659: out = 24'(-51492);
			10660: out = 24'(20928);
			10661: out = 24'(80736);
			10662: out = 24'(36236);
			10663: out = 24'(-7856);
			10664: out = 24'(-3488);
			10665: out = 24'(-34436);
			10666: out = 24'(-77364);
			10667: out = 24'(-31476);
			10668: out = 24'(67924);
			10669: out = 24'(6632);
			10670: out = 24'(-21888);
			10671: out = 24'(-2704);
			10672: out = 24'(41896);
			10673: out = 24'(-3104);
			10674: out = 24'(-16124);
			10675: out = 24'(6284);
			10676: out = 24'(17552);
			10677: out = 24'(-71056);
			10678: out = 24'(-48860);
			10679: out = 24'(20256);
			10680: out = 24'(73164);
			10681: out = 24'(24296);
			10682: out = 24'(21628);
			10683: out = 24'(-11248);
			10684: out = 24'(-5416);
			10685: out = 24'(-3368);
			10686: out = 24'(8436);
			10687: out = 24'(-23868);
			10688: out = 24'(-20912);
			10689: out = 24'(-12140);
			10690: out = 24'(-50020);
			10691: out = 24'(10440);
			10692: out = 24'(74572);
			10693: out = 24'(45180);
			10694: out = 24'(-55368);
			10695: out = 24'(-79716);
			10696: out = 24'(6400);
			10697: out = 24'(48096);
			10698: out = 24'(-27080);
			10699: out = 24'(-3984);
			10700: out = 24'(35716);
			10701: out = 24'(21144);
			10702: out = 24'(-68768);
			10703: out = 24'(-47992);
			10704: out = 24'(1416);
			10705: out = 24'(27724);
			10706: out = 24'(-5804);
			10707: out = 24'(6464);
			10708: out = 24'(5848);
			10709: out = 24'(15572);
			10710: out = 24'(14272);
			10711: out = 24'(43308);
			10712: out = 24'(27796);
			10713: out = 24'(8680);
			10714: out = 24'(-21492);
			10715: out = 24'(-14828);
			10716: out = 24'(-48888);
			10717: out = 24'(-23992);
			10718: out = 24'(2784);
			10719: out = 24'(19348);
			10720: out = 24'(-2184);
			10721: out = 24'(32396);
			10722: out = 24'(34008);
			10723: out = 24'(-208);
			10724: out = 24'(-1248);
			10725: out = 24'(1952);
			10726: out = 24'(-21056);
			10727: out = 24'(-40716);
			10728: out = 24'(26876);
			10729: out = 24'(36492);
			10730: out = 24'(6220);
			10731: out = 24'(-36720);
			10732: out = 24'(-12688);
			10733: out = 24'(-7756);
			10734: out = 24'(7884);
			10735: out = 24'(3404);
			10736: out = 24'(8144);
			10737: out = 24'(-17936);
			10738: out = 24'(-5576);
			10739: out = 24'(-984);
			10740: out = 24'(1736);
			10741: out = 24'(-3644);
			10742: out = 24'(34616);
			10743: out = 24'(32288);
			10744: out = 24'(-5144);
			10745: out = 24'(-27856);
			10746: out = 24'(6676);
			10747: out = 24'(20172);
			10748: out = 24'(-4228);
			10749: out = 24'(-14288);
			10750: out = 24'(6012);
			10751: out = 24'(17212);
			10752: out = 24'(-14236);
			10753: out = 24'(-51608);
			10754: out = 24'(-22292);
			10755: out = 24'(8092);
			10756: out = 24'(6144);
			10757: out = 24'(3000);
			10758: out = 24'(12372);
			10759: out = 24'(21168);
			10760: out = 24'(5456);
			10761: out = 24'(4632);
			10762: out = 24'(9636);
			10763: out = 24'(32172);
			10764: out = 24'(-16972);
			10765: out = 24'(-53316);
			10766: out = 24'(8996);
			10767: out = 24'(37848);
			10768: out = 24'(-11904);
			10769: out = 24'(-44044);
			10770: out = 24'(31892);
			10771: out = 24'(55048);
			10772: out = 24'(5528);
			10773: out = 24'(-37624);
			10774: out = 24'(16080);
			10775: out = 24'(31252);
			10776: out = 24'(9020);
			10777: out = 24'(-35232);
			10778: out = 24'(-20272);
			10779: out = 24'(-3320);
			10780: out = 24'(20056);
			10781: out = 24'(-4416);
			10782: out = 24'(-26096);
			10783: out = 24'(-37888);
			10784: out = 24'(14468);
			10785: out = 24'(22364);
			10786: out = 24'(6228);
			10787: out = 24'(160);
			10788: out = 24'(30264);
			10789: out = 24'(18388);
			10790: out = 24'(-11024);
			10791: out = 24'(-15564);
			10792: out = 24'(5004);
			10793: out = 24'(-3092);
			10794: out = 24'(-36416);
			10795: out = 24'(-51324);
			10796: out = 24'(-27928);
			10797: out = 24'(33940);
			10798: out = 24'(77492);
			10799: out = 24'(69316);
			10800: out = 24'(-804);
			10801: out = 24'(-58148);
			10802: out = 24'(-71208);
			10803: out = 24'(-25444);
			10804: out = 24'(-4144);
			10805: out = 24'(40404);
			10806: out = 24'(16532);
			10807: out = 24'(-2196);
			10808: out = 24'(-1624);
			10809: out = 24'(44420);
			10810: out = 24'(-14184);
			10811: out = 24'(-58672);
			10812: out = 24'(-20868);
			10813: out = 24'(11200);
			10814: out = 24'(-6296);
			10815: out = 24'(-21980);
			10816: out = 24'(7488);
			10817: out = 24'(7784);
			10818: out = 24'(18216);
			10819: out = 24'(20452);
			10820: out = 24'(38188);
			10821: out = 24'(44652);
			10822: out = 24'(16488);
			10823: out = 24'(-24500);
			10824: out = 24'(-50276);
			10825: out = 24'(-67564);
			10826: out = 24'(-9748);
			10827: out = 24'(8284);
			10828: out = 24'(-1968);
			10829: out = 24'(-21396);
			10830: out = 24'(24732);
			10831: out = 24'(5100);
			10832: out = 24'(-26240);
			10833: out = 24'(-33708);
			10834: out = 24'(25748);
			10835: out = 24'(35244);
			10836: out = 24'(34556);
			10837: out = 24'(24960);
			10838: out = 24'(43784);
			10839: out = 24'(14880);
			10840: out = 24'(25772);
			10841: out = 24'(-6048);
			10842: out = 24'(-105396);
			10843: out = 24'(-123360);
			10844: out = 24'(-24140);
			10845: out = 24'(68256);
			10846: out = 24'(31232);
			10847: out = 24'(-51444);
			10848: out = 24'(-43236);
			10849: out = 24'(42072);
			10850: out = 24'(49240);
			10851: out = 24'(15344);
			10852: out = 24'(-76904);
			10853: out = 24'(-61384);
			10854: out = 24'(25888);
			10855: out = 24'(15144);
			10856: out = 24'(20904);
			10857: out = 24'(25564);
			10858: out = 24'(41548);
			10859: out = 24'(32708);
			10860: out = 24'(12024);
			10861: out = 24'(-25828);
			10862: out = 24'(-33484);
			10863: out = 24'(2728);
			10864: out = 24'(10372);
			10865: out = 24'(7232);
			10866: out = 24'(-1320);
			10867: out = 24'(4364);
			10868: out = 24'(27728);
			10869: out = 24'(16304);
			10870: out = 24'(-20116);
			10871: out = 24'(-35572);
			10872: out = 24'(-4320);
			10873: out = 24'(31048);
			10874: out = 24'(24488);
			10875: out = 24'(-1308);
			10876: out = 24'(-17540);
			10877: out = 24'(-2888);
			10878: out = 24'(-14160);
			10879: out = 24'(-25936);
			10880: out = 24'(4312);
			10881: out = 24'(33820);
			10882: out = 24'(44024);
			10883: out = 24'(32380);
			10884: out = 24'(12560);
			10885: out = 24'(1992);
			10886: out = 24'(-23080);
			10887: out = 24'(-20264);
			10888: out = 24'(6356);
			10889: out = 24'(-11760);
			10890: out = 24'(-37244);
			10891: out = 24'(-39132);
			10892: out = 24'(2712);
			10893: out = 24'(36740);
			10894: out = 24'(26624);
			10895: out = 24'(3876);
			10896: out = 24'(1956);
			10897: out = 24'(4356);
			10898: out = 24'(24356);
			10899: out = 24'(15056);
			10900: out = 24'(-6224);
			10901: out = 24'(-30416);
			10902: out = 24'(668);
			10903: out = 24'(1632);
			10904: out = 24'(-1540);
			10905: out = 24'(60);
			10906: out = 24'(20644);
			10907: out = 24'(12816);
			10908: out = 24'(13180);
			10909: out = 24'(7708);
			10910: out = 24'(-32540);
			10911: out = 24'(-33668);
			10912: out = 24'(6936);
			10913: out = 24'(32444);
			10914: out = 24'(-1576);
			10915: out = 24'(-12576);
			10916: out = 24'(7224);
			10917: out = 24'(26808);
			10918: out = 24'(11744);
			10919: out = 24'(-23792);
			10920: out = 24'(-30140);
			10921: out = 24'(-26688);
			10922: out = 24'(-37372);
			10923: out = 24'(-41884);
			10924: out = 24'(1820);
			10925: out = 24'(38696);
			10926: out = 24'(29720);
			10927: out = 24'(3768);
			10928: out = 24'(9220);
			10929: out = 24'(17012);
			10930: out = 24'(6148);
			10931: out = 24'(12);
			10932: out = 24'(-3204);
			10933: out = 24'(2156);
			10934: out = 24'(7552);
			10935: out = 24'(13656);
			10936: out = 24'(-21696);
			10937: out = 24'(-41940);
			10938: out = 24'(-33216);
			10939: out = 24'(-10836);
			10940: out = 24'(12008);
			10941: out = 24'(-20568);
			10942: out = 24'(-32452);
			10943: out = 24'(20976);
			10944: out = 24'(51204);
			10945: out = 24'(44056);
			10946: out = 24'(260);
			10947: out = 24'(-11684);
			10948: out = 24'(5932);
			10949: out = 24'(28960);
			10950: out = 24'(-5876);
			10951: out = 24'(-34604);
			10952: out = 24'(-6100);
			10953: out = 24'(18688);
			10954: out = 24'(8860);
			10955: out = 24'(8144);
			10956: out = 24'(35840);
			10957: out = 24'(37072);
			10958: out = 24'(-5996);
			10959: out = 24'(-34052);
			10960: out = 24'(-18096);
			10961: out = 24'(-30176);
			10962: out = 24'(-41692);
			10963: out = 24'(-11944);
			10964: out = 24'(48716);
			10965: out = 24'(31452);
			10966: out = 24'(30188);
			10967: out = 24'(20972);
			10968: out = 24'(6964);
			10969: out = 24'(-65208);
			10970: out = 24'(-47620);
			10971: out = 24'(-23112);
			10972: out = 24'(17488);
			10973: out = 24'(41648);
			10974: out = 24'(31040);
			10975: out = 24'(14508);
			10976: out = 24'(20456);
			10977: out = 24'(16548);
			10978: out = 24'(-22476);
			10979: out = 24'(-60392);
			10980: out = 24'(-39832);
			10981: out = 24'(1836);
			10982: out = 24'(1204);
			10983: out = 24'(-30984);
			10984: out = 24'(-416);
			10985: out = 24'(55016);
			10986: out = 24'(20984);
			10987: out = 24'(7784);
			10988: out = 24'(-9160);
			10989: out = 24'(-22788);
			10990: out = 24'(-60468);
			10991: out = 24'(3272);
			10992: out = 24'(29276);
			10993: out = 24'(8820);
			10994: out = 24'(-26104);
			10995: out = 24'(27892);
			10996: out = 24'(37184);
			10997: out = 24'(-9400);
			10998: out = 24'(-70040);
			10999: out = 24'(-43988);
			11000: out = 24'(1424);
			11001: out = 24'(16360);
			11002: out = 24'(-6180);
			11003: out = 24'(-25744);
			11004: out = 24'(12704);
			11005: out = 24'(36456);
			11006: out = 24'(20896);
			11007: out = 24'(-10560);
			11008: out = 24'(6668);
			11009: out = 24'(14224);
			11010: out = 24'(-2036);
			11011: out = 24'(-42548);
			11012: out = 24'(9112);
			11013: out = 24'(-13080);
			11014: out = 24'(-24332);
			11015: out = 24'(9312);
			11016: out = 24'(51088);
			11017: out = 24'(20360);
			11018: out = 24'(-12356);
			11019: out = 24'(-16868);
			11020: out = 24'(-17200);
			11021: out = 24'(-5444);
			11022: out = 24'(26636);
			11023: out = 24'(45476);
			11024: out = 24'(1608);
			11025: out = 24'(-3928);
			11026: out = 24'(1328);
			11027: out = 24'(7532);
			11028: out = 24'(-22452);
			11029: out = 24'(-31216);
			11030: out = 24'(-18636);
			11031: out = 24'(10768);
			11032: out = 24'(-2580);
			11033: out = 24'(-8544);
			11034: out = 24'(-15336);
			11035: out = 24'(31304);
			11036: out = 24'(55820);
			11037: out = 24'(72160);
			11038: out = 24'(-32772);
			11039: out = 24'(-43904);
			11040: out = 24'(6284);
			11041: out = 24'(10576);
			11042: out = 24'(-20996);
			11043: out = 24'(11700);
			11044: out = 24'(33580);
			11045: out = 24'(-32612);
			11046: out = 24'(-29472);
			11047: out = 24'(33712);
			11048: out = 24'(57072);
			11049: out = 24'(-19072);
			11050: out = 24'(-47532);
			11051: out = 24'(-29996);
			11052: out = 24'(-2800);
			11053: out = 24'(-20704);
			11054: out = 24'(2592);
			11055: out = 24'(3500);
			11056: out = 24'(3132);
			11057: out = 24'(9632);
			11058: out = 24'(51204);
			11059: out = 24'(51552);
			11060: out = 24'(-4628);
			11061: out = 24'(-56488);
			11062: out = 24'(-8708);
			11063: out = 24'(1956);
			11064: out = 24'(-19484);
			11065: out = 24'(-52144);
			11066: out = 24'(-19372);
			11067: out = 24'(15668);
			11068: out = 24'(35300);
			11069: out = 24'(12808);
			11070: out = 24'(5764);
			11071: out = 24'(29092);
			11072: out = 24'(36288);
			11073: out = 24'(-5332);
			11074: out = 24'(-38872);
			11075: out = 24'(-4636);
			11076: out = 24'(40168);
			11077: out = 24'(22844);
			11078: out = 24'(-35996);
			11079: out = 24'(-63112);
			11080: out = 24'(-34436);
			11081: out = 24'(20500);
			11082: out = 24'(50396);
			11083: out = 24'(45912);
			11084: out = 24'(39020);
			11085: out = 24'(4712);
			11086: out = 24'(-15568);
			11087: out = 24'(-1656);
			11088: out = 24'(-19720);
			11089: out = 24'(-26620);
			11090: out = 24'(-31332);
			11091: out = 24'(-21116);
			11092: out = 24'(-13884);
			11093: out = 24'(18572);
			11094: out = 24'(50272);
			11095: out = 24'(56640);
			11096: out = 24'(-3640);
			11097: out = 24'(-27596);
			11098: out = 24'(-30816);
			11099: out = 24'(5592);
			11100: out = 24'(2764);
			11101: out = 24'(41456);
			11102: out = 24'(-23828);
			11103: out = 24'(-50492);
			11104: out = 24'(10252);
			11105: out = 24'(38384);
			11106: out = 24'(-11536);
			11107: out = 24'(-36604);
			11108: out = 24'(11648);
			11109: out = 24'(12348);
			11110: out = 24'(-10760);
			11111: out = 24'(-16684);
			11112: out = 24'(15512);
			11113: out = 24'(-5472);
			11114: out = 24'(-7948);
			11115: out = 24'(-7872);
			11116: out = 24'(8984);
			11117: out = 24'(-5356);
			11118: out = 24'(-2964);
			11119: out = 24'(-7020);
			11120: out = 24'(7980);
			11121: out = 24'(13428);
			11122: out = 24'(27968);
			11123: out = 24'(628);
			11124: out = 24'(-18856);
			11125: out = 24'(-25828);
			11126: out = 24'(-11424);
			11127: out = 24'(-42260);
			11128: out = 24'(-43404);
			11129: out = 24'(-604);
			11130: out = 24'(23892);
			11131: out = 24'(29392);
			11132: out = 24'(24732);
			11133: out = 24'(32520);
			11134: out = 24'(55788);
			11135: out = 24'(11392);
			11136: out = 24'(-24272);
			11137: out = 24'(-57724);
			11138: out = 24'(-91664);
			11139: out = 24'(-64476);
			11140: out = 24'(-1212);
			11141: out = 24'(52128);
			11142: out = 24'(61848);
			11143: out = 24'(6480);
			11144: out = 24'(-3748);
			11145: out = 24'(3260);
			11146: out = 24'(3156);
			11147: out = 24'(-22720);
			11148: out = 24'(-22960);
			11149: out = 24'(-24708);
			11150: out = 24'(-16876);
			11151: out = 24'(328);
			11152: out = 24'(46692);
			11153: out = 24'(39392);
			11154: out = 24'(3032);
			11155: out = 24'(-29640);
			11156: out = 24'(-2496);
			11157: out = 24'(-18392);
			11158: out = 24'(-30148);
			11159: out = 24'(6548);
			11160: out = 24'(33056);
			11161: out = 24'(17048);
			11162: out = 24'(-6352);
			11163: out = 24'(8432);
			11164: out = 24'(49348);
			11165: out = 24'(20952);
			11166: out = 24'(-25304);
			11167: out = 24'(-32152);
			11168: out = 24'(24492);
			11169: out = 24'(7648);
			11170: out = 24'(7744);
			11171: out = 24'(35732);
			11172: out = 24'(43048);
			11173: out = 24'(6260);
			11174: out = 24'(-28204);
			11175: out = 24'(-22064);
			11176: out = 24'(-1544);
			11177: out = 24'(10844);
			11178: out = 24'(996);
			11179: out = 24'(-1156);
			11180: out = 24'(-2076);
			11181: out = 24'(6200);
			11182: out = 24'(22972);
			11183: out = 24'(53848);
			11184: out = 24'(37880);
			11185: out = 24'(-22744);
			11186: out = 24'(-94136);
			11187: out = 24'(-56628);
			11188: out = 24'(20488);
			11189: out = 24'(12640);
			11190: out = 24'(-51164);
			11191: out = 24'(-34700);
			11192: out = 24'(35748);
			11193: out = 24'(32444);
			11194: out = 24'(15048);
			11195: out = 24'(-3496);
			11196: out = 24'(-372);
			11197: out = 24'(-19176);
			11198: out = 24'(-35772);
			11199: out = 24'(-47412);
			11200: out = 24'(-22176);
			11201: out = 24'(6732);
			11202: out = 24'(-21736);
			11203: out = 24'(5184);
			11204: out = 24'(26348);
			11205: out = 24'(22512);
			11206: out = 24'(1280);
			11207: out = 24'(908);
			11208: out = 24'(-13752);
			11209: out = 24'(-31296);
			11210: out = 24'(-19184);
			11211: out = 24'(140);
			11212: out = 24'(27888);
			11213: out = 24'(30240);
			11214: out = 24'(-3644);
			11215: out = 24'(-6296);
			11216: out = 24'(-26064);
			11217: out = 24'(-17924);
			11218: out = 24'(3840);
			11219: out = 24'(13536);
			11220: out = 24'(-8168);
			11221: out = 24'(-11892);
			11222: out = 24'(6252);
			11223: out = 24'(28276);
			11224: out = 24'(18140);
			11225: out = 24'(27548);
			11226: out = 24'(29792);
			11227: out = 24'(-316);
			11228: out = 24'(-16588);
			11229: out = 24'(-8252);
			11230: out = 24'(-7792);
			11231: out = 24'(-29000);
			11232: out = 24'(-22344);
			11233: out = 24'(24212);
			11234: out = 24'(38572);
			11235: out = 24'(-3312);
			11236: out = 24'(-47756);
			11237: out = 24'(-5448);
			11238: out = 24'(42712);
			11239: out = 24'(25400);
			11240: out = 24'(5952);
			11241: out = 24'(-33572);
			11242: out = 24'(-41364);
			11243: out = 24'(-24768);
			11244: out = 24'(24584);
			11245: out = 24'(40080);
			11246: out = 24'(40528);
			11247: out = 24'(10928);
			11248: out = 24'(-17640);
			11249: out = 24'(-57996);
			11250: out = 24'(-41132);
			11251: out = 24'(-14688);
			11252: out = 24'(-692);
			11253: out = 24'(32744);
			11254: out = 24'(35964);
			11255: out = 24'(6180);
			11256: out = 24'(-24260);
			11257: out = 24'(-24656);
			11258: out = 24'(15376);
			11259: out = 24'(21128);
			11260: out = 24'(8856);
			11261: out = 24'(35824);
			11262: out = 24'(23764);
			11263: out = 24'(-23220);
			11264: out = 24'(-57420);
			11265: out = 24'(5760);
			11266: out = 24'(10492);
			11267: out = 24'(18532);
			11268: out = 24'(3848);
			11269: out = 24'(6092);
			11270: out = 24'(27780);
			11271: out = 24'(42520);
			11272: out = 24'(7520);
			11273: out = 24'(-40140);
			11274: out = 24'(-44012);
			11275: out = 24'(1740);
			11276: out = 24'(24952);
			11277: out = 24'(8892);
			11278: out = 24'(-10844);
			11279: out = 24'(-4572);
			11280: out = 24'(608);
			11281: out = 24'(-292);
			11282: out = 24'(11504);
			11283: out = 24'(6096);
			11284: out = 24'(1632);
			11285: out = 24'(5612);
			11286: out = 24'(26792);
			11287: out = 24'(15556);
			11288: out = 24'(8392);
			11289: out = 24'(192);
			11290: out = 24'(-3392);
			11291: out = 24'(-40108);
			11292: out = 24'(-17344);
			11293: out = 24'(13408);
			11294: out = 24'(13812);
			11295: out = 24'(-20552);
			11296: out = 24'(-28840);
			11297: out = 24'(3708);
			11298: out = 24'(39856);
			11299: out = 24'(21620);
			11300: out = 24'(7972);
			11301: out = 24'(-16280);
			11302: out = 24'(-29332);
			11303: out = 24'(-50088);
			11304: out = 24'(-15064);
			11305: out = 24'(-16080);
			11306: out = 24'(-6064);
			11307: out = 24'(18264);
			11308: out = 24'(28780);
			11309: out = 24'(-10520);
			11310: out = 24'(-15408);
			11311: out = 24'(32476);
			11312: out = 24'(2572);
			11313: out = 24'(4096);
			11314: out = 24'(-3988);
			11315: out = 24'(-4420);
			11316: out = 24'(-49816);
			11317: out = 24'(-17724);
			11318: out = 24'(-11260);
			11319: out = 24'(-3160);
			11320: out = 24'(17700);
			11321: out = 24'(44084);
			11322: out = 24'(22356);
			11323: out = 24'(-9324);
			11324: out = 24'(-22328);
			11325: out = 24'(-472);
			11326: out = 24'(-29028);
			11327: out = 24'(-62436);
			11328: out = 24'(-46860);
			11329: out = 24'(30476);
			11330: out = 24'(48604);
			11331: out = 24'(46728);
			11332: out = 24'(51560);
			11333: out = 24'(46804);
			11334: out = 24'(7428);
			11335: out = 24'(-46784);
			11336: out = 24'(-65712);
			11337: out = 24'(2548);
			11338: out = 24'(20256);
			11339: out = 24'(27636);
			11340: out = 24'(1920);
			11341: out = 24'(-22012);
			11342: out = 24'(-99636);
			11343: out = 24'(-29608);
			11344: out = 24'(71428);
			11345: out = 24'(69936);
			11346: out = 24'(-35268);
			11347: out = 24'(-32740);
			11348: out = 24'(38668);
			11349: out = 24'(51104);
			11350: out = 24'(-42908);
			11351: out = 24'(-23624);
			11352: out = 24'(48492);
			11353: out = 24'(56656);
			11354: out = 24'(-8944);
			11355: out = 24'(-83924);
			11356: out = 24'(-71732);
			11357: out = 24'(2980);
			11358: out = 24'(44468);
			11359: out = 24'(40296);
			11360: out = 24'(30148);
			11361: out = 24'(21684);
			11362: out = 24'(5396);
			11363: out = 24'(-70208);
			11364: out = 24'(-47240);
			11365: out = 24'(14440);
			11366: out = 24'(16552);
			11367: out = 24'(-36376);
			11368: out = 24'(-51948);
			11369: out = 24'(-3200);
			11370: out = 24'(37924);
			11371: out = 24'(8628);
			11372: out = 24'(28396);
			11373: out = 24'(46672);
			11374: out = 24'(29712);
			11375: out = 24'(-23292);
			11376: out = 24'(-31440);
			11377: out = 24'(-26756);
			11378: out = 24'(-40940);
			11379: out = 24'(-58424);
			11380: out = 24'(28640);
			11381: out = 24'(72776);
			11382: out = 24'(32532);
			11383: out = 24'(-24328);
			11384: out = 24'(36600);
			11385: out = 24'(63880);
			11386: out = 24'(2340);
			11387: out = 24'(-103612);
			11388: out = 24'(-111912);
			11389: out = 24'(-44580);
			11390: out = 24'(17012);
			11391: out = 24'(23568);
			11392: out = 24'(30316);
			11393: out = 24'(12788);
			11394: out = 24'(-6360);
			11395: out = 24'(-2576);
			11396: out = 24'(50976);
			11397: out = 24'(45172);
			11398: out = 24'(15980);
			11399: out = 24'(-29168);
			11400: out = 24'(-33612);
			11401: out = 24'(3032);
			11402: out = 24'(19648);
			11403: out = 24'(-10776);
			11404: out = 24'(-34604);
			11405: out = 24'(13752);
			11406: out = 24'(26220);
			11407: out = 24'(-1000);
			11408: out = 24'(-21992);
			11409: out = 24'(39340);
			11410: out = 24'(28336);
			11411: out = 24'(14780);
			11412: out = 24'(-3476);
			11413: out = 24'(6016);
			11414: out = 24'(-42804);
			11415: out = 24'(-39604);
			11416: out = 24'(-19604);
			11417: out = 24'(5628);
			11418: out = 24'(-2396);
			11419: out = 24'(33856);
			11420: out = 24'(33540);
			11421: out = 24'(-864);
			11422: out = 24'(-38236);
			11423: out = 24'(18520);
			11424: out = 24'(46684);
			11425: out = 24'(8012);
			11426: out = 24'(-48800);
			11427: out = 24'(-43044);
			11428: out = 24'(-28884);
			11429: out = 24'(-23036);
			11430: out = 24'(6904);
			11431: out = 24'(55512);
			11432: out = 24'(51888);
			11433: out = 24'(3688);
			11434: out = 24'(-27620);
			11435: out = 24'(-53716);
			11436: out = 24'(-21736);
			11437: out = 24'(20412);
			11438: out = 24'(43164);
			11439: out = 24'(2908);
			11440: out = 24'(-28996);
			11441: out = 24'(-54436);
			11442: out = 24'(-31100);
			11443: out = 24'(11988);
			11444: out = 24'(46988);
			11445: out = 24'(24556);
			11446: out = 24'(13164);
			11447: out = 24'(33080);
			11448: out = 24'(53904);
			11449: out = 24'(-15972);
			11450: out = 24'(-78672);
			11451: out = 24'(-40416);
			11452: out = 24'(-3864);
			11453: out = 24'(-43232);
			11454: out = 24'(-84408);
			11455: out = 24'(-10668);
			11456: out = 24'(45788);
			11457: out = 24'(77700);
			11458: out = 24'(42048);
			11459: out = 24'(16540);
			11460: out = 24'(-14288);
			11461: out = 24'(35720);
			11462: out = 24'(23164);
			11463: out = 24'(-28240);
			11464: out = 24'(-84120);
			11465: out = 24'(-32692);
			11466: out = 24'(4772);
			11467: out = 24'(36344);
			11468: out = 24'(75616);
			11469: out = 24'(56308);
			11470: out = 24'(-6608);
			11471: out = 24'(-57384);
			11472: out = 24'(-46740);
			11473: out = 24'(-21292);
			11474: out = 24'(-4);
			11475: out = 24'(13536);
			11476: out = 24'(16004);
			11477: out = 24'(16352);
			11478: out = 24'(-27644);
			11479: out = 24'(-10668);
			11480: out = 24'(47420);
			11481: out = 24'(40404);
			11482: out = 24'(-16456);
			11483: out = 24'(-41916);
			11484: out = 24'(-13348);
			11485: out = 24'(-27144);
			11486: out = 24'(-1248);
			11487: out = 24'(-4952);
			11488: out = 24'(15612);
			11489: out = 24'(23468);
			11490: out = 24'(34668);
			11491: out = 24'(-28336);
			11492: out = 24'(-54504);
			11493: out = 24'(-20600);
			11494: out = 24'(1972);
			11495: out = 24'(8428);
			11496: out = 24'(40092);
			11497: out = 24'(75456);
			11498: out = 24'(59728);
			11499: out = 24'(7636);
			11500: out = 24'(-28100);
			11501: out = 24'(-38000);
			11502: out = 24'(-45668);
			11503: out = 24'(-53696);
			11504: out = 24'(-20032);
			11505: out = 24'(14096);
			11506: out = 24'(7700);
			11507: out = 24'(16324);
			11508: out = 24'(51128);
			11509: out = 24'(64344);
			11510: out = 24'(18064);
			11511: out = 24'(-35724);
			11512: out = 24'(-53192);
			11513: out = 24'(-42064);
			11514: out = 24'(-45648);
			11515: out = 24'(-11944);
			11516: out = 24'(1484);
			11517: out = 24'(39936);
			11518: out = 24'(57076);
			11519: out = 24'(45480);
			11520: out = 24'(-628);
			11521: out = 24'(-13620);
			11522: out = 24'(-14752);
			11523: out = 24'(-27732);
			11524: out = 24'(-24996);
			11525: out = 24'(2168);
			11526: out = 24'(18324);
			11527: out = 24'(2988);
			11528: out = 24'(-12912);
			11529: out = 24'(-2632);
			11530: out = 24'(14068);
			11531: out = 24'(17552);
			11532: out = 24'(17044);
			11533: out = 24'(15620);
			11534: out = 24'(-7364);
			11535: out = 24'(-30544);
			11536: out = 24'(18640);
			11537: out = 24'(5124);
			11538: out = 24'(-2444);
			11539: out = 24'(680);
			11540: out = 24'(27416);
			11541: out = 24'(-9520);
			11542: out = 24'(-8820);
			11543: out = 24'(17988);
			11544: out = 24'(30876);
			11545: out = 24'(-28012);
			11546: out = 24'(-26044);
			11547: out = 24'(32388);
			11548: out = 24'(52308);
			11549: out = 24'(-37548);
			11550: out = 24'(-75532);
			11551: out = 24'(-13936);
			11552: out = 24'(52788);
			11553: out = 24'(2988);
			11554: out = 24'(-20792);
			11555: out = 24'(7716);
			11556: out = 24'(50000);
			11557: out = 24'(39520);
			11558: out = 24'(-57808);
			11559: out = 24'(-79932);
			11560: out = 24'(-4660);
			11561: out = 24'(56172);
			11562: out = 24'(56820);
			11563: out = 24'(21712);
			11564: out = 24'(-20320);
			11565: out = 24'(-45764);
			11566: out = 24'(-39320);
			11567: out = 24'(22128);
			11568: out = 24'(52732);
			11569: out = 24'(19880);
			11570: out = 24'(-52132);
			11571: out = 24'(-48068);
			11572: out = 24'(-15432);
			11573: out = 24'(2256);
			11574: out = 24'(2096);
			11575: out = 24'(64140);
			11576: out = 24'(66712);
			11577: out = 24'(-588);
			11578: out = 24'(-95416);
			11579: out = 24'(-71716);
			11580: out = 24'(-25692);
			11581: out = 24'(11124);
			11582: out = 24'(41876);
			11583: out = 24'(63036);
			11584: out = 24'(39060);
			11585: out = 24'(-7872);
			11586: out = 24'(-32468);
			11587: out = 24'(-15212);
			11588: out = 24'(-18684);
			11589: out = 24'(-42868);
			11590: out = 24'(-42352);
			11591: out = 24'(40);
			11592: out = 24'(39876);
			11593: out = 24'(36652);
			11594: out = 24'(17248);
			11595: out = 24'(5480);
			11596: out = 24'(16416);
			11597: out = 24'(7092);
			11598: out = 24'(-1912);
			11599: out = 24'(-9048);
			11600: out = 24'(-11036);
			11601: out = 24'(-50948);
			11602: out = 24'(-39536);
			11603: out = 24'(38456);
			11604: out = 24'(45592);
			11605: out = 24'(27560);
			11606: out = 24'(20);
			11607: out = 24'(-9116);
			11608: out = 24'(-46156);
			11609: out = 24'(-12860);
			11610: out = 24'(10448);
			11611: out = 24'(13336);
			11612: out = 24'(30312);
			11613: out = 24'(22208);
			11614: out = 24'(44776);
			11615: out = 24'(37776);
			11616: out = 24'(-10624);
			11617: out = 24'(-71972);
			11618: out = 24'(-39412);
			11619: out = 24'(10936);
			11620: out = 24'(-6848);
			11621: out = 24'(-10640);
			11622: out = 24'(-2908);
			11623: out = 24'(27804);
			11624: out = 24'(29532);
			11625: out = 24'(3952);
			11626: out = 24'(3112);
			11627: out = 24'(27948);
			11628: out = 24'(31188);
			11629: out = 24'(-6236);
			11630: out = 24'(-26916);
			11631: out = 24'(-16744);
			11632: out = 24'(6316);
			11633: out = 24'(10248);
			11634: out = 24'(32508);
			11635: out = 24'(20332);
			11636: out = 24'(-11592);
			11637: out = 24'(-40640);
			11638: out = 24'(-16556);
			11639: out = 24'(-9608);
			11640: out = 24'(-19308);
			11641: out = 24'(-25332);
			11642: out = 24'(4172);
			11643: out = 24'(4048);
			11644: out = 24'(-4972);
			11645: out = 24'(728);
			11646: out = 24'(24888);
			11647: out = 24'(28068);
			11648: out = 24'(15436);
			11649: out = 24'(-1764);
			11650: out = 24'(-31620);
			11651: out = 24'(-26692);
			11652: out = 24'(-40988);
			11653: out = 24'(-37184);
			11654: out = 24'(-4800);
			11655: out = 24'(60508);
			11656: out = 24'(33852);
			11657: out = 24'(-13336);
			11658: out = 24'(-29864);
			11659: out = 24'(13740);
			11660: out = 24'(23784);
			11661: out = 24'(29664);
			11662: out = 24'(12880);
			11663: out = 24'(-46296);
			11664: out = 24'(-57228);
			11665: out = 24'(-2588);
			11666: out = 24'(34168);
			11667: out = 24'(2384);
			11668: out = 24'(-35508);
			11669: out = 24'(4636);
			11670: out = 24'(47668);
			11671: out = 24'(8292);
			11672: out = 24'(-61968);
			11673: out = 24'(-53476);
			11674: out = 24'(12584);
			11675: out = 24'(35508);
			11676: out = 24'(39380);
			11677: out = 24'(38144);
			11678: out = 24'(28388);
			11679: out = 24'(-13180);
			11680: out = 24'(-53444);
			11681: out = 24'(-30764);
			11682: out = 24'(3308);
			11683: out = 24'(-2808);
			11684: out = 24'(7268);
			11685: out = 24'(-3972);
			11686: out = 24'(20268);
			11687: out = 24'(15940);
			11688: out = 24'(-13208);
			11689: out = 24'(-8008);
			11690: out = 24'(37644);
			11691: out = 24'(34604);
			11692: out = 24'(-30860);
			11693: out = 24'(-78748);
			11694: out = 24'(-37820);
			11695: out = 24'(32704);
			11696: out = 24'(53620);
			11697: out = 24'(58632);
			11698: out = 24'(29148);
			11699: out = 24'(-11840);
			11700: out = 24'(-55376);
			11701: out = 24'(-63680);
			11702: out = 24'(-53560);
			11703: out = 24'(-22592);
			11704: out = 24'(25260);
			11705: out = 24'(78760);
			11706: out = 24'(31388);
			11707: out = 24'(-24748);
			11708: out = 24'(-46340);
			11709: out = 24'(2324);
			11710: out = 24'(12044);
			11711: out = 24'(27768);
			11712: out = 24'(19176);
			11713: out = 24'(5788);
			11714: out = 24'(680);
			11715: out = 24'(-12888);
			11716: out = 24'(-29632);
			11717: out = 24'(-17756);
			11718: out = 24'(18808);
			11719: out = 24'(60048);
			11720: out = 24'(41172);
			11721: out = 24'(-9872);
			11722: out = 24'(-37904);
			11723: out = 24'(-39204);
			11724: out = 24'(-17144);
			11725: out = 24'(17028);
			11726: out = 24'(52248);
			11727: out = 24'(7404);
			11728: out = 24'(-23300);
			11729: out = 24'(-34588);
			11730: out = 24'(-16836);
			11731: out = 24'(7976);
			11732: out = 24'(24820);
			11733: out = 24'(23380);
			11734: out = 24'(14640);
			11735: out = 24'(6056);
			11736: out = 24'(-25032);
			11737: out = 24'(-51968);
			11738: out = 24'(-39024);
			11739: out = 24'(10896);
			11740: out = 24'(11580);
			11741: out = 24'(6484);
			11742: out = 24'(22204);
			11743: out = 24'(31084);
			11744: out = 24'(-2032);
			11745: out = 24'(-52068);
			11746: out = 24'(-43184);
			11747: out = 24'(14468);
			11748: out = 24'(6112);
			11749: out = 24'(-38496);
			11750: out = 24'(-36000);
			11751: out = 24'(27884);
			11752: out = 24'(15948);
			11753: out = 24'(16760);
			11754: out = 24'(23528);
			11755: out = 24'(40364);
			11756: out = 24'(-924);
			11757: out = 24'(-860);
			11758: out = 24'(-5468);
			11759: out = 24'(3800);
			11760: out = 24'(-1972);
			11761: out = 24'(17356);
			11762: out = 24'(9992);
			11763: out = 24'(768);
			11764: out = 24'(-19136);
			11765: out = 24'(3440);
			11766: out = 24'(-18440);
			11767: out = 24'(-19992);
			11768: out = 24'(5260);
			11769: out = 24'(36144);
			11770: out = 24'(11752);
			11771: out = 24'(840);
			11772: out = 24'(5400);
			11773: out = 24'(-2856);
			11774: out = 24'(-6608);
			11775: out = 24'(31584);
			11776: out = 24'(39236);
			11777: out = 24'(-65428);
			11778: out = 24'(-75584);
			11779: out = 24'(-21168);
			11780: out = 24'(33864);
			11781: out = 24'(-4160);
			11782: out = 24'(28940);
			11783: out = 24'(28544);
			11784: out = 24'(26684);
			11785: out = 24'(-6836);
			11786: out = 24'(992);
			11787: out = 24'(-43644);
			11788: out = 24'(-45892);
			11789: out = 24'(3248);
			11790: out = 24'(54276);
			11791: out = 24'(14556);
			11792: out = 24'(-36356);
			11793: out = 24'(-40628);
			11794: out = 24'(12172);
			11795: out = 24'(47084);
			11796: out = 24'(44848);
			11797: out = 24'(11260);
			11798: out = 24'(-22096);
			11799: out = 24'(-71152);
			11800: out = 24'(-52796);
			11801: out = 24'(-3692);
			11802: out = 24'(14888);
			11803: out = 24'(52164);
			11804: out = 24'(72816);
			11805: out = 24'(75068);
			11806: out = 24'(27860);
			11807: out = 24'(-1688);
			11808: out = 24'(-82360);
			11809: out = 24'(-95968);
			11810: out = 24'(-43788);
			11811: out = 24'(22048);
			11812: out = 24'(24564);
			11813: out = 24'(45620);
			11814: out = 24'(46648);
			11815: out = 24'(824);
			11816: out = 24'(-52268);
			11817: out = 24'(-6644);
			11818: out = 24'(65244);
			11819: out = 24'(43284);
			11820: out = 24'(-42672);
			11821: out = 24'(-81480);
			11822: out = 24'(-34536);
			11823: out = 24'(22452);
			11824: out = 24'(56588);
			11825: out = 24'(46640);
			11826: out = 24'(20608);
			11827: out = 24'(-23448);
			11828: out = 24'(-48280);
			11829: out = 24'(-77024);
			11830: out = 24'(-62376);
			11831: out = 24'(-16280);
			11832: out = 24'(38952);
			11833: out = 24'(61780);
			11834: out = 24'(46376);
			11835: out = 24'(-27860);
			11836: out = 24'(-110680);
			11837: out = 24'(-43092);
			11838: out = 24'(37160);
			11839: out = 24'(18048);
			11840: out = 24'(-49712);
			11841: out = 24'(-33036);
			11842: out = 24'(23436);
			11843: out = 24'(15908);
			11844: out = 24'(-39324);
			11845: out = 24'(-8984);
			11846: out = 24'(41796);
			11847: out = 24'(33756);
			11848: out = 24'(-27608);
			11849: out = 24'(-31344);
			11850: out = 24'(-9456);
			11851: out = 24'(19844);
			11852: out = 24'(29056);
			11853: out = 24'(46532);
			11854: out = 24'(-8624);
			11855: out = 24'(-35736);
			11856: out = 24'(-21616);
			11857: out = 24'(18176);
			11858: out = 24'(-40736);
			11859: out = 24'(-39264);
			11860: out = 24'(21088);
			11861: out = 24'(72036);
			11862: out = 24'(8516);
			11863: out = 24'(-2328);
			11864: out = 24'(30152);
			11865: out = 24'(57960);
			11866: out = 24'(-5492);
			11867: out = 24'(-27072);
			11868: out = 24'(-12504);
			11869: out = 24'(41800);
			11870: out = 24'(58660);
			11871: out = 24'(19088);
			11872: out = 24'(-44528);
			11873: out = 24'(-48356);
			11874: out = 24'(15060);
			11875: out = 24'(3208);
			11876: out = 24'(4);
			11877: out = 24'(11184);
			11878: out = 24'(22780);
			11879: out = 24'(-28544);
			11880: out = 24'(-17864);
			11881: out = 24'(37756);
			11882: out = 24'(80172);
			11883: out = 24'(49556);
			11884: out = 24'(-5032);
			11885: out = 24'(-59128);
			11886: out = 24'(-62616);
			11887: out = 24'(-4624);
			11888: out = 24'(49328);
			11889: out = 24'(59796);
			11890: out = 24'(10848);
			11891: out = 24'(-82316);
			11892: out = 24'(-65124);
			11893: out = 24'(-47436);
			11894: out = 24'(-28688);
			11895: out = 24'(5852);
			11896: out = 24'(55924);
			11897: out = 24'(63772);
			11898: out = 24'(26292);
			11899: out = 24'(-13780);
			11900: out = 24'(-6904);
			11901: out = 24'(-7396);
			11902: out = 24'(-24404);
			11903: out = 24'(-21704);
			11904: out = 24'(39724);
			11905: out = 24'(25260);
			11906: out = 24'(-16292);
			11907: out = 24'(-49164);
			11908: out = 24'(-29680);
			11909: out = 24'(-1684);
			11910: out = 24'(16500);
			11911: out = 24'(17408);
			11912: out = 24'(17080);
			11913: out = 24'(8104);
			11914: out = 24'(-4192);
			11915: out = 24'(-13248);
			11916: out = 24'(-5348);
			11917: out = 24'(25052);
			11918: out = 24'(21436);
			11919: out = 24'(9856);
			11920: out = 24'(-5352);
			11921: out = 24'(-32908);
			11922: out = 24'(-36160);
			11923: out = 24'(-22356);
			11924: out = 24'(-5488);
			11925: out = 24'(3836);
			11926: out = 24'(18432);
			11927: out = 24'(33244);
			11928: out = 24'(32812);
			11929: out = 24'(17532);
			11930: out = 24'(-48956);
			11931: out = 24'(-30324);
			11932: out = 24'(29008);
			11933: out = 24'(54796);
			11934: out = 24'(29148);
			11935: out = 24'(4040);
			11936: out = 24'(-19108);
			11937: out = 24'(-37836);
			11938: out = 24'(-44600);
			11939: out = 24'(-8172);
			11940: out = 24'(18380);
			11941: out = 24'(11512);
			11942: out = 24'(-2396);
			11943: out = 24'(-1360);
			11944: out = 24'(7192);
			11945: out = 24'(3928);
			11946: out = 24'(4320);
			11947: out = 24'(28556);
			11948: out = 24'(42428);
			11949: out = 24'(9436);
			11950: out = 24'(-40252);
			11951: out = 24'(-16496);
			11952: out = 24'(27956);
			11953: out = 24'(38504);
			11954: out = 24'(4608);
			11955: out = 24'(-36080);
			11956: out = 24'(-32408);
			11957: out = 24'(-10760);
			11958: out = 24'(1608);
			11959: out = 24'(6080);
			11960: out = 24'(6808);
			11961: out = 24'(2228);
			11962: out = 24'(2160);
			11963: out = 24'(11440);
			11964: out = 24'(24344);
			11965: out = 24'(11968);
			11966: out = 24'(-5968);
			11967: out = 24'(-13384);
			11968: out = 24'(-27144);
			11969: out = 24'(-18708);
			11970: out = 24'(12912);
			11971: out = 24'(31804);
			11972: out = 24'(4608);
			11973: out = 24'(-9832);
			11974: out = 24'(20064);
			11975: out = 24'(50264);
			11976: out = 24'(18588);
			11977: out = 24'(-44824);
			11978: out = 24'(-65600);
			11979: out = 24'(-24948);
			11980: out = 24'(3568);
			11981: out = 24'(50672);
			11982: out = 24'(52220);
			11983: out = 24'(27112);
			11984: out = 24'(-18008);
			11985: out = 24'(-46704);
			11986: out = 24'(-68964);
			11987: out = 24'(-61688);
			11988: out = 24'(-15872);
			11989: out = 24'(37356);
			11990: out = 24'(70200);
			11991: out = 24'(46676);
			11992: out = 24'(-7292);
			11993: out = 24'(-36760);
			11994: out = 24'(-3188);
			11995: out = 24'(28564);
			11996: out = 24'(14240);
			11997: out = 24'(-13716);
			11998: out = 24'(4004);
			11999: out = 24'(28632);
			12000: out = 24'(-1012);
			12001: out = 24'(-78000);
			12002: out = 24'(-27856);
			12003: out = 24'(18496);
			12004: out = 24'(11668);
			12005: out = 24'(-26260);
			12006: out = 24'(-51912);
			12007: out = 24'(-12712);
			12008: out = 24'(23116);
			12009: out = 24'(16664);
			12010: out = 24'(-7320);
			12011: out = 24'(6660);
			12012: out = 24'(31844);
			12013: out = 24'(46584);
			12014: out = 24'(44720);
			12015: out = 24'(1292);
			12016: out = 24'(-53600);
			12017: out = 24'(-56356);
			12018: out = 24'(16752);
			12019: out = 24'(5260);
			12020: out = 24'(-23020);
			12021: out = 24'(-19600);
			12022: out = 24'(28916);
			12023: out = 24'(8116);
			12024: out = 24'(-23880);
			12025: out = 24'(-27308);
			12026: out = 24'(31068);
			12027: out = 24'(57232);
			12028: out = 24'(36896);
			12029: out = 24'(-36328);
			12030: out = 24'(-80912);
			12031: out = 24'(-19664);
			12032: out = 24'(11888);
			12033: out = 24'(21052);
			12034: out = 24'(40584);
			12035: out = 24'(78432);
			12036: out = 24'(432);
			12037: out = 24'(-88508);
			12038: out = 24'(-104096);
			12039: out = 24'(3888);
			12040: out = 24'(41432);
			12041: out = 24'(53088);
			12042: out = 24'(27712);
			12043: out = 24'(-6348);
			12044: out = 24'(-79348);
			12045: out = 24'(-35732);
			12046: out = 24'(41544);
			12047: out = 24'(64036);
			12048: out = 24'(2116);
			12049: out = 24'(-14464);
			12050: out = 24'(-8816);
			12051: out = 24'(7848);
			12052: out = 24'(-2780);
			12053: out = 24'(3872);
			12054: out = 24'(1904);
			12055: out = 24'(26696);
			12056: out = 24'(45332);
			12057: out = 24'(-4508);
			12058: out = 24'(-73636);
			12059: out = 24'(-54868);
			12060: out = 24'(46088);
			12061: out = 24'(23684);
			12062: out = 24'(-5560);
			12063: out = 24'(3656);
			12064: out = 24'(52832);
			12065: out = 24'(22812);
			12066: out = 24'(-26540);
			12067: out = 24'(-65328);
			12068: out = 24'(-40176);
			12069: out = 24'(-15900);
			12070: out = 24'(16664);
			12071: out = 24'(10608);
			12072: out = 24'(9620);
			12073: out = 24'(9280);
			12074: out = 24'(6776);
			12075: out = 24'(-15752);
			12076: out = 24'(-9924);
			12077: out = 24'(22948);
			12078: out = 24'(13948);
			12079: out = 24'(-3784);
			12080: out = 24'(-8600);
			12081: out = 24'(-1416);
			12082: out = 24'(-19632);
			12083: out = 24'(-6708);
			12084: out = 24'(35616);
			12085: out = 24'(49832);
			12086: out = 24'(-31608);
			12087: out = 24'(-51412);
			12088: out = 24'(-18456);
			12089: out = 24'(28816);
			12090: out = 24'(7132);
			12091: out = 24'(23624);
			12092: out = 24'(6488);
			12093: out = 24'(-17620);
			12094: out = 24'(-51252);
			12095: out = 24'(-4268);
			12096: out = 24'(1024);
			12097: out = 24'(12132);
			12098: out = 24'(39420);
			12099: out = 24'(42272);
			12100: out = 24'(15624);
			12101: out = 24'(-7536);
			12102: out = 24'(3604);
			12103: out = 24'(-6100);
			12104: out = 24'(-6260);
			12105: out = 24'(-44576);
			12106: out = 24'(-50104);
			12107: out = 24'(16684);
			12108: out = 24'(74072);
			12109: out = 24'(43472);
			12110: out = 24'(-21464);
			12111: out = 24'(-47668);
			12112: out = 24'(-9900);
			12113: out = 24'(5908);
			12114: out = 24'(-5004);
			12115: out = 24'(-8036);
			12116: out = 24'(13792);
			12117: out = 24'(7912);
			12118: out = 24'(-104);
			12119: out = 24'(9164);
			12120: out = 24'(23536);
			12121: out = 24'(9680);
			12122: out = 24'(-14280);
			12123: out = 24'(-28792);
			12124: out = 24'(-14180);
			12125: out = 24'(13304);
			12126: out = 24'(50504);
			12127: out = 24'(56608);
			12128: out = 24'(28912);
			12129: out = 24'(-59780);
			12130: out = 24'(-76124);
			12131: out = 24'(-25436);
			12132: out = 24'(25124);
			12133: out = 24'(-17940);
			12134: out = 24'(4692);
			12135: out = 24'(38660);
			12136: out = 24'(30748);
			12137: out = 24'(-56432);
			12138: out = 24'(-39468);
			12139: out = 24'(8468);
			12140: out = 24'(22460);
			12141: out = 24'(0);
			12142: out = 24'(-20040);
			12143: out = 24'(-44532);
			12144: out = 24'(-48020);
			12145: out = 24'(6044);
			12146: out = 24'(29724);
			12147: out = 24'(39004);
			12148: out = 24'(39756);
			12149: out = 24'(60328);
			12150: out = 24'(13644);
			12151: out = 24'(-17504);
			12152: out = 24'(-57136);
			12153: out = 24'(-55304);
			12154: out = 24'(-22120);
			12155: out = 24'(47024);
			12156: out = 24'(43040);
			12157: out = 24'(2952);
			12158: out = 24'(-34344);
			12159: out = 24'(12700);
			12160: out = 24'(11600);
			12161: out = 24'(-10528);
			12162: out = 24'(10188);
			12163: out = 24'(27500);
			12164: out = 24'(-21824);
			12165: out = 24'(-55324);
			12166: out = 24'(23540);
			12167: out = 24'(26644);
			12168: out = 24'(6108);
			12169: out = 24'(-22724);
			12170: out = 24'(-4276);
			12171: out = 24'(20036);
			12172: out = 24'(12800);
			12173: out = 24'(-4920);
			12174: out = 24'(28);
			12175: out = 24'(-18608);
			12176: out = 24'(-8956);
			12177: out = 24'(2152);
			12178: out = 24'(4636);
			12179: out = 24'(-45500);
			12180: out = 24'(-11912);
			12181: out = 24'(25568);
			12182: out = 24'(41904);
			12183: out = 24'(11276);
			12184: out = 24'(10360);
			12185: out = 24'(-10392);
			12186: out = 24'(-15876);
			12187: out = 24'(-14820);
			12188: out = 24'(-33464);
			12189: out = 24'(-38560);
			12190: out = 24'(5444);
			12191: out = 24'(51156);
			12192: out = 24'(3568);
			12193: out = 24'(-11128);
			12194: out = 24'(10768);
			12195: out = 24'(37148);
			12196: out = 24'(-6912);
			12197: out = 24'(-10224);
			12198: out = 24'(1152);
			12199: out = 24'(13288);
			12200: out = 24'(-24972);
			12201: out = 24'(7736);
			12202: out = 24'(11020);
			12203: out = 24'(11000);
			12204: out = 24'(928);
			12205: out = 24'(-5512);
			12206: out = 24'(-42680);
			12207: out = 24'(-41960);
			12208: out = 24'(16048);
			12209: out = 24'(26224);
			12210: out = 24'(15120);
			12211: out = 24'(-9716);
			12212: out = 24'(5776);
			12213: out = 24'(32240);
			12214: out = 24'(30084);
			12215: out = 24'(-17144);
			12216: out = 24'(-26792);
			12217: out = 24'(20720);
			12218: out = 24'(26404);
			12219: out = 24'(-38160);
			12220: out = 24'(-55884);
			12221: out = 24'(49076);
			12222: out = 24'(47540);
			12223: out = 24'(4348);
			12224: out = 24'(-30348);
			12225: out = 24'(6156);
			12226: out = 24'(5476);
			12227: out = 24'(928);
			12228: out = 24'(-28556);
			12229: out = 24'(-41160);
			12230: out = 24'(-2784);
			12231: out = 24'(8340);
			12232: out = 24'(25252);
			12233: out = 24'(45208);
			12234: out = 24'(35308);
			12235: out = 24'(-2868);
			12236: out = 24'(-32212);
			12237: out = 24'(-29280);
			12238: out = 24'(-12884);
			12239: out = 24'(-23992);
			12240: out = 24'(-27560);
			12241: out = 24'(-9976);
			12242: out = 24'(20188);
			12243: out = 24'(32252);
			12244: out = 24'(34956);
			12245: out = 24'(18200);
			12246: out = 24'(-1964);
			12247: out = 24'(-17140);
			12248: out = 24'(-2388);
			12249: out = 24'(3416);
			12250: out = 24'(-1060);
			12251: out = 24'(-392);
			12252: out = 24'(9544);
			12253: out = 24'(-2204);
			12254: out = 24'(-16760);
			12255: out = 24'(-524);
			12256: out = 24'(1592);
			12257: out = 24'(-17920);
			12258: out = 24'(-29876);
			12259: out = 24'(6028);
			12260: out = 24'(20560);
			12261: out = 24'(20036);
			12262: out = 24'(10512);
			12263: out = 24'(27724);
			12264: out = 24'(-2536);
			12265: out = 24'(2756);
			12266: out = 24'(-9764);
			12267: out = 24'(-8968);
			12268: out = 24'(-22744);
			12269: out = 24'(27240);
			12270: out = 24'(1632);
			12271: out = 24'(-52704);
			12272: out = 24'(-43776);
			12273: out = 24'(-768);
			12274: out = 24'(9672);
			12275: out = 24'(504);
			12276: out = 24'(11724);
			12277: out = 24'(8984);
			12278: out = 24'(-9884);
			12279: out = 24'(-1856);
			12280: out = 24'(33008);
			12281: out = 24'(-8392);
			12282: out = 24'(-46416);
			12283: out = 24'(-13776);
			12284: out = 24'(67944);
			12285: out = 24'(44604);
			12286: out = 24'(-7476);
			12287: out = 24'(-41208);
			12288: out = 24'(-14256);
			12289: out = 24'(-16472);
			12290: out = 24'(2124);
			12291: out = 24'(-1244);
			12292: out = 24'(-3292);
			12293: out = 24'(-28588);
			12294: out = 24'(26664);
			12295: out = 24'(42232);
			12296: out = 24'(37156);
			12297: out = 24'(10432);
			12298: out = 24'(14684);
			12299: out = 24'(-30576);
			12300: out = 24'(-51828);
			12301: out = 24'(-18124);
			12302: out = 24'(37364);
			12303: out = 24'(-5672);
			12304: out = 24'(-69460);
			12305: out = 24'(-66464);
			12306: out = 24'(21700);
			12307: out = 24'(60912);
			12308: out = 24'(57556);
			12309: out = 24'(38596);
			12310: out = 24'(2924);
			12311: out = 24'(2528);
			12312: out = 24'(-20932);
			12313: out = 24'(-34168);
			12314: out = 24'(-20012);
			12315: out = 24'(11560);
			12316: out = 24'(11856);
			12317: out = 24'(2248);
			12318: out = 24'(2064);
			12319: out = 24'(32584);
			12320: out = 24'(12432);
			12321: out = 24'(-14768);
			12322: out = 24'(-32276);
			12323: out = 24'(-37568);
			12324: out = 24'(-39756);
			12325: out = 24'(-1392);
			12326: out = 24'(42736);
			12327: out = 24'(35396);
			12328: out = 24'(-2760);
			12329: out = 24'(-26712);
			12330: out = 24'(-9932);
			12331: out = 24'(20340);
			12332: out = 24'(4244);
			12333: out = 24'(-1628);
			12334: out = 24'(1576);
			12335: out = 24'(1820);
			12336: out = 24'(-35596);
			12337: out = 24'(-17952);
			12338: out = 24'(15024);
			12339: out = 24'(25424);
			12340: out = 24'(26248);
			12341: out = 24'(-3140);
			12342: out = 24'(-35800);
			12343: out = 24'(-45524);
			12344: out = 24'(1904);
			12345: out = 24'(33644);
			12346: out = 24'(55144);
			12347: out = 24'(44420);
			12348: out = 24'(6352);
			12349: out = 24'(-51216);
			12350: out = 24'(-67288);
			12351: out = 24'(-23028);
			12352: out = 24'(37716);
			12353: out = 24'(27704);
			12354: out = 24'(-2836);
			12355: out = 24'(-28952);
			12356: out = 24'(-11948);
			12357: out = 24'(24344);
			12358: out = 24'(45844);
			12359: out = 24'(23224);
			12360: out = 24'(-3168);
			12361: out = 24'(-2328);
			12362: out = 24'(-3200);
			12363: out = 24'(-17440);
			12364: out = 24'(-15344);
			12365: out = 24'(7404);
			12366: out = 24'(-35324);
			12367: out = 24'(-64708);
			12368: out = 24'(-7944);
			12369: out = 24'(80308);
			12370: out = 24'(45876);
			12371: out = 24'(-31240);
			12372: out = 24'(-49444);
			12373: out = 24'(11360);
			12374: out = 24'(-15000);
			12375: out = 24'(-26864);
			12376: out = 24'(7444);
			12377: out = 24'(64852);
			12378: out = 24'(22252);
			12379: out = 24'(9040);
			12380: out = 24'(-2484);
			12381: out = 24'(-9676);
			12382: out = 24'(-63668);
			12383: out = 24'(-5100);
			12384: out = 24'(36520);
			12385: out = 24'(26400);
			12386: out = 24'(-36996);
			12387: out = 24'(-47800);
			12388: out = 24'(-30672);
			12389: out = 24'(12932);
			12390: out = 24'(43984);
			12391: out = 24'(9856);
			12392: out = 24'(18408);
			12393: out = 24'(32464);
			12394: out = 24'(25080);
			12395: out = 24'(-54076);
			12396: out = 24'(-11420);
			12397: out = 24'(25712);
			12398: out = 24'(17912);
			12399: out = 24'(-9896);
			12400: out = 24'(-11544);
			12401: out = 24'(-11372);
			12402: out = 24'(-6108);
			12403: out = 24'(7172);
			12404: out = 24'(24440);
			12405: out = 24'(14764);
			12406: out = 24'(380);
			12407: out = 24'(-5240);
			12408: out = 24'(20556);
			12409: out = 24'(-10132);
			12410: out = 24'(-24512);
			12411: out = 24'(9084);
			12412: out = 24'(43188);
			12413: out = 24'(6652);
			12414: out = 24'(-34876);
			12415: out = 24'(-31012);
			12416: out = 24'(1884);
			12417: out = 24'(-25260);
			12418: out = 24'(-29032);
			12419: out = 24'(26180);
			12420: out = 24'(60500);
			12421: out = 24'(40940);
			12422: out = 24'(-24368);
			12423: out = 24'(-42216);
			12424: out = 24'(1856);
			12425: out = 24'(24968);
			12426: out = 24'(-12140);
			12427: out = 24'(-49672);
			12428: out = 24'(-44788);
			12429: out = 24'(1764);
			12430: out = 24'(4756);
			12431: out = 24'(7248);
			12432: out = 24'(21364);
			12433: out = 24'(44076);
			12434: out = 24'(2216);
			12435: out = 24'(-11864);
			12436: out = 24'(-9848);
			12437: out = 24'(-32684);
			12438: out = 24'(-41380);
			12439: out = 24'(4564);
			12440: out = 24'(55308);
			12441: out = 24'(46880);
			12442: out = 24'(23076);
			12443: out = 24'(568);
			12444: out = 24'(-7184);
			12445: out = 24'(900);
			12446: out = 24'(-14896);
			12447: out = 24'(16520);
			12448: out = 24'(6136);
			12449: out = 24'(-43996);
			12450: out = 24'(-91952);
			12451: out = 24'(-5288);
			12452: out = 24'(50184);
			12453: out = 24'(27300);
			12454: out = 24'(30212);
			12455: out = 24'(23856);
			12456: out = 24'(-592);
			12457: out = 24'(-57912);
			12458: out = 24'(-68564);
			12459: out = 24'(-25676);
			12460: out = 24'(31016);
			12461: out = 24'(19004);
			12462: out = 24'(-9524);
			12463: out = 24'(25108);
			12464: out = 24'(59072);
			12465: out = 24'(17748);
			12466: out = 24'(-54596);
			12467: out = 24'(-36480);
			12468: out = 24'(22340);
			12469: out = 24'(42788);
			12470: out = 24'(19104);
			12471: out = 24'(6296);
			12472: out = 24'(6892);
			12473: out = 24'(-20224);
			12474: out = 24'(-59204);
			12475: out = 24'(-54140);
			12476: out = 24'(-10808);
			12477: out = 24'(17380);
			12478: out = 24'(25608);
			12479: out = 24'(28488);
			12480: out = 24'(-7532);
			12481: out = 24'(-20216);
			12482: out = 24'(18600);
			12483: out = 24'(63492);
			12484: out = 24'(46776);
			12485: out = 24'(-12068);
			12486: out = 24'(-27788);
			12487: out = 24'(4332);
			12488: out = 24'(-724);
			12489: out = 24'(-26104);
			12490: out = 24'(-15248);
			12491: out = 24'(20156);
			12492: out = 24'(-2844);
			12493: out = 24'(-7452);
			12494: out = 24'(-6844);
			12495: out = 24'(-9044);
			12496: out = 24'(-50100);
			12497: out = 24'(30988);
			12498: out = 24'(46240);
			12499: out = 24'(9988);
			12500: out = 24'(-39516);
			12501: out = 24'(-14912);
			12502: out = 24'(5892);
			12503: out = 24'(12828);
			12504: out = 24'(20464);
			12505: out = 24'(30448);
			12506: out = 24'(45976);
			12507: out = 24'(4376);
			12508: out = 24'(-55940);
			12509: out = 24'(-56572);
			12510: out = 24'(-13664);
			12511: out = 24'(-992);
			12512: out = 24'(-21876);
			12513: out = 24'(-17136);
			12514: out = 24'(308);
			12515: out = 24'(23336);
			12516: out = 24'(34328);
			12517: out = 24'(31840);
			12518: out = 24'(11432);
			12519: out = 24'(-31544);
			12520: out = 24'(-49964);
			12521: out = 24'(-19576);
			12522: out = 24'(3168);
			12523: out = 24'(-4580);
			12524: out = 24'(-20336);
			12525: out = 24'(-5808);
			12526: out = 24'(19532);
			12527: out = 24'(42860);
			12528: out = 24'(25040);
			12529: out = 24'(-9460);
			12530: out = 24'(-19644);
			12531: out = 24'(-33860);
			12532: out = 24'(-15820);
			12533: out = 24'(10948);
			12534: out = 24'(26332);
			12535: out = 24'(4440);
			12536: out = 24'(1768);
			12537: out = 24'(-6512);
			12538: out = 24'(-28704);
			12539: out = 24'(-20640);
			12540: out = 24'(-5380);
			12541: out = 24'(3884);
			12542: out = 24'(-5576);
			12543: out = 24'(5664);
			12544: out = 24'(6828);
			12545: out = 24'(30376);
			12546: out = 24'(45232);
			12547: out = 24'(43296);
			12548: out = 24'(7960);
			12549: out = 24'(-3636);
			12550: out = 24'(-15700);
			12551: out = 24'(-45600);
			12552: out = 24'(-37384);
			12553: out = 24'(6748);
			12554: out = 24'(50416);
			12555: out = 24'(48484);
			12556: out = 24'(8496);
			12557: out = 24'(-33388);
			12558: out = 24'(-35048);
			12559: out = 24'(13208);
			12560: out = 24'(44608);
			12561: out = 24'(40840);
			12562: out = 24'(-17140);
			12563: out = 24'(-50236);
			12564: out = 24'(14716);
			12565: out = 24'(33768);
			12566: out = 24'(13404);
			12567: out = 24'(-5456);
			12568: out = 24'(15444);
			12569: out = 24'(7108);
			12570: out = 24'(-10016);
			12571: out = 24'(-14096);
			12572: out = 24'(-2148);
			12573: out = 24'(-18360);
			12574: out = 24'(-33036);
			12575: out = 24'(1580);
			12576: out = 24'(50312);
			12577: out = 24'(8300);
			12578: out = 24'(-26520);
			12579: out = 24'(-10080);
			12580: out = 24'(40320);
			12581: out = 24'(20200);
			12582: out = 24'(-1452);
			12583: out = 24'(-17660);
			12584: out = 24'(-14052);
			12585: out = 24'(-37244);
			12586: out = 24'(-6012);
			12587: out = 24'(320);
			12588: out = 24'(-1572);
			12589: out = 24'(60);
			12590: out = 24'(-908);
			12591: out = 24'(15756);
			12592: out = 24'(28704);
			12593: out = 24'(23472);
			12594: out = 24'(-35624);
			12595: out = 24'(-7184);
			12596: out = 24'(30656);
			12597: out = 24'(19416);
			12598: out = 24'(-59864);
			12599: out = 24'(-44348);
			12600: out = 24'(-9316);
			12601: out = 24'(-2928);
			12602: out = 24'(-19936);
			12603: out = 24'(-944);
			12604: out = 24'(22208);
			12605: out = 24'(27692);
			12606: out = 24'(9400);
			12607: out = 24'(25416);
			12608: out = 24'(-7776);
			12609: out = 24'(-45624);
			12610: out = 24'(-35784);
			12611: out = 24'(25328);
			12612: out = 24'(23820);
			12613: out = 24'(-17504);
			12614: out = 24'(-23904);
			12615: out = 24'(13976);
			12616: out = 24'(33440);
			12617: out = 24'(-11268);
			12618: out = 24'(-46384);
			12619: out = 24'(404);
			12620: out = 24'(29280);
			12621: out = 24'(-2428);
			12622: out = 24'(-38048);
			12623: out = 24'(5052);
			12624: out = 24'(-96);
			12625: out = 24'(2328);
			12626: out = 24'(2880);
			12627: out = 24'(16208);
			12628: out = 24'(52188);
			12629: out = 24'(24804);
			12630: out = 24'(-22504);
			12631: out = 24'(-40912);
			12632: out = 24'(2308);
			12633: out = 24'(21160);
			12634: out = 24'(22280);
			12635: out = 24'(828);
			12636: out = 24'(-23896);
			12637: out = 24'(-34592);
			12638: out = 24'(10240);
			12639: out = 24'(41512);
			12640: out = 24'(9044);
			12641: out = 24'(-4520);
			12642: out = 24'(16080);
			12643: out = 24'(29672);
			12644: out = 24'(-5320);
			12645: out = 24'(-19144);
			12646: out = 24'(-8544);
			12647: out = 24'(8296);
			12648: out = 24'(-5516);
			12649: out = 24'(-24344);
			12650: out = 24'(-2892);
			12651: out = 24'(30036);
			12652: out = 24'(30396);
			12653: out = 24'(31840);
			12654: out = 24'(11504);
			12655: out = 24'(10244);
			12656: out = 24'(5008);
			12657: out = 24'(-76);
			12658: out = 24'(-40220);
			12659: out = 24'(-27484);
			12660: out = 24'(7620);
			12661: out = 24'(7772);
			12662: out = 24'(20440);
			12663: out = 24'(5148);
			12664: out = 24'(-24000);
			12665: out = 24'(-55512);
			12666: out = 24'(18604);
			12667: out = 24'(18696);
			12668: out = 24'(-1176);
			12669: out = 24'(-19888);
			12670: out = 24'(-21052);
			12671: out = 24'(-5776);
			12672: out = 24'(26224);
			12673: out = 24'(37840);
			12674: out = 24'(9692);
			12675: out = 24'(-16272);
			12676: out = 24'(-30716);
			12677: out = 24'(-34212);
			12678: out = 24'(-20264);
			12679: out = 24'(-30088);
			12680: out = 24'(-1532);
			12681: out = 24'(19956);
			12682: out = 24'(13672);
			12683: out = 24'(-23252);
			12684: out = 24'(-23912);
			12685: out = 24'(-29036);
			12686: out = 24'(-39144);
			12687: out = 24'(1424);
			12688: out = 24'(55380);
			12689: out = 24'(49196);
			12690: out = 24'(-6620);
			12691: out = 24'(-27896);
			12692: out = 24'(-7124);
			12693: out = 24'(15680);
			12694: out = 24'(5848);
			12695: out = 24'(-1824);
			12696: out = 24'(18416);
			12697: out = 24'(18992);
			12698: out = 24'(-17628);
			12699: out = 24'(-45236);
			12700: out = 24'(-1460);
			12701: out = 24'(34936);
			12702: out = 24'(16000);
			12703: out = 24'(-20144);
			12704: out = 24'(1824);
			12705: out = 24'(35384);
			12706: out = 24'(25576);
			12707: out = 24'(-15860);
			12708: out = 24'(1352);
			12709: out = 24'(6632);
			12710: out = 24'(4236);
			12711: out = 24'(-15792);
			12712: out = 24'(-1892);
			12713: out = 24'(-15404);
			12714: out = 24'(22396);
			12715: out = 24'(56380);
			12716: out = 24'(45708);
			12717: out = 24'(7320);
			12718: out = 24'(7820);
			12719: out = 24'(24304);
			12720: out = 24'(-6936);
			12721: out = 24'(-25636);
			12722: out = 24'(-54484);
			12723: out = 24'(-15312);
			12724: out = 24'(36360);
			12725: out = 24'(51872);
			12726: out = 24'(1488);
			12727: out = 24'(-12004);
			12728: out = 24'(-7028);
			12729: out = 24'(-16476);
			12730: out = 24'(-70636);
			12731: out = 24'(-44668);
			12732: out = 24'(23724);
			12733: out = 24'(53540);
			12734: out = 24'(5720);
			12735: out = 24'(25872);
			12736: out = 24'(46940);
			12737: out = 24'(17892);
			12738: out = 24'(-22796);
			12739: out = 24'(16124);
			12740: out = 24'(16448);
			12741: out = 24'(-79084);
			12742: out = 24'(-112700);
			12743: out = 24'(-53740);
			12744: out = 24'(41736);
			12745: out = 24'(48664);
			12746: out = 24'(9460);
			12747: out = 24'(-1620);
			12748: out = 24'(-11792);
			12749: out = 24'(-50372);
			12750: out = 24'(-81528);
			12751: out = 24'(12704);
			12752: out = 24'(76164);
			12753: out = 24'(50120);
			12754: out = 24'(-76);
			12755: out = 24'(-28516);
			12756: out = 24'(-14420);
			12757: out = 24'(-8472);
			12758: out = 24'(-16696);
			12759: out = 24'(-22428);
			12760: out = 24'(-13096);
			12761: out = 24'(-7416);
			12762: out = 24'(5348);
			12763: out = 24'(7704);
			12764: out = 24'(17188);
			12765: out = 24'(-10112);
			12766: out = 24'(-17540);
			12767: out = 24'(16764);
			12768: out = 24'(17272);
			12769: out = 24'(-57904);
			12770: out = 24'(-98184);
			12771: out = 24'(752);
			12772: out = 24'(60444);
			12773: out = 24'(48464);
			12774: out = 24'(5292);
			12775: out = 24'(-5304);
			12776: out = 24'(31544);
			12777: out = 24'(-1684);
			12778: out = 24'(-33252);
			12779: out = 24'(-11916);
			12780: out = 24'(13460);
			12781: out = 24'(17704);
			12782: out = 24'(35116);
			12783: out = 24'(65524);
			12784: out = 24'(35220);
			12785: out = 24'(1192);
			12786: out = 24'(-45988);
			12787: out = 24'(-45584);
			12788: out = 24'(-16);
			12789: out = 24'(18856);
			12790: out = 24'(9680);
			12791: out = 24'(-6372);
			12792: out = 24'(-9244);
			12793: out = 24'(2680);
			12794: out = 24'(19524);
			12795: out = 24'(17952);
			12796: out = 24'(-1420);
			12797: out = 24'(20632);
			12798: out = 24'(7544);
			12799: out = 24'(7960);
			12800: out = 24'(15900);
			12801: out = 24'(23464);
			12802: out = 24'(21736);
			12803: out = 24'(18784);
			12804: out = 24'(-11608);
			12805: out = 24'(-77312);
			12806: out = 24'(-77644);
			12807: out = 24'(-32848);
			12808: out = 24'(10532);
			12809: out = 24'(17276);
			12810: out = 24'(54792);
			12811: out = 24'(41300);
			12812: out = 24'(-2736);
			12813: out = 24'(-45496);
			12814: out = 24'(-20168);
			12815: out = 24'(-2384);
			12816: out = 24'(-9420);
			12817: out = 24'(-27764);
			12818: out = 24'(-10040);
			12819: out = 24'(-1100);
			12820: out = 24'(-372);
			12821: out = 24'(-3516);
			12822: out = 24'(8624);
			12823: out = 24'(35848);
			12824: out = 24'(31264);
			12825: out = 24'(-10604);
			12826: out = 24'(-55260);
			12827: out = 24'(-54028);
			12828: out = 24'(-16300);
			12829: out = 24'(15388);
			12830: out = 24'(16912);
			12831: out = 24'(35640);
			12832: out = 24'(33824);
			12833: out = 24'(25448);
			12834: out = 24'(-14020);
			12835: out = 24'(-59300);
			12836: out = 24'(-100640);
			12837: out = 24'(-52468);
			12838: out = 24'(31880);
			12839: out = 24'(58156);
			12840: out = 24'(24096);
			12841: out = 24'(9004);
			12842: out = 24'(12308);
			12843: out = 24'(7456);
			12844: out = 24'(9376);
			12845: out = 24'(31508);
			12846: out = 24'(37128);
			12847: out = 24'(9932);
			12848: out = 24'(-38300);
			12849: out = 24'(-20324);
			12850: out = 24'(8136);
			12851: out = 24'(3884);
			12852: out = 24'(1156);
			12853: out = 24'(8680);
			12854: out = 24'(-3904);
			12855: out = 24'(-40188);
			12856: out = 24'(-45632);
			12857: out = 24'(-5916);
			12858: out = 24'(31160);
			12859: out = 24'(28160);
			12860: out = 24'(7740);
			12861: out = 24'(9172);
			12862: out = 24'(15192);
			12863: out = 24'(12004);
			12864: out = 24'(-468);
			12865: out = 24'(596);
			12866: out = 24'(-13420);
			12867: out = 24'(-27092);
			12868: out = 24'(-30092);
			12869: out = 24'(-64);
			12870: out = 24'(13736);
			12871: out = 24'(32736);
			12872: out = 24'(38652);
			12873: out = 24'(21712);
			12874: out = 24'(-32880);
			12875: out = 24'(-49940);
			12876: out = 24'(-22776);
			12877: out = 24'(-1004);
			12878: out = 24'(2216);
			12879: out = 24'(13056);
			12880: out = 24'(29336);
			12881: out = 24'(21704);
			12882: out = 24'(6260);
			12883: out = 24'(-11556);
			12884: out = 24'(-15188);
			12885: out = 24'(-11772);
			12886: out = 24'(-25524);
			12887: out = 24'(-11212);
			12888: out = 24'(11460);
			12889: out = 24'(22804);
			12890: out = 24'(33964);
			12891: out = 24'(24816);
			12892: out = 24'(4712);
			12893: out = 24'(-23672);
			12894: out = 24'(-29684);
			12895: out = 24'(328);
			12896: out = 24'(31612);
			12897: out = 24'(7000);
			12898: out = 24'(-59108);
			12899: out = 24'(-30476);
			12900: out = 24'(29428);
			12901: out = 24'(43728);
			12902: out = 24'(13476);
			12903: out = 24'(3584);
			12904: out = 24'(19828);
			12905: out = 24'(4660);
			12906: out = 24'(-45024);
			12907: out = 24'(-55836);
			12908: out = 24'(11832);
			12909: out = 24'(63696);
			12910: out = 24'(45016);
			12911: out = 24'(12904);
			12912: out = 24'(-42132);
			12913: out = 24'(-70180);
			12914: out = 24'(-55908);
			12915: out = 24'(2148);
			12916: out = 24'(2520);
			12917: out = 24'(10556);
			12918: out = 24'(29164);
			12919: out = 24'(28648);
			12920: out = 24'(76);
			12921: out = 24'(-41948);
			12922: out = 24'(-31136);
			12923: out = 24'(15300);
			12924: out = 24'(26400);
			12925: out = 24'(6400);
			12926: out = 24'(5224);
			12927: out = 24'(4320);
			12928: out = 24'(-21476);
			12929: out = 24'(-73824);
			12930: out = 24'(-40696);
			12931: out = 24'(28312);
			12932: out = 24'(19800);
			12933: out = 24'(292);
			12934: out = 24'(24396);
			12935: out = 24'(46928);
			12936: out = 24'(-6380);
			12937: out = 24'(-50276);
			12938: out = 24'(-33684);
			12939: out = 24'(21644);
			12940: out = 24'(21448);
			12941: out = 24'(35400);
			12942: out = 24'(20780);
			12943: out = 24'(16908);
			12944: out = 24'(-6700);
			12945: out = 24'(172);
			12946: out = 24'(-1064);
			12947: out = 24'(39316);
			12948: out = 24'(43192);
			12949: out = 24'(-25076);
			12950: out = 24'(-65880);
			12951: out = 24'(-37612);
			12952: out = 24'(11816);
			12953: out = 24'(15340);
			12954: out = 24'(24068);
			12955: out = 24'(29660);
			12956: out = 24'(18760);
			12957: out = 24'(-6860);
			12958: out = 24'(-8508);
			12959: out = 24'(12256);
			12960: out = 24'(13488);
			12961: out = 24'(-5160);
			12962: out = 24'(-34184);
			12963: out = 24'(-8852);
			12964: out = 24'(-5384);
			12965: out = 24'(-13728);
			12966: out = 24'(-2108);
			12967: out = 24'(32164);
			12968: out = 24'(-2832);
			12969: out = 24'(-42552);
			12970: out = 24'(3828);
			12971: out = 24'(44236);
			12972: out = 24'(9704);
			12973: out = 24'(-45988);
			12974: out = 24'(-29516);
			12975: out = 24'(30612);
			12976: out = 24'(24288);
			12977: out = 24'(-11520);
			12978: out = 24'(-4012);
			12979: out = 24'(14804);
			12980: out = 24'(10056);
			12981: out = 24'(-6468);
			12982: out = 24'(3024);
			12983: out = 24'(-2972);
			12984: out = 24'(17532);
			12985: out = 24'(11800);
			12986: out = 24'(-11156);
			12987: out = 24'(-56556);
			12988: out = 24'(-35168);
			12989: out = 24'(-10832);
			12990: out = 24'(8700);
			12991: out = 24'(20896);
			12992: out = 24'(17416);
			12993: out = 24'(12664);
			12994: out = 24'(7884);
			12995: out = 24'(-1656);
			12996: out = 24'(1460);
			12997: out = 24'(8044);
			12998: out = 24'(23456);
			12999: out = 24'(25956);
			13000: out = 24'(21768);
			13001: out = 24'(-17476);
			13002: out = 24'(-20388);
			13003: out = 24'(2220);
			13004: out = 24'(-13900);
			13005: out = 24'(-14936);
			13006: out = 24'(-10256);
			13007: out = 24'(2944);
			13008: out = 24'(-7912);
			13009: out = 24'(15016);
			13010: out = 24'(6024);
			13011: out = 24'(-1060);
			13012: out = 24'(2764);
			13013: out = 24'(38852);
			13014: out = 24'(5068);
			13015: out = 24'(-41348);
			13016: out = 24'(-39132);
			13017: out = 24'(29448);
			13018: out = 24'(36204);
			13019: out = 24'(-9760);
			13020: out = 24'(-49548);
			13021: out = 24'(-5436);
			13022: out = 24'(-484);
			13023: out = 24'(-872);
			13024: out = 24'(-7800);
			13025: out = 24'(-10216);
			13026: out = 24'(-19888);
			13027: out = 24'(-21640);
			13028: out = 24'(-16216);
			13029: out = 24'(6184);
			13030: out = 24'(36136);
			13031: out = 24'(58188);
			13032: out = 24'(39212);
			13033: out = 24'(-11388);
			13034: out = 24'(-69152);
			13035: out = 24'(-30316);
			13036: out = 24'(37740);
			13037: out = 24'(44420);
			13038: out = 24'(4544);
			13039: out = 24'(-18692);
			13040: out = 24'(4620);
			13041: out = 24'(20976);
			13042: out = 24'(-6844);
			13043: out = 24'(-33688);
			13044: out = 24'(-22352);
			13045: out = 24'(18252);
			13046: out = 24'(50012);
			13047: out = 24'(35024);
			13048: out = 24'(20352);
			13049: out = 24'(-8352);
			13050: out = 24'(-39576);
			13051: out = 24'(-21220);
			13052: out = 24'(-2912);
			13053: out = 24'(-6508);
			13054: out = 24'(-12768);
			13055: out = 24'(12260);
			13056: out = 24'(9332);
			13057: out = 24'(-21440);
			13058: out = 24'(-27208);
			13059: out = 24'(27648);
			13060: out = 24'(53840);
			13061: out = 24'(20604);
			13062: out = 24'(-18844);
			13063: out = 24'(-16284);
			13064: out = 24'(7500);
			13065: out = 24'(-19432);
			13066: out = 24'(-51420);
			13067: out = 24'(-38632);
			13068: out = 24'(14844);
			13069: out = 24'(9628);
			13070: out = 24'(11928);
			13071: out = 24'(37672);
			13072: out = 24'(1900);
			13073: out = 24'(-36128);
			13074: out = 24'(-36788);
			13075: out = 24'(10888);
			13076: out = 24'(11556);
			13077: out = 24'(7572);
			13078: out = 24'(-4288);
			13079: out = 24'(4072);
			13080: out = 24'(2404);
			13081: out = 24'(4240);
			13082: out = 24'(-1480);
			13083: out = 24'(3256);
			13084: out = 24'(-2484);
			13085: out = 24'(-15668);
			13086: out = 24'(-19176);
			13087: out = 24'(840);
			13088: out = 24'(2024);
			13089: out = 24'(-3220);
			13090: out = 24'(-24392);
			13091: out = 24'(11404);
			13092: out = 24'(52428);
			13093: out = 24'(35348);
			13094: out = 24'(-1868);
			13095: out = 24'(-4624);
			13096: out = 24'(360);
			13097: out = 24'(-25564);
			13098: out = 24'(-23644);
			13099: out = 24'(26096);
			13100: out = 24'(48072);
			13101: out = 24'(3536);
			13102: out = 24'(-89544);
			13103: out = 24'(-62160);
			13104: out = 24'(11352);
			13105: out = 24'(-664);
			13106: out = 24'(-1820);
			13107: out = 24'(21028);
			13108: out = 24'(68180);
			13109: out = 24'(55684);
			13110: out = 24'(36972);
			13111: out = 24'(-31188);
			13112: out = 24'(-35020);
			13113: out = 24'(-18540);
			13114: out = 24'(-30904);
			13115: out = 24'(-46460);
			13116: out = 24'(4280);
			13117: out = 24'(59852);
			13118: out = 24'(33936);
			13119: out = 24'(-15568);
			13120: out = 24'(-51244);
			13121: out = 24'(-36648);
			13122: out = 24'(-6404);
			13123: out = 24'(32276);
			13124: out = 24'(36252);
			13125: out = 24'(27316);
			13126: out = 24'(8352);
			13127: out = 24'(22296);
			13128: out = 24'(-14308);
			13129: out = 24'(-22380);
			13130: out = 24'(13224);
			13131: out = 24'(53940);
			13132: out = 24'(28912);
			13133: out = 24'(-16756);
			13134: out = 24'(-56280);
			13135: out = 24'(-80044);
			13136: out = 24'(-17492);
			13137: out = 24'(27484);
			13138: out = 24'(26624);
			13139: out = 24'(-268);
			13140: out = 24'(-8464);
			13141: out = 24'(-13696);
			13142: out = 24'(-14920);
			13143: out = 24'(-3320);
			13144: out = 24'(38136);
			13145: out = 24'(46856);
			13146: out = 24'(21544);
			13147: out = 24'(-19892);
			13148: out = 24'(-41208);
			13149: out = 24'(-59660);
			13150: out = 24'(-49164);
			13151: out = 24'(-12476);
			13152: out = 24'(15396);
			13153: out = 24'(17624);
			13154: out = 24'(1064);
			13155: out = 24'(5616);
			13156: out = 24'(29544);
			13157: out = 24'(12896);
			13158: out = 24'(-20108);
			13159: out = 24'(-16940);
			13160: out = 24'(28960);
			13161: out = 24'(8252);
			13162: out = 24'(-13840);
			13163: out = 24'(-24788);
			13164: out = 24'(-4072);
			13165: out = 24'(-360);
			13166: out = 24'(8080);
			13167: out = 24'(7700);
			13168: out = 24'(17864);
			13169: out = 24'(31916);
			13170: out = 24'(-4252);
			13171: out = 24'(-45404);
			13172: out = 24'(-43060);
			13173: out = 24'(9508);
			13174: out = 24'(38420);
			13175: out = 24'(41308);
			13176: out = 24'(24132);
			13177: out = 24'(-3520);
			13178: out = 24'(-12924);
			13179: out = 24'(-26096);
			13180: out = 24'(-16448);
			13181: out = 24'(11388);
			13182: out = 24'(28096);
			13183: out = 24'(27480);
			13184: out = 24'(19096);
			13185: out = 24'(4468);
			13186: out = 24'(-14520);
			13187: out = 24'(-7636);
			13188: out = 24'(16260);
			13189: out = 24'(12008);
			13190: out = 24'(-38060);
			13191: out = 24'(-43444);
			13192: out = 24'(8220);
			13193: out = 24'(50872);
			13194: out = 24'(17088);
			13195: out = 24'(16728);
			13196: out = 24'(-7176);
			13197: out = 24'(-13880);
			13198: out = 24'(-26900);
			13199: out = 24'(-23336);
			13200: out = 24'(-51336);
			13201: out = 24'(-33048);
			13202: out = 24'(26784);
			13203: out = 24'(65240);
			13204: out = 24'(22764);
			13205: out = 24'(-20564);
			13206: out = 24'(-16480);
			13207: out = 24'(23620);
			13208: out = 24'(19240);
			13209: out = 24'(7508);
			13210: out = 24'(4380);
			13211: out = 24'(584);
			13212: out = 24'(-25684);
			13213: out = 24'(-55088);
			13214: out = 24'(-50172);
			13215: out = 24'(-2648);
			13216: out = 24'(16984);
			13217: out = 24'(28432);
			13218: out = 24'(16024);
			13219: out = 24'(-2344);
			13220: out = 24'(-25448);
			13221: out = 24'(9820);
			13222: out = 24'(35768);
			13223: out = 24'(24964);
			13224: out = 24'(-9636);
			13225: out = 24'(-12656);
			13226: out = 24'(-7712);
			13227: out = 24'(-2248);
			13228: out = 24'(13720);
			13229: out = 24'(28976);
			13230: out = 24'(37344);
			13231: out = 24'(21364);
			13232: out = 24'(-4680);
			13233: out = 24'(-36692);
			13234: out = 24'(-30300);
			13235: out = 24'(-18892);
			13236: out = 24'(-15416);
			13237: out = 24'(-11364);
			13238: out = 24'(21516);
			13239: out = 24'(35620);
			13240: out = 24'(13364);
			13241: out = 24'(-24616);
			13242: out = 24'(-9968);
			13243: out = 24'(20328);
			13244: out = 24'(34028);
			13245: out = 24'(26400);
			13246: out = 24'(6076);
			13247: out = 24'(-34536);
			13248: out = 24'(-75804);
			13249: out = 24'(-65512);
			13250: out = 24'(17256);
			13251: out = 24'(52356);
			13252: out = 24'(15196);
			13253: out = 24'(-12184);
			13254: out = 24'(49032);
			13255: out = 24'(46788);
			13256: out = 24'(-41664);
			13257: out = 24'(-110224);
			13258: out = 24'(-17472);
			13259: out = 24'(44544);
			13260: out = 24'(26308);
			13261: out = 24'(-9144);
			13262: out = 24'(-6184);
			13263: out = 24'(5376);
			13264: out = 24'(-40920);
			13265: out = 24'(-61944);
			13266: out = 24'(18368);
			13267: out = 24'(81064);
			13268: out = 24'(42736);
			13269: out = 24'(-23052);
			13270: out = 24'(-34684);
			13271: out = 24'(-40124);
			13272: out = 24'(-26824);
			13273: out = 24'(5404);
			13274: out = 24'(45000);
			13275: out = 24'(220);
			13276: out = 24'(-20000);
			13277: out = 24'(-33040);
			13278: out = 24'(-6484);
			13279: out = 24'(23824);
			13280: out = 24'(15252);
			13281: out = 24'(-172);
			13282: out = 24'(14752);
			13283: out = 24'(38664);
			13284: out = 24'(-36372);
			13285: out = 24'(-64104);
			13286: out = 24'(-14896);
			13287: out = 24'(45292);
			13288: out = 24'(39092);
			13289: out = 24'(19720);
			13290: out = 24'(25296);
			13291: out = 24'(23188);
			13292: out = 24'(-52976);
			13293: out = 24'(-68284);
			13294: out = 24'(-256);
			13295: out = 24'(68308);
			13296: out = 24'(31048);
			13297: out = 24'(10236);
			13298: out = 24'(-12840);
			13299: out = 24'(-26064);
			13300: out = 24'(-34732);
			13301: out = 24'(-9600);
			13302: out = 24'(38760);
			13303: out = 24'(55812);
			13304: out = 24'(26864);
			13305: out = 24'(-51168);
			13306: out = 24'(-31748);
			13307: out = 24'(15376);
			13308: out = 24'(12068);
			13309: out = 24'(19004);
			13310: out = 24'(4240);
			13311: out = 24'(-7548);
			13312: out = 24'(-19780);
			13313: out = 24'(17268);
			13314: out = 24'(-16548);
			13315: out = 24'(-20244);
			13316: out = 24'(18088);
			13317: out = 24'(58248);
			13318: out = 24'(15960);
			13319: out = 24'(-34432);
			13320: out = 24'(-39536);
			13321: out = 24'(2096);
			13322: out = 24'(2720);
			13323: out = 24'(-10560);
			13324: out = 24'(-7852);
			13325: out = 24'(12344);
			13326: out = 24'(12672);
			13327: out = 24'(-21136);
			13328: out = 24'(-35212);
			13329: out = 24'(-7376);
			13330: out = 24'(9108);
			13331: out = 24'(6624);
			13332: out = 24'(3572);
			13333: out = 24'(17632);
			13334: out = 24'(27944);
			13335: out = 24'(456);
			13336: out = 24'(-16000);
			13337: out = 24'(708);
			13338: out = 24'(23188);
			13339: out = 24'(-2692);
			13340: out = 24'(-15504);
			13341: out = 24'(36);
			13342: out = 24'(14016);
			13343: out = 24'(4776);
			13344: out = 24'(-9548);
			13345: out = 24'(-1612);
			13346: out = 24'(5668);
			13347: out = 24'(-38688);
			13348: out = 24'(-53084);
			13349: out = 24'(-21760);
			13350: out = 24'(25532);
			13351: out = 24'(29680);
			13352: out = 24'(46736);
			13353: out = 24'(60360);
			13354: out = 24'(54872);
			13355: out = 24'(3896);
			13356: out = 24'(-42072);
			13357: out = 24'(-80668);
			13358: out = 24'(-59992);
			13359: out = 24'(19652);
			13360: out = 24'(51636);
			13361: out = 24'(50004);
			13362: out = 24'(6452);
			13363: out = 24'(-34584);
			13364: out = 24'(-36724);
			13365: out = 24'(-800);
			13366: out = 24'(5000);
			13367: out = 24'(-9668);
			13368: out = 24'(10432);
			13369: out = 24'(24148);
			13370: out = 24'(2296);
			13371: out = 24'(-27288);
			13372: out = 24'(11008);
			13373: out = 24'(39864);
			13374: out = 24'(39564);
			13375: out = 24'(-7888);
			13376: out = 24'(-41784);
			13377: out = 24'(-72296);
			13378: out = 24'(-19080);
			13379: out = 24'(32628);
			13380: out = 24'(39884);
			13381: out = 24'(17792);
			13382: out = 24'(21280);
			13383: out = 24'(12368);
			13384: out = 24'(-30692);
			13385: out = 24'(-86392);
			13386: out = 24'(-75360);
			13387: out = 24'(-19980);
			13388: out = 24'(19624);
			13389: out = 24'(31944);
			13390: out = 24'(20400);
			13391: out = 24'(12436);
			13392: out = 24'(5200);
			13393: out = 24'(6448);
			13394: out = 24'(-27956);
			13395: out = 24'(-9772);
			13396: out = 24'(27140);
			13397: out = 24'(38408);
			13398: out = 24'(-12964);
			13399: out = 24'(-20356);
			13400: out = 24'(14152);
			13401: out = 24'(54052);
			13402: out = 24'(35404);
			13403: out = 24'(24896);
			13404: out = 24'(-4248);
			13405: out = 24'(-26056);
			13406: out = 24'(-46752);
			13407: out = 24'(-16672);
			13408: out = 24'(-16424);
			13409: out = 24'(-11688);
			13410: out = 24'(21476);
			13411: out = 24'(65620);
			13412: out = 24'(15440);
			13413: out = 24'(-43580);
			13414: out = 24'(-12108);
			13415: out = 24'(23056);
			13416: out = 24'(21196);
			13417: out = 24'(-16556);
			13418: out = 24'(-10732);
			13419: out = 24'(31320);
			13420: out = 24'(45900);
			13421: out = 24'(-9804);
			13422: out = 24'(-62504);
			13423: out = 24'(-19572);
			13424: out = 24'(160);
			13425: out = 24'(-16636);
			13426: out = 24'(-40336);
			13427: out = 24'(-29380);
			13428: out = 24'(18072);
			13429: out = 24'(35144);
			13430: out = 24'(19948);
			13431: out = 24'(-8348);
			13432: out = 24'(-35192);
			13433: out = 24'(-52256);
			13434: out = 24'(-22348);
			13435: out = 24'(36332);
			13436: out = 24'(45772);
			13437: out = 24'(17436);
			13438: out = 24'(-4432);
			13439: out = 24'(6740);
			13440: out = 24'(22424);
			13441: out = 24'(-9344);
			13442: out = 24'(-37948);
			13443: out = 24'(-29144);
			13444: out = 24'(-5436);
			13445: out = 24'(27696);
			13446: out = 24'(36948);
			13447: out = 24'(26396);
			13448: out = 24'(4444);
			13449: out = 24'(-8144);
			13450: out = 24'(-11764);
			13451: out = 24'(-7728);
			13452: out = 24'(996);
			13453: out = 24'(-1336);
			13454: out = 24'(2752);
			13455: out = 24'(-6076);
			13456: out = 24'(-13212);
			13457: out = 24'(-804);
			13458: out = 24'(37388);
			13459: out = 24'(45196);
			13460: out = 24'(13004);
			13461: out = 24'(-47268);
			13462: out = 24'(-15600);
			13463: out = 24'(9800);
			13464: out = 24'(8492);
			13465: out = 24'(12568);
			13466: out = 24'(34036);
			13467: out = 24'(39632);
			13468: out = 24'(17260);
			13469: out = 24'(-16132);
			13470: out = 24'(-46408);
			13471: out = 24'(-32912);
			13472: out = 24'(15460);
			13473: out = 24'(44360);
			13474: out = 24'(3708);
			13475: out = 24'(-22532);
			13476: out = 24'(-19684);
			13477: out = 24'(5100);
			13478: out = 24'(26844);
			13479: out = 24'(13292);
			13480: out = 24'(11720);
			13481: out = 24'(18792);
			13482: out = 24'(15520);
			13483: out = 24'(-37476);
			13484: out = 24'(-45196);
			13485: out = 24'(-2656);
			13486: out = 24'(30536);
			13487: out = 24'(29572);
			13488: out = 24'(14404);
			13489: out = 24'(4360);
			13490: out = 24'(-3592);
			13491: out = 24'(-6680);
			13492: out = 24'(-25552);
			13493: out = 24'(-40052);
			13494: out = 24'(-31340);
			13495: out = 24'(11364);
			13496: out = 24'(30036);
			13497: out = 24'(16868);
			13498: out = 24'(-15304);
			13499: out = 24'(-20108);
			13500: out = 24'(-56504);
			13501: out = 24'(-46248);
			13502: out = 24'(-3140);
			13503: out = 24'(34448);
			13504: out = 24'(40860);
			13505: out = 24'(27724);
			13506: out = 24'(548);
			13507: out = 24'(-23124);
			13508: out = 24'(-33380);
			13509: out = 24'(-12024);
			13510: out = 24'(9248);
			13511: out = 24'(11460);
			13512: out = 24'(-19632);
			13513: out = 24'(-32576);
			13514: out = 24'(-36216);
			13515: out = 24'(-14864);
			13516: out = 24'(13036);
			13517: out = 24'(22740);
			13518: out = 24'(-14220);
			13519: out = 24'(-38548);
			13520: out = 24'(-6864);
			13521: out = 24'(27264);
			13522: out = 24'(2088);
			13523: out = 24'(-22200);
			13524: out = 24'(20652);
			13525: out = 24'(32616);
			13526: out = 24'(26912);
			13527: out = 24'(1612);
			13528: out = 24'(5904);
			13529: out = 24'(-4100);
			13530: out = 24'(9780);
			13531: out = 24'(-11524);
			13532: out = 24'(-28060);
			13533: out = 24'(-1712);
			13534: out = 24'(8436);
			13535: out = 24'(-1608);
			13536: out = 24'(7620);
			13537: out = 24'(48128);
			13538: out = 24'(32792);
			13539: out = 24'(-9792);
			13540: out = 24'(-28636);
			13541: out = 24'(4200);
			13542: out = 24'(25836);
			13543: out = 24'(-1228);
			13544: out = 24'(-37720);
			13545: out = 24'(-29388);
			13546: out = 24'(5080);
			13547: out = 24'(15352);
			13548: out = 24'(8600);
			13549: out = 24'(13356);
			13550: out = 24'(8908);
			13551: out = 24'(12556);
			13552: out = 24'(6688);
			13553: out = 24'(5840);
			13554: out = 24'(-1136);
			13555: out = 24'(9768);
			13556: out = 24'(3700);
			13557: out = 24'(-1292);
			13558: out = 24'(-3272);
			13559: out = 24'(-21480);
			13560: out = 24'(-28588);
			13561: out = 24'(-8344);
			13562: out = 24'(11196);
			13563: out = 24'(34368);
			13564: out = 24'(15952);
			13565: out = 24'(11192);
			13566: out = 24'(4084);
			13567: out = 24'(-5240);
			13568: out = 24'(-49448);
			13569: out = 24'(-23340);
			13570: out = 24'(30916);
			13571: out = 24'(28584);
			13572: out = 24'(2116);
			13573: out = 24'(31008);
			13574: out = 24'(57488);
			13575: out = 24'(1744);
			13576: out = 24'(-77136);
			13577: out = 24'(-91976);
			13578: out = 24'(-40156);
			13579: out = 24'(-6792);
			13580: out = 24'(45048);
			13581: out = 24'(63292);
			13582: out = 24'(41180);
			13583: out = 24'(-20892);
			13584: out = 24'(-38552);
			13585: out = 24'(-18900);
			13586: out = 24'(15912);
			13587: out = 24'(11784);
			13588: out = 24'(-17320);
			13589: out = 24'(-9844);
			13590: out = 24'(11704);
			13591: out = 24'(10996);
			13592: out = 24'(2348);
			13593: out = 24'(-2048);
			13594: out = 24'(-4912);
			13595: out = 24'(-31228);
			13596: out = 24'(-64424);
			13597: out = 24'(-44708);
			13598: out = 24'(6076);
			13599: out = 24'(44460);
			13600: out = 24'(56204);
			13601: out = 24'(26348);
			13602: out = 24'(9904);
			13603: out = 24'(-12452);
			13604: out = 24'(-18336);
			13605: out = 24'(-14876);
			13606: out = 24'(10484);
			13607: out = 24'(-9364);
			13608: out = 24'(-27636);
			13609: out = 24'(-1856);
			13610: out = 24'(45996);
			13611: out = 24'(1408);
			13612: out = 24'(-64140);
			13613: out = 24'(-35016);
			13614: out = 24'(12808);
			13615: out = 24'(19276);
			13616: out = 24'(-1944);
			13617: out = 24'(19104);
			13618: out = 24'(35360);
			13619: out = 24'(30992);
			13620: out = 24'(-1692);
			13621: out = 24'(-11460);
			13622: out = 24'(1156);
			13623: out = 24'(16640);
			13624: out = 24'(-2176);
			13625: out = 24'(-31932);
			13626: out = 24'(-41600);
			13627: out = 24'(-20668);
			13628: out = 24'(13388);
			13629: out = 24'(41212);
			13630: out = 24'(46604);
			13631: out = 24'(23424);
			13632: out = 24'(-12864);
			13633: out = 24'(-43712);
			13634: out = 24'(-62484);
			13635: out = 24'(-61476);
			13636: out = 24'(-26128);
			13637: out = 24'(45772);
			13638: out = 24'(92296);
			13639: out = 24'(67280);
			13640: out = 24'(-6956);
			13641: out = 24'(-70692);
			13642: out = 24'(-74464);
			13643: out = 24'(-3948);
			13644: out = 24'(-11480);
			13645: out = 24'(-20008);
			13646: out = 24'(4576);
			13647: out = 24'(41760);
			13648: out = 24'(41100);
			13649: out = 24'(21444);
			13650: out = 24'(-2504);
			13651: out = 24'(-14340);
			13652: out = 24'(-13528);
			13653: out = 24'(-1384);
			13654: out = 24'(-10024);
			13655: out = 24'(-28968);
			13656: out = 24'(6480);
			13657: out = 24'(40792);
			13658: out = 24'(39340);
			13659: out = 24'(-2940);
			13660: out = 24'(-61140);
			13661: out = 24'(-36796);
			13662: out = 24'(9072);
			13663: out = 24'(17096);
			13664: out = 24'(5072);
			13665: out = 24'(30592);
			13666: out = 24'(52608);
			13667: out = 24'(35372);
			13668: out = 24'(3888);
			13669: out = 24'(-31216);
			13670: out = 24'(-9528);
			13671: out = 24'(11616);
			13672: out = 24'(-7568);
			13673: out = 24'(-59924);
			13674: out = 24'(-32352);
			13675: out = 24'(27480);
			13676: out = 24'(36300);
			13677: out = 24'(34480);
			13678: out = 24'(-4228);
			13679: out = 24'(-2452);
			13680: out = 24'(11184);
			13681: out = 24'(20120);
			13682: out = 24'(-58188);
			13683: out = 24'(-70328);
			13684: out = 24'(-6700);
			13685: out = 24'(39280);
			13686: out = 24'(34984);
			13687: out = 24'(15764);
			13688: out = 24'(12956);
			13689: out = 24'(15884);
			13690: out = 24'(-25536);
			13691: out = 24'(-54332);
			13692: out = 24'(-52316);
			13693: out = 24'(-11920);
			13694: out = 24'(1632);
			13695: out = 24'(31432);
			13696: out = 24'(22612);
			13697: out = 24'(8072);
			13698: out = 24'(18352);
			13699: out = 24'(31128);
			13700: out = 24'(-72);
			13701: out = 24'(-36600);
			13702: out = 24'(-25748);
			13703: out = 24'(-7668);
			13704: out = 24'(-20980);
			13705: out = 24'(-31392);
			13706: out = 24'(7552);
			13707: out = 24'(44200);
			13708: out = 24'(36572);
			13709: out = 24'(9288);
			13710: out = 24'(-868);
			13711: out = 24'(-14800);
			13712: out = 24'(-37572);
			13713: out = 24'(-40588);
			13714: out = 24'(7340);
			13715: out = 24'(52816);
			13716: out = 24'(75728);
			13717: out = 24'(45200);
			13718: out = 24'(-9068);
			13719: out = 24'(-60020);
			13720: out = 24'(-56716);
			13721: out = 24'(-28468);
			13722: out = 24'(-1756);
			13723: out = 24'(13772);
			13724: out = 24'(37752);
			13725: out = 24'(35936);
			13726: out = 24'(4288);
			13727: out = 24'(-33964);
			13728: out = 24'(-28416);
			13729: out = 24'(-13964);
			13730: out = 24'(-17076);
			13731: out = 24'(-24664);
			13732: out = 24'(37140);
			13733: out = 24'(56492);
			13734: out = 24'(49028);
			13735: out = 24'(9868);
			13736: out = 24'(-16980);
			13737: out = 24'(-27688);
			13738: out = 24'(408);
			13739: out = 24'(12308);
			13740: out = 24'(-388);
			13741: out = 24'(-34140);
			13742: out = 24'(-11700);
			13743: out = 24'(17412);
			13744: out = 24'(13232);
			13745: out = 24'(1860);
			13746: out = 24'(616);
			13747: out = 24'(-4588);
			13748: out = 24'(-14684);
			13749: out = 24'(-7040);
			13750: out = 24'(15128);
			13751: out = 24'(9256);
			13752: out = 24'(-11348);
			13753: out = 24'(1260);
			13754: out = 24'(13640);
			13755: out = 24'(1240);
			13756: out = 24'(-11100);
			13757: out = 24'(26548);
			13758: out = 24'(24272);
			13759: out = 24'(1620);
			13760: out = 24'(-31100);
			13761: out = 24'(-28260);
			13762: out = 24'(-12000);
			13763: out = 24'(12928);
			13764: out = 24'(24956);
			13765: out = 24'(31340);
			13766: out = 24'(1368);
			13767: out = 24'(-16972);
			13768: out = 24'(-37328);
			13769: out = 24'(-42560);
			13770: out = 24'(-49696);
			13771: out = 24'(9640);
			13772: out = 24'(42868);
			13773: out = 24'(35228);
			13774: out = 24'(11856);
			13775: out = 24'(17492);
			13776: out = 24'(12544);
			13777: out = 24'(-16892);
			13778: out = 24'(-60148);
			13779: out = 24'(-28144);
			13780: out = 24'(20);
			13781: out = 24'(23380);
			13782: out = 24'(42144);
			13783: out = 24'(21612);
			13784: out = 24'(19468);
			13785: out = 24'(13888);
			13786: out = 24'(-9800);
			13787: out = 24'(-50348);
			13788: out = 24'(-48768);
			13789: out = 24'(-14556);
			13790: out = 24'(11180);
			13791: out = 24'(31700);
			13792: out = 24'(4656);
			13793: out = 24'(17660);
			13794: out = 24'(29936);
			13795: out = 24'(2088);
			13796: out = 24'(-26684);
			13797: out = 24'(-25600);
			13798: out = 24'(-12212);
			13799: out = 24'(-7204);
			13800: out = 24'(19932);
			13801: out = 24'(44332);
			13802: out = 24'(39604);
			13803: out = 24'(15824);
			13804: out = 24'(-2064);
			13805: out = 24'(5268);
			13806: out = 24'(-25120);
			13807: out = 24'(-65756);
			13808: out = 24'(-5124);
			13809: out = 24'(45908);
			13810: out = 24'(50360);
			13811: out = 24'(7300);
			13812: out = 24'(-18244);
			13813: out = 24'(-9668);
			13814: out = 24'(8724);
			13815: out = 24'(5100);
			13816: out = 24'(-168);
			13817: out = 24'(2144);
			13818: out = 24'(3764);
			13819: out = 24'(-14872);
			13820: out = 24'(-36132);
			13821: out = 24'(1536);
			13822: out = 24'(35008);
			13823: out = 24'(51096);
			13824: out = 24'(23556);
			13825: out = 24'(-43372);
			13826: out = 24'(-63860);
			13827: out = 24'(-21172);
			13828: out = 24'(27792);
			13829: out = 24'(35008);
			13830: out = 24'(6844);
			13831: out = 24'(-292);
			13832: out = 24'(208);
			13833: out = 24'(-13668);
			13834: out = 24'(-40980);
			13835: out = 24'(-21344);
			13836: out = 24'(6480);
			13837: out = 24'(-4068);
			13838: out = 24'(-17024);
			13839: out = 24'(-17612);
			13840: out = 24'(-3576);
			13841: out = 24'(-2000);
			13842: out = 24'(-8152);
			13843: out = 24'(-7484);
			13844: out = 24'(-616);
			13845: out = 24'(4756);
			13846: out = 24'(21080);
			13847: out = 24'(20800);
			13848: out = 24'(7568);
			13849: out = 24'(-19652);
			13850: out = 24'(-27840);
			13851: out = 24'(-8080);
			13852: out = 24'(20820);
			13853: out = 24'(13700);
			13854: out = 24'(-17428);
			13855: out = 24'(-46272);
			13856: out = 24'(-25804);
			13857: out = 24'(1628);
			13858: out = 24'(15840);
			13859: out = 24'(27796);
			13860: out = 24'(52684);
			13861: out = 24'(37784);
			13862: out = 24'(-15508);
			13863: out = 24'(-68424);
			13864: out = 24'(-49020);
			13865: out = 24'(7152);
			13866: out = 24'(58616);
			13867: out = 24'(82284);
			13868: out = 24'(32016);
			13869: out = 24'(-26980);
			13870: out = 24'(-41324);
			13871: out = 24'(1044);
			13872: out = 24'(1800);
			13873: out = 24'(-16924);
			13874: out = 24'(-17720);
			13875: out = 24'(18124);
			13876: out = 24'(45596);
			13877: out = 24'(22208);
			13878: out = 24'(-3988);
			13879: out = 24'(6628);
			13880: out = 24'(36112);
			13881: out = 24'(-12336);
			13882: out = 24'(-65772);
			13883: out = 24'(-59472);
			13884: out = 24'(4752);
			13885: out = 24'(36908);
			13886: out = 24'(38448);
			13887: out = 24'(26280);
			13888: out = 24'(7612);
			13889: out = 24'(620);
			13890: out = 24'(-3092);
			13891: out = 24'(3840);
			13892: out = 24'(7260);
			13893: out = 24'(1828);
			13894: out = 24'(-7524);
			13895: out = 24'(3432);
			13896: out = 24'(15832);
			13897: out = 24'(-10460);
			13898: out = 24'(-22196);
			13899: out = 24'(-14032);
			13900: out = 24'(-568);
			13901: out = 24'(-1764);
			13902: out = 24'(-27144);
			13903: out = 24'(-20452);
			13904: out = 24'(9708);
			13905: out = 24'(16432);
			13906: out = 24'(4560);
			13907: out = 24'(-7508);
			13908: out = 24'(-188);
			13909: out = 24'(8980);
			13910: out = 24'(6868);
			13911: out = 24'(-18628);
			13912: out = 24'(-34912);
			13913: out = 24'(-11380);
			13914: out = 24'(26720);
			13915: out = 24'(49960);
			13916: out = 24'(27600);
			13917: out = 24'(-6728);
			13918: out = 24'(-23276);
			13919: out = 24'(-40324);
			13920: out = 24'(-74164);
			13921: out = 24'(-76148);
			13922: out = 24'(4736);
			13923: out = 24'(56528);
			13924: out = 24'(49108);
			13925: out = 24'(11552);
			13926: out = 24'(3708);
			13927: out = 24'(-7704);
			13928: out = 24'(-168);
			13929: out = 24'(-6456);
			13930: out = 24'(-14136);
			13931: out = 24'(-928);
			13932: out = 24'(12260);
			13933: out = 24'(12788);
			13934: out = 24'(5060);
			13935: out = 24'(11096);
			13936: out = 24'(16688);
			13937: out = 24'(13752);
			13938: out = 24'(-14860);
			13939: out = 24'(-52048);
			13940: out = 24'(-43124);
			13941: out = 24'(7236);
			13942: out = 24'(32252);
			13943: out = 24'(4052);
			13944: out = 24'(10924);
			13945: out = 24'(12016);
			13946: out = 24'(88);
			13947: out = 24'(-29064);
			13948: out = 24'(-25724);
			13949: out = 24'(-9948);
			13950: out = 24'(7856);
			13951: out = 24'(14888);
			13952: out = 24'(41860);
			13953: out = 24'(47172);
			13954: out = 24'(35448);
			13955: out = 24'(-10064);
			13956: out = 24'(-68784);
			13957: out = 24'(-42596);
			13958: out = 24'(23988);
			13959: out = 24'(40688);
			13960: out = 24'(-80);
			13961: out = 24'(-2932);
			13962: out = 24'(13624);
			13963: out = 24'(4452);
			13964: out = 24'(-38780);
			13965: out = 24'(-5392);
			13966: out = 24'(4604);
			13967: out = 24'(-19200);
			13968: out = 24'(-55244);
			13969: out = 24'(-27800);
			13970: out = 24'(8024);
			13971: out = 24'(29656);
			13972: out = 24'(38820);
			13973: out = 24'(55380);
			13974: out = 24'(47832);
			13975: out = 24'(1624);
			13976: out = 24'(-45544);
			13977: out = 24'(-29252);
			13978: out = 24'(-8972);
			13979: out = 24'(10984);
			13980: out = 24'(20716);
			13981: out = 24'(35888);
			13982: out = 24'(3264);
			13983: out = 24'(-11744);
			13984: out = 24'(-15844);
			13985: out = 24'(-3348);
			13986: out = 24'(7564);
			13987: out = 24'(-5652);
			13988: out = 24'(-26000);
			13989: out = 24'(-19524);
			13990: out = 24'(12740);
			13991: out = 24'(43160);
			13992: out = 24'(41028);
			13993: out = 24'(19872);
			13994: out = 24'(3320);
			13995: out = 24'(-780);
			13996: out = 24'(-13620);
			13997: out = 24'(-39208);
			13998: out = 24'(-52808);
			13999: out = 24'(-20528);
			14000: out = 24'(18824);
			14001: out = 24'(39100);
			14002: out = 24'(39804);
			14003: out = 24'(-17560);
			14004: out = 24'(-23900);
			14005: out = 24'(-22508);
			14006: out = 24'(-19416);
			14007: out = 24'(-12536);
			14008: out = 24'(25952);
			14009: out = 24'(29488);
			14010: out = 24'(352);
			14011: out = 24'(-18576);
			14012: out = 24'(11332);
			14013: out = 24'(27040);
			14014: out = 24'(-12540);
			14015: out = 24'(-95404);
			14016: out = 24'(-34376);
			14017: out = 24'(20972);
			14018: out = 24'(26632);
			14019: out = 24'(504);
			14020: out = 24'(34748);
			14021: out = 24'(33120);
			14022: out = 24'(17948);
			14023: out = 24'(-4604);
			14024: out = 24'(1212);
			14025: out = 24'(-25720);
			14026: out = 24'(-21812);
			14027: out = 24'(5968);
			14028: out = 24'(8916);
			14029: out = 24'(10376);
			14030: out = 24'(18688);
			14031: out = 24'(23948);
			14032: out = 24'(-10220);
			14033: out = 24'(-39452);
			14034: out = 24'(-42836);
			14035: out = 24'(772);
			14036: out = 24'(28988);
			14037: out = 24'(14168);
			14038: out = 24'(-16852);
			14039: out = 24'(-6796);
			14040: out = 24'(20792);
			14041: out = 24'(34744);
			14042: out = 24'(6504);
			14043: out = 24'(6432);
			14044: out = 24'(14884);
			14045: out = 24'(2944);
			14046: out = 24'(-59344);
			14047: out = 24'(-44400);
			14048: out = 24'(24852);
			14049: out = 24'(28284);
			14050: out = 24'(19628);
			14051: out = 24'(19364);
			14052: out = 24'(18860);
			14053: out = 24'(-25636);
			14054: out = 24'(-4700);
			14055: out = 24'(13408);
			14056: out = 24'(18252);
			14057: out = 24'(-5236);
			14058: out = 24'(-1744);
			14059: out = 24'(18716);
			14060: out = 24'(25048);
			14061: out = 24'(-12864);
			14062: out = 24'(-32804);
			14063: out = 24'(-49996);
			14064: out = 24'(-23840);
			14065: out = 24'(4764);
			14066: out = 24'(19992);
			14067: out = 24'(2820);
			14068: out = 24'(10560);
			14069: out = 24'(27572);
			14070: out = 24'(30352);
			14071: out = 24'(12424);
			14072: out = 24'(2540);
			14073: out = 24'(-12964);
			14074: out = 24'(-39700);
			14075: out = 24'(-25364);
			14076: out = 24'(-9284);
			14077: out = 24'(3532);
			14078: out = 24'(14200);
			14079: out = 24'(44668);
			14080: out = 24'(18688);
			14081: out = 24'(-37212);
			14082: out = 24'(-72984);
			14083: out = 24'(-29956);
			14084: out = 24'(-13392);
			14085: out = 24'(-5376);
			14086: out = 24'(21440);
			14087: out = 24'(60612);
			14088: out = 24'(46408);
			14089: out = 24'(-19476);
			14090: out = 24'(-64724);
			14091: out = 24'(-20416);
			14092: out = 24'(14596);
			14093: out = 24'(15648);
			14094: out = 24'(-14392);
			14095: out = 24'(-25032);
			14096: out = 24'(-24888);
			14097: out = 24'(-8624);
			14098: out = 24'(-4060);
			14099: out = 24'(6732);
			14100: out = 24'(33992);
			14101: out = 24'(29960);
			14102: out = 24'(5924);
			14103: out = 24'(-12564);
			14104: out = 24'(-5872);
			14105: out = 24'(-18244);
			14106: out = 24'(-9236);
			14107: out = 24'(31288);
			14108: out = 24'(66772);
			14109: out = 24'(21380);
			14110: out = 24'(-39788);
			14111: out = 24'(-61972);
			14112: out = 24'(-12472);
			14113: out = 24'(7928);
			14114: out = 24'(19760);
			14115: out = 24'(5296);
			14116: out = 24'(4988);
			14117: out = 24'(27576);
			14118: out = 24'(41336);
			14119: out = 24'(19648);
			14120: out = 24'(-3684);
			14121: out = 24'(-2116);
			14122: out = 24'(3392);
			14123: out = 24'(-13492);
			14124: out = 24'(-30680);
			14125: out = 24'(-26276);
			14126: out = 24'(8080);
			14127: out = 24'(7204);
			14128: out = 24'(-3744);
			14129: out = 24'(3444);
			14130: out = 24'(42752);
			14131: out = 24'(7416);
			14132: out = 24'(-47084);
			14133: out = 24'(-60568);
			14134: out = 24'(-6740);
			14135: out = 24'(12960);
			14136: out = 24'(17760);
			14137: out = 24'(25180);
			14138: out = 24'(25512);
			14139: out = 24'(6728);
			14140: out = 24'(-19092);
			14141: out = 24'(-34732);
			14142: out = 24'(-23476);
			14143: out = 24'(11844);
			14144: out = 24'(37236);
			14145: out = 24'(14168);
			14146: out = 24'(-40160);
			14147: out = 24'(-55460);
			14148: out = 24'(-22620);
			14149: out = 24'(6944);
			14150: out = 24'(208);
			14151: out = 24'(-28256);
			14152: out = 24'(15312);
			14153: out = 24'(51304);
			14154: out = 24'(22344);
			14155: out = 24'(-41068);
			14156: out = 24'(-40440);
			14157: out = 24'(7912);
			14158: out = 24'(27212);
			14159: out = 24'(-10660);
			14160: out = 24'(-15612);
			14161: out = 24'(-1096);
			14162: out = 24'(9076);
			14163: out = 24'(-11064);
			14164: out = 24'(18040);
			14165: out = 24'(17512);
			14166: out = 24'(10872);
			14167: out = 24'(-2884);
			14168: out = 24'(3204);
			14169: out = 24'(-22528);
			14170: out = 24'(-22576);
			14171: out = 24'(11544);
			14172: out = 24'(45076);
			14173: out = 24'(9888);
			14174: out = 24'(-36416);
			14175: out = 24'(-48572);
			14176: out = 24'(-14552);
			14177: out = 24'(-2172);
			14178: out = 24'(9656);
			14179: out = 24'(17728);
			14180: out = 24'(16524);
			14181: out = 24'(37068);
			14182: out = 24'(32312);
			14183: out = 24'(-8624);
			14184: out = 24'(-73176);
			14185: out = 24'(-20444);
			14186: out = 24'(16136);
			14187: out = 24'(44680);
			14188: out = 24'(42920);
			14189: out = 24'(35352);
			14190: out = 24'(-18932);
			14191: out = 24'(-45004);
			14192: out = 24'(-36632);
			14193: out = 24'(476);
			14194: out = 24'(-1192);
			14195: out = 24'(10852);
			14196: out = 24'(7592);
			14197: out = 24'(-12624);
			14198: out = 24'(-20816);
			14199: out = 24'(28744);
			14200: out = 24'(48312);
			14201: out = 24'(5840);
			14202: out = 24'(92);
			14203: out = 24'(25456);
			14204: out = 24'(26548);
			14205: out = 24'(-20564);
			14206: out = 24'(-45116);
			14207: out = 24'(1564);
			14208: out = 24'(45664);
			14209: out = 24'(26316);
			14210: out = 24'(-7216);
			14211: out = 24'(-16036);
			14212: out = 24'(-11024);
			14213: out = 24'(-22940);
			14214: out = 24'(-28612);
			14215: out = 24'(12824);
			14216: out = 24'(33880);
			14217: out = 24'(2640);
			14218: out = 24'(-33268);
			14219: out = 24'(-10544);
			14220: out = 24'(32728);
			14221: out = 24'(30276);
			14222: out = 24'(-5676);
			14223: out = 24'(-26372);
			14224: out = 24'(-10324);
			14225: out = 24'(-3412);
			14226: out = 24'(-9476);
			14227: out = 24'(8456);
			14228: out = 24'(27272);
			14229: out = 24'(22560);
			14230: out = 24'(4952);
			14231: out = 24'(-3312);
			14232: out = 24'(-26976);
			14233: out = 24'(-59196);
			14234: out = 24'(-44176);
			14235: out = 24'(37700);
			14236: out = 24'(23996);
			14237: out = 24'(-3556);
			14238: out = 24'(-7456);
			14239: out = 24'(16284);
			14240: out = 24'(-33384);
			14241: out = 24'(-73400);
			14242: out = 24'(-56388);
			14243: out = 24'(18148);
			14244: out = 24'(37568);
			14245: out = 24'(29944);
			14246: out = 24'(11612);
			14247: out = 24'(1832);
			14248: out = 24'(-13632);
			14249: out = 24'(-17556);
			14250: out = 24'(14536);
			14251: out = 24'(48772);
			14252: out = 24'(26656);
			14253: out = 24'(-20952);
			14254: out = 24'(-39804);
			14255: out = 24'(-12556);
			14256: out = 24'(488);
			14257: out = 24'(40436);
			14258: out = 24'(21256);
			14259: out = 24'(4856);
			14260: out = 24'(-12624);
			14261: out = 24'(-52028);
			14262: out = 24'(-67616);
			14263: out = 24'(-21300);
			14264: out = 24'(47100);
			14265: out = 24'(73376);
			14266: out = 24'(38380);
			14267: out = 24'(10368);
			14268: out = 24'(2040);
			14269: out = 24'(-1900);
			14270: out = 24'(-49580);
			14271: out = 24'(-36776);
			14272: out = 24'(16668);
			14273: out = 24'(19216);
			14274: out = 24'(36916);
			14275: out = 24'(7328);
			14276: out = 24'(-11616);
			14277: out = 24'(-18752);
			14278: out = 24'(37848);
			14279: out = 24'(13440);
			14280: out = 24'(-11160);
			14281: out = 24'(-24648);
			14282: out = 24'(-23360);
			14283: out = 24'(-50752);
			14284: out = 24'(-18768);
			14285: out = 24'(48428);
			14286: out = 24'(57944);
			14287: out = 24'(37984);
			14288: out = 24'(8832);
			14289: out = 24'(-5156);
			14290: out = 24'(-14668);
			14291: out = 24'(-70852);
			14292: out = 24'(-65148);
			14293: out = 24'(4264);
			14294: out = 24'(54804);
			14295: out = 24'(32556);
			14296: out = 24'(22100);
			14297: out = 24'(21288);
			14298: out = 24'(396);
			14299: out = 24'(-25908);
			14300: out = 24'(-50692);
			14301: out = 24'(-19680);
			14302: out = 24'(27128);
			14303: out = 24'(34568);
			14304: out = 24'(8156);
			14305: out = 24'(-7552);
			14306: out = 24'(-18796);
			14307: out = 24'(-48028);
			14308: out = 24'(-36944);
			14309: out = 24'(-5900);
			14310: out = 24'(12440);
			14311: out = 24'(-1336);
			14312: out = 24'(-7760);
			14313: out = 24'(5076);
			14314: out = 24'(24600);
			14315: out = 24'(35240);
			14316: out = 24'(46152);
			14317: out = 24'(35048);
			14318: out = 24'(-13084);
			14319: out = 24'(-74864);
			14320: out = 24'(-69276);
			14321: out = 24'(-22052);
			14322: out = 24'(31452);
			14323: out = 24'(40476);
			14324: out = 24'(20556);
			14325: out = 24'(11188);
			14326: out = 24'(2016);
			14327: out = 24'(-26540);
			14328: out = 24'(-62512);
			14329: out = 24'(-11364);
			14330: out = 24'(19644);
			14331: out = 24'(7560);
			14332: out = 24'(-18188);
			14333: out = 24'(2652);
			14334: out = 24'(26552);
			14335: out = 24'(28860);
			14336: out = 24'(12396);
			14337: out = 24'(11488);
			14338: out = 24'(9536);
			14339: out = 24'(6096);
			14340: out = 24'(-2800);
			14341: out = 24'(-76);
			14342: out = 24'(-9892);
			14343: out = 24'(-6624);
			14344: out = 24'(3080);
			14345: out = 24'(9080);
			14346: out = 24'(-2496);
			14347: out = 24'(-10688);
			14348: out = 24'(-4568);
			14349: out = 24'(11996);
			14350: out = 24'(17908);
			14351: out = 24'(11192);
			14352: out = 24'(656);
			14353: out = 24'(176);
			14354: out = 24'(2304);
			14355: out = 24'(14664);
			14356: out = 24'(19352);
			14357: out = 24'(13292);
			14358: out = 24'(-12192);
			14359: out = 24'(-4740);
			14360: out = 24'(1120);
			14361: out = 24'(5804);
			14362: out = 24'(8408);
			14363: out = 24'(24428);
			14364: out = 24'(12672);
			14365: out = 24'(-19344);
			14366: out = 24'(-55088);
			14367: out = 24'(-7788);
			14368: out = 24'(-10660);
			14369: out = 24'(-30400);
			14370: out = 24'(-31900);
			14371: out = 24'(6628);
			14372: out = 24'(18844);
			14373: out = 24'(12792);
			14374: out = 24'(-2052);
			14375: out = 24'(6608);
			14376: out = 24'(-21728);
			14377: out = 24'(-11164);
			14378: out = 24'(16532);
			14379: out = 24'(22228);
			14380: out = 24'(-788);
			14381: out = 24'(4848);
			14382: out = 24'(19044);
			14383: out = 24'(164);
			14384: out = 24'(6052);
			14385: out = 24'(604);
			14386: out = 24'(-7816);
			14387: out = 24'(-29328);
			14388: out = 24'(-10844);
			14389: out = 24'(-5876);
			14390: out = 24'(2440);
			14391: out = 24'(-864);
			14392: out = 24'(12424);
			14393: out = 24'(-14828);
			14394: out = 24'(-13824);
			14395: out = 24'(6276);
			14396: out = 24'(28072);
			14397: out = 24'(-15608);
			14398: out = 24'(-15188);
			14399: out = 24'(19140);
			14400: out = 24'(37020);
			14401: out = 24'(6240);
			14402: out = 24'(-5196);
			14403: out = 24'(3660);
			14404: out = 24'(7292);
			14405: out = 24'(-9052);
			14406: out = 24'(-5824);
			14407: out = 24'(1824);
			14408: out = 24'(-1632);
			14409: out = 24'(-100);
			14410: out = 24'(5228);
			14411: out = 24'(7848);
			14412: out = 24'(-5716);
			14413: out = 24'(-13544);
			14414: out = 24'(-7432);
			14415: out = 24'(15352);
			14416: out = 24'(15552);
			14417: out = 24'(-11932);
			14418: out = 24'(-26412);
			14419: out = 24'(-12436);
			14420: out = 24'(2576);
			14421: out = 24'(-1620);
			14422: out = 24'(-236);
			14423: out = 24'(19536);
			14424: out = 24'(31724);
			14425: out = 24'(7860);
			14426: out = 24'(-42052);
			14427: out = 24'(-37940);
			14428: out = 24'(6300);
			14429: out = 24'(31952);
			14430: out = 24'(23804);
			14431: out = 24'(10912);
			14432: out = 24'(7272);
			14433: out = 24'(-2340);
			14434: out = 24'(-9952);
			14435: out = 24'(-20144);
			14436: out = 24'(12400);
			14437: out = 24'(35892);
			14438: out = 24'(16452);
			14439: out = 24'(-30184);
			14440: out = 24'(-22900);
			14441: out = 24'(11388);
			14442: out = 24'(13040);
			14443: out = 24'(2444);
			14444: out = 24'(-6556);
			14445: out = 24'(9840);
			14446: out = 24'(21124);
			14447: out = 24'(18552);
			14448: out = 24'(1012);
			14449: out = 24'(8132);
			14450: out = 24'(20968);
			14451: out = 24'(5632);
			14452: out = 24'(-8404);
			14453: out = 24'(-11460);
			14454: out = 24'(3380);
			14455: out = 24'(8928);
			14456: out = 24'(-10648);
			14457: out = 24'(-40924);
			14458: out = 24'(-38740);
			14459: out = 24'(3440);
			14460: out = 24'(-2948);
			14461: out = 24'(908);
			14462: out = 24'(-5564);
			14463: out = 24'(-4132);
			14464: out = 24'(644);
			14465: out = 24'(10136);
			14466: out = 24'(2588);
			14467: out = 24'(1852);
			14468: out = 24'(10708);
			14469: out = 24'(6424);
			14470: out = 24'(-19072);
			14471: out = 24'(-15096);
			14472: out = 24'(26012);
			14473: out = 24'(40716);
			14474: out = 24'(280);
			14475: out = 24'(-32372);
			14476: out = 24'(-21356);
			14477: out = 24'(-11176);
			14478: out = 24'(-46220);
			14479: out = 24'(-57468);
			14480: out = 24'(-3676);
			14481: out = 24'(27312);
			14482: out = 24'(14760);
			14483: out = 24'(-4816);
			14484: out = 24'(5104);
			14485: out = 24'(2768);
			14486: out = 24'(7728);
			14487: out = 24'(1968);
			14488: out = 24'(-680);
			14489: out = 24'(-11296);
			14490: out = 24'(-18384);
			14491: out = 24'(-8664);
			14492: out = 24'(12956);
			14493: out = 24'(12432);
			14494: out = 24'(13480);
			14495: out = 24'(7712);
			14496: out = 24'(10024);
			14497: out = 24'(-4872);
			14498: out = 24'(8348);
			14499: out = 24'(-24020);
			14500: out = 24'(-17228);
			14501: out = 24'(14344);
			14502: out = 24'(24080);
			14503: out = 24'(-6680);
			14504: out = 24'(-3188);
			14505: out = 24'(19856);
			14506: out = 24'(-2816);
			14507: out = 24'(-17452);
			14508: out = 24'(-3100);
			14509: out = 24'(20716);
			14510: out = 24'(-3832);
			14511: out = 24'(29384);
			14512: out = 24'(26828);
			14513: out = 24'(12448);
			14514: out = 24'(-14424);
			14515: out = 24'(-364);
			14516: out = 24'(-632);
			14517: out = 24'(9712);
			14518: out = 24'(14048);
			14519: out = 24'(-10092);
			14520: out = 24'(-28608);
			14521: out = 24'(-27472);
			14522: out = 24'(-480);
			14523: out = 24'(36760);
			14524: out = 24'(34984);
			14525: out = 24'(9628);
			14526: out = 24'(-21328);
			14527: out = 24'(-31388);
			14528: out = 24'(-27108);
			14529: out = 24'(-3468);
			14530: out = 24'(13528);
			14531: out = 24'(18968);
			14532: out = 24'(24472);
			14533: out = 24'(30464);
			14534: out = 24'(18864);
			14535: out = 24'(-4896);
			14536: out = 24'(6952);
			14537: out = 24'(1912);
			14538: out = 24'(-15572);
			14539: out = 24'(-35600);
			14540: out = 24'(-22080);
			14541: out = 24'(15904);
			14542: out = 24'(27996);
			14543: out = 24'(-9084);
			14544: out = 24'(-38228);
			14545: out = 24'(-31300);
			14546: out = 24'(24400);
			14547: out = 24'(41484);
			14548: out = 24'(18828);
			14549: out = 24'(-59272);
			14550: out = 24'(-20532);
			14551: out = 24'(35840);
			14552: out = 24'(12356);
			14553: out = 24'(-69848);
			14554: out = 24'(-63624);
			14555: out = 24'(448);
			14556: out = 24'(17256);
			14557: out = 24'(-4536);
			14558: out = 24'(-13872);
			14559: out = 24'(23480);
			14560: out = 24'(43208);
			14561: out = 24'(9132);
			14562: out = 24'(-16424);
			14563: out = 24'(-12952);
			14564: out = 24'(3264);
			14565: out = 24'(-1716);
			14566: out = 24'(640);
			14567: out = 24'(-12936);
			14568: out = 24'(-24068);
			14569: out = 24'(-15532);
			14570: out = 24'(22140);
			14571: out = 24'(27364);
			14572: out = 24'(4404);
			14573: out = 24'(-6572);
			14574: out = 24'(14192);
			14575: out = 24'(1980);
			14576: out = 24'(-60980);
			14577: out = 24'(-96488);
			14578: out = 24'(6256);
			14579: out = 24'(60012);
			14580: out = 24'(51680);
			14581: out = 24'(11196);
			14582: out = 24'(-2412);
			14583: out = 24'(13632);
			14584: out = 24'(9320);
			14585: out = 24'(-18112);
			14586: out = 24'(-28592);
			14587: out = 24'(-1688);
			14588: out = 24'(11496);
			14589: out = 24'(5804);
			14590: out = 24'(-2300);
			14591: out = 24'(-30008);
			14592: out = 24'(-11568);
			14593: out = 24'(15408);
			14594: out = 24'(14812);
			14595: out = 24'(-39496);
			14596: out = 24'(-25648);
			14597: out = 24'(11828);
			14598: out = 24'(35032);
			14599: out = 24'(23052);
			14600: out = 24'(28088);
			14601: out = 24'(15432);
			14602: out = 24'(-19792);
			14603: out = 24'(-66732);
			14604: out = 24'(-47484);
			14605: out = 24'(-15176);
			14606: out = 24'(10752);
			14607: out = 24'(26196);
			14608: out = 24'(60836);
			14609: out = 24'(60844);
			14610: out = 24'(32808);
			14611: out = 24'(-13920);
			14612: out = 24'(-51364);
			14613: out = 24'(-59108);
			14614: out = 24'(-38964);
			14615: out = 24'(-11368);
			14616: out = 24'(12216);
			14617: out = 24'(32808);
			14618: out = 24'(33352);
			14619: out = 24'(15336);
			14620: out = 24'(1276);
			14621: out = 24'(-11016);
			14622: out = 24'(2872);
			14623: out = 24'(6404);
			14624: out = 24'(-16656);
			14625: out = 24'(-59452);
			14626: out = 24'(-26632);
			14627: out = 24'(39612);
			14628: out = 24'(57196);
			14629: out = 24'(28128);
			14630: out = 24'(2132);
			14631: out = 24'(10152);
			14632: out = 24'(12936);
			14633: out = 24'(-9860);
			14634: out = 24'(-62296);
			14635: out = 24'(-38184);
			14636: out = 24'(36864);
			14637: out = 24'(61072);
			14638: out = 24'(1848);
			14639: out = 24'(-45784);
			14640: out = 24'(-46512);
			14641: out = 24'(-23500);
			14642: out = 24'(-1092);
			14643: out = 24'(12380);
			14644: out = 24'(32012);
			14645: out = 24'(42760);
			14646: out = 24'(28936);
			14647: out = 24'(-9732);
			14648: out = 24'(-40240);
			14649: out = 24'(-50188);
			14650: out = 24'(-64644);
			14651: out = 24'(-896);
			14652: out = 24'(42576);
			14653: out = 24'(30236);
			14654: out = 24'(-24168);
			14655: out = 24'(-1016);
			14656: out = 24'(16768);
			14657: out = 24'(20060);
			14658: out = 24'(21764);
			14659: out = 24'(33376);
			14660: out = 24'(15540);
			14661: out = 24'(-33260);
			14662: out = 24'(-69412);
			14663: out = 24'(-41636);
			14664: out = 24'(9608);
			14665: out = 24'(28600);
			14666: out = 24'(26156);
			14667: out = 24'(31740);
			14668: out = 24'(29484);
			14669: out = 24'(-2504);
			14670: out = 24'(-37476);
			14671: out = 24'(-40624);
			14672: out = 24'(-7768);
			14673: out = 24'(5400);
			14674: out = 24'(14792);
			14675: out = 24'(36376);
			14676: out = 24'(28072);
			14677: out = 24'(-7456);
			14678: out = 24'(-22204);
			14679: out = 24'(3748);
			14680: out = 24'(908);
			14681: out = 24'(-26460);
			14682: out = 24'(-35128);
			14683: out = 24'(9596);
			14684: out = 24'(46636);
			14685: out = 24'(20752);
			14686: out = 24'(-28540);
			14687: out = 24'(-41664);
			14688: out = 24'(-11340);
			14689: out = 24'(-3108);
			14690: out = 24'(-3220);
			14691: out = 24'(12596);
			14692: out = 24'(37096);
			14693: out = 24'(48600);
			14694: out = 24'(26988);
			14695: out = 24'(124);
			14696: out = 24'(-11292);
			14697: out = 24'(-20748);
			14698: out = 24'(-21320);
			14699: out = 24'(-17676);
			14700: out = 24'(-7332);
			14701: out = 24'(-1316);
			14702: out = 24'(26356);
			14703: out = 24'(36956);
			14704: out = 24'(20112);
			14705: out = 24'(1916);
			14706: out = 24'(-1552);
			14707: out = 24'(18192);
			14708: out = 24'(19604);
			14709: out = 24'(-12896);
			14710: out = 24'(-48288);
			14711: out = 24'(-36356);
			14712: out = 24'(6224);
			14713: out = 24'(28800);
			14714: out = 24'(53136);
			14715: out = 24'(41868);
			14716: out = 24'(10196);
			14717: out = 24'(-33744);
			14718: out = 24'(-41152);
			14719: out = 24'(-24288);
			14720: out = 24'(17636);
			14721: out = 24'(37408);
			14722: out = 24'(28024);
			14723: out = 24'(-4612);
			14724: out = 24'(-7576);
			14725: out = 24'(6136);
			14726: out = 24'(6476);
			14727: out = 24'(-42532);
			14728: out = 24'(-41868);
			14729: out = 24'(8232);
			14730: out = 24'(25844);
			14731: out = 24'(9296);
			14732: out = 24'(-20112);
			14733: out = 24'(-4980);
			14734: out = 24'(27148);
			14735: out = 24'(29124);
			14736: out = 24'(-19772);
			14737: out = 24'(-49192);
			14738: out = 24'(-29152);
			14739: out = 24'(6512);
			14740: out = 24'(14568);
			14741: out = 24'(16312);
			14742: out = 24'(14136);
			14743: out = 24'(-11124);
			14744: out = 24'(3824);
			14745: out = 24'(8632);
			14746: out = 24'(-15504);
			14747: out = 24'(-52708);
			14748: out = 24'(-49908);
			14749: out = 24'(2944);
			14750: out = 24'(37916);
			14751: out = 24'(23992);
			14752: out = 24'(3540);
			14753: out = 24'(13460);
			14754: out = 24'(21944);
			14755: out = 24'(3556);
			14756: out = 24'(-13692);
			14757: out = 24'(-4216);
			14758: out = 24'(11872);
			14759: out = 24'(9416);
			14760: out = 24'(-10820);
			14761: out = 24'(-15288);
			14762: out = 24'(-19776);
			14763: out = 24'(-16624);
			14764: out = 24'(2644);
			14765: out = 24'(47196);
			14766: out = 24'(37548);
			14767: out = 24'(-4692);
			14768: out = 24'(-29352);
			14769: out = 24'(-6844);
			14770: out = 24'(-3516);
			14771: out = 24'(-14948);
			14772: out = 24'(-4884);
			14773: out = 24'(9088);
			14774: out = 24'(16900);
			14775: out = 24'(-15528);
			14776: out = 24'(-43440);
			14777: out = 24'(-380);
			14778: out = 24'(22704);
			14779: out = 24'(20560);
			14780: out = 24'(10340);
			14781: out = 24'(26972);
			14782: out = 24'(-3736);
			14783: out = 24'(-24768);
			14784: out = 24'(-28572);
			14785: out = 24'(-7516);
			14786: out = 24'(13244);
			14787: out = 24'(28488);
			14788: out = 24'(24480);
			14789: out = 24'(5640);
			14790: out = 24'(248);
			14791: out = 24'(-10236);
			14792: out = 24'(-7604);
			14793: out = 24'(464);
			14794: out = 24'(4124);
			14795: out = 24'(60);
			14796: out = 24'(-128);
			14797: out = 24'(-4100);
			14798: out = 24'(-15180);
			14799: out = 24'(-22504);
			14800: out = 24'(-1512);
			14801: out = 24'(27660);
			14802: out = 24'(39832);
			14803: out = 24'(5588);
			14804: out = 24'(-8808);
			14805: out = 24'(-18352);
			14806: out = 24'(-32436);
			14807: out = 24'(-23584);
			14808: out = 24'(10164);
			14809: out = 24'(29192);
			14810: out = 24'(11956);
			14811: out = 24'(1972);
			14812: out = 24'(-4684);
			14813: out = 24'(1080);
			14814: out = 24'(-8356);
			14815: out = 24'(-28712);
			14816: out = 24'(-8928);
			14817: out = 24'(26960);
			14818: out = 24'(31356);
			14819: out = 24'(3676);
			14820: out = 24'(-18488);
			14821: out = 24'(-16300);
			14822: out = 24'(-13200);
			14823: out = 24'(-20784);
			14824: out = 24'(-21788);
			14825: out = 24'(4088);
			14826: out = 24'(26704);
			14827: out = 24'(28576);
			14828: out = 24'(5284);
			14829: out = 24'(2696);
			14830: out = 24'(-15624);
			14831: out = 24'(-35720);
			14832: out = 24'(-11068);
			14833: out = 24'(6320);
			14834: out = 24'(1764);
			14835: out = 24'(-10680);
			14836: out = 24'(1708);
			14837: out = 24'(580);
			14838: out = 24'(-636);
			14839: out = 24'(5036);
			14840: out = 24'(17276);
			14841: out = 24'(-308);
			14842: out = 24'(-27036);
			14843: out = 24'(-24004);
			14844: out = 24'(15332);
			14845: out = 24'(21560);
			14846: out = 24'(5292);
			14847: out = 24'(-836);
			14848: out = 24'(25536);
			14849: out = 24'(26616);
			14850: out = 24'(12312);
			14851: out = 24'(-12336);
			14852: out = 24'(-1116);
			14853: out = 24'(17348);
			14854: out = 24'(41840);
			14855: out = 24'(-14968);
			14856: out = 24'(-72344);
			14857: out = 24'(-33252);
			14858: out = 24'(16404);
			14859: out = 24'(44440);
			14860: out = 24'(22584);
			14861: out = 24'(-3128);
			14862: out = 24'(-36504);
			14863: out = 24'(-13220);
			14864: out = 24'(3872);
			14865: out = 24'(5736);
			14866: out = 24'(20760);
			14867: out = 24'(30380);
			14868: out = 24'(9460);
			14869: out = 24'(-29908);
			14870: out = 24'(-28616);
			14871: out = 24'(-11572);
			14872: out = 24'(18328);
			14873: out = 24'(19184);
			14874: out = 24'(-6404);
			14875: out = 24'(-12264);
			14876: out = 24'(680);
			14877: out = 24'(8144);
			14878: out = 24'(-2468);
			14879: out = 24'(-14208);
			14880: out = 24'(-2140);
			14881: out = 24'(13504);
			14882: out = 24'(2200);
			14883: out = 24'(-26348);
			14884: out = 24'(-20192);
			14885: out = 24'(17164);
			14886: out = 24'(28588);
			14887: out = 24'(1312);
			14888: out = 24'(-35860);
			14889: out = 24'(-23104);
			14890: out = 24'(15704);
			14891: out = 24'(28572);
			14892: out = 24'(-5820);
			14893: out = 24'(-18200);
			14894: out = 24'(-872);
			14895: out = 24'(17300);
			14896: out = 24'(-7296);
			14897: out = 24'(-2864);
			14898: out = 24'(6344);
			14899: out = 24'(-4172);
			14900: out = 24'(-27624);
			14901: out = 24'(-13756);
			14902: out = 24'(9032);
			14903: out = 24'(6584);
			14904: out = 24'(3472);
			14905: out = 24'(-2112);
			14906: out = 24'(5604);
			14907: out = 24'(-1036);
			14908: out = 24'(-18044);
			14909: out = 24'(-23528);
			14910: out = 24'(-236);
			14911: out = 24'(17996);
			14912: out = 24'(17644);
			14913: out = 24'(-19400);
			14914: out = 24'(-14400);
			14915: out = 24'(16192);
			14916: out = 24'(41620);
			14917: out = 24'(-7516);
			14918: out = 24'(-12928);
			14919: out = 24'(-23168);
			14920: out = 24'(-25504);
			14921: out = 24'(-4564);
			14922: out = 24'(44808);
			14923: out = 24'(33716);
			14924: out = 24'(-6336);
			14925: out = 24'(-9736);
			14926: out = 24'(10720);
			14927: out = 24'(-8472);
			14928: out = 24'(-36560);
			14929: out = 24'(-6040);
			14930: out = 24'(24960);
			14931: out = 24'(14852);
			14932: out = 24'(-10460);
			14933: out = 24'(2964);
			14934: out = 24'(1404);
			14935: out = 24'(5592);
			14936: out = 24'(11308);
			14937: out = 24'(26152);
			14938: out = 24'(-596);
			14939: out = 24'(-15500);
			14940: out = 24'(-14088);
			14941: out = 24'(11072);
			14942: out = 24'(14960);
			14943: out = 24'(26544);
			14944: out = 24'(20916);
			14945: out = 24'(15484);
			14946: out = 24'(6196);
			14947: out = 24'(1280);
			14948: out = 24'(-17588);
			14949: out = 24'(-25892);
			14950: out = 24'(-9800);
			14951: out = 24'(-4120);
			14952: out = 24'(2888);
			14953: out = 24'(3768);
			14954: out = 24'(3804);
			14955: out = 24'(-1768);
			14956: out = 24'(-780);
			14957: out = 24'(-1072);
			14958: out = 24'(148);
			14959: out = 24'(3200);
			14960: out = 24'(1412);
			14961: out = 24'(-2764);
			14962: out = 24'(5724);
			14963: out = 24'(28464);
			14964: out = 24'(28060);
			14965: out = 24'(5848);
			14966: out = 24'(-20776);
			14967: out = 24'(-33412);
			14968: out = 24'(-36632);
			14969: out = 24'(-44728);
			14970: out = 24'(-36624);
			14971: out = 24'(8388);
			14972: out = 24'(32376);
			14973: out = 24'(44080);
			14974: out = 24'(19284);
			14975: out = 24'(-18820);
			14976: out = 24'(-67748);
			14977: out = 24'(-33024);
			14978: out = 24'(6528);
			14979: out = 24'(4132);
			14980: out = 24'(-16020);
			14981: out = 24'(-7756);
			14982: out = 24'(25956);
			14983: out = 24'(39904);
			14984: out = 24'(11468);
			14985: out = 24'(-8768);
			14986: out = 24'(-22400);
			14987: out = 24'(-9296);
			14988: out = 24'(17856);
			14989: out = 24'(-20136);
			14990: out = 24'(-20848);
			14991: out = 24'(9500);
			14992: out = 24'(37352);
			14993: out = 24'(-7712);
			14994: out = 24'(-12356);
			14995: out = 24'(-2356);
			14996: out = 24'(11160);
			14997: out = 24'(-2588);
			14998: out = 24'(-5040);
			14999: out = 24'(-23348);
			15000: out = 24'(-20356);
			15001: out = 24'(24988);
			15002: out = 24'(66300);
			15003: out = 24'(45796);
			15004: out = 24'(-6372);
			15005: out = 24'(-29612);
			15006: out = 24'(-31204);
			15007: out = 24'(-15288);
			15008: out = 24'(-5884);
			15009: out = 24'(16592);
			15010: out = 24'(36164);
			15011: out = 24'(43768);
			15012: out = 24'(-1356);
			15013: out = 24'(-58996);
			15014: out = 24'(-48168);
			15015: out = 24'(-28312);
			15016: out = 24'(-14732);
			15017: out = 24'(-1660);
			15018: out = 24'(28292);
			15019: out = 24'(50820);
			15020: out = 24'(37600);
			15021: out = 24'(8896);
			15022: out = 24'(-1856);
			15023: out = 24'(-23328);
			15024: out = 24'(-32036);
			15025: out = 24'(-22472);
			15026: out = 24'(1824);
			15027: out = 24'(-9152);
			15028: out = 24'(388);
			15029: out = 24'(26744);
			15030: out = 24'(42012);
			15031: out = 24'(1084);
			15032: out = 24'(-35128);
			15033: out = 24'(-46648);
			15034: out = 24'(-19140);
			15035: out = 24'(16924);
			15036: out = 24'(11196);
			15037: out = 24'(-40);
			15038: out = 24'(10156);
			15039: out = 24'(38128);
			15040: out = 24'(6852);
			15041: out = 24'(-13804);
			15042: out = 24'(-22660);
			15043: out = 24'(-21396);
			15044: out = 24'(-44992);
			15045: out = 24'(-32428);
			15046: out = 24'(-5740);
			15047: out = 24'(11244);
			15048: out = 24'(-8200);
			15049: out = 24'(13564);
			15050: out = 24'(33340);
			15051: out = 24'(26280);
			15052: out = 24'(-34392);
			15053: out = 24'(-8928);
			15054: out = 24'(-828);
			15055: out = 24'(-11684);
			15056: out = 24'(-5344);
			15057: out = 24'(43488);
			15058: out = 24'(47580);
			15059: out = 24'(6072);
			15060: out = 24'(-27688);
			15061: out = 24'(-6184);
			15062: out = 24'(8368);
			15063: out = 24'(-5224);
			15064: out = 24'(-11484);
			15065: out = 24'(-4628);
			15066: out = 24'(28492);
			15067: out = 24'(24404);
			15068: out = 24'(1412);
			15069: out = 24'(-10588);
			15070: out = 24'(30304);
			15071: out = 24'(31896);
			15072: out = 24'(-4160);
			15073: out = 24'(-29732);
			15074: out = 24'(-8456);
			15075: out = 24'(2596);
			15076: out = 24'(2060);
			15077: out = 24'(20420);
			15078: out = 24'(23628);
			15079: out = 24'(12548);
			15080: out = 24'(-18884);
			15081: out = 24'(-42748);
			15082: out = 24'(-33932);
			15083: out = 24'(-12272);
			15084: out = 24'(14456);
			15085: out = 24'(30020);
			15086: out = 24'(9500);
			15087: out = 24'(1740);
			15088: out = 24'(2716);
			15089: out = 24'(7452);
			15090: out = 24'(-13016);
			15091: out = 24'(-9508);
			15092: out = 24'(-22440);
			15093: out = 24'(-26976);
			15094: out = 24'(3164);
			15095: out = 24'(21412);
			15096: out = 24'(28768);
			15097: out = 24'(10428);
			15098: out = 24'(-13216);
			15099: out = 24'(-50432);
			15100: out = 24'(-23236);
			15101: out = 24'(20612);
			15102: out = 24'(45948);
			15103: out = 24'(51176);
			15104: out = 24'(22480);
			15105: out = 24'(-35284);
			15106: out = 24'(-76068);
			15107: out = 24'(-30936);
			15108: out = 24'(17492);
			15109: out = 24'(32448);
			15110: out = 24'(1900);
			15111: out = 24'(-44800);
			15112: out = 24'(-23316);
			15113: out = 24'(1648);
			15114: out = 24'(18108);
			15115: out = 24'(37984);
			15116: out = 24'(47580);
			15117: out = 24'(23312);
			15118: out = 24'(-26268);
			15119: out = 24'(-56940);
			15120: out = 24'(-36232);
			15121: out = 24'(8188);
			15122: out = 24'(30068);
			15123: out = 24'(29516);
			15124: out = 24'(17056);
			15125: out = 24'(-7512);
			15126: out = 24'(-46008);
			15127: out = 24'(-55428);
			15128: out = 24'(720);
			15129: out = 24'(13748);
			15130: out = 24'(12384);
			15131: out = 24'(14640);
			15132: out = 24'(26496);
			15133: out = 24'(13624);
			15134: out = 24'(-9668);
			15135: out = 24'(-20864);
			15136: out = 24'(-17056);
			15137: out = 24'(-42488);
			15138: out = 24'(-28568);
			15139: out = 24'(24112);
			15140: out = 24'(50276);
			15141: out = 24'(-18644);
			15142: out = 24'(-42804);
			15143: out = 24'(-2188);
			15144: out = 24'(43972);
			15145: out = 24'(-6900);
			15146: out = 24'(2984);
			15147: out = 24'(20548);
			15148: out = 24'(35348);
			15149: out = 24'(14572);
			15150: out = 24'(-12756);
			15151: out = 24'(-9820);
			15152: out = 24'(28088);
			15153: out = 24'(43316);
			15154: out = 24'(-1556);
			15155: out = 24'(-39844);
			15156: out = 24'(-37356);
			15157: out = 24'(-7912);
			15158: out = 24'(-15684);
			15159: out = 24'(-4488);
			15160: out = 24'(14604);
			15161: out = 24'(29860);
			15162: out = 24'(-7208);
			15163: out = 24'(21028);
			15164: out = 24'(22068);
			15165: out = 24'(6940);
			15166: out = 24'(-16580);
			15167: out = 24'(20716);
			15168: out = 24'(3752);
			15169: out = 24'(-31244);
			15170: out = 24'(-26128);
			15171: out = 24'(17060);
			15172: out = 24'(22368);
			15173: out = 24'(-8948);
			15174: out = 24'(-29556);
			15175: out = 24'(-14696);
			15176: out = 24'(-1084);
			15177: out = 24'(-5884);
			15178: out = 24'(-5772);
			15179: out = 24'(17056);
			15180: out = 24'(38580);
			15181: out = 24'(29500);
			15182: out = 24'(-2168);
			15183: out = 24'(-24340);
			15184: out = 24'(-13864);
			15185: out = 24'(9664);
			15186: out = 24'(14388);
			15187: out = 24'(-744);
			15188: out = 24'(6716);
			15189: out = 24'(17276);
			15190: out = 24'(16264);
			15191: out = 24'(-7320);
			15192: out = 24'(-23112);
			15193: out = 24'(-22148);
			15194: out = 24'(6256);
			15195: out = 24'(26744);
			15196: out = 24'(31036);
			15197: out = 24'(-1744);
			15198: out = 24'(-11476);
			15199: out = 24'(1544);
			15200: out = 24'(12060);
			15201: out = 24'(-3600);
			15202: out = 24'(-5492);
			15203: out = 24'(-1192);
			15204: out = 24'(-3628);
			15205: out = 24'(-42128);
			15206: out = 24'(-32920);
			15207: out = 24'(5712);
			15208: out = 24'(31712);
			15209: out = 24'(36740);
			15210: out = 24'(21804);
			15211: out = 24'(-13628);
			15212: out = 24'(-41924);
			15213: out = 24'(-20332);
			15214: out = 24'(7584);
			15215: out = 24'(4176);
			15216: out = 24'(-11404);
			15217: out = 24'(-1312);
			15218: out = 24'(1860);
			15219: out = 24'(-22420);
			15220: out = 24'(-37712);
			15221: out = 24'(-3464);
			15222: out = 24'(33640);
			15223: out = 24'(10960);
			15224: out = 24'(-34140);
			15225: out = 24'(-35468);
			15226: out = 24'(1668);
			15227: out = 24'(15000);
			15228: out = 24'(10456);
			15229: out = 24'(21176);
			15230: out = 24'(8304);
			15231: out = 24'(1460);
			15232: out = 24'(-9272);
			15233: out = 24'(-2140);
			15234: out = 24'(-3464);
			15235: out = 24'(3260);
			15236: out = 24'(-3228);
			15237: out = 24'(11240);
			15238: out = 24'(38692);
			15239: out = 24'(13180);
			15240: out = 24'(-34096);
			15241: out = 24'(-45688);
			15242: out = 24'(-9620);
			15243: out = 24'(468);
			15244: out = 24'(-3440);
			15245: out = 24'(22952);
			15246: out = 24'(61008);
			15247: out = 24'(31616);
			15248: out = 24'(-35688);
			15249: out = 24'(-58488);
			15250: out = 24'(-4680);
			15251: out = 24'(-5072);
			15252: out = 24'(14436);
			15253: out = 24'(11316);
			15254: out = 24'(5072);
			15255: out = 24'(-27436);
			15256: out = 24'(-20652);
			15257: out = 24'(-13196);
			15258: out = 24'(16432);
			15259: out = 24'(54484);
			15260: out = 24'(57904);
			15261: out = 24'(24956);
			15262: out = 24'(-23644);
			15263: out = 24'(-53804);
			15264: out = 24'(-51676);
			15265: out = 24'(-17104);
			15266: out = 24'(11628);
			15267: out = 24'(15148);
			15268: out = 24'(-17680);
			15269: out = 24'(7920);
			15270: out = 24'(34868);
			15271: out = 24'(20848);
			15272: out = 24'(-43828);
			15273: out = 24'(-24248);
			15274: out = 24'(15700);
			15275: out = 24'(26752);
			15276: out = 24'(-332);
			15277: out = 24'(2828);
			15278: out = 24'(14352);
			15279: out = 24'(21448);
			15280: out = 24'(6792);
			15281: out = 24'(22748);
			15282: out = 24'(1088);
			15283: out = 24'(-19952);
			15284: out = 24'(-25160);
			15285: out = 24'(-1928);
			15286: out = 24'(-264);
			15287: out = 24'(-96);
			15288: out = 24'(-3624);
			15289: out = 24'(-9360);
			15290: out = 24'(1768);
			15291: out = 24'(21452);
			15292: out = 24'(19820);
			15293: out = 24'(400);
			15294: out = 24'(-2332);
			15295: out = 24'(27384);
			15296: out = 24'(33332);
			15297: out = 24'(184);
			15298: out = 24'(-34356);
			15299: out = 24'(-7104);
			15300: out = 24'(18208);
			15301: out = 24'(-9676);
			15302: out = 24'(-27712);
			15303: out = 24'(-9940);
			15304: out = 24'(19700);
			15305: out = 24'(10424);
			15306: out = 24'(2712);
			15307: out = 24'(-28728);
			15308: out = 24'(-17948);
			15309: out = 24'(7376);
			15310: out = 24'(7208);
			15311: out = 24'(-17556);
			15312: out = 24'(-29124);
			15313: out = 24'(-6820);
			15314: out = 24'(26160);
			15315: out = 24'(13604);
			15316: out = 24'(-4800);
			15317: out = 24'(-6060);
			15318: out = 24'(9204);
			15319: out = 24'(-4300);
			15320: out = 24'(-26372);
			15321: out = 24'(-28288);
			15322: out = 24'(9712);
			15323: out = 24'(17088);
			15324: out = 24'(26168);
			15325: out = 24'(-6496);
			15326: out = 24'(-30096);
			15327: out = 24'(-17216);
			15328: out = 24'(11460);
			15329: out = 24'(-160);
			15330: out = 24'(-11564);
			15331: out = 24'(10464);
			15332: out = 24'(27472);
			15333: out = 24'(-9784);
			15334: out = 24'(-45768);
			15335: out = 24'(-19760);
			15336: out = 24'(-9372);
			15337: out = 24'(6304);
			15338: out = 24'(24660);
			15339: out = 24'(51172);
			15340: out = 24'(13636);
			15341: out = 24'(8376);
			15342: out = 24'(880);
			15343: out = 24'(-3836);
			15344: out = 24'(-31780);
			15345: out = 24'(-1656);
			15346: out = 24'(24912);
			15347: out = 24'(30832);
			15348: out = 24'(5468);
			15349: out = 24'(-34440);
			15350: out = 24'(-55908);
			15351: out = 24'(-26300);
			15352: out = 24'(19096);
			15353: out = 24'(14124);
			15354: out = 24'(1184);
			15355: out = 24'(13460);
			15356: out = 24'(35356);
			15357: out = 24'(36300);
			15358: out = 24'(2240);
			15359: out = 24'(-6776);
			15360: out = 24'(9188);
			15361: out = 24'(-11240);
			15362: out = 24'(-30728);
			15363: out = 24'(-16372);
			15364: out = 24'(29852);
			15365: out = 24'(28516);
			15366: out = 24'(26044);
			15367: out = 24'(-6684);
			15368: out = 24'(-24936);
			15369: out = 24'(-33488);
			15370: out = 24'(-11948);
			15371: out = 24'(-15932);
			15372: out = 24'(-2140);
			15373: out = 24'(28336);
			15374: out = 24'(27588);
			15375: out = 24'(1232);
			15376: out = 24'(-7852);
			15377: out = 24'(10460);
			15378: out = 24'(-7564);
			15379: out = 24'(-3664);
			15380: out = 24'(9412);
			15381: out = 24'(28000);
			15382: out = 24'(13584);
			15383: out = 24'(-6000);
			15384: out = 24'(-32072);
			15385: out = 24'(-33936);
			15386: out = 24'(-25808);
			15387: out = 24'(33324);
			15388: out = 24'(34544);
			15389: out = 24'(10004);
			15390: out = 24'(-11248);
			15391: out = 24'(15064);
			15392: out = 24'(744);
			15393: out = 24'(-18716);
			15394: out = 24'(-17400);
			15395: out = 24'(15180);
			15396: out = 24'(12224);
			15397: out = 24'(5864);
			15398: out = 24'(-1624);
			15399: out = 24'(-20020);
			15400: out = 24'(-24964);
			15401: out = 24'(80);
			15402: out = 24'(22124);
			15403: out = 24'(2496);
			15404: out = 24'(-8980);
			15405: out = 24'(5972);
			15406: out = 24'(33420);
			15407: out = 24'(26512);
			15408: out = 24'(-20668);
			15409: out = 24'(-41468);
			15410: out = 24'(-12008);
			15411: out = 24'(20412);
			15412: out = 24'(1756);
			15413: out = 24'(-24252);
			15414: out = 24'(-23916);
			15415: out = 24'(4016);
			15416: out = 24'(6484);
			15417: out = 24'(4572);
			15418: out = 24'(-9248);
			15419: out = 24'(-4348);
			15420: out = 24'(15180);
			15421: out = 24'(-196);
			15422: out = 24'(-39904);
			15423: out = 24'(-48600);
			15424: out = 24'(3804);
			15425: out = 24'(16628);
			15426: out = 24'(18452);
			15427: out = 24'(29000);
			15428: out = 24'(51028);
			15429: out = 24'(5024);
			15430: out = 24'(-32392);
			15431: out = 24'(-45160);
			15432: out = 24'(-14260);
			15433: out = 24'(-15172);
			15434: out = 24'(19956);
			15435: out = 24'(19740);
			15436: out = 24'(804);
			15437: out = 24'(-4420);
			15438: out = 24'(17616);
			15439: out = 24'(26544);
			15440: out = 24'(2240);
			15441: out = 24'(-39984);
			15442: out = 24'(-23228);
			15443: out = 24'(1960);
			15444: out = 24'(3784);
			15445: out = 24'(-13712);
			15446: out = 24'(21804);
			15447: out = 24'(19336);
			15448: out = 24'(-5700);
			15449: out = 24'(-25380);
			15450: out = 24'(-22200);
			15451: out = 24'(12676);
			15452: out = 24'(31076);
			15453: out = 24'(16672);
			15454: out = 24'(-28564);
			15455: out = 24'(-14552);
			15456: out = 24'(4396);
			15457: out = 24'(8540);
			15458: out = 24'(4628);
			15459: out = 24'(8532);
			15460: out = 24'(2072);
			15461: out = 24'(-10436);
			15462: out = 24'(-15656);
			15463: out = 24'(-24520);
			15464: out = 24'(-11936);
			15465: out = 24'(15128);
			15466: out = 24'(32928);
			15467: out = 24'(20068);
			15468: out = 24'(-11348);
			15469: out = 24'(-31832);
			15470: out = 24'(-27948);
			15471: out = 24'(-20300);
			15472: out = 24'(1324);
			15473: out = 24'(32128);
			15474: out = 24'(52664);
			15475: out = 24'(26464);
			15476: out = 24'(14964);
			15477: out = 24'(-4444);
			15478: out = 24'(-18904);
			15479: out = 24'(-50820);
			15480: out = 24'(-43764);
			15481: out = 24'(-34824);
			15482: out = 24'(18268);
			15483: out = 24'(62160);
			15484: out = 24'(38068);
			15485: out = 24'(-27580);
			15486: out = 24'(-39740);
			15487: out = 24'(8040);
			15488: out = 24'(7512);
			15489: out = 24'(-10328);
			15490: out = 24'(-13212);
			15491: out = 24'(13124);
			15492: out = 24'(20312);
			15493: out = 24'(13548);
			15494: out = 24'(10076);
			15495: out = 24'(10904);
			15496: out = 24'(-7604);
			15497: out = 24'(-10064);
			15498: out = 24'(444);
			15499: out = 24'(4264);
			15500: out = 24'(-22700);
			15501: out = 24'(472);
			15502: out = 24'(1776);
			15503: out = 24'(4384);
			15504: out = 24'(-1668);
			15505: out = 24'(2132);
			15506: out = 24'(-8992);
			15507: out = 24'(-4508);
			15508: out = 24'(4244);
			15509: out = 24'(336);
			15510: out = 24'(-15484);
			15511: out = 24'(-13808);
			15512: out = 24'(8612);
			15513: out = 24'(25032);
			15514: out = 24'(17448);
			15515: out = 24'(4376);
			15516: out = 24'(-2788);
			15517: out = 24'(-13364);
			15518: out = 24'(-27000);
			15519: out = 24'(-28096);
			15520: out = 24'(-5364);
			15521: out = 24'(16052);
			15522: out = 24'(27756);
			15523: out = 24'(19176);
			15524: out = 24'(19660);
			15525: out = 24'(12016);
			15526: out = 24'(1984);
			15527: out = 24'(-75324);
			15528: out = 24'(-81788);
			15529: out = 24'(-8140);
			15530: out = 24'(39244);
			15531: out = 24'(27864);
			15532: out = 24'(14292);
			15533: out = 24'(24824);
			15534: out = 24'(21784);
			15535: out = 24'(-796);
			15536: out = 24'(-36080);
			15537: out = 24'(-35024);
			15538: out = 24'(2888);
			15539: out = 24'(38308);
			15540: out = 24'(37424);
			15541: out = 24'(18644);
			15542: out = 24'(824);
			15543: out = 24'(-4988);
			15544: out = 24'(4012);
			15545: out = 24'(11560);
			15546: out = 24'(2884);
			15547: out = 24'(-14224);
			15548: out = 24'(-21948);
			15549: out = 24'(-9084);
			15550: out = 24'(1092);
			15551: out = 24'(1204);
			15552: out = 24'(-2560);
			15553: out = 24'(24616);
			15554: out = 24'(39044);
			15555: out = 24'(8880);
			15556: out = 24'(-32752);
			15557: out = 24'(-32324);
			15558: out = 24'(3064);
			15559: out = 24'(12612);
			15560: out = 24'(-5496);
			15561: out = 24'(-23144);
			15562: out = 24'(3192);
			15563: out = 24'(29360);
			15564: out = 24'(4400);
			15565: out = 24'(-8428);
			15566: out = 24'(212);
			15567: out = 24'(13332);
			15568: out = 24'(-3676);
			15569: out = 24'(-45428);
			15570: out = 24'(-46264);
			15571: out = 24'(9960);
			15572: out = 24'(54100);
			15573: out = 24'(36108);
			15574: out = 24'(2420);
			15575: out = 24'(-15652);
			15576: out = 24'(-21944);
			15577: out = 24'(-18008);
			15578: out = 24'(-29904);
			15579: out = 24'(-8176);
			15580: out = 24'(35816);
			15581: out = 24'(45936);
			15582: out = 24'(21404);
			15583: out = 24'(-4624);
			15584: out = 24'(-12112);
			15585: out = 24'(-21980);
			15586: out = 24'(-11568);
			15587: out = 24'(-6260);
			15588: out = 24'(3752);
			15589: out = 24'(10448);
			15590: out = 24'(48400);
			15591: out = 24'(28448);
			15592: out = 24'(-6380);
			15593: out = 24'(-17052);
			15594: out = 24'(20184);
			15595: out = 24'(11348);
			15596: out = 24'(-18204);
			15597: out = 24'(-28972);
			15598: out = 24'(-14096);
			15599: out = 24'(-1896);
			15600: out = 24'(-3188);
			15601: out = 24'(9412);
			15602: out = 24'(42016);
			15603: out = 24'(50436);
			15604: out = 24'(4312);
			15605: out = 24'(-65328);
			15606: out = 24'(-98944);
			15607: out = 24'(-23168);
			15608: out = 24'(35256);
			15609: out = 24'(33260);
			15610: out = 24'(20860);
			15611: out = 24'(35672);
			15612: out = 24'(21944);
			15613: out = 24'(-47948);
			15614: out = 24'(-111152);
			15615: out = 24'(-49040);
			15616: out = 24'(12936);
			15617: out = 24'(27100);
			15618: out = 24'(22832);
			15619: out = 24'(44216);
			15620: out = 24'(28628);
			15621: out = 24'(-20704);
			15622: out = 24'(-56544);
			15623: out = 24'(-15620);
			15624: out = 24'(18400);
			15625: out = 24'(22256);
			15626: out = 24'(2856);
			15627: out = 24'(1888);
			15628: out = 24'(-1704);
			15629: out = 24'(9992);
			15630: out = 24'(11760);
			15631: out = 24'(2756);
			15632: out = 24'(580);
			15633: out = 24'(-8856);
			15634: out = 24'(-10248);
			15635: out = 24'(-10460);
			15636: out = 24'(1012);
			15637: out = 24'(-3696);
			15638: out = 24'(13976);
			15639: out = 24'(26236);
			15640: out = 24'(26600);
			15641: out = 24'(-11064);
			15642: out = 24'(-3120);
			15643: out = 24'(3060);
			15644: out = 24'(-22524);
			15645: out = 24'(-55292);
			15646: out = 24'(-9764);
			15647: out = 24'(35836);
			15648: out = 24'(16672);
			15649: out = 24'(17456);
			15650: out = 24'(14192);
			15651: out = 24'(13572);
			15652: out = 24'(-11108);
			15653: out = 24'(-53320);
			15654: out = 24'(-28132);
			15655: out = 24'(5892);
			15656: out = 24'(6704);
			15657: out = 24'(3964);
			15658: out = 24'(27852);
			15659: out = 24'(39060);
			15660: out = 24'(5908);
			15661: out = 24'(-40144);
			15662: out = 24'(-68840);
			15663: out = 24'(-42856);
			15664: out = 24'(-5800);
			15665: out = 24'(14004);
			15666: out = 24'(32236);
			15667: out = 24'(47016);
			15668: out = 24'(39156);
			15669: out = 24'(9304);
			15670: out = 24'(-32048);
			15671: out = 24'(-41008);
			15672: out = 24'(-39188);
			15673: out = 24'(-26848);
			15674: out = 24'(5528);
			15675: out = 24'(28432);
			15676: out = 24'(18944);
			15677: out = 24'(-2756);
			15678: out = 24'(2380);
			15679: out = 24'(-360);
			15680: out = 24'(2668);
			15681: out = 24'(-8148);
			15682: out = 24'(-29524);
			15683: out = 24'(-10932);
			15684: out = 24'(5876);
			15685: out = 24'(20620);
			15686: out = 24'(14588);
			15687: out = 24'(6212);
			15688: out = 24'(-14244);
			15689: out = 24'(4472);
			15690: out = 24'(25888);
			15691: out = 24'(12100);
			15692: out = 24'(-38340);
			15693: out = 24'(-24760);
			15694: out = 24'(33548);
			15695: out = 24'(37048);
			15696: out = 24'(18924);
			15697: out = 24'(632);
			15698: out = 24'(-2680);
			15699: out = 24'(-22940);
			15700: out = 24'(-18620);
			15701: out = 24'(-4880);
			15702: out = 24'(18372);
			15703: out = 24'(14092);
			15704: out = 24'(22476);
			15705: out = 24'(-17480);
			15706: out = 24'(-23328);
			15707: out = 24'(5652);
			15708: out = 24'(20428);
			15709: out = 24'(7064);
			15710: out = 24'(-7952);
			15711: out = 24'(-8292);
			15712: out = 24'(544);
			15713: out = 24'(10560);
			15714: out = 24'(18916);
			15715: out = 24'(23528);
			15716: out = 24'(29028);
			15717: out = 24'(2604);
			15718: out = 24'(-11620);
			15719: out = 24'(-33744);
			15720: out = 24'(-47796);
			15721: out = 24'(-9516);
			15722: out = 24'(44316);
			15723: out = 24'(44728);
			15724: out = 24'(1520);
			15725: out = 24'(788);
			15726: out = 24'(15876);
			15727: out = 24'(17536);
			15728: out = 24'(-22596);
			15729: out = 24'(-58156);
			15730: out = 24'(-38912);
			15731: out = 24'(21704);
			15732: out = 24'(47228);
			15733: out = 24'(27036);
			15734: out = 24'(-21640);
			15735: out = 24'(-20652);
			15736: out = 24'(12132);
			15737: out = 24'(20532);
			15738: out = 24'(-12940);
			15739: out = 24'(-30272);
			15740: out = 24'(-7532);
			15741: out = 24'(22156);
			15742: out = 24'(4352);
			15743: out = 24'(-7264);
			15744: out = 24'(-10244);
			15745: out = 24'(-3084);
			15746: out = 24'(7928);
			15747: out = 24'(-11404);
			15748: out = 24'(-37916);
			15749: out = 24'(-46076);
			15750: out = 24'(-548);
			15751: out = 24'(18556);
			15752: out = 24'(41064);
			15753: out = 24'(31100);
			15754: out = 24'(8392);
			15755: out = 24'(-29096);
			15756: out = 24'(-14256);
			15757: out = 24'(-15240);
			15758: out = 24'(-38760);
			15759: out = 24'(-13604);
			15760: out = 24'(39072);
			15761: out = 24'(50080);
			15762: out = 24'(18452);
			15763: out = 24'(704);
			15764: out = 24'(-7252);
			15765: out = 24'(-27612);
			15766: out = 24'(-42212);
			15767: out = 24'(-8960);
			15768: out = 24'(12180);
			15769: out = 24'(-1808);
			15770: out = 24'(-15876);
			15771: out = 24'(14092);
			15772: out = 24'(28256);
			15773: out = 24'(14828);
			15774: out = 24'(-4328);
			15775: out = 24'(4200);
			15776: out = 24'(23828);
			15777: out = 24'(-7336);
			15778: out = 24'(-39388);
			15779: out = 24'(-18432);
			15780: out = 24'(24968);
			15781: out = 24'(7872);
			15782: out = 24'(-27440);
			15783: out = 24'(-14384);
			15784: out = 24'(38352);
			15785: out = 24'(34884);
			15786: out = 24'(3412);
			15787: out = 24'(-7648);
			15788: out = 24'(3444);
			15789: out = 24'(25768);
			15790: out = 24'(-3600);
			15791: out = 24'(-26444);
			15792: out = 24'(-404);
			15793: out = 24'(28204);
			15794: out = 24'(20712);
			15795: out = 24'(580);
			15796: out = 24'(-1296);
			15797: out = 24'(-12536);
			15798: out = 24'(-4152);
			15799: out = 24'(1004);
			15800: out = 24'(2876);
			15801: out = 24'(-10832);
			15802: out = 24'(21832);
			15803: out = 24'(34840);
			15804: out = 24'(7836);
			15805: out = 24'(-41028);
			15806: out = 24'(-68192);
			15807: out = 24'(-41700);
			15808: out = 24'(7836);
			15809: out = 24'(30356);
			15810: out = 24'(38132);
			15811: out = 24'(21396);
			15812: out = 24'(-6824);
			15813: out = 24'(-30268);
			15814: out = 24'(-8532);
			15815: out = 24'(904);
			15816: out = 24'(-12996);
			15817: out = 24'(-34160);
			15818: out = 24'(492);
			15819: out = 24'(6508);
			15820: out = 24'(13872);
			15821: out = 24'(10460);
			15822: out = 24'(1036);
			15823: out = 24'(-13020);
			15824: out = 24'(-7968);
			15825: out = 24'(4588);
			15826: out = 24'(8516);
			15827: out = 24'(2500);
			15828: out = 24'(-6336);
			15829: out = 24'(-8768);
			15830: out = 24'(2224);
			15831: out = 24'(6648);
			15832: out = 24'(25720);
			15833: out = 24'(16068);
			15834: out = 24'(-21088);
			15835: out = 24'(-17316);
			15836: out = 24'(3000);
			15837: out = 24'(33124);
			15838: out = 24'(28108);
			15839: out = 24'(1468);
			15840: out = 24'(-21300);
			15841: out = 24'(-4668);
			15842: out = 24'(3532);
			15843: out = 24'(-21396);
			15844: out = 24'(-58584);
			15845: out = 24'(-23028);
			15846: out = 24'(37464);
			15847: out = 24'(38696);
			15848: out = 24'(17068);
			15849: out = 24'(2860);
			15850: out = 24'(19972);
			15851: out = 24'(24004);
			15852: out = 24'(3132);
			15853: out = 24'(-33224);
			15854: out = 24'(-28308);
			15855: out = 24'(6820);
			15856: out = 24'(15000);
			15857: out = 24'(24836);
			15858: out = 24'(19596);
			15859: out = 24'(7768);
			15860: out = 24'(-1544);
			15861: out = 24'(-18268);
			15862: out = 24'(-27544);
			15863: out = 24'(-34256);
			15864: out = 24'(-32980);
			15865: out = 24'(-16460);
			15866: out = 24'(21540);
			15867: out = 24'(38124);
			15868: out = 24'(21824);
			15869: out = 24'(10664);
			15870: out = 24'(1660);
			15871: out = 24'(-12988);
			15872: out = 24'(-30804);
			15873: out = 24'(-876);
			15874: out = 24'(-1024);
			15875: out = 24'(4184);
			15876: out = 24'(10636);
			15877: out = 24'(16920);
			15878: out = 24'(2920);
			15879: out = 24'(-4704);
			15880: out = 24'(-9980);
			15881: out = 24'(-22372);
			15882: out = 24'(-24916);
			15883: out = 24'(-13636);
			15884: out = 24'(13480);
			15885: out = 24'(28396);
			15886: out = 24'(24860);
			15887: out = 24'(4780);
			15888: out = 24'(-252);
			15889: out = 24'(-7228);
			15890: out = 24'(-36076);
			15891: out = 24'(-77540);
			15892: out = 24'(-56092);
			15893: out = 24'(19600);
			15894: out = 24'(48880);
			15895: out = 24'(37236);
			15896: out = 24'(11440);
			15897: out = 24'(8112);
			15898: out = 24'(14164);
			15899: out = 24'(-41164);
			15900: out = 24'(-73224);
			15901: out = 24'(-47156);
			15902: out = 24'(10592);
			15903: out = 24'(40240);
			15904: out = 24'(35796);
			15905: out = 24'(17932);
			15906: out = 24'(2944);
			15907: out = 24'(28);
			15908: out = 24'(2856);
			15909: out = 24'(5128);
			15910: out = 24'(-7824);
			15911: out = 24'(-48404);
			15912: out = 24'(-24216);
			15913: out = 24'(12500);
			15914: out = 24'(19196);
			15915: out = 24'(3448);
			15916: out = 24'(20224);
			15917: out = 24'(30888);
			15918: out = 24'(3912);
			15919: out = 24'(-31920);
			15920: out = 24'(-19000);
			15921: out = 24'(37228);
			15922: out = 24'(42148);
			15923: out = 24'(-7116);
			15924: out = 24'(-28216);
			15925: out = 24'(-1380);
			15926: out = 24'(4920);
			15927: out = 24'(-30764);
			15928: out = 24'(-11396);
			15929: out = 24'(-6672);
			15930: out = 24'(6908);
			15931: out = 24'(17048);
			15932: out = 24'(54376);
			15933: out = 24'(35968);
			15934: out = 24'(12512);
			15935: out = 24'(-29148);
			15936: out = 24'(-54816);
			15937: out = 24'(-40184);
			15938: out = 24'(7752);
			15939: out = 24'(27608);
			15940: out = 24'(16284);
			15941: out = 24'(4492);
			15942: out = 24'(13644);
			15943: out = 24'(12140);
			15944: out = 24'(-96);
			15945: out = 24'(17128);
			15946: out = 24'(23664);
			15947: out = 24'(14884);
			15948: out = 24'(-8188);
			15949: out = 24'(-9764);
			15950: out = 24'(-21940);
			15951: out = 24'(-3664);
			15952: out = 24'(30588);
			15953: out = 24'(50868);
			15954: out = 24'(17156);
			15955: out = 24'(-35800);
			15956: out = 24'(-75020);
			15957: out = 24'(-66092);
			15958: out = 24'(-47544);
			15959: out = 24'(-5792);
			15960: out = 24'(20256);
			15961: out = 24'(27004);
			15962: out = 24'(18856);
			15963: out = 24'(18784);
			15964: out = 24'(12948);
			15965: out = 24'(-3836);
			15966: out = 24'(-34272);
			15967: out = 24'(-40892);
			15968: out = 24'(-20560);
			15969: out = 24'(23080);
			15970: out = 24'(45124);
			15971: out = 24'(22596);
			15972: out = 24'(-37948);
			15973: out = 24'(-62432);
			15974: out = 24'(-11752);
			15975: out = 24'(14656);
			15976: out = 24'(3424);
			15977: out = 24'(-17260);
			15978: out = 24'(6284);
			15979: out = 24'(28628);
			15980: out = 24'(26620);
			15981: out = 24'(-20384);
			15982: out = 24'(-41536);
			15983: out = 24'(7068);
			15984: out = 24'(36416);
			15985: out = 24'(1072);
			15986: out = 24'(-41080);
			15987: out = 24'(-9092);
			15988: out = 24'(19756);
			15989: out = 24'(27480);
			15990: out = 24'(16404);
			15991: out = 24'(19820);
			15992: out = 24'(-2548);
			15993: out = 24'(-8408);
			15994: out = 24'(-6576);
			15995: out = 24'(2300);
			15996: out = 24'(196);
			15997: out = 24'(148);
			15998: out = 24'(9392);
			15999: out = 24'(23404);
			16000: out = 24'(8732);
			16001: out = 24'(13224);
			16002: out = 24'(8644);
			16003: out = 24'(-7460);
			16004: out = 24'(-33776);
			16005: out = 24'(-17352);
			16006: out = 24'(1784);
			16007: out = 24'(2780);
			16008: out = 24'(-3160);
			16009: out = 24'(-7108);
			16010: out = 24'(22152);
			16011: out = 24'(36728);
			16012: out = 24'(11964);
			16013: out = 24'(-14372);
			16014: out = 24'(-17500);
			16015: out = 24'(-3052);
			16016: out = 24'(244);
			16017: out = 24'(11076);
			16018: out = 24'(1408);
			16019: out = 24'(-332);
			16020: out = 24'(-1544);
			16021: out = 24'(836);
			16022: out = 24'(5508);
			16023: out = 24'(13296);
			16024: out = 24'(-4936);
			16025: out = 24'(-48200);
			16026: out = 24'(-5052);
			16027: out = 24'(46540);
			16028: out = 24'(48828);
			16029: out = 24'(4168);
			16030: out = 24'(-8488);
			16031: out = 24'(-5592);
			16032: out = 24'(-2452);
			16033: out = 24'(-10344);
			16034: out = 24'(7788);
			16035: out = 24'(21024);
			16036: out = 24'(20020);
			16037: out = 24'(7648);
			16038: out = 24'(25532);
			16039: out = 24'(4620);
			16040: out = 24'(-17816);
			16041: out = 24'(-31476);
			16042: out = 24'(-9656);
			16043: out = 24'(-20784);
			16044: out = 24'(-10064);
			16045: out = 24'(6196);
			16046: out = 24'(17768);
			16047: out = 24'(13528);
			16048: out = 24'(10456);
			16049: out = 24'(4928);
			16050: out = 24'(-3800);
			16051: out = 24'(-28744);
			16052: out = 24'(-32804);
			16053: out = 24'(-23596);
			16054: out = 24'(-6180);
			16055: out = 24'(-1236);
			16056: out = 24'(9776);
			16057: out = 24'(2004);
			16058: out = 24'(2480);
			16059: out = 24'(40392);
			16060: out = 24'(11292);
			16061: out = 24'(-30092);
			16062: out = 24'(-45572);
			16063: out = 24'(4620);
			16064: out = 24'(19904);
			16065: out = 24'(32792);
			16066: out = 24'(18876);
			16067: out = 24'(-3696);
			16068: out = 24'(-20336);
			16069: out = 24'(-20420);
			16070: out = 24'(-26560);
			16071: out = 24'(-32980);
			16072: out = 24'(-11228);
			16073: out = 24'(17488);
			16074: out = 24'(27556);
			16075: out = 24'(12632);
			16076: out = 24'(2644);
			16077: out = 24'(-9660);
			16078: out = 24'(-5260);
			16079: out = 24'(120);
			16080: out = 24'(1156);
			16081: out = 24'(-1124);
			16082: out = 24'(5644);
			16083: out = 24'(10144);
			16084: out = 24'(8424);
			16085: out = 24'(-8500);
			16086: out = 24'(3016);
			16087: out = 24'(21584);
			16088: out = 24'(20196);
			16089: out = 24'(-21124);
			16090: out = 24'(-35192);
			16091: out = 24'(-22600);
			16092: out = 24'(6988);
			16093: out = 24'(15776);
			16094: out = 24'(33380);
			16095: out = 24'(21652);
			16096: out = 24'(8832);
			16097: out = 24'(16296);
			16098: out = 24'(3604);
			16099: out = 24'(-20800);
			16100: out = 24'(-21396);
			16101: out = 24'(19348);
			16102: out = 24'(192);
			16103: out = 24'(-6116);
			16104: out = 24'(3032);
			16105: out = 24'(27104);
			16106: out = 24'(11500);
			16107: out = 24'(10308);
			16108: out = 24'(-100);
			16109: out = 24'(-17980);
			16110: out = 24'(-49760);
			16111: out = 24'(552);
			16112: out = 24'(43908);
			16113: out = 24'(25720);
			16114: out = 24'(-27420);
			16115: out = 24'(-37728);
			16116: out = 24'(-1840);
			16117: out = 24'(9080);
			16118: out = 24'(-25020);
			16119: out = 24'(-20592);
			16120: out = 24'(31564);
			16121: out = 24'(54600);
			16122: out = 24'(11296);
			16123: out = 24'(-10360);
			16124: out = 24'(-4792);
			16125: out = 24'(8456);
			16126: out = 24'(-14480);
			16127: out = 24'(-15740);
			16128: out = 24'(-26512);
			16129: out = 24'(-1484);
			16130: out = 24'(19660);
			16131: out = 24'(32952);
			16132: out = 24'(-14940);
			16133: out = 24'(-18756);
			16134: out = 24'(6172);
			16135: out = 24'(12836);
			16136: out = 24'(-28996);
			16137: out = 24'(-52848);
			16138: out = 24'(-36548);
			16139: out = 24'(4712);
			16140: out = 24'(15160);
			16141: out = 24'(18164);
			16142: out = 24'(6524);
			16143: out = 24'(2800);
			16144: out = 24'(5660);
			16145: out = 24'(19784);
			16146: out = 24'(-9000);
			16147: out = 24'(-44352);
			16148: out = 24'(-5348);
			16149: out = 24'(8252);
			16150: out = 24'(-7788);
			16151: out = 24'(-27456);
			16152: out = 24'(7804);
			16153: out = 24'(8268);
			16154: out = 24'(-816);
			16155: out = 24'(-14840);
			16156: out = 24'(6868);
			16157: out = 24'(12248);
			16158: out = 24'(30616);
			16159: out = 24'(16864);
			16160: out = 24'(-6408);
			16161: out = 24'(-11564);
			16162: out = 24'(10004);
			16163: out = 24'(14120);
			16164: out = 24'(-252);
			16165: out = 24'(-9900);
			16166: out = 24'(-10348);
			16167: out = 24'(-9652);
			16168: out = 24'(2128);
			16169: out = 24'(24588);
			16170: out = 24'(33836);
			16171: out = 24'(15448);
			16172: out = 24'(4768);
			16173: out = 24'(19344);
			16174: out = 24'(-5324);
			16175: out = 24'(-41372);
			16176: out = 24'(-45956);
			16177: out = 24'(9852);
			16178: out = 24'(33648);
			16179: out = 24'(24784);
			16180: out = 24'(-8012);
			16181: out = 24'(-9600);
			16182: out = 24'(2848);
			16183: out = 24'(26188);
			16184: out = 24'(-1368);
			16185: out = 24'(-30296);
			16186: out = 24'(-960);
			16187: out = 24'(32080);
			16188: out = 24'(22332);
			16189: out = 24'(-13916);
			16190: out = 24'(-16252);
			16191: out = 24'(10080);
			16192: out = 24'(30908);
			16193: out = 24'(13600);
			16194: out = 24'(-12912);
			16195: out = 24'(-27584);
			16196: out = 24'(-3908);
			16197: out = 24'(4696);
			16198: out = 24'(-19424);
			16199: out = 24'(-58112);
			16200: out = 24'(-12748);
			16201: out = 24'(45352);
			16202: out = 24'(37672);
			16203: out = 24'(-25652);
			16204: out = 24'(-37744);
			16205: out = 24'(2060);
			16206: out = 24'(26680);
			16207: out = 24'(-3860);
			16208: out = 24'(-25984);
			16209: out = 24'(-14860);
			16210: out = 24'(10344);
			16211: out = 24'(5360);
			16212: out = 24'(-1632);
			16213: out = 24'(-11456);
			16214: out = 24'(-5592);
			16215: out = 24'(444);
			16216: out = 24'(5324);
			16217: out = 24'(9232);
			16218: out = 24'(17068);
			16219: out = 24'(11584);
			16220: out = 24'(-8820);
			16221: out = 24'(-35024);
			16222: out = 24'(-27468);
			16223: out = 24'(2776);
			16224: out = 24'(6992);
			16225: out = 24'(15336);
			16226: out = 24'(4668);
			16227: out = 24'(-1196);
			16228: out = 24'(-712);
			16229: out = 24'(16240);
			16230: out = 24'(7128);
			16231: out = 24'(-2228);
			16232: out = 24'(-672);
			16233: out = 24'(-556);
			16234: out = 24'(4968);
			16235: out = 24'(9880);
			16236: out = 24'(7488);
			16237: out = 24'(17832);
			16238: out = 24'(1328);
			16239: out = 24'(-1624);
			16240: out = 24'(-404);
			16241: out = 24'(13376);
			16242: out = 24'(-36328);
			16243: out = 24'(-32508);
			16244: out = 24'(340);
			16245: out = 24'(15568);
			16246: out = 24'(-31880);
			16247: out = 24'(-11760);
			16248: out = 24'(33620);
			16249: out = 24'(34052);
			16250: out = 24'(5408);
			16251: out = 24'(-11472);
			16252: out = 24'(-5624);
			16253: out = 24'(-1856);
			16254: out = 24'(-14072);
			16255: out = 24'(-6272);
			16256: out = 24'(4552);
			16257: out = 24'(12076);
			16258: out = 24'(24232);
			16259: out = 24'(17344);
			16260: out = 24'(-12996);
			16261: out = 24'(-46568);
			16262: out = 24'(-35484);
			16263: out = 24'(-10988);
			16264: out = 24'(19592);
			16265: out = 24'(23328);
			16266: out = 24'(17200);
			16267: out = 24'(232);
			16268: out = 24'(916);
			16269: out = 24'(-4680);
			16270: out = 24'(-11728);
			16271: out = 24'(-39976);
			16272: out = 24'(-8624);
			16273: out = 24'(6776);
			16274: out = 24'(1848);
			16275: out = 24'(17800);
			16276: out = 24'(33072);
			16277: out = 24'(25660);
			16278: out = 24'(-320);
			16279: out = 24'(-19704);
			16280: out = 24'(-16204);
			16281: out = 24'(-23084);
			16282: out = 24'(-22420);
			16283: out = 24'(13868);
			16284: out = 24'(28560);
			16285: out = 24'(26876);
			16286: out = 24'(7652);
			16287: out = 24'(-400);
			16288: out = 24'(-2288);
			16289: out = 24'(1192);
			16290: out = 24'(-7000);
			16291: out = 24'(-16424);
			16292: out = 24'(-20264);
			16293: out = 24'(-9536);
			16294: out = 24'(-2552);
			16295: out = 24'(312);
			16296: out = 24'(4136);
			16297: out = 24'(21616);
			16298: out = 24'(17432);
			16299: out = 24'(-4948);
			16300: out = 24'(-12676);
			16301: out = 24'(-13804);
			16302: out = 24'(3188);
			16303: out = 24'(9108);
			16304: out = 24'(9660);
			16305: out = 24'(-1380);
			16306: out = 24'(12856);
			16307: out = 24'(8520);
			16308: out = 24'(-16312);
			16309: out = 24'(-48732);
			16310: out = 24'(-24200);
			16311: out = 24'(-1680);
			16312: out = 24'(-56);
			16313: out = 24'(1772);
			16314: out = 24'(35168);
			16315: out = 24'(29592);
			16316: out = 24'(-20012);
			16317: out = 24'(-62548);
			16318: out = 24'(-41668);
			16319: out = 24'(2852);
			16320: out = 24'(20180);
			16321: out = 24'(15992);
			16322: out = 24'(31532);
			16323: out = 24'(31356);
			16324: out = 24'(18584);
			16325: out = 24'(8148);
			16326: out = 24'(-1128);
			16327: out = 24'(-9920);
			16328: out = 24'(-16828);
			16329: out = 24'(-3776);
			16330: out = 24'(13500);
			16331: out = 24'(15708);
			16332: out = 24'(-12688);
			16333: out = 24'(-25212);
			16334: out = 24'(2464);
			16335: out = 24'(14912);
			16336: out = 24'(-9872);
			16337: out = 24'(-29840);
			16338: out = 24'(-12004);
			16339: out = 24'(14916);
			16340: out = 24'(7752);
			16341: out = 24'(10764);
			16342: out = 24'(44696);
			16343: out = 24'(48936);
			16344: out = 24'(32);
			16345: out = 24'(-46340);
			16346: out = 24'(-28556);
			16347: out = 24'(10148);
			16348: out = 24'(28572);
			16349: out = 24'(11972);
			16350: out = 24'(9212);
			16351: out = 24'(29152);
			16352: out = 24'(22436);
			16353: out = 24'(-12848);
			16354: out = 24'(-39932);
			16355: out = 24'(-29392);
			16356: out = 24'(-7068);
			16357: out = 24'(-4628);
			16358: out = 24'(-11028);
			16359: out = 24'(4336);
			16360: out = 24'(16292);
			16361: out = 24'(29440);
			16362: out = 24'(19580);
			16363: out = 24'(5144);
			16364: out = 24'(-12560);
			16365: out = 24'(-816);
			16366: out = 24'(-10556);
			16367: out = 24'(-38124);
			16368: out = 24'(-49000);
			16369: out = 24'(4172);
			16370: out = 24'(50852);
			16371: out = 24'(49020);
			16372: out = 24'(13136);
			16373: out = 24'(-23020);
			16374: out = 24'(-46068);
			16375: out = 24'(-54428);
			16376: out = 24'(-53744);
			16377: out = 24'(-6820);
			16378: out = 24'(14080);
			16379: out = 24'(20316);
			16380: out = 24'(14072);
			16381: out = 24'(-10524);
			16382: out = 24'(-30536);
			16383: out = 24'(-20944);
			16384: out = 24'(5544);
			16385: out = 24'(12);
			16386: out = 24'(2848);
			16387: out = 24'(4300);
			16388: out = 24'(15744);
			16389: out = 24'(25088);
			16390: out = 24'(14496);
			16391: out = 24'(-2592);
			16392: out = 24'(-9648);
			16393: out = 24'(-5820);
			16394: out = 24'(-26164);
			16395: out = 24'(-14916);
			16396: out = 24'(14188);
			16397: out = 24'(22740);
			16398: out = 24'(-100);
			16399: out = 24'(-6348);
			16400: out = 24'(12396);
			16401: out = 24'(17784);
			16402: out = 24'(3856);
			16403: out = 24'(-25656);
			16404: out = 24'(-14460);
			16405: out = 24'(3836);
			16406: out = 24'(-8264);
			16407: out = 24'(-5648);
			16408: out = 24'(32532);
			16409: out = 24'(49844);
			16410: out = 24'(11716);
			16411: out = 24'(-31724);
			16412: out = 24'(-21832);
			16413: out = 24'(9828);
			16414: out = 24'(2556);
			16415: out = 24'(-33088);
			16416: out = 24'(-16624);
			16417: out = 24'(26904);
			16418: out = 24'(34596);
			16419: out = 24'(3680);
			16420: out = 24'(8872);
			16421: out = 24'(22304);
			16422: out = 24'(3160);
			16423: out = 24'(-42512);
			16424: out = 24'(-42876);
			16425: out = 24'(-5256);
			16426: out = 24'(21432);
			16427: out = 24'(16888);
			16428: out = 24'(10048);
			16429: out = 24'(14316);
			16430: out = 24'(9616);
			16431: out = 24'(-18520);
			16432: out = 24'(-22372);
			16433: out = 24'(-9300);
			16434: out = 24'(22320);
			16435: out = 24'(38988);
			16436: out = 24'(26620);
			16437: out = 24'(4996);
			16438: out = 24'(-1624);
			16439: out = 24'(4136);
			16440: out = 24'(-2316);
			16441: out = 24'(-14784);
			16442: out = 24'(-24440);
			16443: out = 24'(-10952);
			16444: out = 24'(14664);
			16445: out = 24'(-27280);
			16446: out = 24'(-41292);
			16447: out = 24'(3608);
			16448: out = 24'(51436);
			16449: out = 24'(25804);
			16450: out = 24'(-31260);
			16451: out = 24'(-52644);
			16452: out = 24'(-18364);
			16453: out = 24'(-2692);
			16454: out = 24'(6952);
			16455: out = 24'(23100);
			16456: out = 24'(41576);
			16457: out = 24'(28848);
			16458: out = 24'(-12);
			16459: out = 24'(-13960);
			16460: out = 24'(-11412);
			16461: out = 24'(-26120);
			16462: out = 24'(-39876);
			16463: out = 24'(-35092);
			16464: out = 24'(-1724);
			16465: out = 24'(31476);
			16466: out = 24'(31652);
			16467: out = 24'(16384);
			16468: out = 24'(-6116);
			16469: out = 24'(-19088);
			16470: out = 24'(-30280);
			16471: out = 24'(-2496);
			16472: out = 24'(11868);
			16473: out = 24'(500);
			16474: out = 24'(-22116);
			16475: out = 24'(12172);
			16476: out = 24'(28908);
			16477: out = 24'(11664);
			16478: out = 24'(2880);
			16479: out = 24'(-660);
			16480: out = 24'(-6724);
			16481: out = 24'(-23584);
			16482: out = 24'(-13980);
			16483: out = 24'(5008);
			16484: out = 24'(37668);
			16485: out = 24'(32348);
			16486: out = 24'(-4704);
			16487: out = 24'(-26964);
			16488: out = 24'(-16172);
			16489: out = 24'(408);
			16490: out = 24'(-332);
			16491: out = 24'(1632);
			16492: out = 24'(-3040);
			16493: out = 24'(-6892);
			16494: out = 24'(-8684);
			16495: out = 24'(-3968);
			16496: out = 24'(24564);
			16497: out = 24'(37780);
			16498: out = 24'(26000);
			16499: out = 24'(8252);
			16500: out = 24'(-35476);
			16501: out = 24'(-40212);
			16502: out = 24'(-6512);
			16503: out = 24'(24780);
			16504: out = 24'(5764);
			16505: out = 24'(-1436);
			16506: out = 24'(22288);
			16507: out = 24'(41232);
			16508: out = 24'(-22628);
			16509: out = 24'(-56388);
			16510: out = 24'(-43168);
			16511: out = 24'(3996);
			16512: out = 24'(7552);
			16513: out = 24'(35036);
			16514: out = 24'(42972);
			16515: out = 24'(33744);
			16516: out = 24'(6544);
			16517: out = 24'(-21408);
			16518: out = 24'(-43064);
			16519: out = 24'(-35388);
			16520: out = 24'(4736);
			16521: out = 24'(34296);
			16522: out = 24'(40080);
			16523: out = 24'(20556);
			16524: out = 24'(16);
			16525: out = 24'(-33640);
			16526: out = 24'(-20684);
			16527: out = 24'(-4764);
			16528: out = 24'(332);
			16529: out = 24'(-6264);
			16530: out = 24'(14928);
			16531: out = 24'(16476);
			16532: out = 24'(-7388);
			16533: out = 24'(-49476);
			16534: out = 24'(-13344);
			16535: out = 24'(9000);
			16536: out = 24'(7160);
			16537: out = 24'(296);
			16538: out = 24'(5616);
			16539: out = 24'(-8800);
			16540: out = 24'(-19156);
			16541: out = 24'(-5748);
			16542: out = 24'(22836);
			16543: out = 24'(17244);
			16544: out = 24'(6912);
			16545: out = 24'(8364);
			16546: out = 24'(-4976);
			16547: out = 24'(-16568);
			16548: out = 24'(-13696);
			16549: out = 24'(1836);
			16550: out = 24'(-1712);
			16551: out = 24'(684);
			16552: out = 24'(2040);
			16553: out = 24'(3580);
			16554: out = 24'(448);
			16555: out = 24'(-4860);
			16556: out = 24'(-2304);
			16557: out = 24'(-4100);
			16558: out = 24'(-14224);
			16559: out = 24'(-11364);
			16560: out = 24'(13008);
			16561: out = 24'(29844);
			16562: out = 24'(21412);
			16563: out = 24'(-2752);
			16564: out = 24'(-3212);
			16565: out = 24'(-452);
			16566: out = 24'(-8816);
			16567: out = 24'(-18288);
			16568: out = 24'(84);
			16569: out = 24'(20428);
			16570: out = 24'(21072);
			16571: out = 24'(-696);
			16572: out = 24'(260);
			16573: out = 24'(-3608);
			16574: out = 24'(-4132);
			16575: out = 24'(3984);
			16576: out = 24'(19308);
			16577: out = 24'(8964);
			16578: out = 24'(-3888);
			16579: out = 24'(1048);
			16580: out = 24'(6220);
			16581: out = 24'(-2716);
			16582: out = 24'(-15540);
			16583: out = 24'(-3856);
			16584: out = 24'(21028);
			16585: out = 24'(39048);
			16586: out = 24'(21036);
			16587: out = 24'(-8616);
			16588: out = 24'(-10564);
			16589: out = 24'(-1568);
			16590: out = 24'(2648);
			16591: out = 24'(-4088);
			16592: out = 24'(-172);
			16593: out = 24'(6876);
			16594: out = 24'(18048);
			16595: out = 24'(-1896);
			16596: out = 24'(-41524);
			16597: out = 24'(-12312);
			16598: out = 24'(25004);
			16599: out = 24'(29776);
			16600: out = 24'(-10892);
			16601: out = 24'(-16220);
			16602: out = 24'(-13724);
			16603: out = 24'(12932);
			16604: out = 24'(4392);
			16605: out = 24'(-25144);
			16606: out = 24'(-36780);
			16607: out = 24'(16224);
			16608: out = 24'(40016);
			16609: out = 24'(6436);
			16610: out = 24'(-77436);
			16611: out = 24'(-41020);
			16612: out = 24'(41172);
			16613: out = 24'(39976);
			16614: out = 24'(-35844);
			16615: out = 24'(-34952);
			16616: out = 24'(18152);
			16617: out = 24'(22236);
			16618: out = 24'(-30940);
			16619: out = 24'(-44564);
			16620: out = 24'(-12708);
			16621: out = 24'(10500);
			16622: out = 24'(10660);
			16623: out = 24'(1724);
			16624: out = 24'(2392);
			16625: out = 24'(4716);
			16626: out = 24'(9244);
			16627: out = 24'(-10076);
			16628: out = 24'(-21328);
			16629: out = 24'(-21752);
			16630: out = 24'(-7336);
			16631: out = 24'(-10312);
			16632: out = 24'(7880);
			16633: out = 24'(28380);
			16634: out = 24'(40196);
			16635: out = 24'(14452);
			16636: out = 24'(16416);
			16637: out = 24'(11104);
			16638: out = 24'(-9740);
			16639: out = 24'(-59428);
			16640: out = 24'(-13628);
			16641: out = 24'(27444);
			16642: out = 24'(20168);
			16643: out = 24'(-12876);
			16644: out = 24'(-9564);
			16645: out = 24'(2164);
			16646: out = 24'(3272);
			16647: out = 24'(-624);
			16648: out = 24'(-13744);
			16649: out = 24'(2820);
			16650: out = 24'(22752);
			16651: out = 24'(10452);
			16652: out = 24'(-21084);
			16653: out = 24'(-44140);
			16654: out = 24'(-8656);
			16655: out = 24'(47364);
			16656: out = 24'(45840);
			16657: out = 24'(14624);
			16658: out = 24'(-16784);
			16659: out = 24'(-23468);
			16660: out = 24'(-10572);
			16661: out = 24'(688);
			16662: out = 24'(12536);
			16663: out = 24'(14648);
			16664: out = 24'(4024);
			16665: out = 24'(3096);
			16666: out = 24'(3076);
			16667: out = 24'(-11456);
			16668: out = 24'(-30428);
			16669: out = 24'(-46464);
			16670: out = 24'(8120);
			16671: out = 24'(55648);
			16672: out = 24'(45464);
			16673: out = 24'(7968);
			16674: out = 24'(-92);
			16675: out = 24'(4624);
			16676: out = 24'(-7744);
			16677: out = 24'(-27816);
			16678: out = 24'(-12136);
			16679: out = 24'(20300);
			16680: out = 24'(24636);
			16681: out = 24'(-11564);
			16682: out = 24'(272);
			16683: out = 24'(7256);
			16684: out = 24'(4760);
			16685: out = 24'(-456);
			16686: out = 24'(27144);
			16687: out = 24'(20516);
			16688: out = 24'(-10636);
			16689: out = 24'(-38876);
			16690: out = 24'(-57564);
			16691: out = 24'(-22052);
			16692: out = 24'(18308);
			16693: out = 24'(30092);
			16694: out = 24'(4700);
			16695: out = 24'(1264);
			16696: out = 24'(-5360);
			16697: out = 24'(-11684);
			16698: out = 24'(-15452);
			16699: out = 24'(-1428);
			16700: out = 24'(-9344);
			16701: out = 24'(-17776);
			16702: out = 24'(1684);
			16703: out = 24'(-236);
			16704: out = 24'(3368);
			16705: out = 24'(9044);
			16706: out = 24'(16356);
			16707: out = 24'(-12300);
			16708: out = 24'(-15608);
			16709: out = 24'(-16928);
			16710: out = 24'(-25892);
			16711: out = 24'(-21492);
			16712: out = 24'(-9036);
			16713: out = 24'(23912);
			16714: out = 24'(37436);
			16715: out = 24'(9792);
			16716: out = 24'(-44712);
			16717: out = 24'(-57456);
			16718: out = 24'(-25116);
			16719: out = 24'(-2968);
			16720: out = 24'(37896);
			16721: out = 24'(38768);
			16722: out = 24'(23472);
			16723: out = 24'(9328);
			16724: out = 24'(1832);
			16725: out = 24'(-9872);
			16726: out = 24'(-25660);
			16727: out = 24'(-23172);
			16728: out = 24'(-2452);
			16729: out = 24'(23728);
			16730: out = 24'(16800);
			16731: out = 24'(1792);
			16732: out = 24'(9128);
			16733: out = 24'(25316);
			16734: out = 24'(6484);
			16735: out = 24'(-27752);
			16736: out = 24'(-42484);
			16737: out = 24'(-7032);
			16738: out = 24'(4540);
			16739: out = 24'(4672);
			16740: out = 24'(15564);
			16741: out = 24'(19720);
			16742: out = 24'(6264);
			16743: out = 24'(5552);
			16744: out = 24'(16892);
			16745: out = 24'(4264);
			16746: out = 24'(-28432);
			16747: out = 24'(-23584);
			16748: out = 24'(16512);
			16749: out = 24'(16816);
			16750: out = 24'(5828);
			16751: out = 24'(6996);
			16752: out = 24'(17892);
			16753: out = 24'(2204);
			16754: out = 24'(-29572);
			16755: out = 24'(-38992);
			16756: out = 24'(-17636);
			16757: out = 24'(13968);
			16758: out = 24'(41268);
			16759: out = 24'(54448);
			16760: out = 24'(20940);
			16761: out = 24'(-36308);
			16762: out = 24'(-33684);
			16763: out = 24'(16312);
			16764: out = 24'(26840);
			16765: out = 24'(-20884);
			16766: out = 24'(-50496);
			16767: out = 24'(-2700);
			16768: out = 24'(42728);
			16769: out = 24'(25980);
			16770: out = 24'(5104);
			16771: out = 24'(2168);
			16772: out = 24'(14664);
			16773: out = 24'(-6912);
			16774: out = 24'(-47860);
			16775: out = 24'(-42580);
			16776: out = 24'(2368);
			16777: out = 24'(30984);
			16778: out = 24'(23480);
			16779: out = 24'(7624);
			16780: out = 24'(1252);
			16781: out = 24'(-3040);
			16782: out = 24'(-10424);
			16783: out = 24'(-9824);
			16784: out = 24'(-2376);
			16785: out = 24'(1260);
			16786: out = 24'(-2412);
			16787: out = 24'(-13992);
			16788: out = 24'(-3592);
			16789: out = 24'(3840);
			16790: out = 24'(18328);
			16791: out = 24'(44872);
			16792: out = 24'(24436);
			16793: out = 24'(-15224);
			16794: out = 24'(-42412);
			16795: out = 24'(-25032);
			16796: out = 24'(-4884);
			16797: out = 24'(6332);
			16798: out = 24'(-1444);
			16799: out = 24'(-8324);
			16800: out = 24'(-1568);
			16801: out = 24'(7700);
			16802: out = 24'(3848);
			16803: out = 24'(-14336);
			16804: out = 24'(-25268);
			16805: out = 24'(4852);
			16806: out = 24'(42428);
			16807: out = 24'(30736);
			16808: out = 24'(-26088);
			16809: out = 24'(-30700);
			16810: out = 24'(6572);
			16811: out = 24'(17636);
			16812: out = 24'(-20516);
			16813: out = 24'(-37648);
			16814: out = 24'(4976);
			16815: out = 24'(47012);
			16816: out = 24'(31332);
			16817: out = 24'(-11476);
			16818: out = 24'(-11580);
			16819: out = 24'(10224);
			16820: out = 24'(9248);
			16821: out = 24'(1896);
			16822: out = 24'(-9720);
			16823: out = 24'(-5308);
			16824: out = 24'(-2516);
			16825: out = 24'(-13708);
			16826: out = 24'(496);
			16827: out = 24'(12796);
			16828: out = 24'(18336);
			16829: out = 24'(15092);
			16830: out = 24'(-11812);
			16831: out = 24'(-24112);
			16832: out = 24'(-3680);
			16833: out = 24'(25460);
			16834: out = 24'(19732);
			16835: out = 24'(-10300);
			16836: out = 24'(-20520);
			16837: out = 24'(6244);
			16838: out = 24'(21780);
			16839: out = 24'(18824);
			16840: out = 24'(4468);
			16841: out = 24'(-3380);
			16842: out = 24'(-15780);
			16843: out = 24'(-3372);
			16844: out = 24'(2064);
			16845: out = 24'(2528);
			16846: out = 24'(-1220);
			16847: out = 24'(-12084);
			16848: out = 24'(-10512);
			16849: out = 24'(10728);
			16850: out = 24'(30740);
			16851: out = 24'(19088);
			16852: out = 24'(-2544);
			16853: out = 24'(-7680);
			16854: out = 24'(11232);
			16855: out = 24'(13168);
			16856: out = 24'(17196);
			16857: out = 24'(7592);
			16858: out = 24'(-6708);
			16859: out = 24'(-30872);
			16860: out = 24'(-27456);
			16861: out = 24'(-23520);
			16862: out = 24'(-16432);
			16863: out = 24'(-4520);
			16864: out = 24'(37772);
			16865: out = 24'(34800);
			16866: out = 24'(-1968);
			16867: out = 24'(-32304);
			16868: out = 24'(-3960);
			16869: out = 24'(-472);
			16870: out = 24'(-21704);
			16871: out = 24'(-22692);
			16872: out = 24'(9976);
			16873: out = 24'(23660);
			16874: out = 24'(-4984);
			16875: out = 24'(-25808);
			16876: out = 24'(-4388);
			16877: out = 24'(28900);
			16878: out = 24'(11724);
			16879: out = 24'(-20800);
			16880: out = 24'(-33384);
			16881: out = 24'(9772);
			16882: out = 24'(3504);
			16883: out = 24'(-16108);
			16884: out = 24'(-7400);
			16885: out = 24'(22904);
			16886: out = 24'(10340);
			16887: out = 24'(4668);
			16888: out = 24'(13468);
			16889: out = 24'(-11508);
			16890: out = 24'(-49172);
			16891: out = 24'(-22204);
			16892: out = 24'(36036);
			16893: out = 24'(19980);
			16894: out = 24'(-33244);
			16895: out = 24'(-18476);
			16896: out = 24'(41176);
			16897: out = 24'(21376);
			16898: out = 24'(-30688);
			16899: out = 24'(-33272);
			16900: out = 24'(16124);
			16901: out = 24'(21092);
			16902: out = 24'(6972);
			16903: out = 24'(11324);
			16904: out = 24'(24020);
			16905: out = 24'(-7512);
			16906: out = 24'(-35432);
			16907: out = 24'(-34596);
			16908: out = 24'(-5248);
			16909: out = 24'(916);
			16910: out = 24'(28236);
			16911: out = 24'(14716);
			16912: out = 24'(19348);
			16913: out = 24'(23460);
			16914: out = 24'(17644);
			16915: out = 24'(4880);
			16916: out = 24'(1864);
			16917: out = 24'(-10700);
			16918: out = 24'(-42552);
			16919: out = 24'(-11768);
			16920: out = 24'(18852);
			16921: out = 24'(16236);
			16922: out = 24'(-8820);
			16923: out = 24'(11816);
			16924: out = 24'(29920);
			16925: out = 24'(15432);
			16926: out = 24'(-21908);
			16927: out = 24'(-2796);
			16928: out = 24'(6260);
			16929: out = 24'(-1588);
			16930: out = 24'(-20356);
			16931: out = 24'(716);
			16932: out = 24'(10968);
			16933: out = 24'(18924);
			16934: out = 24'(12844);
			16935: out = 24'(7620);
			16936: out = 24'(-33204);
			16937: out = 24'(-52896);
			16938: out = 24'(-34960);
			16939: out = 24'(12104);
			16940: out = 24'(22548);
			16941: out = 24'(26764);
			16942: out = 24'(19440);
			16943: out = 24'(5268);
			16944: out = 24'(-16352);
			16945: out = 24'(-27624);
			16946: out = 24'(-23364);
			16947: out = 24'(-4360);
			16948: out = 24'(11472);
			16949: out = 24'(33820);
			16950: out = 24'(32832);
			16951: out = 24'(4812);
			16952: out = 24'(-31744);
			16953: out = 24'(-52116);
			16954: out = 24'(-50676);
			16955: out = 24'(-35912);
			16956: out = 24'(-9984);
			16957: out = 24'(5804);
			16958: out = 24'(26696);
			16959: out = 24'(32952);
			16960: out = 24'(24436);
			16961: out = 24'(2240);
			16962: out = 24'(-36);
			16963: out = 24'(-7928);
			16964: out = 24'(-23532);
			16965: out = 24'(-9708);
			16966: out = 24'(4728);
			16967: out = 24'(11500);
			16968: out = 24'(8844);
			16969: out = 24'(4828);
			16970: out = 24'(20512);
			16971: out = 24'(23844);
			16972: out = 24'(10184);
			16973: out = 24'(-10092);
			16974: out = 24'(-6248);
			16975: out = 24'(-8208);
			16976: out = 24'(-5624);
			16977: out = 24'(11452);
			16978: out = 24'(28840);
			16979: out = 24'(24616);
			16980: out = 24'(7104);
			16981: out = 24'(-6996);
			16982: out = 24'(-1612);
			16983: out = 24'(-22940);
			16984: out = 24'(-32620);
			16985: out = 24'(-680);
			16986: out = 24'(48036);
			16987: out = 24'(41464);
			16988: out = 24'(8148);
			16989: out = 24'(-12968);
			16990: out = 24'(-11712);
			16991: out = 24'(-2032);
			16992: out = 24'(-1876);
			16993: out = 24'(-1044);
			16994: out = 24'(-3408);
			16995: out = 24'(4128);
			16996: out = 24'(-2516);
			16997: out = 24'(12408);
			16998: out = 24'(35880);
			16999: out = 24'(11160);
			17000: out = 24'(-20380);
			17001: out = 24'(-26400);
			17002: out = 24'(-11912);
			17003: out = 24'(-28908);
			17004: out = 24'(-19836);
			17005: out = 24'(14596);
			17006: out = 24'(37300);
			17007: out = 24'(16020);
			17008: out = 24'(-584);
			17009: out = 24'(11292);
			17010: out = 24'(14984);
			17011: out = 24'(-27940);
			17012: out = 24'(-39192);
			17013: out = 24'(-10664);
			17014: out = 24'(25584);
			17015: out = 24'(18944);
			17016: out = 24'(3644);
			17017: out = 24'(-4032);
			17018: out = 24'(480);
			17019: out = 24'(-5580);
			17020: out = 24'(-18428);
			17021: out = 24'(-15844);
			17022: out = 24'(-1776);
			17023: out = 24'(10700);
			17024: out = 24'(14908);
			17025: out = 24'(4632);
			17026: out = 24'(-13852);
			17027: out = 24'(-14332);
			17028: out = 24'(7104);
			17029: out = 24'(10624);
			17030: out = 24'(-15728);
			17031: out = 24'(-32892);
			17032: out = 24'(-6176);
			17033: out = 24'(5028);
			17034: out = 24'(17116);
			17035: out = 24'(24920);
			17036: out = 24'(28308);
			17037: out = 24'(1716);
			17038: out = 24'(-30692);
			17039: out = 24'(-48352);
			17040: out = 24'(-28792);
			17041: out = 24'(14128);
			17042: out = 24'(13708);
			17043: out = 24'(6240);
			17044: out = 24'(12176);
			17045: out = 24'(14092);
			17046: out = 24'(-5680);
			17047: out = 24'(-29148);
			17048: out = 24'(-28660);
			17049: out = 24'(-14948);
			17050: out = 24'(-8048);
			17051: out = 24'(-6204);
			17052: out = 24'(16348);
			17053: out = 24'(38368);
			17054: out = 24'(24840);
			17055: out = 24'(-4888);
			17056: out = 24'(-11196);
			17057: out = 24'(-2136);
			17058: out = 24'(-12432);
			17059: out = 24'(-28216);
			17060: out = 24'(-5312);
			17061: out = 24'(28004);
			17062: out = 24'(7456);
			17063: out = 24'(8772);
			17064: out = 24'(17212);
			17065: out = 24'(20608);
			17066: out = 24'(-2764);
			17067: out = 24'(-20592);
			17068: out = 24'(-18604);
			17069: out = 24'(-5260);
			17070: out = 24'(1040);
			17071: out = 24'(1904);
			17072: out = 24'(31744);
			17073: out = 24'(42712);
			17074: out = 24'(14776);
			17075: out = 24'(-16220);
			17076: out = 24'(-10396);
			17077: out = 24'(3536);
			17078: out = 24'(-8852);
			17079: out = 24'(-30960);
			17080: out = 24'(-12664);
			17081: out = 24'(23880);
			17082: out = 24'(35244);
			17083: out = 24'(14376);
			17084: out = 24'(1620);
			17085: out = 24'(-5108);
			17086: out = 24'(-8516);
			17087: out = 24'(-11960);
			17088: out = 24'(-19760);
			17089: out = 24'(-6652);
			17090: out = 24'(8396);
			17091: out = 24'(7504);
			17092: out = 24'(24652);
			17093: out = 24'(22272);
			17094: out = 24'(16848);
			17095: out = 24'(-14852);
			17096: out = 24'(-49380);
			17097: out = 24'(-77652);
			17098: out = 24'(-23548);
			17099: out = 24'(44376);
			17100: out = 24'(41932);
			17101: out = 24'(-1944);
			17102: out = 24'(-14160);
			17103: out = 24'(5596);
			17104: out = 24'(3716);
			17105: out = 24'(-25956);
			17106: out = 24'(-34128);
			17107: out = 24'(-7704);
			17108: out = 24'(16872);
			17109: out = 24'(-3108);
			17110: out = 24'(13212);
			17111: out = 24'(30008);
			17112: out = 24'(14976);
			17113: out = 24'(-24836);
			17114: out = 24'(-17708);
			17115: out = 24'(13804);
			17116: out = 24'(15704);
			17117: out = 24'(-23012);
			17118: out = 24'(-38752);
			17119: out = 24'(-19552);
			17120: out = 24'(7840);
			17121: out = 24'(12368);
			17122: out = 24'(6948);
			17123: out = 24'(1992);
			17124: out = 24'(-7100);
			17125: out = 24'(-23744);
			17126: out = 24'(-5892);
			17127: out = 24'(84);
			17128: out = 24'(1344);
			17129: out = 24'(4184);
			17130: out = 24'(24560);
			17131: out = 24'(16208);
			17132: out = 24'(-4476);
			17133: out = 24'(-17616);
			17134: out = 24'(1012);
			17135: out = 24'(-6508);
			17136: out = 24'(-12864);
			17137: out = 24'(-9804);
			17138: out = 24'(4960);
			17139: out = 24'(2016);
			17140: out = 24'(2428);
			17141: out = 24'(10004);
			17142: out = 24'(15564);
			17143: out = 24'(-4888);
			17144: out = 24'(-24284);
			17145: out = 24'(-17164);
			17146: out = 24'(14596);
			17147: out = 24'(15372);
			17148: out = 24'(19276);
			17149: out = 24'(15940);
			17150: out = 24'(17236);
			17151: out = 24'(6896);
			17152: out = 24'(3868);
			17153: out = 24'(-14436);
			17154: out = 24'(-20300);
			17155: out = 24'(584);
			17156: out = 24'(8352);
			17157: out = 24'(3828);
			17158: out = 24'(3816);
			17159: out = 24'(16660);
			17160: out = 24'(5628);
			17161: out = 24'(-9004);
			17162: out = 24'(-11888);
			17163: out = 24'(1976);
			17164: out = 24'(7552);
			17165: out = 24'(-5684);
			17166: out = 24'(-16424);
			17167: out = 24'(-5796);
			17168: out = 24'(-1468);
			17169: out = 24'(13780);
			17170: out = 24'(20968);
			17171: out = 24'(21852);
			17172: out = 24'(-2336);
			17173: out = 24'(4664);
			17174: out = 24'(-11796);
			17175: out = 24'(-25980);
			17176: out = 24'(-16076);
			17177: out = 24'(23556);
			17178: out = 24'(43236);
			17179: out = 24'(38572);
			17180: out = 24'(12780);
			17181: out = 24'(-22524);
			17182: out = 24'(-54916);
			17183: out = 24'(-45928);
			17184: out = 24'(-2296);
			17185: out = 24'(14448);
			17186: out = 24'(18308);
			17187: out = 24'(16256);
			17188: out = 24'(14024);
			17189: out = 24'(-620);
			17190: out = 24'(-22860);
			17191: out = 24'(-20384);
			17192: out = 24'(9888);
			17193: out = 24'(20788);
			17194: out = 24'(6684);
			17195: out = 24'(-14444);
			17196: out = 24'(-2712);
			17197: out = 24'(21560);
			17198: out = 24'(-16584);
			17199: out = 24'(-23432);
			17200: out = 24'(14388);
			17201: out = 24'(40500);
			17202: out = 24'(5200);
			17203: out = 24'(-46708);
			17204: out = 24'(-42500);
			17205: out = 24'(8248);
			17206: out = 24'(14852);
			17207: out = 24'(1600);
			17208: out = 24'(1916);
			17209: out = 24'(21124);
			17210: out = 24'(13444);
			17211: out = 24'(-6132);
			17212: out = 24'(-23984);
			17213: out = 24'(-17904);
			17214: out = 24'(-384);
			17215: out = 24'(-8720);
			17216: out = 24'(5216);
			17217: out = 24'(23312);
			17218: out = 24'(21248);
			17219: out = 24'(3124);
			17220: out = 24'(-5844);
			17221: out = 24'(-2308);
			17222: out = 24'(2176);
			17223: out = 24'(-10252);
			17224: out = 24'(-3576);
			17225: out = 24'(-984);
			17226: out = 24'(2088);
			17227: out = 24'(16300);
			17228: out = 24'(20480);
			17229: out = 24'(9968);
			17230: out = 24'(-3348);
			17231: out = 24'(-1480);
			17232: out = 24'(-18088);
			17233: out = 24'(-12380);
			17234: out = 24'(8916);
			17235: out = 24'(22788);
			17236: out = 24'(18140);
			17237: out = 24'(7616);
			17238: out = 24'(16040);
			17239: out = 24'(28068);
			17240: out = 24'(8596);
			17241: out = 24'(-14912);
			17242: out = 24'(-16212);
			17243: out = 24'(-1648);
			17244: out = 24'(-7944);
			17245: out = 24'(-14736);
			17246: out = 24'(-6292);
			17247: out = 24'(11368);
			17248: out = 24'(9608);
			17249: out = 24'(12164);
			17250: out = 24'(3772);
			17251: out = 24'(-6036);
			17252: out = 24'(-12416);
			17253: out = 24'(-25556);
			17254: out = 24'(-9896);
			17255: out = 24'(9492);
			17256: out = 24'(13924);
			17257: out = 24'(-1892);
			17258: out = 24'(4076);
			17259: out = 24'(1024);
			17260: out = 24'(-17232);
			17261: out = 24'(-33596);
			17262: out = 24'(488);
			17263: out = 24'(25596);
			17264: out = 24'(14284);
			17265: out = 24'(-10028);
			17266: out = 24'(-3104);
			17267: out = 24'(7488);
			17268: out = 24'(3048);
			17269: out = 24'(-1772);
			17270: out = 24'(-8928);
			17271: out = 24'(7648);
			17272: out = 24'(11448);
			17273: out = 24'(-6156);
			17274: out = 24'(-19316);
			17275: out = 24'(-7500);
			17276: out = 24'(4712);
			17277: out = 24'(-5284);
			17278: out = 24'(-8616);
			17279: out = 24'(-6732);
			17280: out = 24'(6244);
			17281: out = 24'(3756);
			17282: out = 24'(1012);
			17283: out = 24'(1276);
			17284: out = 24'(27480);
			17285: out = 24'(30248);
			17286: out = 24'(4124);
			17287: out = 24'(-58956);
			17288: out = 24'(-41792);
			17289: out = 24'(4920);
			17290: out = 24'(11720);
			17291: out = 24'(-20252);
			17292: out = 24'(-2040);
			17293: out = 24'(26048);
			17294: out = 24'(15616);
			17295: out = 24'(-15804);
			17296: out = 24'(-11168);
			17297: out = 24'(11336);
			17298: out = 24'(8496);
			17299: out = 24'(-17864);
			17300: out = 24'(-13572);
			17301: out = 24'(15736);
			17302: out = 24'(27448);
			17303: out = 24'(84);
			17304: out = 24'(-19660);
			17305: out = 24'(-22332);
			17306: out = 24'(4660);
			17307: out = 24'(29904);
			17308: out = 24'(18956);
			17309: out = 24'(-12076);
			17310: out = 24'(-22104);
			17311: out = 24'(3348);
			17312: out = 24'(-4464);
			17313: out = 24'(18736);
			17314: out = 24'(15204);
			17315: out = 24'(-11964);
			17316: out = 24'(-54336);
			17317: out = 24'(-54356);
			17318: out = 24'(-32620);
			17319: out = 24'(7200);
			17320: out = 24'(46564);
			17321: out = 24'(58212);
			17322: out = 24'(31564);
			17323: out = 24'(-12404);
			17324: out = 24'(-51636);
			17325: out = 24'(-36908);
			17326: out = 24'(-31632);
			17327: out = 24'(-18640);
			17328: out = 24'(11736);
			17329: out = 24'(46924);
			17330: out = 24'(39872);
			17331: out = 24'(20308);
			17332: out = 24'(2560);
			17333: out = 24'(-19304);
			17334: out = 24'(-39624);
			17335: out = 24'(-34280);
			17336: out = 24'(-6144);
			17337: out = 24'(-1888);
			17338: out = 24'(11124);
			17339: out = 24'(-1732);
			17340: out = 24'(-5388);
			17341: out = 24'(10812);
			17342: out = 24'(16972);
			17343: out = 24'(7556);
			17344: out = 24'(-3052);
			17345: out = 24'(2132);
			17346: out = 24'(14824);
			17347: out = 24'(10948);
			17348: out = 24'(-3520);
			17349: out = 24'(-7128);
			17350: out = 24'(6732);
			17351: out = 24'(16352);
			17352: out = 24'(4008);
			17353: out = 24'(-24620);
			17354: out = 24'(-52708);
			17355: out = 24'(-29568);
			17356: out = 24'(-528);
			17357: out = 24'(12664);
			17358: out = 24'(19156);
			17359: out = 24'(30104);
			17360: out = 24'(17952);
			17361: out = 24'(-17360);
			17362: out = 24'(-43144);
			17363: out = 24'(-56556);
			17364: out = 24'(-18240);
			17365: out = 24'(12288);
			17366: out = 24'(17868);
			17367: out = 24'(1840);
			17368: out = 24'(34488);
			17369: out = 24'(47132);
			17370: out = 24'(27428);
			17371: out = 24'(-376);
			17372: out = 24'(-14540);
			17373: out = 24'(-35188);
			17374: out = 24'(-44080);
			17375: out = 24'(-6108);
			17376: out = 24'(6088);
			17377: out = 24'(19720);
			17378: out = 24'(31360);
			17379: out = 24'(35944);
			17380: out = 24'(-9964);
			17381: out = 24'(-39164);
			17382: out = 24'(-30080);
			17383: out = 24'(3536);
			17384: out = 24'(-8364);
			17385: out = 24'(-4264);
			17386: out = 24'(14816);
			17387: out = 24'(31188);
			17388: out = 24'(724);
			17389: out = 24'(2712);
			17390: out = 24'(7316);
			17391: out = 24'(6292);
			17392: out = 24'(-4624);
			17393: out = 24'(-10336);
			17394: out = 24'(4420);
			17395: out = 24'(19848);
			17396: out = 24'(14892);
			17397: out = 24'(1800);
			17398: out = 24'(704);
			17399: out = 24'(2888);
			17400: out = 24'(-11224);
			17401: out = 24'(-54012);
			17402: out = 24'(-39956);
			17403: out = 24'(7572);
			17404: out = 24'(32844);
			17405: out = 24'(27064);
			17406: out = 24'(11632);
			17407: out = 24'(15352);
			17408: out = 24'(23564);
			17409: out = 24'(6352);
			17410: out = 24'(-26380);
			17411: out = 24'(-50284);
			17412: out = 24'(-36916);
			17413: out = 24'(1628);
			17414: out = 24'(22988);
			17415: out = 24'(33952);
			17416: out = 24'(44072);
			17417: out = 24'(40736);
			17418: out = 24'(14528);
			17419: out = 24'(-34480);
			17420: out = 24'(-58520);
			17421: out = 24'(-39076);
			17422: out = 24'(-22104);
			17423: out = 24'(-4668);
			17424: out = 24'(8360);
			17425: out = 24'(19636);
			17426: out = 24'(16916);
			17427: out = 24'(11604);
			17428: out = 24'(8176);
			17429: out = 24'(6080);
			17430: out = 24'(-11796);
			17431: out = 24'(-24448);
			17432: out = 24'(-27068);
			17433: out = 24'(-7904);
			17434: out = 24'(10880);
			17435: out = 24'(39180);
			17436: out = 24'(16448);
			17437: out = 24'(-4580);
			17438: out = 24'(4328);
			17439: out = 24'(28760);
			17440: out = 24'(7188);
			17441: out = 24'(-28280);
			17442: out = 24'(-31392);
			17443: out = 24'(5456);
			17444: out = 24'(6336);
			17445: out = 24'(-19120);
			17446: out = 24'(-26168);
			17447: out = 24'(9888);
			17448: out = 24'(24672);
			17449: out = 24'(72);
			17450: out = 24'(-39644);
			17451: out = 24'(-40244);
			17452: out = 24'(5364);
			17453: out = 24'(42444);
			17454: out = 24'(36108);
			17455: out = 24'(15468);
			17456: out = 24'(-4);
			17457: out = 24'(12788);
			17458: out = 24'(5344);
			17459: out = 24'(-27064);
			17460: out = 24'(-60448);
			17461: out = 24'(-14740);
			17462: out = 24'(29408);
			17463: out = 24'(26576);
			17464: out = 24'(20560);
			17465: out = 24'(13164);
			17466: out = 24'(21412);
			17467: out = 24'(1052);
			17468: out = 24'(-37036);
			17469: out = 24'(-59632);
			17470: out = 24'(-24144);
			17471: out = 24'(7232);
			17472: out = 24'(404);
			17473: out = 24'(1132);
			17474: out = 24'(25440);
			17475: out = 24'(44044);
			17476: out = 24'(32432);
			17477: out = 24'(6056);
			17478: out = 24'(2256);
			17479: out = 24'(3232);
			17480: out = 24'(-6536);
			17481: out = 24'(-28192);
			17482: out = 24'(-21352);
			17483: out = 24'(-10188);
			17484: out = 24'(11976);
			17485: out = 24'(36720);
			17486: out = 24'(29892);
			17487: out = 24'(-9724);
			17488: out = 24'(-32188);
			17489: out = 24'(-5464);
			17490: out = 24'(5552);
			17491: out = 24'(4972);
			17492: out = 24'(-1328);
			17493: out = 24'(-1004);
			17494: out = 24'(-17116);
			17495: out = 24'(-23392);
			17496: out = 24'(-13384);
			17497: out = 24'(3076);
			17498: out = 24'(1112);
			17499: out = 24'(-564);
			17500: out = 24'(14704);
			17501: out = 24'(36772);
			17502: out = 24'(35496);
			17503: out = 24'(8028);
			17504: out = 24'(-9252);
			17505: out = 24'(-9408);
			17506: out = 24'(-12448);
			17507: out = 24'(-29000);
			17508: out = 24'(-30888);
			17509: out = 24'(-9284);
			17510: out = 24'(14632);
			17511: out = 24'(9540);
			17512: out = 24'(3364);
			17513: out = 24'(-1340);
			17514: out = 24'(4204);
			17515: out = 24'(14964);
			17516: out = 24'(10380);
			17517: out = 24'(-14560);
			17518: out = 24'(-31360);
			17519: out = 24'(-12428);
			17520: out = 24'(-1240);
			17521: out = 24'(1340);
			17522: out = 24'(4136);
			17523: out = 24'(18792);
			17524: out = 24'(24312);
			17525: out = 24'(2412);
			17526: out = 24'(-31456);
			17527: out = 24'(-35344);
			17528: out = 24'(9540);
			17529: out = 24'(19436);
			17530: out = 24'(-11140);
			17531: out = 24'(-32604);
			17532: out = 24'(-2892);
			17533: out = 24'(22516);
			17534: out = 24'(15656);
			17535: out = 24'(-1564);
			17536: out = 24'(-8544);
			17537: out = 24'(13244);
			17538: out = 24'(10284);
			17539: out = 24'(1072);
			17540: out = 24'(8984);
			17541: out = 24'(2956);
			17542: out = 24'(-17816);
			17543: out = 24'(-19512);
			17544: out = 24'(13032);
			17545: out = 24'(16160);
			17546: out = 24'(9520);
			17547: out = 24'(6384);
			17548: out = 24'(21136);
			17549: out = 24'(36200);
			17550: out = 24'(18728);
			17551: out = 24'(-6012);
			17552: out = 24'(-21488);
			17553: out = 24'(-18232);
			17554: out = 24'(-31600);
			17555: out = 24'(-18432);
			17556: out = 24'(4160);
			17557: out = 24'(5244);
			17558: out = 24'(20404);
			17559: out = 24'(34900);
			17560: out = 24'(28072);
			17561: out = 24'(-5356);
			17562: out = 24'(-34024);
			17563: out = 24'(-24060);
			17564: out = 24'(228);
			17565: out = 24'(8860);
			17566: out = 24'(8532);
			17567: out = 24'(26996);
			17568: out = 24'(27592);
			17569: out = 24'(-1548);
			17570: out = 24'(-25388);
			17571: out = 24'(-18636);
			17572: out = 24'(2064);
			17573: out = 24'(7844);
			17574: out = 24'(9100);
			17575: out = 24'(88);
			17576: out = 24'(212);
			17577: out = 24'(-4504);
			17578: out = 24'(-12936);
			17579: out = 24'(10880);
			17580: out = 24'(19800);
			17581: out = 24'(-16);
			17582: out = 24'(-35784);
			17583: out = 24'(-28860);
			17584: out = 24'(-532);
			17585: out = 24'(28424);
			17586: out = 24'(24188);
			17587: out = 24'(3412);
			17588: out = 24'(-24612);
			17589: out = 24'(-19756);
			17590: out = 24'(-2876);
			17591: out = 24'(-160);
			17592: out = 24'(-26312);
			17593: out = 24'(-22736);
			17594: out = 24'(7972);
			17595: out = 24'(29956);
			17596: out = 24'(5728);
			17597: out = 24'(-2632);
			17598: out = 24'(1724);
			17599: out = 24'(464);
			17600: out = 24'(-32424);
			17601: out = 24'(-31368);
			17602: out = 24'(-10116);
			17603: out = 24'(9292);
			17604: out = 24'(24376);
			17605: out = 24'(21268);
			17606: out = 24'(8928);
			17607: out = 24'(-832);
			17608: out = 24'(612);
			17609: out = 24'(1556);
			17610: out = 24'(-7940);
			17611: out = 24'(-22424);
			17612: out = 24'(-30084);
			17613: out = 24'(2528);
			17614: out = 24'(11120);
			17615: out = 24'(2420);
			17616: out = 24'(4168);
			17617: out = 24'(21628);
			17618: out = 24'(16008);
			17619: out = 24'(-3676);
			17620: out = 24'(-7372);
			17621: out = 24'(-20168);
			17622: out = 24'(3120);
			17623: out = 24'(6960);
			17624: out = 24'(2176);
			17625: out = 24'(8016);
			17626: out = 24'(11804);
			17627: out = 24'(-4700);
			17628: out = 24'(-14328);
			17629: out = 24'(9432);
			17630: out = 24'(10428);
			17631: out = 24'(2824);
			17632: out = 24'(2552);
			17633: out = 24'(8668);
			17634: out = 24'(30868);
			17635: out = 24'(11280);
			17636: out = 24'(2716);
			17637: out = 24'(15200);
			17638: out = 24'(10400);
			17639: out = 24'(-34116);
			17640: out = 24'(-42572);
			17641: out = 24'(12412);
			17642: out = 24'(38948);
			17643: out = 24'(22344);
			17644: out = 24'(-4816);
			17645: out = 24'(-1300);
			17646: out = 24'(4592);
			17647: out = 24'(10392);
			17648: out = 24'(-7484);
			17649: out = 24'(-20820);
			17650: out = 24'(-13308);
			17651: out = 24'(3968);
			17652: out = 24'(5552);
			17653: out = 24'(-3624);
			17654: out = 24'(1500);
			17655: out = 24'(-3880);
			17656: out = 24'(22584);
			17657: out = 24'(18276);
			17658: out = 24'(-16696);
			17659: out = 24'(-36080);
			17660: out = 24'(-7936);
			17661: out = 24'(11136);
			17662: out = 24'(-8028);
			17663: out = 24'(-19036);
			17664: out = 24'(1856);
			17665: out = 24'(37564);
			17666: out = 24'(29500);
			17667: out = 24'(-23548);
			17668: out = 24'(-27200);
			17669: out = 24'(-916);
			17670: out = 24'(15748);
			17671: out = 24'(-3632);
			17672: out = 24'(-10912);
			17673: out = 24'(-9520);
			17674: out = 24'(8028);
			17675: out = 24'(13480);
			17676: out = 24'(2932);
			17677: out = 24'(-9580);
			17678: out = 24'(-2080);
			17679: out = 24'(7324);
			17680: out = 24'(752);
			17681: out = 24'(-21956);
			17682: out = 24'(-23272);
			17683: out = 24'(-912);
			17684: out = 24'(23648);
			17685: out = 24'(7632);
			17686: out = 24'(4248);
			17687: out = 24'(7648);
			17688: out = 24'(-3820);
			17689: out = 24'(-39852);
			17690: out = 24'(-48428);
			17691: out = 24'(-17980);
			17692: out = 24'(20932);
			17693: out = 24'(30436);
			17694: out = 24'(19068);
			17695: out = 24'(-4404);
			17696: out = 24'(-16428);
			17697: out = 24'(1836);
			17698: out = 24'(3760);
			17699: out = 24'(-7940);
			17700: out = 24'(-7092);
			17701: out = 24'(23804);
			17702: out = 24'(31784);
			17703: out = 24'(14648);
			17704: out = 24'(-3892);
			17705: out = 24'(2512);
			17706: out = 24'(-19676);
			17707: out = 24'(-32000);
			17708: out = 24'(-21736);
			17709: out = 24'(12220);
			17710: out = 24'(14768);
			17711: out = 24'(17452);
			17712: out = 24'(15544);
			17713: out = 24'(16040);
			17714: out = 24'(15304);
			17715: out = 24'(3588);
			17716: out = 24'(-4212);
			17717: out = 24'(-720);
			17718: out = 24'(-2092);
			17719: out = 24'(-17792);
			17720: out = 24'(-22184);
			17721: out = 24'(-244);
			17722: out = 24'(13676);
			17723: out = 24'(25892);
			17724: out = 24'(7396);
			17725: out = 24'(28);
			17726: out = 24'(6112);
			17727: out = 24'(6452);
			17728: out = 24'(-27788);
			17729: out = 24'(-35428);
			17730: out = 24'(7400);
			17731: out = 24'(26308);
			17732: out = 24'(23516);
			17733: out = 24'(5520);
			17734: out = 24'(-4236);
			17735: out = 24'(-20632);
			17736: out = 24'(-9416);
			17737: out = 24'(-7040);
			17738: out = 24'(-12296);
			17739: out = 24'(-12880);
			17740: out = 24'(5884);
			17741: out = 24'(22160);
			17742: out = 24'(16316);
			17743: out = 24'(-1704);
			17744: out = 24'(-3804);
			17745: out = 24'(14896);
			17746: out = 24'(17332);
			17747: out = 24'(-7308);
			17748: out = 24'(-26748);
			17749: out = 24'(-13340);
			17750: out = 24'(9784);
			17751: out = 24'(12032);
			17752: out = 24'(-4716);
			17753: out = 24'(2124);
			17754: out = 24'(10468);
			17755: out = 24'(-2972);
			17756: out = 24'(-42452);
			17757: out = 24'(-9628);
			17758: out = 24'(15604);
			17759: out = 24'(4208);
			17760: out = 24'(-27468);
			17761: out = 24'(8380);
			17762: out = 24'(24688);
			17763: out = 24'(14796);
			17764: out = 24'(-1336);
			17765: out = 24'(-1884);
			17766: out = 24'(-2220);
			17767: out = 24'(-18048);
			17768: out = 24'(-28736);
			17769: out = 24'(14036);
			17770: out = 24'(31508);
			17771: out = 24'(20628);
			17772: out = 24'(-6140);
			17773: out = 24'(852);
			17774: out = 24'(-12056);
			17775: out = 24'(-204);
			17776: out = 24'(6368);
			17777: out = 24'(-1880);
			17778: out = 24'(-21132);
			17779: out = 24'(-18588);
			17780: out = 24'(-2924);
			17781: out = 24'(8164);
			17782: out = 24'(504);
			17783: out = 24'(-2636);
			17784: out = 24'(-12352);
			17785: out = 24'(-22376);
			17786: out = 24'(-5760);
			17787: out = 24'(5900);
			17788: out = 24'(8008);
			17789: out = 24'(3720);
			17790: out = 24'(8880);
			17791: out = 24'(-7652);
			17792: out = 24'(-21180);
			17793: out = 24'(-14464);
			17794: out = 24'(17824);
			17795: out = 24'(10780);
			17796: out = 24'(3648);
			17797: out = 24'(2060);
			17798: out = 24'(8380);
			17799: out = 24'(-7204);
			17800: out = 24'(-13048);
			17801: out = 24'(-11020);
			17802: out = 24'(-1840);
			17803: out = 24'(15628);
			17804: out = 24'(7244);
			17805: out = 24'(-5772);
			17806: out = 24'(-4372);
			17807: out = 24'(23252);
			17808: out = 24'(7728);
			17809: out = 24'(-7396);
			17810: out = 24'(-4240);
			17811: out = 24'(16376);
			17812: out = 24'(16648);
			17813: out = 24'(11804);
			17814: out = 24'(5660);
			17815: out = 24'(1472);
			17816: out = 24'(-20732);
			17817: out = 24'(-18444);
			17818: out = 24'(-1852);
			17819: out = 24'(7100);
			17820: out = 24'(-3456);
			17821: out = 24'(-4092);
			17822: out = 24'(10448);
			17823: out = 24'(21480);
			17824: out = 24'(-5040);
			17825: out = 24'(-12716);
			17826: out = 24'(-9904);
			17827: out = 24'(6336);
			17828: out = 24'(21384);
			17829: out = 24'(6584);
			17830: out = 24'(-16892);
			17831: out = 24'(-17168);
			17832: out = 24'(9280);
			17833: out = 24'(21680);
			17834: out = 24'(15204);
			17835: out = 24'(3236);
			17836: out = 24'(-2412);
			17837: out = 24'(-17472);
			17838: out = 24'(-17096);
			17839: out = 24'(5748);
			17840: out = 24'(29224);
			17841: out = 24'(40);
			17842: out = 24'(-3268);
			17843: out = 24'(8288);
			17844: out = 24'(21804);
			17845: out = 24'(-4608);
			17846: out = 24'(-10168);
			17847: out = 24'(-31080);
			17848: out = 24'(-43732);
			17849: out = 24'(-30912);
			17850: out = 24'(7744);
			17851: out = 24'(16740);
			17852: out = 24'(2560);
			17853: out = 24'(2472);
			17854: out = 24'(4024);
			17855: out = 24'(18012);
			17856: out = 24'(-3676);
			17857: out = 24'(-43660);
			17858: out = 24'(-20736);
			17859: out = 24'(16436);
			17860: out = 24'(33992);
			17861: out = 24'(17236);
			17862: out = 24'(2468);
			17863: out = 24'(-12872);
			17864: out = 24'(-8340);
			17865: out = 24'(1752);
			17866: out = 24'(-1348);
			17867: out = 24'(-3056);
			17868: out = 24'(-9588);
			17869: out = 24'(-6348);
			17870: out = 24'(16);
			17871: out = 24'(15836);
			17872: out = 24'(5868);
			17873: out = 24'(2452);
			17874: out = 24'(11108);
			17875: out = 24'(-3408);
			17876: out = 24'(-28524);
			17877: out = 24'(-31776);
			17878: out = 24'(-1236);
			17879: out = 24'(21168);
			17880: out = 24'(11900);
			17881: out = 24'(-2520);
			17882: out = 24'(8708);
			17883: out = 24'(35192);
			17884: out = 24'(6440);
			17885: out = 24'(-25216);
			17886: out = 24'(-26152);
			17887: out = 24'(336);
			17888: out = 24'(748);
			17889: out = 24'(928);
			17890: out = 24'(8312);
			17891: out = 24'(14916);
			17892: out = 24'(2276);
			17893: out = 24'(-3112);
			17894: out = 24'(6116);
			17895: out = 24'(13316);
			17896: out = 24'(-8096);
			17897: out = 24'(-10268);
			17898: out = 24'(8372);
			17899: out = 24'(21156);
			17900: out = 24'(-1780);
			17901: out = 24'(-13284);
			17902: out = 24'(-5040);
			17903: out = 24'(8952);
			17904: out = 24'(-3284);
			17905: out = 24'(-10936);
			17906: out = 24'(-15420);
			17907: out = 24'(-3152);
			17908: out = 24'(7428);
			17909: out = 24'(9268);
			17910: out = 24'(-1000);
			17911: out = 24'(-6920);
			17912: out = 24'(-2936);
			17913: out = 24'(22392);
			17914: out = 24'(-3592);
			17915: out = 24'(-29228);
			17916: out = 24'(-19992);
			17917: out = 24'(13252);
			17918: out = 24'(10284);
			17919: out = 24'(-7268);
			17920: out = 24'(-40);
			17921: out = 24'(28868);
			17922: out = 24'(28672);
			17923: out = 24'(-8244);
			17924: out = 24'(-35480);
			17925: out = 24'(-14556);
			17926: out = 24'(23712);
			17927: out = 24'(11488);
			17928: out = 24'(-24044);
			17929: out = 24'(-19900);
			17930: out = 24'(22072);
			17931: out = 24'(38152);
			17932: out = 24'(4424);
			17933: out = 24'(-29484);
			17934: out = 24'(-16576);
			17935: out = 24'(25888);
			17936: out = 24'(25336);
			17937: out = 24'(-13828);
			17938: out = 24'(-28856);
			17939: out = 24'(800);
			17940: out = 24'(31784);
			17941: out = 24'(12760);
			17942: out = 24'(-32860);
			17943: out = 24'(-41988);
			17944: out = 24'(-1696);
			17945: out = 24'(29980);
			17946: out = 24'(19840);
			17947: out = 24'(10628);
			17948: out = 24'(932);
			17949: out = 24'(-11072);
			17950: out = 24'(-29532);
			17951: out = 24'(-416);
			17952: out = 24'(3168);
			17953: out = 24'(20352);
			17954: out = 24'(25832);
			17955: out = 24'(-1432);
			17956: out = 24'(-13712);
			17957: out = 24'(-4896);
			17958: out = 24'(10648);
			17959: out = 24'(4792);
			17960: out = 24'(-13124);
			17961: out = 24'(-28616);
			17962: out = 24'(-20936);
			17963: out = 24'(608);
			17964: out = 24'(7564);
			17965: out = 24'(11028);
			17966: out = 24'(11464);
			17967: out = 24'(7496);
			17968: out = 24'(16196);
			17969: out = 24'(-7992);
			17970: out = 24'(-28948);
			17971: out = 24'(-27376);
			17972: out = 24'(7808);
			17973: out = 24'(8488);
			17974: out = 24'(8564);
			17975: out = 24'(5964);
			17976: out = 24'(136);
			17977: out = 24'(-1864);
			17978: out = 24'(9156);
			17979: out = 24'(13892);
			17980: out = 24'(-128);
			17981: out = 24'(-25012);
			17982: out = 24'(-15332);
			17983: out = 24'(12372);
			17984: out = 24'(19408);
			17985: out = 24'(-10440);
			17986: out = 24'(-15060);
			17987: out = 24'(-2072);
			17988: out = 24'(2884);
			17989: out = 24'(1380);
			17990: out = 24'(-2032);
			17991: out = 24'(5340);
			17992: out = 24'(5636);
			17993: out = 24'(988);
			17994: out = 24'(-25220);
			17995: out = 24'(-7096);
			17996: out = 24'(24144);
			17997: out = 24'(19472);
			17998: out = 24'(-6460);
			17999: out = 24'(-24492);
			18000: out = 24'(-15908);
			18001: out = 24'(-4);
			18002: out = 24'(3384);
			18003: out = 24'(11260);
			18004: out = 24'(21236);
			18005: out = 24'(19996);
			18006: out = 24'(1028);
			18007: out = 24'(-3356);
			18008: out = 24'(6440);
			18009: out = 24'(14612);
			18010: out = 24'(1036);
			18011: out = 24'(3600);
			18012: out = 24'(-5732);
			18013: out = 24'(-21856);
			18014: out = 24'(-31216);
			18015: out = 24'(6304);
			18016: out = 24'(28700);
			18017: out = 24'(21536);
			18018: out = 24'(0);
			18019: out = 24'(-10448);
			18020: out = 24'(-8208);
			18021: out = 24'(-12092);
			18022: out = 24'(-25308);
			18023: out = 24'(-9892);
			18024: out = 24'(-4300);
			18025: out = 24'(7768);
			18026: out = 24'(17820);
			18027: out = 24'(22780);
			18028: out = 24'(-8508);
			18029: out = 24'(-26908);
			18030: out = 24'(-16584);
			18031: out = 24'(2764);
			18032: out = 24'(-1928);
			18033: out = 24'(-13264);
			18034: out = 24'(-5764);
			18035: out = 24'(17736);
			18036: out = 24'(23528);
			18037: out = 24'(1484);
			18038: out = 24'(-23164);
			18039: out = 24'(-17904);
			18040: out = 24'(11616);
			18041: out = 24'(25108);
			18042: out = 24'(11528);
			18043: out = 24'(-11204);
			18044: out = 24'(-28060);
			18045: out = 24'(-22620);
			18046: out = 24'(-9784);
			18047: out = 24'(1980);
			18048: out = 24'(92);
			18049: out = 24'(21680);
			18050: out = 24'(13428);
			18051: out = 24'(-7532);
			18052: out = 24'(-16596);
			18053: out = 24'(4064);
			18054: out = 24'(11772);
			18055: out = 24'(-2028);
			18056: out = 24'(-22656);
			18057: out = 24'(6908);
			18058: out = 24'(9540);
			18059: out = 24'(4236);
			18060: out = 24'(-7136);
			18061: out = 24'(1484);
			18062: out = 24'(-10204);
			18063: out = 24'(7964);
			18064: out = 24'(28572);
			18065: out = 24'(15256);
			18066: out = 24'(-1892);
			18067: out = 24'(3552);
			18068: out = 24'(15220);
			18069: out = 24'(-3328);
			18070: out = 24'(304);
			18071: out = 24'(304);
			18072: out = 24'(5616);
			18073: out = 24'(6304);
			18074: out = 24'(72);
			18075: out = 24'(-1412);
			18076: out = 24'(-3752);
			18077: out = 24'(-12516);
			18078: out = 24'(-18372);
			18079: out = 24'(-11132);
			18080: out = 24'(1360);
			18081: out = 24'(11716);
			18082: out = 24'(26384);
			18083: out = 24'(3348);
			18084: out = 24'(-18368);
			18085: out = 24'(-19440);
			18086: out = 24'(-588);
			18087: out = 24'(-10964);
			18088: out = 24'(-12548);
			18089: out = 24'(5480);
			18090: out = 24'(23376);
			18091: out = 24'(25692);
			18092: out = 24'(6580);
			18093: out = 24'(-2768);
			18094: out = 24'(-3416);
			18095: out = 24'(-3960);
			18096: out = 24'(-15880);
			18097: out = 24'(5108);
			18098: out = 24'(34320);
			18099: out = 24'(14796);
			18100: out = 24'(-18440);
			18101: out = 24'(-21988);
			18102: out = 24'(8680);
			18103: out = 24'(19796);
			18104: out = 24'(12388);
			18105: out = 24'(-4452);
			18106: out = 24'(-14488);
			18107: out = 24'(-19768);
			18108: out = 24'(-13284);
			18109: out = 24'(5464);
			18110: out = 24'(15308);
			18111: out = 24'(6088);
			18112: out = 24'(14824);
			18113: out = 24'(5748);
			18114: out = 24'(-18048);
			18115: out = 24'(-44092);
			18116: out = 24'(-14872);
			18117: out = 24'(-5896);
			18118: out = 24'(7784);
			18119: out = 24'(18532);
			18120: out = 24'(22064);
			18121: out = 24'(1680);
			18122: out = 24'(-15280);
			18123: out = 24'(-16380);
			18124: out = 24'(-10988);
			18125: out = 24'(-15120);
			18126: out = 24'(-21388);
			18127: out = 24'(-4048);
			18128: out = 24'(24780);
			18129: out = 24'(24976);
			18130: out = 24'(-5992);
			18131: out = 24'(-25608);
			18132: out = 24'(-6792);
			18133: out = 24'(19672);
			18134: out = 24'(20716);
			18135: out = 24'(6656);
			18136: out = 24'(216);
			18137: out = 24'(6916);
			18138: out = 24'(7808);
			18139: out = 24'(-2052);
			18140: out = 24'(-23508);
			18141: out = 24'(-39416);
			18142: out = 24'(-11564);
			18143: out = 24'(23324);
			18144: out = 24'(14284);
			18145: out = 24'(-32356);
			18146: out = 24'(-6564);
			18147: out = 24'(29988);
			18148: out = 24'(33404);
			18149: out = 24'(-8772);
			18150: out = 24'(-18464);
			18151: out = 24'(-24916);
			18152: out = 24'(-5164);
			18153: out = 24'(7832);
			18154: out = 24'(964);
			18155: out = 24'(7908);
			18156: out = 24'(13072);
			18157: out = 24'(1436);
			18158: out = 24'(-11724);
			18159: out = 24'(-5768);
			18160: out = 24'(12280);
			18161: out = 24'(8720);
			18162: out = 24'(-10416);
			18163: out = 24'(-40200);
			18164: out = 24'(-13204);
			18165: out = 24'(16720);
			18166: out = 24'(14884);
			18167: out = 24'(16604);
			18168: out = 24'(17076);
			18169: out = 24'(600);
			18170: out = 24'(-32644);
			18171: out = 24'(-24872);
			18172: out = 24'(-19792);
			18173: out = 24'(2516);
			18174: out = 24'(20144);
			18175: out = 24'(23172);
			18176: out = 24'(12228);
			18177: out = 24'(828);
			18178: out = 24'(-13268);
			18179: out = 24'(-42856);
			18180: out = 24'(-15824);
			18181: out = 24'(-5684);
			18182: out = 24'(11300);
			18183: out = 24'(23088);
			18184: out = 24'(27472);
			18185: out = 24'(-11712);
			18186: out = 24'(-21464);
			18187: out = 24'(2364);
			18188: out = 24'(-468);
			18189: out = 24'(-29688);
			18190: out = 24'(-30836);
			18191: out = 24'(8564);
			18192: out = 24'(28692);
			18193: out = 24'(28160);
			18194: out = 24'(18692);
			18195: out = 24'(14560);
			18196: out = 24'(6812);
			18197: out = 24'(-10572);
			18198: out = 24'(-8584);
			18199: out = 24'(1540);
			18200: out = 24'(-2488);
			18201: out = 24'(-3800);
			18202: out = 24'(2296);
			18203: out = 24'(13120);
			18204: out = 24'(16412);
			18205: out = 24'(26652);
			18206: out = 24'(13840);
			18207: out = 24'(-4352);
			18208: out = 24'(-24036);
			18209: out = 24'(-36144);
			18210: out = 24'(-28008);
			18211: out = 24'(-12712);
			18212: out = 24'(-608);
			18213: out = 24'(10048);
			18214: out = 24'(21224);
			18215: out = 24'(21836);
			18216: out = 24'(9704);
			18217: out = 24'(-384);
			18218: out = 24'(-21528);
			18219: out = 24'(-10000);
			18220: out = 24'(2296);
			18221: out = 24'(-512);
			18222: out = 24'(232);
			18223: out = 24'(5172);
			18224: out = 24'(10088);
			18225: out = 24'(6200);
			18226: out = 24'(904);
			18227: out = 24'(-7612);
			18228: out = 24'(-8080);
			18229: out = 24'(-3520);
			18230: out = 24'(-628);
			18231: out = 24'(3888);
			18232: out = 24'(7200);
			18233: out = 24'(4296);
			18234: out = 24'(-15236);
			18235: out = 24'(-104);
			18236: out = 24'(-11708);
			18237: out = 24'(-12580);
			18238: out = 24'(7840);
			18239: out = 24'(22088);
			18240: out = 24'(10084);
			18241: out = 24'(-6716);
			18242: out = 24'(-4752);
			18243: out = 24'(14348);
			18244: out = 24'(22764);
			18245: out = 24'(15116);
			18246: out = 24'(-4984);
			18247: out = 24'(-26384);
			18248: out = 24'(-15512);
			18249: out = 24'(-1224);
			18250: out = 24'(-3888);
			18251: out = 24'(-10600);
			18252: out = 24'(9220);
			18253: out = 24'(31568);
			18254: out = 24'(18072);
			18255: out = 24'(-20472);
			18256: out = 24'(-19608);
			18257: out = 24'(-2728);
			18258: out = 24'(-4180);
			18259: out = 24'(-21196);
			18260: out = 24'(8112);
			18261: out = 24'(40880);
			18262: out = 24'(50740);
			18263: out = 24'(25516);
			18264: out = 24'(1164);
			18265: out = 24'(-4168);
			18266: out = 24'(-6548);
			18267: out = 24'(-19580);
			18268: out = 24'(-15724);
			18269: out = 24'(-636);
			18270: out = 24'(22836);
			18271: out = 24'(15288);
			18272: out = 24'(-12804);
			18273: out = 24'(-40592);
			18274: out = 24'(-18168);
			18275: out = 24'(6104);
			18276: out = 24'(2036);
			18277: out = 24'(5004);
			18278: out = 24'(11044);
			18279: out = 24'(11656);
			18280: out = 24'(-6808);
			18281: out = 24'(-6564);
			18282: out = 24'(-6812);
			18283: out = 24'(17236);
			18284: out = 24'(24144);
			18285: out = 24'(-1740);
			18286: out = 24'(-35240);
			18287: out = 24'(-28016);
			18288: out = 24'(11068);
			18289: out = 24'(35676);
			18290: out = 24'(37564);
			18291: out = 24'(13748);
			18292: out = 24'(-17260);
			18293: out = 24'(-37404);
			18294: out = 24'(-21840);
			18295: out = 24'(-11400);
			18296: out = 24'(-13244);
			18297: out = 24'(-16168);
			18298: out = 24'(-172);
			18299: out = 24'(22628);
			18300: out = 24'(30236);
			18301: out = 24'(16392);
			18302: out = 24'(224);
			18303: out = 24'(-9156);
			18304: out = 24'(-12192);
			18305: out = 24'(-15316);
			18306: out = 24'(-13904);
			18307: out = 24'(-29844);
			18308: out = 24'(-15876);
			18309: out = 24'(16160);
			18310: out = 24'(35088);
			18311: out = 24'(12068);
			18312: out = 24'(-18268);
			18313: out = 24'(-36028);
			18314: out = 24'(-27052);
			18315: out = 24'(-11348);
			18316: out = 24'(-9204);
			18317: out = 24'(-13984);
			18318: out = 24'(-916);
			18319: out = 24'(14352);
			18320: out = 24'(32584);
			18321: out = 24'(5444);
			18322: out = 24'(-30700);
			18323: out = 24'(-37720);
			18324: out = 24'(7400);
			18325: out = 24'(17720);
			18326: out = 24'(6332);
			18327: out = 24'(12480);
			18328: out = 24'(21372);
			18329: out = 24'(17060);
			18330: out = 24'(2344);
			18331: out = 24'(2192);
			18332: out = 24'(-2000);
			18333: out = 24'(2680);
			18334: out = 24'(-14268);
			18335: out = 24'(-30720);
			18336: out = 24'(-12644);
			18337: out = 24'(9384);
			18338: out = 24'(23372);
			18339: out = 24'(19176);
			18340: out = 24'(260);
			18341: out = 24'(7116);
			18342: out = 24'(-720);
			18343: out = 24'(-27008);
			18344: out = 24'(-53716);
			18345: out = 24'(-7884);
			18346: out = 24'(23892);
			18347: out = 24'(28476);
			18348: out = 24'(14352);
			18349: out = 24'(10188);
			18350: out = 24'(4896);
			18351: out = 24'(3220);
			18352: out = 24'(-3208);
			18353: out = 24'(-7884);
			18354: out = 24'(-10876);
			18355: out = 24'(-3500);
			18356: out = 24'(-3128);
			18357: out = 24'(-11472);
			18358: out = 24'(-12312);
			18359: out = 24'(13940);
			18360: out = 24'(29364);
			18361: out = 24'(5932);
			18362: out = 24'(1796);
			18363: out = 24'(-1684);
			18364: out = 24'(-2448);
			18365: out = 24'(-9548);
			18366: out = 24'(-1036);
			18367: out = 24'(5628);
			18368: out = 24'(6740);
			18369: out = 24'(-384);
			18370: out = 24'(9084);
			18371: out = 24'(1644);
			18372: out = 24'(-1660);
			18373: out = 24'(2176);
			18374: out = 24'(16112);
			18375: out = 24'(15692);
			18376: out = 24'(12156);
			18377: out = 24'(4352);
			18378: out = 24'(-2196);
			18379: out = 24'(-24316);
			18380: out = 24'(-23260);
			18381: out = 24'(-3244);
			18382: out = 24'(16100);
			18383: out = 24'(9084);
			18384: out = 24'(2008);
			18385: out = 24'(-1760);
			18386: out = 24'(240);
			18387: out = 24'(-1616);
			18388: out = 24'(-164);
			18389: out = 24'(2216);
			18390: out = 24'(10552);
			18391: out = 24'(13212);
			18392: out = 24'(2292);
			18393: out = 24'(-22700);
			18394: out = 24'(-22008);
			18395: out = 24'(24648);
			18396: out = 24'(43008);
			18397: out = 24'(24916);
			18398: out = 24'(-13236);
			18399: out = 24'(-31124);
			18400: out = 24'(-23484);
			18401: out = 24'(-6340);
			18402: out = 24'(4520);
			18403: out = 24'(17148);
			18404: out = 24'(13204);
			18405: out = 24'(11988);
			18406: out = 24'(-3632);
			18407: out = 24'(-16024);
			18408: out = 24'(-24780);
			18409: out = 24'(6352);
			18410: out = 24'(14304);
			18411: out = 24'(4564);
			18412: out = 24'(-656);
			18413: out = 24'(12800);
			18414: out = 24'(1056);
			18415: out = 24'(-20132);
			18416: out = 24'(-16464);
			18417: out = 24'(-5624);
			18418: out = 24'(5884);
			18419: out = 24'(7636);
			18420: out = 24'(6980);
			18421: out = 24'(-100);
			18422: out = 24'(-1740);
			18423: out = 24'(-1612);
			18424: out = 24'(-1856);
			18425: out = 24'(3004);
			18426: out = 24'(-2064);
			18427: out = 24'(6220);
			18428: out = 24'(13356);
			18429: out = 24'(-1748);
			18430: out = 24'(-25936);
			18431: out = 24'(-25576);
			18432: out = 24'(-1216);
			18433: out = 24'(6884);
			18434: out = 24'(28832);
			18435: out = 24'(17320);
			18436: out = 24'(1508);
			18437: out = 24'(-6024);
			18438: out = 24'(-1284);
			18439: out = 24'(-8880);
			18440: out = 24'(-18160);
			18441: out = 24'(-15948);
			18442: out = 24'(-1960);
			18443: out = 24'(3592);
			18444: out = 24'(604);
			18445: out = 24'(4044);
			18446: out = 24'(21688);
			18447: out = 24'(24524);
			18448: out = 24'(1220);
			18449: out = 24'(-35152);
			18450: out = 24'(-48808);
			18451: out = 24'(-13732);
			18452: out = 24'(19204);
			18453: out = 24'(16168);
			18454: out = 24'(2092);
			18455: out = 24'(18288);
			18456: out = 24'(27608);
			18457: out = 24'(3416);
			18458: out = 24'(-27328);
			18459: out = 24'(-3840);
			18460: out = 24'(27816);
			18461: out = 24'(23972);
			18462: out = 24'(-8784);
			18463: out = 24'(-12540);
			18464: out = 24'(-236);
			18465: out = 24'(10344);
			18466: out = 24'(3228);
			18467: out = 24'(-984);
			18468: out = 24'(-10616);
			18469: out = 24'(-5644);
			18470: out = 24'(1904);
			18471: out = 24'(6152);
			18472: out = 24'(-7756);
			18473: out = 24'(-12296);
			18474: out = 24'(-6396);
			18475: out = 24'(-832);
			18476: out = 24'(124);
			18477: out = 24'(-1828);
			18478: out = 24'(896);
			18479: out = 24'(-7160);
			18480: out = 24'(-28656);
			18481: out = 24'(-40180);
			18482: out = 24'(-8728);
			18483: out = 24'(30472);
			18484: out = 24'(28144);
			18485: out = 24'(3100);
			18486: out = 24'(-6976);
			18487: out = 24'(3260);
			18488: out = 24'(5900);
			18489: out = 24'(-13724);
			18490: out = 24'(-11808);
			18491: out = 24'(13732);
			18492: out = 24'(30932);
			18493: out = 24'(6412);
			18494: out = 24'(-16324);
			18495: out = 24'(-19184);
			18496: out = 24'(5936);
			18497: out = 24'(22232);
			18498: out = 24'(28156);
			18499: out = 24'(3416);
			18500: out = 24'(-13984);
			18501: out = 24'(-4224);
			18502: out = 24'(3168);
			18503: out = 24'(-25808);
			18504: out = 24'(-38840);
			18505: out = 24'(11948);
			18506: out = 24'(41336);
			18507: out = 24'(24844);
			18508: out = 24'(-5580);
			18509: out = 24'(2780);
			18510: out = 24'(17304);
			18511: out = 24'(9068);
			18512: out = 24'(-24144);
			18513: out = 24'(-38492);
			18514: out = 24'(-9952);
			18515: out = 24'(6736);
			18516: out = 24'(3992);
			18517: out = 24'(904);
			18518: out = 24'(7012);
			18519: out = 24'(8572);
			18520: out = 24'(3140);
			18521: out = 24'(-1104);
			18522: out = 24'(-1316);
			18523: out = 24'(12492);
			18524: out = 24'(8260);
			18525: out = 24'(-6944);
			18526: out = 24'(-12144);
			18527: out = 24'(9996);
			18528: out = 24'(13800);
			18529: out = 24'(-1648);
			18530: out = 24'(-8372);
			18531: out = 24'(-5452);
			18532: out = 24'(19744);
			18533: out = 24'(15316);
			18534: out = 24'(-14380);
			18535: out = 24'(-45228);
			18536: out = 24'(-10292);
			18537: out = 24'(20928);
			18538: out = 24'(15828);
			18539: out = 24'(-4708);
			18540: out = 24'(-3280);
			18541: out = 24'(-1140);
			18542: out = 24'(-14580);
			18543: out = 24'(-35400);
			18544: out = 24'(-3520);
			18545: out = 24'(18144);
			18546: out = 24'(21372);
			18547: out = 24'(14448);
			18548: out = 24'(15192);
			18549: out = 24'(4740);
			18550: out = 24'(-9964);
			18551: out = 24'(-19084);
			18552: out = 24'(-10288);
			18553: out = 24'(1576);
			18554: out = 24'(16136);
			18555: out = 24'(20248);
			18556: out = 24'(7116);
			18557: out = 24'(-13428);
			18558: out = 24'(-16144);
			18559: out = 24'(1448);
			18560: out = 24'(13236);
			18561: out = 24'(2732);
			18562: out = 24'(-11140);
			18563: out = 24'(-14404);
			18564: out = 24'(-16132);
			18565: out = 24'(-28604);
			18566: out = 24'(-19940);
			18567: out = 24'(16704);
			18568: out = 24'(43204);
			18569: out = 24'(41792);
			18570: out = 24'(900);
			18571: out = 24'(-16168);
			18572: out = 24'(-3476);
			18573: out = 24'(-2136);
			18574: out = 24'(-17408);
			18575: out = 24'(-20984);
			18576: out = 24'(-2460);
			18577: out = 24'(14056);
			18578: out = 24'(5972);
			18579: out = 24'(-584);
			18580: out = 24'(-464);
			18581: out = 24'(-1024);
			18582: out = 24'(-1500);
			18583: out = 24'(-916);
			18584: out = 24'(-800);
			18585: out = 24'(-1428);
			18586: out = 24'(-18140);
			18587: out = 24'(-7940);
			18588: out = 24'(120);
			18589: out = 24'(-1428);
			18590: out = 24'(-596);
			18591: out = 24'(11860);
			18592: out = 24'(9604);
			18593: out = 24'(-412);
			18594: out = 24'(16284);
			18595: out = 24'(8196);
			18596: out = 24'(2508);
			18597: out = 24'(-3212);
			18598: out = 24'(-716);
			18599: out = 24'(-1376);
			18600: out = 24'(-12680);
			18601: out = 24'(-29560);
			18602: out = 24'(-21620);
			18603: out = 24'(21784);
			18604: out = 24'(39832);
			18605: out = 24'(20360);
			18606: out = 24'(-5088);
			18607: out = 24'(-15836);
			18608: out = 24'(-19800);
			18609: out = 24'(-31244);
			18610: out = 24'(-24076);
			18611: out = 24'(5136);
			18612: out = 24'(28008);
			18613: out = 24'(-2612);
			18614: out = 24'(-30188);
			18615: out = 24'(7256);
			18616: out = 24'(34084);
			18617: out = 24'(23036);
			18618: out = 24'(-7480);
			18619: out = 24'(-7356);
			18620: out = 24'(-8972);
			18621: out = 24'(-1528);
			18622: out = 24'(36);
			18623: out = 24'(10480);
			18624: out = 24'(12756);
			18625: out = 24'(9196);
			18626: out = 24'(-5300);
			18627: out = 24'(-10072);
			18628: out = 24'(-16476);
			18629: out = 24'(9952);
			18630: out = 24'(8884);
			18631: out = 24'(-3028);
			18632: out = 24'(-692);
			18633: out = 24'(17808);
			18634: out = 24'(16656);
			18635: out = 24'(-3868);
			18636: out = 24'(-24688);
			18637: out = 24'(-20804);
			18638: out = 24'(-9428);
			18639: out = 24'(5832);
			18640: out = 24'(15884);
			18641: out = 24'(22736);
			18642: out = 24'(11212);
			18643: out = 24'(6076);
			18644: out = 24'(2276);
			18645: out = 24'(-23164);
			18646: out = 24'(-23376);
			18647: out = 24'(-8928);
			18648: out = 24'(-5572);
			18649: out = 24'(-32032);
			18650: out = 24'(-33992);
			18651: out = 24'(-10604);
			18652: out = 24'(15120);
			18653: out = 24'(16180);
			18654: out = 24'(32080);
			18655: out = 24'(32960);
			18656: out = 24'(17392);
			18657: out = 24'(-17368);
			18658: out = 24'(-57172);
			18659: out = 24'(-52032);
			18660: out = 24'(-15264);
			18661: out = 24'(14272);
			18662: out = 24'(37540);
			18663: out = 24'(22568);
			18664: out = 24'(7824);
			18665: out = 24'(-1696);
			18666: out = 24'(-468);
			18667: out = 24'(-19032);
			18668: out = 24'(-21548);
			18669: out = 24'(-17896);
			18670: out = 24'(-21620);
			18671: out = 24'(-2152);
			18672: out = 24'(7392);
			18673: out = 24'(9652);
			18674: out = 24'(8400);
			18675: out = 24'(-7180);
			18676: out = 24'(-3912);
			18677: out = 24'(4604);
			18678: out = 24'(7220);
			18679: out = 24'(-16616);
			18680: out = 24'(-5428);
			18681: out = 24'(3856);
			18682: out = 24'(7316);
			18683: out = 24'(16908);
			18684: out = 24'(17032);
			18685: out = 24'(12756);
			18686: out = 24'(3676);
			18687: out = 24'(-14244);
			18688: out = 24'(-1532);
			18689: out = 24'(3476);
			18690: out = 24'(17040);
			18691: out = 24'(28244);
			18692: out = 24'(23616);
			18693: out = 24'(-20144);
			18694: out = 24'(-40556);
			18695: out = 24'(-8664);
			18696: out = 24'(25964);
			18697: out = 24'(18120);
			18698: out = 24'(3588);
			18699: out = 24'(11756);
			18700: out = 24'(12804);
			18701: out = 24'(5896);
			18702: out = 24'(-6720);
			18703: out = 24'(-892);
			18704: out = 24'(5420);
			18705: out = 24'(10372);
			18706: out = 24'(-4448);
			18707: out = 24'(-3784);
			18708: out = 24'(14172);
			18709: out = 24'(3172);
			18710: out = 24'(-27272);
			18711: out = 24'(-37148);
			18712: out = 24'(-720);
			18713: out = 24'(30960);
			18714: out = 24'(27320);
			18715: out = 24'(-2528);
			18716: out = 24'(-16628);
			18717: out = 24'(-2740);
			18718: out = 24'(12984);
			18719: out = 24'(7828);
			18720: out = 24'(-3128);
			18721: out = 24'(-1224);
			18722: out = 24'(-18028);
			18723: out = 24'(-29436);
			18724: out = 24'(-18456);
			18725: out = 24'(9544);
			18726: out = 24'(28036);
			18727: out = 24'(13532);
			18728: out = 24'(-5796);
			18729: out = 24'(-4784);
			18730: out = 24'(-14848);
			18731: out = 24'(-16304);
			18732: out = 24'(-18552);
			18733: out = 24'(-10884);
			18734: out = 24'(-10932);
			18735: out = 24'(23340);
			18736: out = 24'(27812);
			18737: out = 24'(-4824);
			18738: out = 24'(-41704);
			18739: out = 24'(-3492);
			18740: out = 24'(34596);
			18741: out = 24'(4608);
			18742: out = 24'(-73352);
			18743: out = 24'(-71544);
			18744: out = 24'(-9232);
			18745: out = 24'(32272);
			18746: out = 24'(22828);
			18747: out = 24'(3952);
			18748: out = 24'(16420);
			18749: out = 24'(18196);
			18750: out = 24'(-10644);
			18751: out = 24'(-41736);
			18752: out = 24'(-5848);
			18753: out = 24'(33124);
			18754: out = 24'(27396);
			18755: out = 24'(2844);
			18756: out = 24'(412);
			18757: out = 24'(8688);
			18758: out = 24'(3532);
			18759: out = 24'(-17392);
			18760: out = 24'(-10676);
			18761: out = 24'(504);
			18762: out = 24'(17484);
			18763: out = 24'(28092);
			18764: out = 24'(7028);
			18765: out = 24'(-27340);
			18766: out = 24'(-34768);
			18767: out = 24'(-1772);
			18768: out = 24'(27740);
			18769: out = 24'(13456);
			18770: out = 24'(-5616);
			18771: out = 24'(-2524);
			18772: out = 24'(-6180);
			18773: out = 24'(-9728);
			18774: out = 24'(-6852);
			18775: out = 24'(19316);
			18776: out = 24'(36656);
			18777: out = 24'(19120);
			18778: out = 24'(-17588);
			18779: out = 24'(-28420);
			18780: out = 24'(-8976);
			18781: out = 24'(7552);
			18782: out = 24'(6948);
			18783: out = 24'(16420);
			18784: out = 24'(27828);
			18785: out = 24'(19676);
			18786: out = 24'(-29812);
			18787: out = 24'(-48456);
			18788: out = 24'(-6376);
			18789: out = 24'(28764);
			18790: out = 24'(19560);
			18791: out = 24'(-1484);
			18792: out = 24'(6184);
			18793: out = 24'(26016);
			18794: out = 24'(15016);
			18795: out = 24'(-9232);
			18796: out = 24'(-16012);
			18797: out = 24'(-1736);
			18798: out = 24'(140);
			18799: out = 24'(-6372);
			18800: out = 24'(-8076);
			18801: out = 24'(1932);
			18802: out = 24'(19524);
			18803: out = 24'(10328);
			18804: out = 24'(-10488);
			18805: out = 24'(-16836);
			18806: out = 24'(-16132);
			18807: out = 24'(3176);
			18808: out = 24'(5216);
			18809: out = 24'(-424);
			18810: out = 24'(-1128);
			18811: out = 24'(22360);
			18812: out = 24'(25004);
			18813: out = 24'(4876);
			18814: out = 24'(-22904);
			18815: out = 24'(-4740);
			18816: out = 24'(-10212);
			18817: out = 24'(-27024);
			18818: out = 24'(-18204);
			18819: out = 24'(1756);
			18820: out = 24'(24188);
			18821: out = 24'(27404);
			18822: out = 24'(18964);
			18823: out = 24'(-8236);
			18824: out = 24'(-5784);
			18825: out = 24'(300);
			18826: out = 24'(-6808);
			18827: out = 24'(-44288);
			18828: out = 24'(-27848);
			18829: out = 24'(-3216);
			18830: out = 24'(13512);
			18831: out = 24'(29848);
			18832: out = 24'(29128);
			18833: out = 24'(15332);
			18834: out = 24'(-12600);
			18835: out = 24'(-30684);
			18836: out = 24'(-51060);
			18837: out = 24'(-26976);
			18838: out = 24'(672);
			18839: out = 24'(10544);
			18840: out = 24'(21848);
			18841: out = 24'(35548);
			18842: out = 24'(32308);
			18843: out = 24'(4836);
			18844: out = 24'(-46564);
			18845: out = 24'(-37944);
			18846: out = 24'(-11084);
			18847: out = 24'(468);
			18848: out = 24'(-8064);
			18849: out = 24'(-944);
			18850: out = 24'(5260);
			18851: out = 24'(11764);
			18852: out = 24'(16128);
			18853: out = 24'(28872);
			18854: out = 24'(13788);
			18855: out = 24'(-12644);
			18856: out = 24'(-31108);
			18857: out = 24'(-23164);
			18858: out = 24'(-9600);
			18859: out = 24'(11520);
			18860: out = 24'(20688);
			18861: out = 24'(3332);
			18862: out = 24'(-12384);
			18863: out = 24'(4904);
			18864: out = 24'(31324);
			18865: out = 24'(13584);
			18866: out = 24'(-25504);
			18867: out = 24'(-43308);
			18868: out = 24'(-18064);
			18869: out = 24'(2792);
			18870: out = 24'(4796);
			18871: out = 24'(1920);
			18872: out = 24'(18832);
			18873: out = 24'(25316);
			18874: out = 24'(68);
			18875: out = 24'(-36428);
			18876: out = 24'(-30088);
			18877: out = 24'(7996);
			18878: out = 24'(9296);
			18879: out = 24'(2128);
			18880: out = 24'(9496);
			18881: out = 24'(24404);
			18882: out = 24'(15948);
			18883: out = 24'(-9308);
			18884: out = 24'(-12100);
			18885: out = 24'(4044);
			18886: out = 24'(-1372);
			18887: out = 24'(-8792);
			18888: out = 24'(-8444);
			18889: out = 24'(10512);
			18890: out = 24'(26056);
			18891: out = 24'(21424);
			18892: out = 24'(2724);
			18893: out = 24'(-19016);
			18894: out = 24'(-29208);
			18895: out = 24'(-15740);
			18896: out = 24'(3352);
			18897: out = 24'(8164);
			18898: out = 24'(2600);
			18899: out = 24'(-4504);
			18900: out = 24'(5948);
			18901: out = 24'(8332);
			18902: out = 24'(11848);
			18903: out = 24'(21412);
			18904: out = 24'(31100);
			18905: out = 24'(-3104);
			18906: out = 24'(-46780);
			18907: out = 24'(-45280);
			18908: out = 24'(-2508);
			18909: out = 24'(18768);
			18910: out = 24'(11648);
			18911: out = 24'(9840);
			18912: out = 24'(2592);
			18913: out = 24'(-5056);
			18914: out = 24'(-18600);
			18915: out = 24'(-11232);
			18916: out = 24'(4732);
			18917: out = 24'(24096);
			18918: out = 24'(5500);
			18919: out = 24'(-19160);
			18920: out = 24'(-11904);
			18921: out = 24'(21580);
			18922: out = 24'(20096);
			18923: out = 24'(-13188);
			18924: out = 24'(-36000);
			18925: out = 24'(10456);
			18926: out = 24'(37736);
			18927: out = 24'(24316);
			18928: out = 24'(-4276);
			18929: out = 24'(-36500);
			18930: out = 24'(-36932);
			18931: out = 24'(-21420);
			18932: out = 24'(-4720);
			18933: out = 24'(8528);
			18934: out = 24'(35372);
			18935: out = 24'(48928);
			18936: out = 24'(26668);
			18937: out = 24'(-13852);
			18938: out = 24'(-33432);
			18939: out = 24'(-7656);
			18940: out = 24'(15988);
			18941: out = 24'(-2576);
			18942: out = 24'(-25604);
			18943: out = 24'(-17460);
			18944: out = 24'(7232);
			18945: out = 24'(6312);
			18946: out = 24'(3328);
			18947: out = 24'(13468);
			18948: out = 24'(38340);
			18949: out = 24'(37552);
			18950: out = 24'(-3524);
			18951: out = 24'(-29464);
			18952: out = 24'(-19128);
			18953: out = 24'(1852);
			18954: out = 24'(-648);
			18955: out = 24'(-10840);
			18956: out = 24'(-4456);
			18957: out = 24'(11052);
			18958: out = 24'(6564);
			18959: out = 24'(2064);
			18960: out = 24'(-2088);
			18961: out = 24'(3108);
			18962: out = 24'(6688);
			18963: out = 24'(1084);
			18964: out = 24'(-2880);
			18965: out = 24'(2952);
			18966: out = 24'(6560);
			18967: out = 24'(1544);
			18968: out = 24'(-10132);
			18969: out = 24'(-9344);
			18970: out = 24'(2384);
			18971: out = 24'(7036);
			18972: out = 24'(2124);
			18973: out = 24'(-1944);
			18974: out = 24'(2240);
			18975: out = 24'(6680);
			18976: out = 24'(-848);
			18977: out = 24'(-15124);
			18978: out = 24'(-20484);
			18979: out = 24'(-7328);
			18980: out = 24'(-1396);
			18981: out = 24'(5820);
			18982: out = 24'(10652);
			18983: out = 24'(16384);
			18984: out = 24'(14796);
			18985: out = 24'(7212);
			18986: out = 24'(-9152);
			18987: out = 24'(-16268);
			18988: out = 24'(-11512);
			18989: out = 24'(10360);
			18990: out = 24'(9936);
			18991: out = 24'(-3524);
			18992: out = 24'(-9368);
			18993: out = 24'(5440);
			18994: out = 24'(-4748);
			18995: out = 24'(-24256);
			18996: out = 24'(-8964);
			18997: out = 24'(28848);
			18998: out = 24'(39996);
			18999: out = 24'(13528);
			19000: out = 24'(-13004);
			19001: out = 24'(-12320);
			19002: out = 24'(-76);
			19003: out = 24'(-1144);
			19004: out = 24'(-9876);
			19005: out = 24'(-9680);
			19006: out = 24'(-3248);
			19007: out = 24'(-368);
			19008: out = 24'(-976);
			19009: out = 24'(-4640);
			19010: out = 24'(25084);
			19011: out = 24'(40324);
			19012: out = 24'(22528);
			19013: out = 24'(-23320);
			19014: out = 24'(-37792);
			19015: out = 24'(-43032);
			19016: out = 24'(-31756);
			19017: out = 24'(-84);
			19018: out = 24'(32904);
			19019: out = 24'(50028);
			19020: out = 24'(41840);
			19021: out = 24'(16000);
			19022: out = 24'(-14288);
			19023: out = 24'(-19908);
			19024: out = 24'(-4172);
			19025: out = 24'(4104);
			19026: out = 24'(-16520);
			19027: out = 24'(-21300);
			19028: out = 24'(-3200);
			19029: out = 24'(18308);
			19030: out = 24'(17684);
			19031: out = 24'(15356);
			19032: out = 24'(15804);
			19033: out = 24'(14832);
			19034: out = 24'(-812);
			19035: out = 24'(-26080);
			19036: out = 24'(-36120);
			19037: out = 24'(-24548);
			19038: out = 24'(-8532);
			19039: out = 24'(-936);
			19040: out = 24'(13460);
			19041: out = 24'(27208);
			19042: out = 24'(18000);
			19043: out = 24'(-22440);
			19044: out = 24'(-30072);
			19045: out = 24'(-1356);
			19046: out = 24'(21200);
			19047: out = 24'(-1172);
			19048: out = 24'(-2352);
			19049: out = 24'(10960);
			19050: out = 24'(19260);
			19051: out = 24'(-4320);
			19052: out = 24'(-15216);
			19053: out = 24'(-18796);
			19054: out = 24'(-11300);
			19055: out = 24'(-11132);
			19056: out = 24'(-11988);
			19057: out = 24'(-10672);
			19058: out = 24'(4004);
			19059: out = 24'(15576);
			19060: out = 24'(16212);
			19061: out = 24'(5840);
			19062: out = 24'(1812);
			19063: out = 24'(-5416);
			19064: out = 24'(-29404);
			19065: out = 24'(-51364);
			19066: out = 24'(-37568);
			19067: out = 24'(5704);
			19068: out = 24'(24856);
			19069: out = 24'(27432);
			19070: out = 24'(16896);
			19071: out = 24'(18508);
			19072: out = 24'(15520);
			19073: out = 24'(5388);
			19074: out = 24'(-38676);
			19075: out = 24'(-60924);
			19076: out = 24'(-30748);
			19077: out = 24'(17680);
			19078: out = 24'(23808);
			19079: out = 24'(7576);
			19080: out = 24'(4196);
			19081: out = 24'(25664);
			19082: out = 24'(20612);
			19083: out = 24'(5528);
			19084: out = 24'(-8556);
			19085: out = 24'(-17152);
			19086: out = 24'(-14796);
			19087: out = 24'(-6212);
			19088: out = 24'(2848);
			19089: out = 24'(10580);
			19090: out = 24'(34872);
			19091: out = 24'(38532);
			19092: out = 24'(20036);
			19093: out = 24'(-2748);
			19094: out = 24'(-14088);
			19095: out = 24'(-9028);
			19096: out = 24'(-5600);
			19097: out = 24'(-6024);
			19098: out = 24'(-14524);
			19099: out = 24'(7684);
			19100: out = 24'(14424);
			19101: out = 24'(1488);
			19102: out = 24'(-22184);
			19103: out = 24'(1080);
			19104: out = 24'(6220);
			19105: out = 24'(-3124);
			19106: out = 24'(-4296);
			19107: out = 24'(5700);
			19108: out = 24'(3852);
			19109: out = 24'(364);
			19110: out = 24'(9408);
			19111: out = 24'(20328);
			19112: out = 24'(9116);
			19113: out = 24'(-10180);
			19114: out = 24'(-17336);
			19115: out = 24'(-2728);
			19116: out = 24'(4272);
			19117: out = 24'(16672);
			19118: out = 24'(28952);
			19119: out = 24'(19888);
			19120: out = 24'(1060);
			19121: out = 24'(-19460);
			19122: out = 24'(-32404);
			19123: out = 24'(-40944);
			19124: out = 24'(-23772);
			19125: out = 24'(1884);
			19126: out = 24'(20716);
			19127: out = 24'(21540);
			19128: out = 24'(23116);
			19129: out = 24'(7852);
			19130: out = 24'(-10236);
			19131: out = 24'(-16956);
			19132: out = 24'(-3824);
			19133: out = 24'(11288);
			19134: out = 24'(9676);
			19135: out = 24'(-3572);
			19136: out = 24'(-4616);
			19137: out = 24'(-2860);
			19138: out = 24'(3884);
			19139: out = 24'(6068);
			19140: out = 24'(-1080);
			19141: out = 24'(-1008);
			19142: out = 24'(-3924);
			19143: out = 24'(-7828);
			19144: out = 24'(-14844);
			19145: out = 24'(-16952);
			19146: out = 24'(-5488);
			19147: out = 24'(24472);
			19148: out = 24'(40224);
			19149: out = 24'(3980);
			19150: out = 24'(-31420);
			19151: out = 24'(-34020);
			19152: out = 24'(-10200);
			19153: out = 24'(-9684);
			19154: out = 24'(-3092);
			19155: out = 24'(18336);
			19156: out = 24'(41356);
			19157: out = 24'(25640);
			19158: out = 24'(7300);
			19159: out = 24'(-12664);
			19160: out = 24'(-23216);
			19161: out = 24'(-41624);
			19162: out = 24'(-9580);
			19163: out = 24'(3260);
			19164: out = 24'(12028);
			19165: out = 24'(15220);
			19166: out = 24'(29712);
			19167: out = 24'(1372);
			19168: out = 24'(-17324);
			19169: out = 24'(-5356);
			19170: out = 24'(5148);
			19171: out = 24'(-10812);
			19172: out = 24'(-29964);
			19173: out = 24'(-17848);
			19174: out = 24'(5236);
			19175: out = 24'(23556);
			19176: out = 24'(10300);
			19177: out = 24'(2512);
			19178: out = 24'(14452);
			19179: out = 24'(17520);
			19180: out = 24'(-10860);
			19181: out = 24'(-33720);
			19182: out = 24'(-18408);
			19183: out = 24'(-404);
			19184: out = 24'(-1864);
			19185: out = 24'(-8936);
			19186: out = 24'(6168);
			19187: out = 24'(22556);
			19188: out = 24'(24968);
			19189: out = 24'(4004);
			19190: out = 24'(-16472);
			19191: out = 24'(-22356);
			19192: out = 24'(-12788);
			19193: out = 24'(-4348);
			19194: out = 24'(500);
			19195: out = 24'(1212);
			19196: out = 24'(29880);
			19197: out = 24'(29288);
			19198: out = 24'(-2176);
			19199: out = 24'(-39284);
			19200: out = 24'(-8068);
			19201: out = 24'(8496);
			19202: out = 24'(2836);
			19203: out = 24'(-3032);
			19204: out = 24'(5412);
			19205: out = 24'(19980);
			19206: out = 24'(14296);
			19207: out = 24'(-3632);
			19208: out = 24'(-12920);
			19209: out = 24'(11416);
			19210: out = 24'(26420);
			19211: out = 24'(12160);
			19212: out = 24'(-22004);
			19213: out = 24'(-11412);
			19214: out = 24'(-1192);
			19215: out = 24'(-5456);
			19216: out = 24'(-12556);
			19217: out = 24'(3224);
			19218: out = 24'(16088);
			19219: out = 24'(13420);
			19220: out = 24'(-3144);
			19221: out = 24'(-12276);
			19222: out = 24'(-10788);
			19223: out = 24'(-2120);
			19224: out = 24'(-3192);
			19225: out = 24'(412);
			19226: out = 24'(1856);
			19227: out = 24'(19568);
			19228: out = 24'(24128);
			19229: out = 24'(8648);
			19230: out = 24'(-23332);
			19231: out = 24'(-8996);
			19232: out = 24'(17556);
			19233: out = 24'(2784);
			19234: out = 24'(-48188);
			19235: out = 24'(-49312);
			19236: out = 24'(-2964);
			19237: out = 24'(11556);
			19238: out = 24'(6572);
			19239: out = 24'(-1324);
			19240: out = 24'(28456);
			19241: out = 24'(44760);
			19242: out = 24'(13772);
			19243: out = 24'(-56356);
			19244: out = 24'(-66508);
			19245: out = 24'(-3116);
			19246: out = 24'(2496);
			19247: out = 24'(14628);
			19248: out = 24'(-24);
			19249: out = 24'(10220);
			19250: out = 24'(25760);
			19251: out = 24'(33012);
			19252: out = 24'(-12616);
			19253: out = 24'(-35808);
			19254: out = 24'(2764);
			19255: out = 24'(13988);
			19256: out = 24'(-728);
			19257: out = 24'(-10760);
			19258: out = 24'(14544);
			19259: out = 24'(34660);
			19260: out = 24'(28436);
			19261: out = 24'(4300);
			19262: out = 24'(-12760);
			19263: out = 24'(-22912);
			19264: out = 24'(-29972);
			19265: out = 24'(-23720);
			19266: out = 24'(-1496);
			19267: out = 24'(14456);
			19268: out = 24'(16764);
			19269: out = 24'(10800);
			19270: out = 24'(5432);
			19271: out = 24'(-1012);
			19272: out = 24'(-568);
			19273: out = 24'(-732);
			19274: out = 24'(-3024);
			19275: out = 24'(-10172);
			19276: out = 24'(-1692);
			19277: out = 24'(-696);
			19278: out = 24'(-328);
			19279: out = 24'(124);
			19280: out = 24'(14976);
			19281: out = 24'(4176);
			19282: out = 24'(-5500);
			19283: out = 24'(-9968);
			19284: out = 24'(-4768);
			19285: out = 24'(-9584);
			19286: out = 24'(-1064);
			19287: out = 24'(11228);
			19288: out = 24'(15288);
			19289: out = 24'(26700);
			19290: out = 24'(19004);
			19291: out = 24'(-7108);
			19292: out = 24'(-31320);
			19293: out = 24'(-26176);
			19294: out = 24'(-6576);
			19295: out = 24'(-3464);
			19296: out = 24'(-14604);
			19297: out = 24'(-22212);
			19298: out = 24'(11696);
			19299: out = 24'(27908);
			19300: out = 24'(4132);
			19301: out = 24'(-36900);
			19302: out = 24'(-14200);
			19303: out = 24'(10460);
			19304: out = 24'(-212);
			19305: out = 24'(-19196);
			19306: out = 24'(-28708);
			19307: out = 24'(-5672);
			19308: out = 24'(12132);
			19309: out = 24'(7380);
			19310: out = 24'(-9076);
			19311: out = 24'(-13400);
			19312: out = 24'(-10272);
			19313: out = 24'(-6372);
			19314: out = 24'(1108);
			19315: out = 24'(7724);
			19316: out = 24'(9936);
			19317: out = 24'(10600);
			19318: out = 24'(16084);
			19319: out = 24'(11960);
			19320: out = 24'(1792);
			19321: out = 24'(-3384);
			19322: out = 24'(3580);
			19323: out = 24'(2212);
			19324: out = 24'(-1056);
			19325: out = 24'(3068);
			19326: out = 24'(8664);
			19327: out = 24'(28560);
			19328: out = 24'(12220);
			19329: out = 24'(-6596);
			19330: out = 24'(-9428);
			19331: out = 24'(-8752);
			19332: out = 24'(-19020);
			19333: out = 24'(-9960);
			19334: out = 24'(22336);
			19335: out = 24'(30148);
			19336: out = 24'(26836);
			19337: out = 24'(18156);
			19338: out = 24'(17052);
			19339: out = 24'(4804);
			19340: out = 24'(-5720);
			19341: out = 24'(-13928);
			19342: out = 24'(-5976);
			19343: out = 24'(240);
			19344: out = 24'(260);
			19345: out = 24'(3428);
			19346: out = 24'(29132);
			19347: out = 24'(44464);
			19348: out = 24'(13464);
			19349: out = 24'(-38108);
			19350: out = 24'(-53808);
			19351: out = 24'(-20940);
			19352: out = 24'(3988);
			19353: out = 24'(2352);
			19354: out = 24'(6224);
			19355: out = 24'(26068);
			19356: out = 24'(25184);
			19357: out = 24'(7132);
			19358: out = 24'(-11960);
			19359: out = 24'(-15956);
			19360: out = 24'(-25504);
			19361: out = 24'(-14868);
			19362: out = 24'(-13436);
			19363: out = 24'(-3784);
			19364: out = 24'(8100);
			19365: out = 24'(24584);
			19366: out = 24'(14212);
			19367: out = 24'(2304);
			19368: out = 24'(-3944);
			19369: out = 24'(-13496);
			19370: out = 24'(-27004);
			19371: out = 24'(-31728);
			19372: out = 24'(-23892);
			19373: out = 24'(-9012);
			19374: out = 24'(-2392);
			19375: out = 24'(13624);
			19376: out = 24'(27172);
			19377: out = 24'(13308);
			19378: out = 24'(60);
			19379: out = 24'(-12128);
			19380: out = 24'(-13036);
			19381: out = 24'(-14020);
			19382: out = 24'(-4588);
			19383: out = 24'(-3220);
			19384: out = 24'(12552);
			19385: out = 24'(38904);
			19386: out = 24'(43324);
			19387: out = 24'(3900);
			19388: out = 24'(-51228);
			19389: out = 24'(-68532);
			19390: out = 24'(-22944);
			19391: out = 24'(1892);
			19392: out = 24'(-19320);
			19393: out = 24'(-41440);
			19394: out = 24'(-5152);
			19395: out = 24'(26280);
			19396: out = 24'(33740);
			19397: out = 24'(15644);
			19398: out = 24'(704);
			19399: out = 24'(-26004);
			19400: out = 24'(-24624);
			19401: out = 24'(-4692);
			19402: out = 24'(14300);
			19403: out = 24'(11012);
			19404: out = 24'(3784);
			19405: out = 24'(7040);
			19406: out = 24'(16864);
			19407: out = 24'(884);
			19408: out = 24'(6068);
			19409: out = 24'(13848);
			19410: out = 24'(11936);
			19411: out = 24'(-11852);
			19412: out = 24'(-23588);
			19413: out = 24'(-14376);
			19414: out = 24'(10272);
			19415: out = 24'(22516);
			19416: out = 24'(22060);
			19417: out = 24'(18200);
			19418: out = 24'(20056);
			19419: out = 24'(10808);
			19420: out = 24'(-22568);
			19421: out = 24'(-31780);
			19422: out = 24'(-996);
			19423: out = 24'(25692);
			19424: out = 24'(19016);
			19425: out = 24'(-4544);
			19426: out = 24'(4392);
			19427: out = 24'(29804);
			19428: out = 24'(38124);
			19429: out = 24'(-10860);
			19430: out = 24'(-26228);
			19431: out = 24'(360);
			19432: out = 24'(19792);
			19433: out = 24'(-5892);
			19434: out = 24'(-11656);
			19435: out = 24'(4068);
			19436: out = 24'(4928);
			19437: out = 24'(-6224);
			19438: out = 24'(-6924);
			19439: out = 24'(6184);
			19440: out = 24'(13668);
			19441: out = 24'(7896);
			19442: out = 24'(1192);
			19443: out = 24'(-7528);
			19444: out = 24'(-14100);
			19445: out = 24'(-6392);
			19446: out = 24'(9036);
			19447: out = 24'(16132);
			19448: out = 24'(11036);
			19449: out = 24'(-2424);
			19450: out = 24'(-1480);
			19451: out = 24'(-10888);
			19452: out = 24'(-16968);
			19453: out = 24'(176);
			19454: out = 24'(17756);
			19455: out = 24'(11832);
			19456: out = 24'(-11132);
			19457: out = 24'(-20588);
			19458: out = 24'(-4960);
			19459: out = 24'(6788);
			19460: out = 24'(3668);
			19461: out = 24'(-2128);
			19462: out = 24'(-9604);
			19463: out = 24'(-19640);
			19464: out = 24'(-28336);
			19465: out = 24'(-11472);
			19466: out = 24'(18804);
			19467: out = 24'(38408);
			19468: out = 24'(16820);
			19469: out = 24'(-10744);
			19470: out = 24'(-17392);
			19471: out = 24'(4132);
			19472: out = 24'(-8864);
			19473: out = 24'(-28412);
			19474: out = 24'(-12528);
			19475: out = 24'(19420);
			19476: out = 24'(16192);
			19477: out = 24'(-2128);
			19478: out = 24'(2588);
			19479: out = 24'(-2588);
			19480: out = 24'(-2980);
			19481: out = 24'(-18316);
			19482: out = 24'(-22484);
			19483: out = 24'(-11024);
			19484: out = 24'(3176);
			19485: out = 24'(-9456);
			19486: out = 24'(-24508);
			19487: out = 24'(-2068);
			19488: out = 24'(24040);
			19489: out = 24'(36504);
			19490: out = 24'(21916);
			19491: out = 24'(-1816);
			19492: out = 24'(-20072);
			19493: out = 24'(-13544);
			19494: out = 24'(-1312);
			19495: out = 24'(-88);
			19496: out = 24'(7484);
			19497: out = 24'(13860);
			19498: out = 24'(19332);
			19499: out = 24'(8504);
			19500: out = 24'(-14108);
			19501: out = 24'(-33996);
			19502: out = 24'(-15196);
			19503: out = 24'(23772);
			19504: out = 24'(31404);
			19505: out = 24'(9628);
			19506: out = 24'(-18636);
			19507: out = 24'(-21616);
			19508: out = 24'(-896);
			19509: out = 24'(144);
			19510: out = 24'(3144);
			19511: out = 24'(11160);
			19512: out = 24'(12580);
			19513: out = 24'(2056);
			19514: out = 24'(992);
			19515: out = 24'(15824);
			19516: out = 24'(21076);
			19517: out = 24'(9336);
			19518: out = 24'(-16852);
			19519: out = 24'(-15604);
			19520: out = 24'(424);
			19521: out = 24'(-1896);
			19522: out = 24'(-19148);
			19523: out = 24'(-7240);
			19524: out = 24'(20096);
			19525: out = 24'(14172);
			19526: out = 24'(484);
			19527: out = 24'(-15832);
			19528: out = 24'(-15872);
			19529: out = 24'(-9168);
			19530: out = 24'(-1156);
			19531: out = 24'(-144);
			19532: out = 24'(-732);
			19533: out = 24'(580);
			19534: out = 24'(6204);
			19535: out = 24'(19280);
			19536: out = 24'(27224);
			19537: out = 24'(23700);
			19538: out = 24'(5332);
			19539: out = 24'(-20272);
			19540: out = 24'(-47956);
			19541: out = 24'(-45228);
			19542: out = 24'(-512);
			19543: out = 24'(8400);
			19544: out = 24'(-3980);
			19545: out = 24'(-9484);
			19546: out = 24'(9280);
			19547: out = 24'(14896);
			19548: out = 24'(-10112);
			19549: out = 24'(-34552);
			19550: out = 24'(-13284);
			19551: out = 24'(8944);
			19552: out = 24'(32108);
			19553: out = 24'(18660);
			19554: out = 24'(-1944);
			19555: out = 24'(-5884);
			19556: out = 24'(-2952);
			19557: out = 24'(-19016);
			19558: out = 24'(-31260);
			19559: out = 24'(792);
			19560: out = 24'(1076);
			19561: out = 24'(-3668);
			19562: out = 24'(-5404);
			19563: out = 24'(10284);
			19564: out = 24'(7756);
			19565: out = 24'(6648);
			19566: out = 24'(1440);
			19567: out = 24'(1412);
			19568: out = 24'(-944);
			19569: out = 24'(2572);
			19570: out = 24'(-13420);
			19571: out = 24'(-40816);
			19572: out = 24'(-23524);
			19573: out = 24'(13800);
			19574: out = 24'(52384);
			19575: out = 24'(47860);
			19576: out = 24'(20660);
			19577: out = 24'(-37156);
			19578: out = 24'(-40364);
			19579: out = 24'(-13252);
			19580: out = 24'(-52);
			19581: out = 24'(-4864);
			19582: out = 24'(27604);
			19583: out = 24'(58064);
			19584: out = 24'(41536);
			19585: out = 24'(6820);
			19586: out = 24'(-18576);
			19587: out = 24'(-22588);
			19588: out = 24'(-22444);
			19589: out = 24'(-17196);
			19590: out = 24'(-12016);
			19591: out = 24'(-5796);
			19592: out = 24'(-3752);
			19593: out = 24'(1688);
			19594: out = 24'(26372);
			19595: out = 24'(37816);
			19596: out = 24'(21436);
			19597: out = 24'(-600);
			19598: out = 24'(-14252);
			19599: out = 24'(-6300);
			19600: out = 24'(-5592);
			19601: out = 24'(-17760);
			19602: out = 24'(-11272);
			19603: out = 24'(6584);
			19604: out = 24'(14468);
			19605: out = 24'(5088);
			19606: out = 24'(564);
			19607: out = 24'(-3436);
			19608: out = 24'(-12112);
			19609: out = 24'(-20028);
			19610: out = 24'(4096);
			19611: out = 24'(6684);
			19612: out = 24'(4804);
			19613: out = 24'(-544);
			19614: out = 24'(8624);
			19615: out = 24'(56);
			19616: out = 24'(164);
			19617: out = 24'(-1328);
			19618: out = 24'(-856);
			19619: out = 24'(-20296);
			19620: out = 24'(-9696);
			19621: out = 24'(4936);
			19622: out = 24'(6988);
			19623: out = 24'(140);
			19624: out = 24'(1192);
			19625: out = 24'(5288);
			19626: out = 24'(7520);
			19627: out = 24'(-908);
			19628: out = 24'(1648);
			19629: out = 24'(-11896);
			19630: out = 24'(-23356);
			19631: out = 24'(4432);
			19632: out = 24'(12716);
			19633: out = 24'(12764);
			19634: out = 24'(6096);
			19635: out = 24'(6648);
			19636: out = 24'(-31236);
			19637: out = 24'(-43820);
			19638: out = 24'(-26048);
			19639: out = 24'(3296);
			19640: out = 24'(12332);
			19641: out = 24'(168);
			19642: out = 24'(-4900);
			19643: out = 24'(14236);
			19644: out = 24'(26312);
			19645: out = 24'(17524);
			19646: out = 24'(132);
			19647: out = 24'(4472);
			19648: out = 24'(11148);
			19649: out = 24'(-2992);
			19650: out = 24'(-51364);
			19651: out = 24'(-63632);
			19652: out = 24'(11940);
			19653: out = 24'(35840);
			19654: out = 24'(18848);
			19655: out = 24'(-13036);
			19656: out = 24'(-12488);
			19657: out = 24'(-4080);
			19658: out = 24'(5720);
			19659: out = 24'(1168);
			19660: out = 24'(3640);
			19661: out = 24'(16824);
			19662: out = 24'(26352);
			19663: out = 24'(18448);
			19664: out = 24'(5420);
			19665: out = 24'(-4388);
			19666: out = 24'(14724);
			19667: out = 24'(21840);
			19668: out = 24'(5660);
			19669: out = 24'(-20024);
			19670: out = 24'(4780);
			19671: out = 24'(24660);
			19672: out = 24'(14572);
			19673: out = 24'(-9456);
			19674: out = 24'(-4732);
			19675: out = 24'(19640);
			19676: out = 24'(23776);
			19677: out = 24'(-8436);
			19678: out = 24'(-34976);
			19679: out = 24'(-20964);
			19680: out = 24'(21444);
			19681: out = 24'(30864);
			19682: out = 24'(11048);
			19683: out = 24'(-31612);
			19684: out = 24'(-26524);
			19685: out = 24'(2504);
			19686: out = 24'(-2036);
			19687: out = 24'(-20780);
			19688: out = 24'(-16900);
			19689: out = 24'(9328);
			19690: out = 24'(20464);
			19691: out = 24'(28200);
			19692: out = 24'(16612);
			19693: out = 24'(-6092);
			19694: out = 24'(-31412);
			19695: out = 24'(-16356);
			19696: out = 24'(-4204);
			19697: out = 24'(-7676);
			19698: out = 24'(-22204);
			19699: out = 24'(-4992);
			19700: out = 24'(-7056);
			19701: out = 24'(-12788);
			19702: out = 24'(-13440);
			19703: out = 24'(8464);
			19704: out = 24'(2952);
			19705: out = 24'(-2164);
			19706: out = 24'(-3028);
			19707: out = 24'(752);
			19708: out = 24'(456);
			19709: out = 24'(1088);
			19710: out = 24'(6472);
			19711: out = 24'(6828);
			19712: out = 24'(3484);
			19713: out = 24'(-14560);
			19714: out = 24'(-15068);
			19715: out = 24'(2792);
			19716: out = 24'(708);
			19717: out = 24'(-13020);
			19718: out = 24'(-18956);
			19719: out = 24'(1684);
			19720: out = 24'(33600);
			19721: out = 24'(18468);
			19722: out = 24'(-8472);
			19723: out = 24'(-17860);
			19724: out = 24'(1172);
			19725: out = 24'(-15824);
			19726: out = 24'(-20844);
			19727: out = 24'(-4628);
			19728: out = 24'(24668);
			19729: out = 24'(10028);
			19730: out = 24'(8956);
			19731: out = 24'(5980);
			19732: out = 24'(-1136);
			19733: out = 24'(-11748);
			19734: out = 24'(-3428);
			19735: out = 24'(2048);
			19736: out = 24'(124);
			19737: out = 24'(1044);
			19738: out = 24'(17428);
			19739: out = 24'(18884);
			19740: out = 24'(3112);
			19741: out = 24'(-2856);
			19742: out = 24'(-6004);
			19743: out = 24'(-872);
			19744: out = 24'(1844);
			19745: out = 24'(8312);
			19746: out = 24'(-13732);
			19747: out = 24'(-15320);
			19748: out = 24'(-9576);
			19749: out = 24'(-1060);
			19750: out = 24'(19848);
			19751: out = 24'(34600);
			19752: out = 24'(34600);
			19753: out = 24'(20872);
			19754: out = 24'(8396);
			19755: out = 24'(-11600);
			19756: out = 24'(-17904);
			19757: out = 24'(-4208);
			19758: out = 24'(5080);
			19759: out = 24'(23244);
			19760: out = 24'(12076);
			19761: out = 24'(-3792);
			19762: out = 24'(-1180);
			19763: out = 24'(5324);
			19764: out = 24'(2128);
			19765: out = 24'(1580);
			19766: out = 24'(16176);
			19767: out = 24'(33788);
			19768: out = 24'(7312);
			19769: out = 24'(-31948);
			19770: out = 24'(-33736);
			19771: out = 24'(3588);
			19772: out = 24'(29080);
			19773: out = 24'(15916);
			19774: out = 24'(-5068);
			19775: out = 24'(-3064);
			19776: out = 24'(9984);
			19777: out = 24'(3444);
			19778: out = 24'(-18396);
			19779: out = 24'(-30232);
			19780: out = 24'(-9232);
			19781: out = 24'(5168);
			19782: out = 24'(6492);
			19783: out = 24'(9684);
			19784: out = 24'(-8620);
			19785: out = 24'(-13464);
			19786: out = 24'(-13800);
			19787: out = 24'(-9696);
			19788: out = 24'(-18628);
			19789: out = 24'(-3992);
			19790: out = 24'(2992);
			19791: out = 24'(-2356);
			19792: out = 24'(3336);
			19793: out = 24'(1708);
			19794: out = 24'(1508);
			19795: out = 24'(-2312);
			19796: out = 24'(3676);
			19797: out = 24'(-5376);
			19798: out = 24'(-4260);
			19799: out = 24'(-8708);
			19800: out = 24'(-10488);
			19801: out = 24'(1600);
			19802: out = 24'(32908);
			19803: out = 24'(34168);
			19804: out = 24'(1380);
			19805: out = 24'(-15712);
			19806: out = 24'(-24400);
			19807: out = 24'(-32964);
			19808: out = 24'(-34176);
			19809: out = 24'(5500);
			19810: out = 24'(21164);
			19811: out = 24'(12136);
			19812: out = 24'(-1236);
			19813: out = 24'(7972);
			19814: out = 24'(21988);
			19815: out = 24'(16856);
			19816: out = 24'(3004);
			19817: out = 24'(-1516);
			19818: out = 24'(-7372);
			19819: out = 24'(-19576);
			19820: out = 24'(-12056);
			19821: out = 24'(16812);
			19822: out = 24'(21316);
			19823: out = 24'(-852);
			19824: out = 24'(-16172);
			19825: out = 24'(-8208);
			19826: out = 24'(-9800);
			19827: out = 24'(-24348);
			19828: out = 24'(-18404);
			19829: out = 24'(20112);
			19830: out = 24'(42860);
			19831: out = 24'(32824);
			19832: out = 24'(8076);
			19833: out = 24'(-3792);
			19834: out = 24'(-7164);
			19835: out = 24'(-2184);
			19836: out = 24'(-3524);
			19837: out = 24'(2552);
			19838: out = 24'(13788);
			19839: out = 24'(13564);
			19840: out = 24'(956);
			19841: out = 24'(-8464);
			19842: out = 24'(152);
			19843: out = 24'(3364);
			19844: out = 24'(8004);
			19845: out = 24'(-1208);
			19846: out = 24'(-4428);
			19847: out = 24'(4184);
			19848: out = 24'(28584);
			19849: out = 24'(17800);
			19850: out = 24'(-11644);
			19851: out = 24'(-21564);
			19852: out = 24'(4920);
			19853: out = 24'(9364);
			19854: out = 24'(-13412);
			19855: out = 24'(-29744);
			19856: out = 24'(-15352);
			19857: out = 24'(-2124);
			19858: out = 24'(-316);
			19859: out = 24'(10652);
			19860: out = 24'(19728);
			19861: out = 24'(32048);
			19862: out = 24'(9036);
			19863: out = 24'(-30088);
			19864: out = 24'(-43856);
			19865: out = 24'(-15248);
			19866: out = 24'(10136);
			19867: out = 24'(14428);
			19868: out = 24'(24524);
			19869: out = 24'(2896);
			19870: out = 24'(-15820);
			19871: out = 24'(-29660);
			19872: out = 24'(-19800);
			19873: out = 24'(-17552);
			19874: out = 24'(1188);
			19875: out = 24'(5600);
			19876: out = 24'(376);
			19877: out = 24'(1052);
			19878: out = 24'(18456);
			19879: out = 24'(20124);
			19880: out = 24'(3052);
			19881: out = 24'(-8700);
			19882: out = 24'(-7020);
			19883: out = 24'(-13236);
			19884: out = 24'(-28680);
			19885: out = 24'(-20120);
			19886: out = 24'(-16508);
			19887: out = 24'(1044);
			19888: out = 24'(24216);
			19889: out = 24'(41740);
			19890: out = 24'(21212);
			19891: out = 24'(-11544);
			19892: out = 24'(-38040);
			19893: out = 24'(-41256);
			19894: out = 24'(-10384);
			19895: out = 24'(9908);
			19896: out = 24'(19020);
			19897: out = 24'(19940);
			19898: out = 24'(1040);
			19899: out = 24'(-7952);
			19900: out = 24'(-5424);
			19901: out = 24'(-1136);
			19902: out = 24'(-12236);
			19903: out = 24'(-26012);
			19904: out = 24'(-18544);
			19905: out = 24'(10312);
			19906: out = 24'(23176);
			19907: out = 24'(14432);
			19908: out = 24'(-76);
			19909: out = 24'(6756);
			19910: out = 24'(16228);
			19911: out = 24'(18824);
			19912: out = 24'(-20304);
			19913: out = 24'(-46148);
			19914: out = 24'(-22228);
			19915: out = 24'(9620);
			19916: out = 24'(29904);
			19917: out = 24'(27492);
			19918: out = 24'(14260);
			19919: out = 24'(-3320);
			19920: out = 24'(-23652);
			19921: out = 24'(-27548);
			19922: out = 24'(-11248);
			19923: out = 24'(-532);
			19924: out = 24'(18964);
			19925: out = 24'(19888);
			19926: out = 24'(13464);
			19927: out = 24'(15500);
			19928: out = 24'(13280);
			19929: out = 24'(15336);
			19930: out = 24'(8860);
			19931: out = 24'(-4140);
			19932: out = 24'(-32536);
			19933: out = 24'(-24344);
			19934: out = 24'(-8988);
			19935: out = 24'(-9788);
			19936: out = 24'(820);
			19937: out = 24'(15480);
			19938: out = 24'(34320);
			19939: out = 24'(31120);
			19940: out = 24'(11800);
			19941: out = 24'(-10988);
			19942: out = 24'(-11720);
			19943: out = 24'(-6320);
			19944: out = 24'(-5488);
			19945: out = 24'(-3940);
			19946: out = 24'(12008);
			19947: out = 24'(18220);
			19948: out = 24'(3916);
			19949: out = 24'(-12332);
			19950: out = 24'(-15480);
			19951: out = 24'(-13800);
			19952: out = 24'(-7768);
			19953: out = 24'(-3668);
			19954: out = 24'(12304);
			19955: out = 24'(408);
			19956: out = 24'(-27188);
			19957: out = 24'(-39384);
			19958: out = 24'(2592);
			19959: out = 24'(26616);
			19960: out = 24'(22080);
			19961: out = 24'(13024);
			19962: out = 24'(-5488);
			19963: out = 24'(-41200);
			19964: out = 24'(-49964);
			19965: out = 24'(4912);
			19966: out = 24'(29884);
			19967: out = 24'(26344);
			19968: out = 24'(8716);
			19969: out = 24'(8332);
			19970: out = 24'(6120);
			19971: out = 24'(-7952);
			19972: out = 24'(-20856);
			19973: out = 24'(-6608);
			19974: out = 24'(14676);
			19975: out = 24'(23624);
			19976: out = 24'(8600);
			19977: out = 24'(-8104);
			19978: out = 24'(-5252);
			19979: out = 24'(-9696);
			19980: out = 24'(-7940);
			19981: out = 24'(-2600);
			19982: out = 24'(7152);
			19983: out = 24'(-18388);
			19984: out = 24'(-12192);
			19985: out = 24'(9504);
			19986: out = 24'(20056);
			19987: out = 24'(2036);
			19988: out = 24'(-2200);
			19989: out = 24'(2732);
			19990: out = 24'(6380);
			19991: out = 24'(-592);
			19992: out = 24'(-4056);
			19993: out = 24'(-8148);
			19994: out = 24'(-10640);
			19995: out = 24'(-18204);
			19996: out = 24'(-1408);
			19997: out = 24'(2740);
			19998: out = 24'(-684);
			19999: out = 24'(60);
			20000: out = 24'(372);
			20001: out = 24'(2876);
			20002: out = 24'(15924);
			20003: out = 24'(30724);
			20004: out = 24'(23252);
			20005: out = 24'(3508);
			20006: out = 24'(-11944);
			20007: out = 24'(-19916);
			20008: out = 24'(-20820);
			20009: out = 24'(-22360);
			20010: out = 24'(1692);
			20011: out = 24'(24496);
			20012: out = 24'(-512);
			20013: out = 24'(-7976);
			20014: out = 24'(-1660);
			20015: out = 24'(6080);
			20016: out = 24'(-9856);
			20017: out = 24'(-2332);
			20018: out = 24'(9220);
			20019: out = 24'(7896);
			20020: out = 24'(-20616);
			20021: out = 24'(-28412);
			20022: out = 24'(-9724);
			20023: out = 24'(17484);
			20024: out = 24'(15688);
			20025: out = 24'(24956);
			20026: out = 24'(-3968);
			20027: out = 24'(-14184);
			20028: out = 24'(-5368);
			20029: out = 24'(18204);
			20030: out = 24'(-2328);
			20031: out = 24'(-10240);
			20032: out = 24'(292);
			20033: out = 24'(18012);
			20034: out = 24'(2300);
			20035: out = 24'(-2412);
			20036: out = 24'(3064);
			20037: out = 24'(14184);
			20038: out = 24'(-10928);
			20039: out = 24'(-7680);
			20040: out = 24'(2236);
			20041: out = 24'(5496);
			20042: out = 24'(-28592);
			20043: out = 24'(-11952);
			20044: out = 24'(2136);
			20045: out = 24'(840);
			20046: out = 24'(6504);
			20047: out = 24'(20548);
			20048: out = 24'(788);
			20049: out = 24'(-35308);
			20050: out = 24'(-22644);
			20051: out = 24'(10236);
			20052: out = 24'(23200);
			20053: out = 24'(2148);
			20054: out = 24'(-5192);
			20055: out = 24'(-5112);
			20056: out = 24'(14388);
			20057: out = 24'(10576);
			20058: out = 24'(-10584);
			20059: out = 24'(-21348);
			20060: out = 24'(-8920);
			20061: out = 24'(2592);
			20062: out = 24'(2676);
			20063: out = 24'(708);
			20064: out = 24'(16976);
			20065: out = 24'(33120);
			20066: out = 24'(34980);
			20067: out = 24'(23484);
			20068: out = 24'(5004);
			20069: out = 24'(-20596);
			20070: out = 24'(-34956);
			20071: out = 24'(-11872);
			20072: out = 24'(-15276);
			20073: out = 24'(-2096);
			20074: out = 24'(15260);
			20075: out = 24'(30156);
			20076: out = 24'(2132);
			20077: out = 24'(-2532);
			20078: out = 24'(-4108);
			20079: out = 24'(-11596);
			20080: out = 24'(-17108);
			20081: out = 24'(-7840);
			20082: out = 24'(9032);
			20083: out = 24'(15832);
			20084: out = 24'(-1164);
			20085: out = 24'(3716);
			20086: out = 24'(10980);
			20087: out = 24'(11756);
			20088: out = 24'(1264);
			20089: out = 24'(1756);
			20090: out = 24'(-4220);
			20091: out = 24'(-14776);
			20092: out = 24'(-21596);
			20093: out = 24'(-5144);
			20094: out = 24'(-32);
			20095: out = 24'(-568);
			20096: out = 24'(10660);
			20097: out = 24'(20768);
			20098: out = 24'(21224);
			20099: out = 24'(-2824);
			20100: out = 24'(-23524);
			20101: out = 24'(-24380);
			20102: out = 24'(10444);
			20103: out = 24'(17920);
			20104: out = 24'(1464);
			20105: out = 24'(-9432);
			20106: out = 24'(-2768);
			20107: out = 24'(-8568);
			20108: out = 24'(-21120);
			20109: out = 24'(-19960);
			20110: out = 24'(14800);
			20111: out = 24'(16968);
			20112: out = 24'(-480);
			20113: out = 24'(-7380);
			20114: out = 24'(11480);
			20115: out = 24'(10996);
			20116: out = 24'(5076);
			20117: out = 24'(7872);
			20118: out = 24'(12888);
			20119: out = 24'(-23768);
			20120: out = 24'(-64360);
			20121: out = 24'(-61884);
			20122: out = 24'(-2680);
			20123: out = 24'(20380);
			20124: out = 24'(20384);
			20125: out = 24'(13420);
			20126: out = 24'(8212);
			20127: out = 24'(13956);
			20128: out = 24'(8356);
			20129: out = 24'(-8096);
			20130: out = 24'(-19660);
			20131: out = 24'(-4184);
			20132: out = 24'(12348);
			20133: out = 24'(2792);
			20134: out = 24'(-27652);
			20135: out = 24'(-15316);
			20136: out = 24'(-1800);
			20137: out = 24'(23508);
			20138: out = 24'(34820);
			20139: out = 24'(14408);
			20140: out = 24'(-11064);
			20141: out = 24'(-34296);
			20142: out = 24'(-38500);
			20143: out = 24'(-10132);
			20144: out = 24'(3396);
			20145: out = 24'(21208);
			20146: out = 24'(28440);
			20147: out = 24'(23008);
			20148: out = 24'(-4108);
			20149: out = 24'(-10588);
			20150: out = 24'(-5264);
			20151: out = 24'(816);
			20152: out = 24'(-980);
			20153: out = 24'(5176);
			20154: out = 24'(8364);
			20155: out = 24'(4492);
			20156: out = 24'(-20148);
			20157: out = 24'(-9552);
			20158: out = 24'(4520);
			20159: out = 24'(20360);
			20160: out = 24'(27840);
			20161: out = 24'(21264);
			20162: out = 24'(-13388);
			20163: out = 24'(-31088);
			20164: out = 24'(-2260);
			20165: out = 24'(20584);
			20166: out = 24'(12012);
			20167: out = 24'(-6112);
			20168: out = 24'(-8464);
			20169: out = 24'(-5164);
			20170: out = 24'(-25292);
			20171: out = 24'(-38568);
			20172: out = 24'(-16368);
			20173: out = 24'(11588);
			20174: out = 24'(29432);
			20175: out = 24'(27640);
			20176: out = 24'(17504);
			20177: out = 24'(2756);
			20178: out = 24'(-12624);
			20179: out = 24'(-20368);
			20180: out = 24'(-18440);
			20181: out = 24'(-7164);
			20182: out = 24'(-5916);
			20183: out = 24'(3820);
			20184: out = 24'(8432);
			20185: out = 24'(7844);
			20186: out = 24'(-7660);
			20187: out = 24'(2140);
			20188: out = 24'(6864);
			20189: out = 24'(-3332);
			20190: out = 24'(-35472);
			20191: out = 24'(-16144);
			20192: out = 24'(4876);
			20193: out = 24'(7756);
			20194: out = 24'(212);
			20195: out = 24'(29268);
			20196: out = 24'(27712);
			20197: out = 24'(-5600);
			20198: out = 24'(-35640);
			20199: out = 24'(-19252);
			20200: out = 24'(-2540);
			20201: out = 24'(5132);
			20202: out = 24'(21480);
			20203: out = 24'(34208);
			20204: out = 24'(22496);
			20205: out = 24'(-8804);
			20206: out = 24'(-28464);
			20207: out = 24'(-23324);
			20208: out = 24'(3916);
			20209: out = 24'(20428);
			20210: out = 24'(19140);
			20211: out = 24'(8004);
			20212: out = 24'(11948);
			20213: out = 24'(9420);
			20214: out = 24'(-7152);
			20215: out = 24'(-19452);
			20216: out = 24'(-23916);
			20217: out = 24'(-8456);
			20218: out = 24'(268);
			20219: out = 24'(-5036);
			20220: out = 24'(-33852);
			20221: out = 24'(-8568);
			20222: out = 24'(39060);
			20223: out = 24'(54084);
			20224: out = 24'(34080);
			20225: out = 24'(7940);
			20226: out = 24'(-13084);
			20227: out = 24'(-36592);
			20228: out = 24'(-62044);
			20229: out = 24'(-42640);
			20230: out = 24'(8548);
			20231: out = 24'(40472);
			20232: out = 24'(36604);
			20233: out = 24'(18760);
			20234: out = 24'(6784);
			20235: out = 24'(-9988);
			20236: out = 24'(-29084);
			20237: out = 24'(-51308);
			20238: out = 24'(-22768);
			20239: out = 24'(16540);
			20240: out = 24'(24272);
			20241: out = 24'(26112);
			20242: out = 24'(18340);
			20243: out = 24'(8356);
			20244: out = 24'(-2208);
			20245: out = 24'(-12716);
			20246: out = 24'(-9564);
			20247: out = 24'(-13588);
			20248: out = 24'(-24048);
			20249: out = 24'(-41988);
			20250: out = 24'(-8724);
			20251: out = 24'(4720);
			20252: out = 24'(808);
			20253: out = 24'(3112);
			20254: out = 24'(37756);
			20255: out = 24'(24560);
			20256: out = 24'(-20636);
			20257: out = 24'(-53268);
			20258: out = 24'(-6860);
			20259: out = 24'(5452);
			20260: out = 24'(-1644);
			20261: out = 24'(3764);
			20262: out = 24'(7468);
			20263: out = 24'(5400);
			20264: out = 24'(-1668);
			20265: out = 24'(3856);
			20266: out = 24'(6984);
			20267: out = 24'(6272);
			20268: out = 24'(-13852);
			20269: out = 24'(-24512);
			20270: out = 24'(2752);
			20271: out = 24'(18240);
			20272: out = 24'(28064);
			20273: out = 24'(27240);
			20274: out = 24'(22640);
			20275: out = 24'(-25364);
			20276: out = 24'(-30508);
			20277: out = 24'(-5844);
			20278: out = 24'(16660);
			20279: out = 24'(19032);
			20280: out = 24'(6780);
			20281: out = 24'(-1736);
			20282: out = 24'(1912);
			20283: out = 24'(10248);
			20284: out = 24'(4768);
			20285: out = 24'(-8752);
			20286: out = 24'(-15916);
			20287: out = 24'(-7636);
			20288: out = 24'(10388);
			20289: out = 24'(11788);
			20290: out = 24'(-3504);
			20291: out = 24'(-9116);
			20292: out = 24'(14152);
			20293: out = 24'(36752);
			20294: out = 24'(29520);
			20295: out = 24'(3272);
			20296: out = 24'(-19496);
			20297: out = 24'(-14656);
			20298: out = 24'(-7488);
			20299: out = 24'(-9244);
			20300: out = 24'(-12180);
			20301: out = 24'(13376);
			20302: out = 24'(33220);
			20303: out = 24'(33156);
			20304: out = 24'(19236);
			20305: out = 24'(-1292);
			20306: out = 24'(-29416);
			20307: out = 24'(-39932);
			20308: out = 24'(-10972);
			20309: out = 24'(3868);
			20310: out = 24'(5220);
			20311: out = 24'(-3880);
			20312: out = 24'(-7980);
			20313: out = 24'(-5392);
			20314: out = 24'(-2000);
			20315: out = 24'(108);
			20316: out = 24'(1084);
			20317: out = 24'(14404);
			20318: out = 24'(6272);
			20319: out = 24'(1216);
			20320: out = 24'(-1136);
			20321: out = 24'(924);
			20322: out = 24'(-14196);
			20323: out = 24'(-6688);
			20324: out = 24'(11944);
			20325: out = 24'(16700);
			20326: out = 24'(2744);
			20327: out = 24'(-6328);
			20328: out = 24'(-8488);
			20329: out = 24'(996);
			20330: out = 24'(-2904);
			20331: out = 24'(9340);
			20332: out = 24'(2468);
			20333: out = 24'(-15184);
			20334: out = 24'(-63512);
			20335: out = 24'(-13804);
			20336: out = 24'(23772);
			20337: out = 24'(8112);
			20338: out = 24'(-21284);
			20339: out = 24'(10320);
			20340: out = 24'(27076);
			20341: out = 24'(5248);
			20342: out = 24'(-22608);
			20343: out = 24'(-9432);
			20344: out = 24'(-3808);
			20345: out = 24'(-6828);
			20346: out = 24'(80);
			20347: out = 24'(2348);
			20348: out = 24'(-21276);
			20349: out = 24'(-30584);
			20350: out = 24'(8080);
			20351: out = 24'(38292);
			20352: out = 24'(39412);
			20353: out = 24'(18540);
			20354: out = 24'(-2364);
			20355: out = 24'(1544);
			20356: out = 24'(-36916);
			20357: out = 24'(-45088);
			20358: out = 24'(-5712);
			20359: out = 24'(35076);
			20360: out = 24'(17876);
			20361: out = 24'(1072);
			20362: out = 24'(1064);
			20363: out = 24'(500);
			20364: out = 24'(-640);
			20365: out = 24'(16180);
			20366: out = 24'(33528);
			20367: out = 24'(19368);
			20368: out = 24'(-5724);
			20369: out = 24'(-22392);
			20370: out = 24'(-13008);
			20371: out = 24'(48);
			20372: out = 24'(-3388);
			20373: out = 24'(-2240);
			20374: out = 24'(4488);
			20375: out = 24'(6360);
			20376: out = 24'(308);
			20377: out = 24'(-1056);
			20378: out = 24'(3956);
			20379: out = 24'(9120);
			20380: out = 24'(18036);
			20381: out = 24'(2632);
			20382: out = 24'(-5032);
			20383: out = 24'(-13544);
			20384: out = 24'(-20164);
			20385: out = 24'(-12632);
			20386: out = 24'(8304);
			20387: out = 24'(21048);
			20388: out = 24'(23144);
			20389: out = 24'(-236);
			20390: out = 24'(13492);
			20391: out = 24'(14552);
			20392: out = 24'(-5620);
			20393: out = 24'(-16864);
			20394: out = 24'(-14992);
			20395: out = 24'(-20132);
			20396: out = 24'(-28480);
			20397: out = 24'(-7784);
			20398: out = 24'(12124);
			20399: out = 24'(19784);
			20400: out = 24'(19368);
			20401: out = 24'(30804);
			20402: out = 24'(29660);
			20403: out = 24'(3048);
			20404: out = 24'(-40788);
			20405: out = 24'(-59820);
			20406: out = 24'(-36804);
			20407: out = 24'(-2324);
			20408: out = 24'(12672);
			20409: out = 24'(21648);
			20410: out = 24'(28016);
			20411: out = 24'(23456);
			20412: out = 24'(-12316);
			20413: out = 24'(-42400);
			20414: out = 24'(-12164);
			20415: out = 24'(14540);
			20416: out = 24'(18028);
			20417: out = 24'(2788);
			20418: out = 24'(616);
			20419: out = 24'(-24900);
			20420: out = 24'(-21492);
			20421: out = 24'(6224);
			20422: out = 24'(29228);
			20423: out = 24'(5316);
			20424: out = 24'(-13796);
			20425: out = 24'(-8336);
			20426: out = 24'(4652);
			20427: out = 24'(-33728);
			20428: out = 24'(-31368);
			20429: out = 24'(9420);
			20430: out = 24'(44712);
			20431: out = 24'(24132);
			20432: out = 24'(-14664);
			20433: out = 24'(-34224);
			20434: out = 24'(-26760);
			20435: out = 24'(-33876);
			20436: out = 24'(-21600);
			20437: out = 24'(6736);
			20438: out = 24'(47104);
			20439: out = 24'(49664);
			20440: out = 24'(25596);
			20441: out = 24'(-29928);
			20442: out = 24'(-47488);
			20443: out = 24'(-13992);
			20444: out = 24'(5920);
			20445: out = 24'(-2304);
			20446: out = 24'(-10952);
			20447: out = 24'(8048);
			20448: out = 24'(22632);
			20449: out = 24'(26960);
			20450: out = 24'(9796);
			20451: out = 24'(3096);
			20452: out = 24'(13584);
			20453: out = 24'(11340);
			20454: out = 24'(-10188);
			20455: out = 24'(-30380);
			20456: out = 24'(-36744);
			20457: out = 24'(-11532);
			20458: out = 24'(2016);
			20459: out = 24'(20076);
			20460: out = 24'(37944);
			20461: out = 24'(38980);
			20462: out = 24'(-992);
			20463: out = 24'(-25832);
			20464: out = 24'(-9120);
			20465: out = 24'(15200);
			20466: out = 24'(10068);
			20467: out = 24'(-6260);
			20468: out = 24'(-11976);
			20469: out = 24'(-8364);
			20470: out = 24'(-5544);
			20471: out = 24'(3716);
			20472: out = 24'(16248);
			20473: out = 24'(24616);
			20474: out = 24'(21704);
			20475: out = 24'(9944);
			20476: out = 24'(-9928);
			20477: out = 24'(-20388);
			20478: out = 24'(-28140);
			20479: out = 24'(2168);
			20480: out = 24'(12496);
			20481: out = 24'(-2140);
			20482: out = 24'(-4208);
			20483: out = 24'(292);
			20484: out = 24'(-10060);
			20485: out = 24'(-24460);
			20486: out = 24'(-11092);
			20487: out = 24'(29776);
			20488: out = 24'(29768);
			20489: out = 24'(-4240);
			20490: out = 24'(-17040);
			20491: out = 24'(-6088);
			20492: out = 24'(8296);
			20493: out = 24'(4040);
			20494: out = 24'(1788);
			20495: out = 24'(-1684);
			20496: out = 24'(11076);
			20497: out = 24'(9152);
			20498: out = 24'(-8544);
			20499: out = 24'(-26812);
			20500: out = 24'(-6408);
			20501: out = 24'(21444);
			20502: out = 24'(22512);
			20503: out = 24'(1896);
			20504: out = 24'(-17344);
			20505: out = 24'(-17572);
			20506: out = 24'(-10368);
			20507: out = 24'(-2972);
			20508: out = 24'(-2060);
			20509: out = 24'(21520);
			20510: out = 24'(36752);
			20511: out = 24'(16756);
			20512: out = 24'(-6836);
			20513: out = 24'(-10088);
			20514: out = 24'(5756);
			20515: out = 24'(1996);
			20516: out = 24'(-15672);
			20517: out = 24'(-36972);
			20518: out = 24'(-23420);
			20519: out = 24'(4920);
			20520: out = 24'(14680);
			20521: out = 24'(3860);
			20522: out = 24'(-904);
			20523: out = 24'(1604);
			20524: out = 24'(8116);
			20525: out = 24'(-15608);
			20526: out = 24'(-12256);
			20527: out = 24'(3028);
			20528: out = 24'(-556);
			20529: out = 24'(-6084);
			20530: out = 24'(1624);
			20531: out = 24'(20408);
			20532: out = 24'(28972);
			20533: out = 24'(9740);
			20534: out = 24'(1284);
			20535: out = 24'(-4656);
			20536: out = 24'(-7844);
			20537: out = 24'(1724);
			20538: out = 24'(23016);
			20539: out = 24'(26408);
			20540: out = 24'(4828);
			20541: out = 24'(-19720);
			20542: out = 24'(-17856);
			20543: out = 24'(-5156);
			20544: out = 24'(-476);
			20545: out = 24'(152);
			20546: out = 24'(19060);
			20547: out = 24'(22076);
			20548: out = 24'(-788);
			20549: out = 24'(-29352);
			20550: out = 24'(-13128);
			20551: out = 24'(3156);
			20552: out = 24'(4696);
			20553: out = 24'(-2688);
			20554: out = 24'(-12816);
			20555: out = 24'(-4616);
			20556: out = 24'(-376);
			20557: out = 24'(4396);
			20558: out = 24'(29144);
			20559: out = 24'(26852);
			20560: out = 24'(10728);
			20561: out = 24'(-5092);
			20562: out = 24'(-6248);
			20563: out = 24'(-14988);
			20564: out = 24'(-22652);
			20565: out = 24'(-9864);
			20566: out = 24'(25900);
			20567: out = 24'(23368);
			20568: out = 24'(9084);
			20569: out = 24'(-9364);
			20570: out = 24'(-14356);
			20571: out = 24'(-30192);
			20572: out = 24'(-11856);
			20573: out = 24'(10828);
			20574: out = 24'(18404);
			20575: out = 24'(56);
			20576: out = 24'(-1760);
			20577: out = 24'(84);
			20578: out = 24'(-3252);
			20579: out = 24'(-8720);
			20580: out = 24'(-30236);
			20581: out = 24'(-22096);
			20582: out = 24'(6696);
			20583: out = 24'(22876);
			20584: out = 24'(4200);
			20585: out = 24'(-6604);
			20586: out = 24'(2800);
			20587: out = 24'(18112);
			20588: out = 24'(14136);
			20589: out = 24'(9152);
			20590: out = 24'(3224);
			20591: out = 24'(-5844);
			20592: out = 24'(-32672);
			20593: out = 24'(-12904);
			20594: out = 24'(14500);
			20595: out = 24'(21468);
			20596: out = 24'(7032);
			20597: out = 24'(-208);
			20598: out = 24'(2704);
			20599: out = 24'(4948);
			20600: out = 24'(-7116);
			20601: out = 24'(-8204);
			20602: out = 24'(-13048);
			20603: out = 24'(-8004);
			20604: out = 24'(8820);
			20605: out = 24'(12228);
			20606: out = 24'(16808);
			20607: out = 24'(13144);
			20608: out = 24'(4520);
			20609: out = 24'(-1700);
			20610: out = 24'(-2516);
			20611: out = 24'(-6236);
			20612: out = 24'(-16704);
			20613: out = 24'(-20424);
			20614: out = 24'(-5604);
			20615: out = 24'(11716);
			20616: out = 24'(9688);
			20617: out = 24'(784);
			20618: out = 24'(-3536);
			20619: out = 24'(14520);
			20620: out = 24'(18508);
			20621: out = 24'(-3108);
			20622: out = 24'(-9276);
			20623: out = 24'(1672);
			20624: out = 24'(9492);
			20625: out = 24'(-752);
			20626: out = 24'(-1288);
			20627: out = 24'(10744);
			20628: out = 24'(28804);
			20629: out = 24'(30180);
			20630: out = 24'(5356);
			20631: out = 24'(-4348);
			20632: out = 24'(-13952);
			20633: out = 24'(-19540);
			20634: out = 24'(-14064);
			20635: out = 24'(6852);
			20636: out = 24'(14660);
			20637: out = 24'(9160);
			20638: out = 24'(4696);
			20639: out = 24'(-5828);
			20640: out = 24'(-10108);
			20641: out = 24'(-10188);
			20642: out = 24'(-6560);
			20643: out = 24'(-7052);
			20644: out = 24'(-6888);
			20645: out = 24'(-2444);
			20646: out = 24'(7156);
			20647: out = 24'(4452);
			20648: out = 24'(-4564);
			20649: out = 24'(-14148);
			20650: out = 24'(-3504);
			20651: out = 24'(13580);
			20652: out = 24'(5560);
			20653: out = 24'(-20088);
			20654: out = 24'(-27684);
			20655: out = 24'(-13404);
			20656: out = 24'(20416);
			20657: out = 24'(9836);
			20658: out = 24'(-1268);
			20659: out = 24'(6256);
			20660: out = 24'(7504);
			20661: out = 24'(-23408);
			20662: out = 24'(-37288);
			20663: out = 24'(-11916);
			20664: out = 24'(-2768);
			20665: out = 24'(-7628);
			20666: out = 24'(-10476);
			20667: out = 24'(3212);
			20668: out = 24'(5960);
			20669: out = 24'(2484);
			20670: out = 24'(-4200);
			20671: out = 24'(-3692);
			20672: out = 24'(-164);
			20673: out = 24'(11552);
			20674: out = 24'(18216);
			20675: out = 24'(11980);
			20676: out = 24'(-1676);
			20677: out = 24'(-20144);
			20678: out = 24'(-712);
			20679: out = 24'(21932);
			20680: out = 24'(17924);
			20681: out = 24'(-25828);
			20682: out = 24'(-21400);
			20683: out = 24'(-5068);
			20684: out = 24'(-624);
			20685: out = 24'(-4216);
			20686: out = 24'(21336);
			20687: out = 24'(31584);
			20688: out = 24'(14476);
			20689: out = 24'(-8864);
			20690: out = 24'(-4148);
			20691: out = 24'(-3348);
			20692: out = 24'(-15872);
			20693: out = 24'(-16504);
			20694: out = 24'(31112);
			20695: out = 24'(50852);
			20696: out = 24'(13816);
			20697: out = 24'(-47692);
			20698: out = 24'(-24308);
			20699: out = 24'(1768);
			20700: out = 24'(14736);
			20701: out = 24'(2920);
			20702: out = 24'(8652);
			20703: out = 24'(28);
			20704: out = 24'(8360);
			20705: out = 24'(9776);
			20706: out = 24'(-908);
			20707: out = 24'(-16964);
			20708: out = 24'(-6232);
			20709: out = 24'(6948);
			20710: out = 24'(-3580);
			20711: out = 24'(-18764);
			20712: out = 24'(-8764);
			20713: out = 24'(18272);
			20714: out = 24'(25640);
			20715: out = 24'(2744);
			20716: out = 24'(-5268);
			20717: out = 24'(112);
			20718: out = 24'(-8536);
			20719: out = 24'(-30640);
			20720: out = 24'(-36908);
			20721: out = 24'(-3096);
			20722: out = 24'(33796);
			20723: out = 24'(42980);
			20724: out = 24'(2240);
			20725: out = 24'(-16708);
			20726: out = 24'(-9996);
			20727: out = 24'(-2716);
			20728: out = 24'(-32664);
			20729: out = 24'(-33468);
			20730: out = 24'(-9680);
			20731: out = 24'(6140);
			20732: out = 24'(-13504);
			20733: out = 24'(-8368);
			20734: out = 24'(9544);
			20735: out = 24'(16948);
			20736: out = 24'(8360);
			20737: out = 24'(1704);
			20738: out = 24'(-7584);
			20739: out = 24'(-18904);
			20740: out = 24'(-19564);
			20741: out = 24'(-21252);
			20742: out = 24'(-10780);
			20743: out = 24'(10040);
			20744: out = 24'(30416);
			20745: out = 24'(16672);
			20746: out = 24'(-4912);
			20747: out = 24'(-19456);
			20748: out = 24'(-20068);
			20749: out = 24'(-19928);
			20750: out = 24'(-13780);
			20751: out = 24'(5428);
			20752: out = 24'(28224);
			20753: out = 24'(31088);
			20754: out = 24'(3784);
			20755: out = 24'(-20928);
			20756: out = 24'(-13032);
			20757: out = 24'(8940);
			20758: out = 24'(22636);
			20759: out = 24'(11040);
			20760: out = 24'(-1372);
			20761: out = 24'(156);
			20762: out = 24'(1524);
			20763: out = 24'(-7000);
			20764: out = 24'(-6424);
			20765: out = 24'(16436);
			20766: out = 24'(11664);
			20767: out = 24'(-1176);
			20768: out = 24'(-20304);
			20769: out = 24'(-26388);
			20770: out = 24'(-14476);
			20771: out = 24'(11320);
			20772: out = 24'(30528);
			20773: out = 24'(35744);
			20774: out = 24'(24440);
			20775: out = 24'(19616);
			20776: out = 24'(3480);
			20777: out = 24'(-28732);
			20778: out = 24'(-58436);
			20779: out = 24'(-29692);
			20780: out = 24'(23016);
			20781: out = 24'(36684);
			20782: out = 24'(6900);
			20783: out = 24'(1860);
			20784: out = 24'(19144);
			20785: out = 24'(25964);
			20786: out = 24'(3048);
			20787: out = 24'(-3504);
			20788: out = 24'(-11128);
			20789: out = 24'(-16952);
			20790: out = 24'(-20404);
			20791: out = 24'(-14260);
			20792: out = 24'(13508);
			20793: out = 24'(28512);
			20794: out = 24'(22448);
			20795: out = 24'(1936);
			20796: out = 24'(728);
			20797: out = 24'(-11236);
			20798: out = 24'(-23064);
			20799: out = 24'(-20576);
			20800: out = 24'(7916);
			20801: out = 24'(18852);
			20802: out = 24'(20236);
			20803: out = 24'(12256);
			20804: out = 24'(-5424);
			20805: out = 24'(-41140);
			20806: out = 24'(-35076);
			20807: out = 24'(13052);
			20808: out = 24'(33548);
			20809: out = 24'(4180);
			20810: out = 24'(-16212);
			20811: out = 24'(-5940);
			20812: out = 24'(-1656);
			20813: out = 24'(-21196);
			20814: out = 24'(-18724);
			20815: out = 24'(5628);
			20816: out = 24'(5576);
			20817: out = 24'(-6968);
			20818: out = 24'(-7812);
			20819: out = 24'(4088);
			20820: out = 24'(6620);
			20821: out = 24'(-9476);
			20822: out = 24'(7296);
			20823: out = 24'(26280);
			20824: out = 24'(8064);
			20825: out = 24'(-10504);
			20826: out = 24'(-22640);
			20827: out = 24'(-11940);
			20828: out = 24'(492);
			20829: out = 24'(588);
			20830: out = 24'(12088);
			20831: out = 24'(18732);
			20832: out = 24'(7228);
			20833: out = 24'(-18596);
			20834: out = 24'(-21908);
			20835: out = 24'(-9152);
			20836: out = 24'(9048);
			20837: out = 24'(16752);
			20838: out = 24'(24520);
			20839: out = 24'(4728);
			20840: out = 24'(-20908);
			20841: out = 24'(-25268);
			20842: out = 24'(4980);
			20843: out = 24'(7672);
			20844: out = 24'(-8776);
			20845: out = 24'(-5764);
			20846: out = 24'(27184);
			20847: out = 24'(31704);
			20848: out = 24'(644);
			20849: out = 24'(-22728);
			20850: out = 24'(5028);
			20851: out = 24'(16636);
			20852: out = 24'(2788);
			20853: out = 24'(-14232);
			20854: out = 24'(-3928);
			20855: out = 24'(15380);
			20856: out = 24'(16264);
			20857: out = 24'(6888);
			20858: out = 24'(6964);
			20859: out = 24'(17540);
			20860: out = 24'(1920);
			20861: out = 24'(-27028);
			20862: out = 24'(-39456);
			20863: out = 24'(-4932);
			20864: out = 24'(6268);
			20865: out = 24'(6116);
			20866: out = 24'(8444);
			20867: out = 24'(19264);
			20868: out = 24'(14944);
			20869: out = 24'(6508);
			20870: out = 24'(-3936);
			20871: out = 24'(-284);
			20872: out = 24'(-14228);
			20873: out = 24'(-2008);
			20874: out = 24'(684);
			20875: out = 24'(-22416);
			20876: out = 24'(-41048);
			20877: out = 24'(-11844);
			20878: out = 24'(23108);
			20879: out = 24'(15408);
			20880: out = 24'(2908);
			20881: out = 24'(-4004);
			20882: out = 24'(1672);
			20883: out = 24'(-4064);
			20884: out = 24'(-10324);
			20885: out = 24'(-6900);
			20886: out = 24'(9140);
			20887: out = 24'(8892);
			20888: out = 24'(-7216);
			20889: out = 24'(-17432);
			20890: out = 24'(-7052);
			20891: out = 24'(-612);
			20892: out = 24'(-3128);
			20893: out = 24'(-2600);
			20894: out = 24'(16124);
			20895: out = 24'(17104);
			20896: out = 24'(-7616);
			20897: out = 24'(-22976);
			20898: out = 24'(-10424);
			20899: out = 24'(2304);
			20900: out = 24'(444);
			20901: out = 24'(6676);
			20902: out = 24'(13796);
			20903: out = 24'(836);
			20904: out = 24'(-24400);
			20905: out = 24'(-22924);
			20906: out = 24'(-12332);
			20907: out = 24'(-6248);
			20908: out = 24'(-3564);
			20909: out = 24'(15832);
			20910: out = 24'(-280);
			20911: out = 24'(-4252);
			20912: out = 24'(11392);
			20913: out = 24'(35700);
			20914: out = 24'(17392);
			20915: out = 24'(-8096);
			20916: out = 24'(-22524);
			20917: out = 24'(-14128);
			20918: out = 24'(-12804);
			20919: out = 24'(-11656);
			20920: out = 24'(-3260);
			20921: out = 24'(16652);
			20922: out = 24'(22452);
			20923: out = 24'(13780);
			20924: out = 24'(-708);
			20925: out = 24'(-2800);
			20926: out = 24'(-1188);
			20927: out = 24'(-11088);
			20928: out = 24'(-18128);
			20929: out = 24'(3776);
			20930: out = 24'(39624);
			20931: out = 24'(41752);
			20932: out = 24'(15620);
			20933: out = 24'(-12472);
			20934: out = 24'(-19028);
			20935: out = 24'(-420);
			20936: out = 24'(1912);
			20937: out = 24'(-3336);
			20938: out = 24'(-4624);
			20939: out = 24'(-1336);
			20940: out = 24'(-796);
			20941: out = 24'(5608);
			20942: out = 24'(14980);
			20943: out = 24'(11800);
			20944: out = 24'(-628);
			20945: out = 24'(-11516);
			20946: out = 24'(-12700);
			20947: out = 24'(-12220);
			20948: out = 24'(10132);
			20949: out = 24'(16548);
			20950: out = 24'(12536);
			20951: out = 24'(388);
			20952: out = 24'(6840);
			20953: out = 24'(180);
			20954: out = 24'(-1072);
			20955: out = 24'(-4572);
			20956: out = 24'(-11368);
			20957: out = 24'(-24548);
			20958: out = 24'(-9676);
			20959: out = 24'(19880);
			20960: out = 24'(26752);
			20961: out = 24'(6232);
			20962: out = 24'(-6084);
			20963: out = 24'(3860);
			20964: out = 24'(13548);
			20965: out = 24'(-13220);
			20966: out = 24'(-34396);
			20967: out = 24'(-33272);
			20968: out = 24'(-17876);
			20969: out = 24'(10920);
			20970: out = 24'(11688);
			20971: out = 24'(2080);
			20972: out = 24'(-4408);
			20973: out = 24'(-164);
			20974: out = 24'(16);
			20975: out = 24'(104);
			20976: out = 24'(-2144);
			20977: out = 24'(-15792);
			20978: out = 24'(1068);
			20979: out = 24'(7360);
			20980: out = 24'(-7928);
			20981: out = 24'(-25248);
			20982: out = 24'(-8184);
			20983: out = 24'(21080);
			20984: out = 24'(23060);
			20985: out = 24'(-3088);
			20986: out = 24'(-25304);
			20987: out = 24'(-13408);
			20988: out = 24'(5916);
			20989: out = 24'(5920);
			20990: out = 24'(-2476);
			20991: out = 24'(8916);
			20992: out = 24'(23600);
			20993: out = 24'(17668);
			20994: out = 24'(-10388);
			20995: out = 24'(-22884);
			20996: out = 24'(-20176);
			20997: out = 24'(-6740);
			20998: out = 24'(7352);
			20999: out = 24'(13908);
			21000: out = 24'(10816);
			21001: out = 24'(5180);
			21002: out = 24'(-2480);
			21003: out = 24'(-15888);
			21004: out = 24'(-27528);
			21005: out = 24'(-17016);
			21006: out = 24'(11328);
			21007: out = 24'(22920);
			21008: out = 24'(16800);
			21009: out = 24'(5780);
			21010: out = 24'(-732);
			21011: out = 24'(812);
			21012: out = 24'(-15008);
			21013: out = 24'(-13600);
			21014: out = 24'(5748);
			21015: out = 24'(12044);
			21016: out = 24'(-18500);
			21017: out = 24'(-42568);
			21018: out = 24'(-28892);
			21019: out = 24'(4812);
			21020: out = 24'(23036);
			21021: out = 24'(34296);
			21022: out = 24'(44288);
			21023: out = 24'(32064);
			21024: out = 24'(7532);
			21025: out = 24'(-28768);
			21026: out = 24'(-27232);
			21027: out = 24'(2536);
			21028: out = 24'(13472);
			21029: out = 24'(7688);
			21030: out = 24'(14216);
			21031: out = 24'(19732);
			21032: out = 24'(-516);
			21033: out = 24'(-31392);
			21034: out = 24'(-20348);
			21035: out = 24'(15396);
			21036: out = 24'(17188);
			21037: out = 24'(4492);
			21038: out = 24'(244);
			21039: out = 24'(10336);
			21040: out = 24'(11720);
			21041: out = 24'(10576);
			21042: out = 24'(2976);
			21043: out = 24'(-9880);
			21044: out = 24'(-17980);
			21045: out = 24'(18720);
			21046: out = 24'(26288);
			21047: out = 24'(4176);
			21048: out = 24'(-21260);
			21049: out = 24'(5320);
			21050: out = 24'(2108);
			21051: out = 24'(-16628);
			21052: out = 24'(-33348);
			21053: out = 24'(-11456);
			21054: out = 24'(-3312);
			21055: out = 24'(-1100);
			21056: out = 24'(-7280);
			21057: out = 24'(-6808);
			21058: out = 24'(9824);
			21059: out = 24'(16360);
			21060: out = 24'(4148);
			21061: out = 24'(-18688);
			21062: out = 24'(-11892);
			21063: out = 24'(-22992);
			21064: out = 24'(-29564);
			21065: out = 24'(-24448);
			21066: out = 24'(-504);
			21067: out = 24'(0);
			21068: out = 24'(7004);
			21069: out = 24'(16184);
			21070: out = 24'(14588);
			21071: out = 24'(11520);
			21072: out = 24'(7240);
			21073: out = 24'(-13148);
			21074: out = 24'(-49200);
			21075: out = 24'(-45472);
			21076: out = 24'(1104);
			21077: out = 24'(41080);
			21078: out = 24'(30032);
			21079: out = 24'(-10476);
			21080: out = 24'(-17688);
			21081: out = 24'(5696);
			21082: out = 24'(10904);
			21083: out = 24'(-6612);
			21084: out = 24'(-15808);
			21085: out = 24'(8984);
			21086: out = 24'(31420);
			21087: out = 24'(21488);
			21088: out = 24'(-1896);
			21089: out = 24'(-2636);
			21090: out = 24'(9384);
			21091: out = 24'(1256);
			21092: out = 24'(-8496);
			21093: out = 24'(-7792);
			21094: out = 24'(7900);
			21095: out = 24'(14908);
			21096: out = 24'(-14136);
			21097: out = 24'(-13212);
			21098: out = 24'(16536);
			21099: out = 24'(33656);
			21100: out = 24'(23352);
			21101: out = 24'(-9176);
			21102: out = 24'(-20920);
			21103: out = 24'(-9248);
			21104: out = 24'(-1676);
			21105: out = 24'(-9156);
			21106: out = 24'(-1324);
			21107: out = 24'(29408);
			21108: out = 24'(49416);
			21109: out = 24'(31500);
			21110: out = 24'(-7432);
			21111: out = 24'(-34984);
			21112: out = 24'(-33192);
			21113: out = 24'(-49840);
			21114: out = 24'(-29260);
			21115: out = 24'(14620);
			21116: out = 24'(43484);
			21117: out = 24'(26272);
			21118: out = 24'(6060);
			21119: out = 24'(2596);
			21120: out = 24'(15864);
			21121: out = 24'(14420);
			21122: out = 24'(-2484);
			21123: out = 24'(-30312);
			21124: out = 24'(-38244);
			21125: out = 24'(-12536);
			21126: out = 24'(3896);
			21127: out = 24'(4832);
			21128: out = 24'(-1508);
			21129: out = 24'(-136);
			21130: out = 24'(-552);
			21131: out = 24'(16);
			21132: out = 24'(-604);
			21133: out = 24'(3932);
			21134: out = 24'(6112);
			21135: out = 24'(3484);
			21136: out = 24'(-1364);
			21137: out = 24'(5964);
			21138: out = 24'(10932);
			21139: out = 24'(12532);
			21140: out = 24'(-12028);
			21141: out = 24'(-35564);
			21142: out = 24'(-36992);
			21143: out = 24'(-1332);
			21144: out = 24'(7636);
			21145: out = 24'(-2388);
			21146: out = 24'(-5916);
			21147: out = 24'(24908);
			21148: out = 24'(20704);
			21149: out = 24'(-2200);
			21150: out = 24'(-15068);
			21151: out = 24'(-1884);
			21152: out = 24'(-11184);
			21153: out = 24'(-22624);
			21154: out = 24'(-14516);
			21155: out = 24'(13048);
			21156: out = 24'(11528);
			21157: out = 24'(7184);
			21158: out = 24'(8056);
			21159: out = 24'(7676);
			21160: out = 24'(-28044);
			21161: out = 24'(-41960);
			21162: out = 24'(-21368);
			21163: out = 24'(-40);
			21164: out = 24'(3496);
			21165: out = 24'(4776);
			21166: out = 24'(11404);
			21167: out = 24'(7452);
			21168: out = 24'(10464);
			21169: out = 24'(3136);
			21170: out = 24'(1684);
			21171: out = 24'(-648);
			21172: out = 24'(1716);
			21173: out = 24'(-6228);
			21174: out = 24'(-2436);
			21175: out = 24'(3908);
			21176: out = 24'(1424);
			21177: out = 24'(4756);
			21178: out = 24'(18576);
			21179: out = 24'(18396);
			21180: out = 24'(-11072);
			21181: out = 24'(-20132);
			21182: out = 24'(3468);
			21183: out = 24'(28560);
			21184: out = 24'(14864);
			21185: out = 24'(22768);
			21186: out = 24'(6228);
			21187: out = 24'(-17200);
			21188: out = 24'(-40444);
			21189: out = 24'(-6440);
			21190: out = 24'(11016);
			21191: out = 24'(23036);
			21192: out = 24'(22764);
			21193: out = 24'(24996);
			21194: out = 24'(-3364);
			21195: out = 24'(-12948);
			21196: out = 24'(4044);
			21197: out = 24'(33780);
			21198: out = 24'(4352);
			21199: out = 24'(-15564);
			21200: out = 24'(-12536);
			21201: out = 24'(-1072);
			21202: out = 24'(-3292);
			21203: out = 24'(-14180);
			21204: out = 24'(-19908);
			21205: out = 24'(-7496);
			21206: out = 24'(16444);
			21207: out = 24'(26288);
			21208: out = 24'(11196);
			21209: out = 24'(-9992);
			21210: out = 24'(-4992);
			21211: out = 24'(-14104);
			21212: out = 24'(-28020);
			21213: out = 24'(-24420);
			21214: out = 24'(10248);
			21215: out = 24'(28448);
			21216: out = 24'(16328);
			21217: out = 24'(-5644);
			21218: out = 24'(-6756);
			21219: out = 24'(-5656);
			21220: out = 24'(-1384);
			21221: out = 24'(4640);
			21222: out = 24'(13504);
			21223: out = 24'(2372);
			21224: out = 24'(-25392);
			21225: out = 24'(-40772);
			21226: out = 24'(-14972);
			21227: out = 24'(9592);
			21228: out = 24'(26576);
			21229: out = 24'(13336);
			21230: out = 24'(764);
			21231: out = 24'(6640);
			21232: out = 24'(15172);
			21233: out = 24'(520);
			21234: out = 24'(-16368);
			21235: out = 24'(-2524);
			21236: out = 24'(7952);
			21237: out = 24'(10908);
			21238: out = 24'(4788);
			21239: out = 24'(-264);
			21240: out = 24'(-13308);
			21241: out = 24'(-13236);
			21242: out = 24'(864);
			21243: out = 24'(15332);
			21244: out = 24'(21064);
			21245: out = 24'(11400);
			21246: out = 24'(6040);
			21247: out = 24'(8212);
			21248: out = 24'(23092);
			21249: out = 24'(-5132);
			21250: out = 24'(-25532);
			21251: out = 24'(-24936);
			21252: out = 24'(-276);
			21253: out = 24'(-11568);
			21254: out = 24'(5192);
			21255: out = 24'(27308);
			21256: out = 24'(20796);
			21257: out = 24'(2876);
			21258: out = 24'(832);
			21259: out = 24'(6292);
			21260: out = 24'(-5536);
			21261: out = 24'(-32648);
			21262: out = 24'(-19352);
			21263: out = 24'(12932);
			21264: out = 24'(16056);
			21265: out = 24'(6560);
			21266: out = 24'(-11792);
			21267: out = 24'(-1308);
			21268: out = 24'(13900);
			21269: out = 24'(6700);
			21270: out = 24'(-5724);
			21271: out = 24'(-5844);
			21272: out = 24'(-860);
			21273: out = 24'(-9480);
			21274: out = 24'(-11872);
			21275: out = 24'(-340);
			21276: out = 24'(25084);
			21277: out = 24'(40860);
			21278: out = 24'(23224);
			21279: out = 24'(-1044);
			21280: out = 24'(-25140);
			21281: out = 24'(-43152);
			21282: out = 24'(-33760);
			21283: out = 24'(-8260);
			21284: out = 24'(23104);
			21285: out = 24'(30908);
			21286: out = 24'(8708);
			21287: out = 24'(-13008);
			21288: out = 24'(-11244);
			21289: out = 24'(-3680);
			21290: out = 24'(-25448);
			21291: out = 24'(-12956);
			21292: out = 24'(5540);
			21293: out = 24'(19808);
			21294: out = 24'(15096);
			21295: out = 24'(9012);
			21296: out = 24'(808);
			21297: out = 24'(-4792);
			21298: out = 24'(-15100);
			21299: out = 24'(-18912);
			21300: out = 24'(-18060);
			21301: out = 24'(-876);
			21302: out = 24'(14652);
			21303: out = 24'(14332);
			21304: out = 24'(-5636);
			21305: out = 24'(-7800);
			21306: out = 24'(15468);
			21307: out = 24'(35020);
			21308: out = 24'(21056);
			21309: out = 24'(-4964);
			21310: out = 24'(-19920);
			21311: out = 24'(-22276);
			21312: out = 24'(-26812);
			21313: out = 24'(-31372);
			21314: out = 24'(-15004);
			21315: out = 24'(21816);
			21316: out = 24'(35824);
			21317: out = 24'(21276);
			21318: out = 24'(-4996);
			21319: out = 24'(-9740);
			21320: out = 24'(-3812);
			21321: out = 24'(3372);
			21322: out = 24'(-14520);
			21323: out = 24'(-23228);
			21324: out = 24'(9012);
			21325: out = 24'(28240);
			21326: out = 24'(10108);
			21327: out = 24'(-17432);
			21328: out = 24'(-9960);
			21329: out = 24'(16344);
			21330: out = 24'(15144);
			21331: out = 24'(-14172);
			21332: out = 24'(-29012);
			21333: out = 24'(-864);
			21334: out = 24'(28956);
			21335: out = 24'(26648);
			21336: out = 24'(2884);
			21337: out = 24'(-308);
			21338: out = 24'(-2440);
			21339: out = 24'(784);
			21340: out = 24'(2616);
			21341: out = 24'(13580);
			21342: out = 24'(3648);
			21343: out = 24'(-132);
			21344: out = 24'(-5568);
			21345: out = 24'(-12780);
			21346: out = 24'(-21772);
			21347: out = 24'(-9868);
			21348: out = 24'(0);
			21349: out = 24'(-6008);
			21350: out = 24'(-23304);
			21351: out = 24'(-4508);
			21352: out = 24'(12240);
			21353: out = 24'(-4440);
			21354: out = 24'(-8972);
			21355: out = 24'(1544);
			21356: out = 24'(25484);
			21357: out = 24'(23580);
			21358: out = 24'(9736);
			21359: out = 24'(-17040);
			21360: out = 24'(-17592);
			21361: out = 24'(-14360);
			21362: out = 24'(-14308);
			21363: out = 24'(-23420);
			21364: out = 24'(9332);
			21365: out = 24'(31768);
			21366: out = 24'(3284);
			21367: out = 24'(-15472);
			21368: out = 24'(-9768);
			21369: out = 24'(6756);
			21370: out = 24'(-2204);
			21371: out = 24'(9008);
			21372: out = 24'(1196);
			21373: out = 24'(-3336);
			21374: out = 24'(-8004);
			21375: out = 24'(7956);
			21376: out = 24'(1484);
			21377: out = 24'(-1596);
			21378: out = 24'(-5956);
			21379: out = 24'(-3448);
			21380: out = 24'(-18100);
			21381: out = 24'(-10824);
			21382: out = 24'(5480);
			21383: out = 24'(10508);
			21384: out = 24'(8652);
			21385: out = 24'(10656);
			21386: out = 24'(15556);
			21387: out = 24'(11508);
			21388: out = 24'(2480);
			21389: out = 24'(-16420);
			21390: out = 24'(-25596);
			21391: out = 24'(-16176);
			21392: out = 24'(-1524);
			21393: out = 24'(2120);
			21394: out = 24'(-3612);
			21395: out = 24'(2376);
			21396: out = 24'(28344);
			21397: out = 24'(18008);
			21398: out = 24'(-7016);
			21399: out = 24'(-16320);
			21400: out = 24'(8204);
			21401: out = 24'(13372);
			21402: out = 24'(6420);
			21403: out = 24'(-192);
			21404: out = 24'(9332);
			21405: out = 24'(25900);
			21406: out = 24'(15624);
			21407: out = 24'(-13320);
			21408: out = 24'(-32640);
			21409: out = 24'(-22452);
			21410: out = 24'(-18780);
			21411: out = 24'(-21620);
			21412: out = 24'(-12340);
			21413: out = 24'(22592);
			21414: out = 24'(30824);
			21415: out = 24'(16440);
			21416: out = 24'(-3648);
			21417: out = 24'(1708);
			21418: out = 24'(236);
			21419: out = 24'(6500);
			21420: out = 24'(4592);
			21421: out = 24'(3364);
			21422: out = 24'(-6372);
			21423: out = 24'(10872);
			21424: out = 24'(17880);
			21425: out = 24'(1756);
			21426: out = 24'(-33412);
			21427: out = 24'(-15124);
			21428: out = 24'(13232);
			21429: out = 24'(5964);
			21430: out = 24'(-27828);
			21431: out = 24'(-17948);
			21432: out = 24'(18608);
			21433: out = 24'(32868);
			21434: out = 24'(17512);
			21435: out = 24'(1468);
			21436: out = 24'(-64);
			21437: out = 24'(-10796);
			21438: out = 24'(-42312);
			21439: out = 24'(-50500);
			21440: out = 24'(-29504);
			21441: out = 24'(-4004);
			21442: out = 24'(-3312);
			21443: out = 24'(15148);
			21444: out = 24'(21088);
			21445: out = 24'(24660);
			21446: out = 24'(14088);
			21447: out = 24'(10252);
			21448: out = 24'(-23772);
			21449: out = 24'(-40616);
			21450: out = 24'(-28052);
			21451: out = 24'(8000);
			21452: out = 24'(21768);
			21453: out = 24'(23920);
			21454: out = 24'(12172);
			21455: out = 24'(776);
			21456: out = 24'(-18420);
			21457: out = 24'(-8304);
			21458: out = 24'(-356);
			21459: out = 24'(-12256);
			21460: out = 24'(-18680);
			21461: out = 24'(6600);
			21462: out = 24'(35320);
			21463: out = 24'(33848);
			21464: out = 24'(4228);
			21465: out = 24'(-192);
			21466: out = 24'(3692);
			21467: out = 24'(-4216);
			21468: out = 24'(-9744);
			21469: out = 24'(-8984);
			21470: out = 24'(7944);
			21471: out = 24'(16576);
			21472: out = 24'(7132);
			21473: out = 24'(-8992);
			21474: out = 24'(-8628);
			21475: out = 24'(2032);
			21476: out = 24'(-2076);
			21477: out = 24'(-5296);
			21478: out = 24'(-18008);
			21479: out = 24'(-15164);
			21480: out = 24'(2796);
			21481: out = 24'(20372);
			21482: out = 24'(22200);
			21483: out = 24'(22488);
			21484: out = 24'(25128);
			21485: out = 24'(32688);
			21486: out = 24'(-13076);
			21487: out = 24'(-57632);
			21488: out = 24'(-64680);
			21489: out = 24'(-20620);
			21490: out = 24'(5128);
			21491: out = 24'(24348);
			21492: out = 24'(31232);
			21493: out = 24'(23744);
			21494: out = 24'(9972);
			21495: out = 24'(2472);
			21496: out = 24'(-6564);
			21497: out = 24'(-21316);
			21498: out = 24'(236);
			21499: out = 24'(1860);
			21500: out = 24'(-6448);
			21501: out = 24'(-8948);
			21502: out = 24'(22776);
			21503: out = 24'(9876);
			21504: out = 24'(-12816);
			21505: out = 24'(-14904);
			21506: out = 24'(16272);
			21507: out = 24'(12564);
			21508: out = 24'(-8412);
			21509: out = 24'(-19684);
			21510: out = 24'(-3236);
			21511: out = 24'(19896);
			21512: out = 24'(26524);
			21513: out = 24'(19340);
			21514: out = 24'(4316);
			21515: out = 24'(1652);
			21516: out = 24'(-15940);
			21517: out = 24'(-16464);
			21518: out = 24'(2120);
			21519: out = 24'(13028);
			21520: out = 24'(832);
			21521: out = 24'(-5736);
			21522: out = 24'(-3588);
			21523: out = 24'(-21256);
			21524: out = 24'(-23152);
			21525: out = 24'(-8052);
			21526: out = 24'(12300);
			21527: out = 24'(17172);
			21528: out = 24'(9448);
			21529: out = 24'(3380);
			21530: out = 24'(-6648);
			21531: out = 24'(-19584);
			21532: out = 24'(1128);
			21533: out = 24'(22432);
			21534: out = 24'(6844);
			21535: out = 24'(-36620);
			21536: out = 24'(-22740);
			21537: out = 24'(-756);
			21538: out = 24'(3088);
			21539: out = 24'(-13412);
			21540: out = 24'(1572);
			21541: out = 24'(15516);
			21542: out = 24'(21564);
			21543: out = 24'(10940);
			21544: out = 24'(8432);
			21545: out = 24'(220);
			21546: out = 24'(-2664);
			21547: out = 24'(-5276);
			21548: out = 24'(-464);
			21549: out = 24'(-1124);
			21550: out = 24'(4144);
			21551: out = 24'(5708);
			21552: out = 24'(-2988);
			21553: out = 24'(-52);
			21554: out = 24'(-2868);
			21555: out = 24'(8248);
			21556: out = 24'(21484);
			21557: out = 24'(24216);
			21558: out = 24'(4412);
			21559: out = 24'(-5436);
			21560: out = 24'(-8952);
			21561: out = 24'(-16936);
			21562: out = 24'(-27532);
			21563: out = 24'(-2092);
			21564: out = 24'(31000);
			21565: out = 24'(25344);
			21566: out = 24'(-21328);
			21567: out = 24'(-44780);
			21568: out = 24'(-24264);
			21569: out = 24'(9912);
			21570: out = 24'(19604);
			21571: out = 24'(28416);
			21572: out = 24'(21228);
			21573: out = 24'(-6004);
			21574: out = 24'(-10836);
			21575: out = 24'(-16424);
			21576: out = 24'(-6692);
			21577: out = 24'(140);
			21578: out = 24'(7808);
			21579: out = 24'(-620);
			21580: out = 24'(2712);
			21581: out = 24'(7488);
			21582: out = 24'(10516);
			21583: out = 24'(-13592);
			21584: out = 24'(-10620);
			21585: out = 24'(-1040);
			21586: out = 24'(-11176);
			21587: out = 24'(-11752);
			21588: out = 24'(-9408);
			21589: out = 24'(-1908);
			21590: out = 24'(2752);
			21591: out = 24'(34952);
			21592: out = 24'(18512);
			21593: out = 24'(-7824);
			21594: out = 24'(-20256);
			21595: out = 24'(-1656);
			21596: out = 24'(-2784);
			21597: out = 24'(-13480);
			21598: out = 24'(-21172);
			21599: out = 24'(-11920);
			21600: out = 24'(-2608);
			21601: out = 24'(3200);
			21602: out = 24'(2120);
			21603: out = 24'(-144);
			21604: out = 24'(6748);
			21605: out = 24'(32);
			21606: out = 24'(-17140);
			21607: out = 24'(-25124);
			21608: out = 24'(14120);
			21609: out = 24'(15812);
			21610: out = 24'(-4932);
			21611: out = 24'(-18420);
			21612: out = 24'(-296);
			21613: out = 24'(23892);
			21614: out = 24'(29824);
			21615: out = 24'(4288);
			21616: out = 24'(-50400);
			21617: out = 24'(-44460);
			21618: out = 24'(-16872);
			21619: out = 24'(10660);
			21620: out = 24'(26132);
			21621: out = 24'(26852);
			21622: out = 24'(12836);
			21623: out = 24'(-11048);
			21624: out = 24'(-32900);
			21625: out = 24'(-21524);
			21626: out = 24'(-1764);
			21627: out = 24'(18652);
			21628: out = 24'(24108);
			21629: out = 24'(10360);
			21630: out = 24'(1884);
			21631: out = 24'(1252);
			21632: out = 24'(-76);
			21633: out = 24'(2296);
			21634: out = 24'(4136);
			21635: out = 24'(19104);
			21636: out = 24'(19844);
			21637: out = 24'(-276);
			21638: out = 24'(-19124);
			21639: out = 24'(-4584);
			21640: out = 24'(17688);
			21641: out = 24'(19336);
			21642: out = 24'(2128);
			21643: out = 24'(-1420);
			21644: out = 24'(-6564);
			21645: out = 24'(-18004);
			21646: out = 24'(-13516);
			21647: out = 24'(1844);
			21648: out = 24'(6268);
			21649: out = 24'(-112);
			21650: out = 24'(7660);
			21651: out = 24'(16064);
			21652: out = 24'(10540);
			21653: out = 24'(-2592);
			21654: out = 24'(556);
			21655: out = 24'(-4232);
			21656: out = 24'(-3496);
			21657: out = 24'(7112);
			21658: out = 24'(23108);
			21659: out = 24'(4236);
			21660: out = 24'(-22136);
			21661: out = 24'(-33416);
			21662: out = 24'(-16588);
			21663: out = 24'(4848);
			21664: out = 24'(11680);
			21665: out = 24'(10224);
			21666: out = 24'(4396);
			21667: out = 24'(-10684);
			21668: out = 24'(-20448);
			21669: out = 24'(-8504);
			21670: out = 24'(13736);
			21671: out = 24'(24008);
			21672: out = 24'(5932);
			21673: out = 24'(-5352);
			21674: out = 24'(-14320);
			21675: out = 24'(-33052);
			21676: out = 24'(-16712);
			21677: out = 24'(7920);
			21678: out = 24'(15436);
			21679: out = 24'(-6260);
			21680: out = 24'(4516);
			21681: out = 24'(1692);
			21682: out = 24'(-716);
			21683: out = 24'(-492);
			21684: out = 24'(33104);
			21685: out = 24'(12716);
			21686: out = 24'(-17084);
			21687: out = 24'(-30400);
			21688: out = 24'(-336);
			21689: out = 24'(200);
			21690: out = 24'(-1856);
			21691: out = 24'(-3968);
			21692: out = 24'(1092);
			21693: out = 24'(5808);
			21694: out = 24'(13972);
			21695: out = 24'(7464);
			21696: out = 24'(-17092);
			21697: out = 24'(-2076);
			21698: out = 24'(5488);
			21699: out = 24'(5456);
			21700: out = 24'(-6604);
			21701: out = 24'(-6280);
			21702: out = 24'(-7912);
			21703: out = 24'(5288);
			21704: out = 24'(12488);
			21705: out = 24'(-6596);
			21706: out = 24'(-13456);
			21707: out = 24'(920);
			21708: out = 24'(14784);
			21709: out = 24'(-1016);
			21710: out = 24'(0);
			21711: out = 24'(8012);
			21712: out = 24'(13256);
			21713: out = 24'(-1528);
			21714: out = 24'(3384);
			21715: out = 24'(5140);
			21716: out = 24'(5368);
			21717: out = 24'(-8316);
			21718: out = 24'(-17632);
			21719: out = 24'(-14704);
			21720: out = 24'(14100);
			21721: out = 24'(38772);
			21722: out = 24'(45272);
			21723: out = 24'(11844);
			21724: out = 24'(-8592);
			21725: out = 24'(-9136);
			21726: out = 24'(-5972);
			21727: out = 24'(-2904);
			21728: out = 24'(6860);
			21729: out = 24'(11308);
			21730: out = 24'(-1680);
			21731: out = 24'(-2516);
			21732: out = 24'(4748);
			21733: out = 24'(7636);
			21734: out = 24'(-3184);
			21735: out = 24'(712);
			21736: out = 24'(916);
			21737: out = 24'(-13116);
			21738: out = 24'(-34804);
			21739: out = 24'(-3872);
			21740: out = 24'(14132);
			21741: out = 24'(20012);
			21742: out = 24'(9888);
			21743: out = 24'(7236);
			21744: out = 24'(-4260);
			21745: out = 24'(-10668);
			21746: out = 24'(-13856);
			21747: out = 24'(-704);
			21748: out = 24'(2776);
			21749: out = 24'(12020);
			21750: out = 24'(8324);
			21751: out = 24'(-2328);
			21752: out = 24'(-25420);
			21753: out = 24'(-13212);
			21754: out = 24'(872);
			21755: out = 24'(-1992);
			21756: out = 24'(-1716);
			21757: out = 24'(3836);
			21758: out = 24'(4476);
			21759: out = 24'(-3536);
			21760: out = 24'(-13216);
			21761: out = 24'(892);
			21762: out = 24'(5768);
			21763: out = 24'(-6468);
			21764: out = 24'(-20776);
			21765: out = 24'(-6780);
			21766: out = 24'(2784);
			21767: out = 24'(876);
			21768: out = 24'(704);
			21769: out = 24'(5000);
			21770: out = 24'(14028);
			21771: out = 24'(15276);
			21772: out = 24'(3784);
			21773: out = 24'(-3172);
			21774: out = 24'(-23064);
			21775: out = 24'(-29380);
			21776: out = 24'(-17716);
			21777: out = 24'(-868);
			21778: out = 24'(-32);
			21779: out = 24'(8820);
			21780: out = 24'(24332);
			21781: out = 24'(18848);
			21782: out = 24'(6196);
			21783: out = 24'(-17304);
			21784: out = 24'(-32160);
			21785: out = 24'(-27780);
			21786: out = 24'(-5408);
			21787: out = 24'(11012);
			21788: out = 24'(14248);
			21789: out = 24'(12056);
			21790: out = 24'(23056);
			21791: out = 24'(11024);
			21792: out = 24'(-14792);
			21793: out = 24'(-26196);
			21794: out = 24'(3968);
			21795: out = 24'(5260);
			21796: out = 24'(-14884);
			21797: out = 24'(-17532);
			21798: out = 24'(23616);
			21799: out = 24'(35032);
			21800: out = 24'(11128);
			21801: out = 24'(-20028);
			21802: out = 24'(-19292);
			21803: out = 24'(1568);
			21804: out = 24'(5972);
			21805: out = 24'(-3088);
			21806: out = 24'(1620);
			21807: out = 24'(10972);
			21808: out = 24'(18668);
			21809: out = 24'(9184);
			21810: out = 24'(-7800);
			21811: out = 24'(-8880);
			21812: out = 24'(-8032);
			21813: out = 24'(-2564);
			21814: out = 24'(-3988);
			21815: out = 24'(-11460);
			21816: out = 24'(-6984);
			21817: out = 24'(16420);
			21818: out = 24'(29540);
			21819: out = 24'(16352);
			21820: out = 24'(548);
			21821: out = 24'(2008);
			21822: out = 24'(2148);
			21823: out = 24'(-16680);
			21824: out = 24'(-36860);
			21825: out = 24'(-19572);
			21826: out = 24'(7316);
			21827: out = 24'(6012);
			21828: out = 24'(25980);
			21829: out = 24'(8084);
			21830: out = 24'(-364);
			21831: out = 24'(-1088);
			21832: out = 24'(11076);
			21833: out = 24'(-5588);
			21834: out = 24'(-3844);
			21835: out = 24'(9584);
			21836: out = 24'(8724);
			21837: out = 24'(2120);
			21838: out = 24'(-2848);
			21839: out = 24'(1084);
			21840: out = 24'(384);
			21841: out = 24'(-3068);
			21842: out = 24'(-17036);
			21843: out = 24'(-15972);
			21844: out = 24'(5904);
			21845: out = 24'(12148);
			21846: out = 24'(11048);
			21847: out = 24'(1608);
			21848: out = 24'(180);
			21849: out = 24'(5008);
			21850: out = 24'(15704);
			21851: out = 24'(10368);
			21852: out = 24'(-512);
			21853: out = 24'(-2068);
			21854: out = 24'(12488);
			21855: out = 24'(14360);
			21856: out = 24'(4184);
			21857: out = 24'(-7184);
			21858: out = 24'(-3404);
			21859: out = 24'(-9516);
			21860: out = 24'(-12820);
			21861: out = 24'(1428);
			21862: out = 24'(10028);
			21863: out = 24'(11148);
			21864: out = 24'(-6208);
			21865: out = 24'(-21868);
			21866: out = 24'(-2880);
			21867: out = 24'(4544);
			21868: out = 24'(3116);
			21869: out = 24'(-544);
			21870: out = 24'(13272);
			21871: out = 24'(-1708);
			21872: out = 24'(-15268);
			21873: out = 24'(-22844);
			21874: out = 24'(-12304);
			21875: out = 24'(-22612);
			21876: out = 24'(-892);
			21877: out = 24'(27824);
			21878: out = 24'(35704);
			21879: out = 24'(4160);
			21880: out = 24'(-17972);
			21881: out = 24'(-33124);
			21882: out = 24'(-35256);
			21883: out = 24'(-4056);
			21884: out = 24'(23584);
			21885: out = 24'(21556);
			21886: out = 24'(-8296);
			21887: out = 24'(-22192);
			21888: out = 24'(-14376);
			21889: out = 24'(10272);
			21890: out = 24'(13180);
			21891: out = 24'(-3636);
			21892: out = 24'(-7608);
			21893: out = 24'(9048);
			21894: out = 24'(13512);
			21895: out = 24'(-7004);
			21896: out = 24'(-19868);
			21897: out = 24'(-8632);
			21898: out = 24'(7440);
			21899: out = 24'(6060);
			21900: out = 24'(7600);
			21901: out = 24'(7260);
			21902: out = 24'(-2028);
			21903: out = 24'(-27244);
			21904: out = 24'(-35188);
			21905: out = 24'(-23948);
			21906: out = 24'(13048);
			21907: out = 24'(36296);
			21908: out = 24'(30288);
			21909: out = 24'(2608);
			21910: out = 24'(-7744);
			21911: out = 24'(-4608);
			21912: out = 24'(-9880);
			21913: out = 24'(-11808);
			21914: out = 24'(-656);
			21915: out = 24'(17544);
			21916: out = 24'(14648);
			21917: out = 24'(11044);
			21918: out = 24'(460);
			21919: out = 24'(10296);
			21920: out = 24'(13012);
			21921: out = 24'(-1332);
			21922: out = 24'(-36676);
			21923: out = 24'(-28308);
			21924: out = 24'(6268);
			21925: out = 24'(13536);
			21926: out = 24'(2368);
			21927: out = 24'(9472);
			21928: out = 24'(17956);
			21929: out = 24'(-7652);
			21930: out = 24'(-26056);
			21931: out = 24'(-12632);
			21932: out = 24'(15896);
			21933: out = 24'(15036);
			21934: out = 24'(19600);
			21935: out = 24'(9488);
			21936: out = 24'(2488);
			21937: out = 24'(-5732);
			21938: out = 24'(13316);
			21939: out = 24'(5464);
			21940: out = 24'(-2636);
			21941: out = 24'(-5960);
			21942: out = 24'(-1256);
			21943: out = 24'(-1936);
			21944: out = 24'(-2468);
			21945: out = 24'(3664);
			21946: out = 24'(23852);
			21947: out = 24'(23104);
			21948: out = 24'(14368);
			21949: out = 24'(-1148);
			21950: out = 24'(-11680);
			21951: out = 24'(-33152);
			21952: out = 24'(-34716);
			21953: out = 24'(-21524);
			21954: out = 24'(3960);
			21955: out = 24'(10436);
			21956: out = 24'(32088);
			21957: out = 24'(23240);
			21958: out = 24'(-7304);
			21959: out = 24'(-16344);
			21960: out = 24'(-22388);
			21961: out = 24'(-19312);
			21962: out = 24'(-4460);
			21963: out = 24'(30096);
			21964: out = 24'(23764);
			21965: out = 24'(4316);
			21966: out = 24'(-11724);
			21967: out = 24'(-1036);
			21968: out = 24'(-24348);
			21969: out = 24'(-20456);
			21970: out = 24'(-5780);
			21971: out = 24'(8180);
			21972: out = 24'(6416);
			21973: out = 24'(7724);
			21974: out = 24'(2160);
			21975: out = 24'(-5832);
			21976: out = 24'(-696);
			21977: out = 24'(9552);
			21978: out = 24'(9920);
			21979: out = 24'(-6560);
			21980: out = 24'(-11176);
			21981: out = 24'(-29392);
			21982: out = 24'(-16140);
			21983: out = 24'(7836);
			21984: out = 24'(24680);
			21985: out = 24'(14960);
			21986: out = 24'(7148);
			21987: out = 24'(-12776);
			21988: out = 24'(-34776);
			21989: out = 24'(-45472);
			21990: out = 24'(-10420);
			21991: out = 24'(10288);
			21992: out = 24'(-2756);
			21993: out = 24'(-10432);
			21994: out = 24'(8324);
			21995: out = 24'(21596);
			21996: out = 24'(8028);
			21997: out = 24'(-14896);
			21998: out = 24'(-20848);
			21999: out = 24'(-18928);
			22000: out = 24'(-11112);
			22001: out = 24'(4028);
			22002: out = 24'(9888);
			22003: out = 24'(-6732);
			22004: out = 24'(-18084);
			22005: out = 24'(6292);
			22006: out = 24'(40372);
			22007: out = 24'(29512);
			22008: out = 24'(-18948);
			22009: out = 24'(-52824);
			22010: out = 24'(-5032);
			22011: out = 24'(18220);
			22012: out = 24'(7500);
			22013: out = 24'(-11440);
			22014: out = 24'(9704);
			22015: out = 24'(2724);
			22016: out = 24'(752);
			22017: out = 24'(148);
			22018: out = 24'(1876);
			22019: out = 24'(-92);
			22020: out = 24'(9320);
			22021: out = 24'(13164);
			22022: out = 24'(-1600);
			22023: out = 24'(80);
			22024: out = 24'(4348);
			22025: out = 24'(7232);
			22026: out = 24'(-2604);
			22027: out = 24'(2164);
			22028: out = 24'(-4676);
			22029: out = 24'(968);
			22030: out = 24'(8464);
			22031: out = 24'(15572);
			22032: out = 24'(1840);
			22033: out = 24'(6824);
			22034: out = 24'(17912);
			22035: out = 24'(5492);
			22036: out = 24'(-17916);
			22037: out = 24'(-27808);
			22038: out = 24'(-12488);
			22039: out = 24'(7664);
			22040: out = 24'(8232);
			22041: out = 24'(7056);
			22042: out = 24'(8728);
			22043: out = 24'(10888);
			22044: out = 24'(7176);
			22045: out = 24'(7304);
			22046: out = 24'(4012);
			22047: out = 24'(-2516);
			22048: out = 24'(-5388);
			22049: out = 24'(-7668);
			22050: out = 24'(-12188);
			22051: out = 24'(-6496);
			22052: out = 24'(23740);
			22053: out = 24'(16044);
			22054: out = 24'(-8688);
			22055: out = 24'(-22060);
			22056: out = 24'(13728);
			22057: out = 24'(-292);
			22058: out = 24'(-5376);
			22059: out = 24'(-19720);
			22060: out = 24'(-21520);
			22061: out = 24'(-6952);
			22062: out = 24'(27656);
			22063: out = 24'(28984);
			22064: out = 24'(1468);
			22065: out = 24'(-27288);
			22066: out = 24'(-8860);
			22067: out = 24'(5740);
			22068: out = 24'(-1964);
			22069: out = 24'(1448);
			22070: out = 24'(17932);
			22071: out = 24'(20688);
			22072: out = 24'(-5876);
			22073: out = 24'(-37044);
			22074: out = 24'(-37944);
			22075: out = 24'(-14896);
			22076: out = 24'(10060);
			22077: out = 24'(25556);
			22078: out = 24'(19388);
			22079: out = 24'(9712);
			22080: out = 24'(-4960);
			22081: out = 24'(-17060);
			22082: out = 24'(-9240);
			22083: out = 24'(-2400);
			22084: out = 24'(1412);
			22085: out = 24'(-360);
			22086: out = 24'(1144);
			22087: out = 24'(-960);
			22088: out = 24'(380);
			22089: out = 24'(-2272);
			22090: out = 24'(-2916);
			22091: out = 24'(-2448);
			22092: out = 24'(11872);
			22093: out = 24'(14740);
			22094: out = 24'(-1572);
			22095: out = 24'(-29356);
			22096: out = 24'(-19316);
			22097: out = 24'(4052);
			22098: out = 24'(6688);
			22099: out = 24'(2332);
			22100: out = 24'(10960);
			22101: out = 24'(21712);
			22102: out = 24'(14936);
			22103: out = 24'(13228);
			22104: out = 24'(92);
			22105: out = 24'(2624);
			22106: out = 24'(7508);
			22107: out = 24'(10696);
			22108: out = 24'(-15200);
			22109: out = 24'(-17608);
			22110: out = 24'(-7772);
			22111: out = 24'(-18620);
			22112: out = 24'(-18552);
			22113: out = 24'(-7640);
			22114: out = 24'(24824);
			22115: out = 24'(42548);
			22116: out = 24'(23440);
			22117: out = 24'(-5384);
			22118: out = 24'(-8216);
			22119: out = 24'(668);
			22120: out = 24'(-14412);
			22121: out = 24'(-37380);
			22122: out = 24'(-28256);
			22123: out = 24'(10976);
			22124: out = 24'(38456);
			22125: out = 24'(24720);
			22126: out = 24'(10700);
			22127: out = 24'(6496);
			22128: out = 24'(6748);
			22129: out = 24'(-13796);
			22130: out = 24'(-13860);
			22131: out = 24'(-10220);
			22132: out = 24'(-15412);
			22133: out = 24'(3120);
			22134: out = 24'(24892);
			22135: out = 24'(19504);
			22136: out = 24'(-13628);
			22137: out = 24'(-23924);
			22138: out = 24'(-5148);
			22139: out = 24'(12992);
			22140: out = 24'(8668);
			22141: out = 24'(8188);
			22142: out = 24'(6696);
			22143: out = 24'(-1072);
			22144: out = 24'(-13432);
			22145: out = 24'(1592);
			22146: out = 24'(-2004);
			22147: out = 24'(-648);
			22148: out = 24'(-11228);
			22149: out = 24'(-23032);
			22150: out = 24'(-9368);
			22151: out = 24'(10924);
			22152: out = 24'(15748);
			22153: out = 24'(6604);
			22154: out = 24'(10264);
			22155: out = 24'(15016);
			22156: out = 24'(12260);
			22157: out = 24'(-6400);
			22158: out = 24'(-25400);
			22159: out = 24'(-40488);
			22160: out = 24'(-28936);
			22161: out = 24'(2916);
			22162: out = 24'(32388);
			22163: out = 24'(48608);
			22164: out = 24'(39276);
			22165: out = 24'(11232);
			22166: out = 24'(-13392);
			22167: out = 24'(-54128);
			22168: out = 24'(-54912);
			22169: out = 24'(-27340);
			22170: out = 24'(3828);
			22171: out = 24'(12760);
			22172: out = 24'(28176);
			22173: out = 24'(29748);
			22174: out = 24'(13688);
			22175: out = 24'(1884);
			22176: out = 24'(-7004);
			22177: out = 24'(-6384);
			22178: out = 24'(-120);
			22179: out = 24'(-5952);
			22180: out = 24'(-92);
			22181: out = 24'(-5712);
			22182: out = 24'(-3592);
			22183: out = 24'(13384);
			22184: out = 24'(15856);
			22185: out = 24'(4284);
			22186: out = 24'(5416);
			22187: out = 24'(21612);
			22188: out = 24'(4280);
			22189: out = 24'(-29116);
			22190: out = 24'(-31132);
			22191: out = 24'(12892);
			22192: out = 24'(20564);
			22193: out = 24'(9180);
			22194: out = 24'(-8696);
			22195: out = 24'(-7444);
			22196: out = 24'(-7076);
			22197: out = 24'(-1384);
			22198: out = 24'(-3784);
			22199: out = 24'(-2888);
			22200: out = 24'(11080);
			22201: out = 24'(14228);
			22202: out = 24'(21760);
			22203: out = 24'(15916);
			22204: out = 24'(-7980);
			22205: out = 24'(-45332);
			22206: out = 24'(-45644);
			22207: out = 24'(-23996);
			22208: out = 24'(-10896);
			22209: out = 24'(-292);
			22210: out = 24'(12556);
			22211: out = 24'(16544);
			22212: out = 24'(6796);
			22213: out = 24'(18360);
			22214: out = 24'(10124);
			22215: out = 24'(-896);
			22216: out = 24'(-16192);
			22217: out = 24'(-18732);
			22218: out = 24'(-25512);
			22219: out = 24'(-8840);
			22220: out = 24'(13976);
			22221: out = 24'(16140);
			22222: out = 24'(11192);
			22223: out = 24'(-812);
			22224: out = 24'(-4300);
			22225: out = 24'(-5092);
			22226: out = 24'(3660);
			22227: out = 24'(-7424);
			22228: out = 24'(-9064);
			22229: out = 24'(212);
			22230: out = 24'(0);
			22231: out = 24'(-1160);
			22232: out = 24'(10900);
			22233: out = 24'(24864);
			22234: out = 24'(16968);
			22235: out = 24'(5856);
			22236: out = 24'(52);
			22237: out = 24'(-5020);
			22238: out = 24'(-16552);
			22239: out = 24'(-28052);
			22240: out = 24'(-10348);
			22241: out = 24'(16120);
			22242: out = 24'(22032);
			22243: out = 24'(3188);
			22244: out = 24'(-1584);
			22245: out = 24'(-6484);
			22246: out = 24'(-20920);
			22247: out = 24'(-1228);
			22248: out = 24'(9356);
			22249: out = 24'(15028);
			22250: out = 24'(7692);
			22251: out = 24'(1320);
			22252: out = 24'(10976);
			22253: out = 24'(20516);
			22254: out = 24'(8884);
			22255: out = 24'(-11884);
			22256: out = 24'(-28500);
			22257: out = 24'(-14976);
			22258: out = 24'(6868);
			22259: out = 24'(17056);
			22260: out = 24'(13692);
			22261: out = 24'(19152);
			22262: out = 24'(21124);
			22263: out = 24'(9284);
			22264: out = 24'(-7352);
			22265: out = 24'(-14116);
			22266: out = 24'(-13184);
			22267: out = 24'(-16148);
			22268: out = 24'(-32284);
			22269: out = 24'(-1548);
			22270: out = 24'(29596);
			22271: out = 24'(28040);
			22272: out = 24'(-180);
			22273: out = 24'(-6292);
			22274: out = 24'(-4268);
			22275: out = 24'(-12012);
			22276: out = 24'(-28512);
			22277: out = 24'(-24140);
			22278: out = 24'(5296);
			22279: out = 24'(32816);
			22280: out = 24'(34380);
			22281: out = 24'(9936);
			22282: out = 24'(-896);
			22283: out = 24'(-1088);
			22284: out = 24'(-4524);
			22285: out = 24'(-16712);
			22286: out = 24'(-15216);
			22287: out = 24'(-17200);
			22288: out = 24'(-24844);
			22289: out = 24'(-2220);
			22290: out = 24'(4304);
			22291: out = 24'(25296);
			22292: out = 24'(27232);
			22293: out = 24'(8988);
			22294: out = 24'(-31556);
			22295: out = 24'(-22828);
			22296: out = 24'(1448);
			22297: out = 24'(-3020);
			22298: out = 24'(-13104);
			22299: out = 24'(-4380);
			22300: out = 24'(15820);
			22301: out = 24'(12164);
			22302: out = 24'(-7908);
			22303: out = 24'(-32136);
			22304: out = 24'(-31112);
			22305: out = 24'(-15800);
			22306: out = 24'(-3516);
			22307: out = 24'(-18096);
			22308: out = 24'(-11564);
			22309: out = 24'(23748);
			22310: out = 24'(49388);
			22311: out = 24'(38024);
			22312: out = 24'(2788);
			22313: out = 24'(-18372);
			22314: out = 24'(-10032);
			22315: out = 24'(5300);
			22316: out = 24'(60);
			22317: out = 24'(-10736);
			22318: out = 24'(-3208);
			22319: out = 24'(20848);
			22320: out = 24'(12436);
			22321: out = 24'(-19016);
			22322: out = 24'(-38400);
			22323: out = 24'(-8916);
			22324: out = 24'(876);
			22325: out = 24'(-3964);
			22326: out = 24'(-9932);
			22327: out = 24'(2608);
			22328: out = 24'(11868);
			22329: out = 24'(17232);
			22330: out = 24'(12168);
			22331: out = 24'(8236);
			22332: out = 24'(-3320);
			22333: out = 24'(-5116);
			22334: out = 24'(-15708);
			22335: out = 24'(-30564);
			22336: out = 24'(-10296);
			22337: out = 24'(11364);
			22338: out = 24'(20432);
			22339: out = 24'(18080);
			22340: out = 24'(18112);
			22341: out = 24'(33000);
			22342: out = 24'(32872);
			22343: out = 24'(2640);
			22344: out = 24'(-47928);
			22345: out = 24'(-29384);
			22346: out = 24'(8960);
			22347: out = 24'(20920);
			22348: out = 24'(-608);
			22349: out = 24'(6012);
			22350: out = 24'(4288);
			22351: out = 24'(-9724);
			22352: out = 24'(-26576);
			22353: out = 24'(6228);
			22354: out = 24'(17768);
			22355: out = 24'(11324);
			22356: out = 24'(-512);
			22357: out = 24'(7120);
			22358: out = 24'(1872);
			22359: out = 24'(-1856);
			22360: out = 24'(2872);
			22361: out = 24'(12676);
			22362: out = 24'(17580);
			22363: out = 24'(8524);
			22364: out = 24'(-2416);
			22365: out = 24'(-596);
			22366: out = 24'(-10372);
			22367: out = 24'(-18288);
			22368: out = 24'(-16276);
			22369: out = 24'(1932);
			22370: out = 24'(-1128);
			22371: out = 24'(10728);
			22372: out = 24'(19252);
			22373: out = 24'(12444);
			22374: out = 24'(-20556);
			22375: out = 24'(-20960);
			22376: out = 24'(6156);
			22377: out = 24'(31796);
			22378: out = 24'(27920);
			22379: out = 24'(7780);
			22380: out = 24'(-10532);
			22381: out = 24'(-9884);
			22382: out = 24'(4292);
			22383: out = 24'(-10472);
			22384: out = 24'(-35848);
			22385: out = 24'(-39340);
			22386: out = 24'(3588);
			22387: out = 24'(-2068);
			22388: out = 24'(7948);
			22389: out = 24'(10308);
			22390: out = 24'(10940);
			22391: out = 24'(-1960);
			22392: out = 24'(9844);
			22393: out = 24'(9208);
			22394: out = 24'(-4208);
			22395: out = 24'(-28556);
			22396: out = 24'(-16392);
			22397: out = 24'(-18192);
			22398: out = 24'(-24604);
			22399: out = 24'(1316);
			22400: out = 24'(15544);
			22401: out = 24'(10332);
			22402: out = 24'(-744);
			22403: out = 24'(8796);
			22404: out = 24'(8028);
			22405: out = 24'(-7088);
			22406: out = 24'(-22564);
			22407: out = 24'(-12300);
			22408: out = 24'(88);
			22409: out = 24'(8344);
			22410: out = 24'(7404);
			22411: out = 24'(7556);
			22412: out = 24'(592);
			22413: out = 24'(-12448);
			22414: out = 24'(-25324);
			22415: out = 24'(-24404);
			22416: out = 24'(-11188);
			22417: out = 24'(-568);
			22418: out = 24'(5996);
			22419: out = 24'(9788);
			22420: out = 24'(8496);
			22421: out = 24'(3124);
			22422: out = 24'(684);
			22423: out = 24'(3580);
			22424: out = 24'(9264);
			22425: out = 24'(10888);
			22426: out = 24'(19892);
			22427: out = 24'(24220);
			22428: out = 24'(12324);
			22429: out = 24'(-20200);
			22430: out = 24'(-20016);
			22431: out = 24'(-960);
			22432: out = 24'(5616);
			22433: out = 24'(-2124);
			22434: out = 24'(-3556);
			22435: out = 24'(13780);
			22436: out = 24'(20284);
			22437: out = 24'(552);
			22438: out = 24'(3128);
			22439: out = 24'(25404);
			22440: out = 24'(32504);
			22441: out = 24'(2804);
			22442: out = 24'(-3716);
			22443: out = 24'(-8624);
			22444: out = 24'(-16644);
			22445: out = 24'(-34004);
			22446: out = 24'(-14264);
			22447: out = 24'(592);
			22448: out = 24'(11364);
			22449: out = 24'(15676);
			22450: out = 24'(28824);
			22451: out = 24'(20908);
			22452: out = 24'(4252);
			22453: out = 24'(-14852);
			22454: out = 24'(-24868);
			22455: out = 24'(-11248);
			22456: out = 24'(2836);
			22457: out = 24'(5256);
			22458: out = 24'(-1216);
			22459: out = 24'(-512);
			22460: out = 24'(-776);
			22461: out = 24'(-2396);
			22462: out = 24'(-9248);
			22463: out = 24'(6680);
			22464: out = 24'(-3216);
			22465: out = 24'(-12796);
			22466: out = 24'(-15436);
			22467: out = 24'(7484);
			22468: out = 24'(8);
			22469: out = 24'(10124);
			22470: out = 24'(24584);
			22471: out = 24'(22480);
			22472: out = 24'(-33388);
			22473: out = 24'(-55796);
			22474: out = 24'(-26072);
			22475: out = 24'(13808);
			22476: out = 24'(3960);
			22477: out = 24'(4064);
			22478: out = 24'(17128);
			22479: out = 24'(20912);
			22480: out = 24'(-14716);
			22481: out = 24'(-19564);
			22482: out = 24'(-2856);
			22483: out = 24'(4348);
			22484: out = 24'(-25028);
			22485: out = 24'(-24924);
			22486: out = 24'(-7340);
			22487: out = 24'(13328);
			22488: out = 24'(23660);
			22489: out = 24'(37416);
			22490: out = 24'(24408);
			22491: out = 24'(-13308);
			22492: out = 24'(-59160);
			22493: out = 24'(-40628);
			22494: out = 24'(-18016);
			22495: out = 24'(-7400);
			22496: out = 24'(3344);
			22497: out = 24'(13324);
			22498: out = 24'(23592);
			22499: out = 24'(22596);
			22500: out = 24'(12600);
			22501: out = 24'(-5584);
			22502: out = 24'(-17948);
			22503: out = 24'(-31412);
			22504: out = 24'(-37408);
			22505: out = 24'(-10516);
			22506: out = 24'(9356);
			22507: out = 24'(23772);
			22508: out = 24'(22440);
			22509: out = 24'(8792);
			22510: out = 24'(-9956);
			22511: out = 24'(-18628);
			22512: out = 24'(-15888);
			22513: out = 24'(-4784);
			22514: out = 24'(6392);
			22515: out = 24'(20072);
			22516: out = 24'(26932);
			22517: out = 24'(22732);
			22518: out = 24'(3208);
			22519: out = 24'(-3188);
			22520: out = 24'(-2624);
			22521: out = 24'(3704);
			22522: out = 24'(16528);
			22523: out = 24'(8156);
			22524: out = 24'(-16244);
			22525: out = 24'(-27412);
			22526: out = 24'(9456);
			22527: out = 24'(40576);
			22528: out = 24'(41476);
			22529: out = 24'(9116);
			22530: out = 24'(-14332);
			22531: out = 24'(-24232);
			22532: out = 24'(-808);
			22533: out = 24'(9048);
			22534: out = 24'(-2060);
			22535: out = 24'(-12400);
			22536: out = 24'(6516);
			22537: out = 24'(19048);
			22538: out = 24'(11920);
			22539: out = 24'(10516);
			22540: out = 24'(10712);
			22541: out = 24'(-3444);
			22542: out = 24'(-30788);
			22543: out = 24'(-30428);
			22544: out = 24'(-11688);
			22545: out = 24'(15900);
			22546: out = 24'(21144);
			22547: out = 24'(10816);
			22548: out = 24'(0);
			22549: out = 24'(7176);
			22550: out = 24'(11240);
			22551: out = 24'(-3572);
			22552: out = 24'(-14088);
			22553: out = 24'(-17336);
			22554: out = 24'(-4716);
			22555: out = 24'(6496);
			22556: out = 24'(120);
			22557: out = 24'(-7564);
			22558: out = 24'(-2328);
			22559: out = 24'(7840);
			22560: out = 24'(-304);
			22561: out = 24'(-8592);
			22562: out = 24'(-8972);
			22563: out = 24'(3708);
			22564: out = 24'(5652);
			22565: out = 24'(9684);
			22566: out = 24'(-3980);
			22567: out = 24'(-12292);
			22568: out = 24'(-7736);
			22569: out = 24'(2464);
			22570: out = 24'(-3528);
			22571: out = 24'(-5800);
			22572: out = 24'(4488);
			22573: out = 24'(544);
			22574: out = 24'(-56);
			22575: out = 24'(6872);
			22576: out = 24'(17568);
			22577: out = 24'(-104);
			22578: out = 24'(16784);
			22579: out = 24'(26912);
			22580: out = 24'(12612);
			22581: out = 24'(-32060);
			22582: out = 24'(-35372);
			22583: out = 24'(-16196);
			22584: out = 24'(5588);
			22585: out = 24'(5984);
			22586: out = 24'(2508);
			22587: out = 24'(-4620);
			22588: out = 24'(796);
			22589: out = 24'(11472);
			22590: out = 24'(14392);
			22591: out = 24'(-3412);
			22592: out = 24'(-26896);
			22593: out = 24'(-31844);
			22594: out = 24'(4892);
			22595: out = 24'(17412);
			22596: out = 24'(14124);
			22597: out = 24'(5864);
			22598: out = 24'(404);
			22599: out = 24'(-2680);
			22600: out = 24'(-10060);
			22601: out = 24'(-16344);
			22602: out = 24'(-10392);
			22603: out = 24'(-2156);
			22604: out = 24'(6152);
			22605: out = 24'(6284);
			22606: out = 24'(1076);
			22607: out = 24'(6656);
			22608: out = 24'(10776);
			22609: out = 24'(7804);
			22610: out = 24'(120);
			22611: out = 24'(7188);
			22612: out = 24'(3396);
			22613: out = 24'(-5308);
			22614: out = 24'(-10252);
			22615: out = 24'(7308);
			22616: out = 24'(7708);
			22617: out = 24'(4292);
			22618: out = 24'(-2868);
			22619: out = 24'(-3428);
			22620: out = 24'(-5788);
			22621: out = 24'(472);
			22622: out = 24'(1204);
			22623: out = 24'(-5008);
			22624: out = 24'(-28892);
			22625: out = 24'(-12240);
			22626: out = 24'(23096);
			22627: out = 24'(35688);
			22628: out = 24'(14876);
			22629: out = 24'(-12740);
			22630: out = 24'(-31776);
			22631: out = 24'(-33872);
			22632: out = 24'(-12916);
			22633: out = 24'(5852);
			22634: out = 24'(16788);
			22635: out = 24'(17120);
			22636: out = 24'(11608);
			22637: out = 24'(-380);
			22638: out = 24'(-5360);
			22639: out = 24'(-3052);
			22640: out = 24'(-4796);
			22641: out = 24'(-6308);
			22642: out = 24'(-5932);
			22643: out = 24'(8584);
			22644: out = 24'(23720);
			22645: out = 24'(19676);
			22646: out = 24'(2320);
			22647: out = 24'(-4772);
			22648: out = 24'(-3324);
			22649: out = 24'(-22368);
			22650: out = 24'(-32736);
			22651: out = 24'(-16800);
			22652: out = 24'(12304);
			22653: out = 24'(6476);
			22654: out = 24'(8680);
			22655: out = 24'(11596);
			22656: out = 24'(18404);
			22657: out = 24'(8864);
			22658: out = 24'(5636);
			22659: out = 24'(-1096);
			22660: out = 24'(2848);
			22661: out = 24'(5148);
			22662: out = 24'(1920);
			22663: out = 24'(-15924);
			22664: out = 24'(-10236);
			22665: out = 24'(21316);
			22666: out = 24'(21488);
			22667: out = 24'(9408);
			22668: out = 24'(-9620);
			22669: out = 24'(-9836);
			22670: out = 24'(-2960);
			22671: out = 24'(4204);
			22672: out = 24'(-3656);
			22673: out = 24'(1440);
			22674: out = 24'(21924);
			22675: out = 24'(28020);
			22676: out = 24'(7512);
			22677: out = 24'(-5252);
			22678: out = 24'(5304);
			22679: out = 24'(1064);
			22680: out = 24'(-27164);
			22681: out = 24'(-38344);
			22682: out = 24'(-3016);
			22683: out = 24'(2908);
			22684: out = 24'(9488);
			22685: out = 24'(2304);
			22686: out = 24'(104);
			22687: out = 24'(-1548);
			22688: out = 24'(140);
			22689: out = 24'(1036);
			22690: out = 24'(10344);
			22691: out = 24'(14548);
			22692: out = 24'(10900);
			22693: out = 24'(-11752);
			22694: out = 24'(-26440);
			22695: out = 24'(-15084);
			22696: out = 24'(5720);
			22697: out = 24'(8384);
			22698: out = 24'(-4152);
			22699: out = 24'(-12592);
			22700: out = 24'(-13552);
			22701: out = 24'(-4228);
			22702: out = 24'(2156);
			22703: out = 24'(2256);
			22704: out = 24'(-420);
			22705: out = 24'(8708);
			22706: out = 24'(20212);
			22707: out = 24'(20712);
			22708: out = 24'(9664);
			22709: out = 24'(-29968);
			22710: out = 24'(-48572);
			22711: out = 24'(-30536);
			22712: out = 24'(216);
			22713: out = 24'(2316);
			22714: out = 24'(-3004);
			22715: out = 24'(876);
			22716: out = 24'(12512);
			22717: out = 24'(17712);
			22718: out = 24'(7768);
			22719: out = 24'(-5700);
			22720: out = 24'(-12176);
			22721: out = 24'(-12292);
			22722: out = 24'(-6556);
			22723: out = 24'(-1416);
			22724: out = 24'(2396);
			22725: out = 24'(11320);
			22726: out = 24'(8676);
			22727: out = 24'(2520);
			22728: out = 24'(-7904);
			22729: out = 24'(-10108);
			22730: out = 24'(-3764);
			22731: out = 24'(12764);
			22732: out = 24'(13368);
			22733: out = 24'(-808);
			22734: out = 24'(-5352);
			22735: out = 24'(15576);
			22736: out = 24'(26952);
			22737: out = 24'(12552);
			22738: out = 24'(-6340);
			22739: out = 24'(-516);
			22740: out = 24'(11240);
			22741: out = 24'(1980);
			22742: out = 24'(-39696);
			22743: out = 24'(-15348);
			22744: out = 24'(19980);
			22745: out = 24'(29264);
			22746: out = 24'(9208);
			22747: out = 24'(868);
			22748: out = 24'(-3316);
			22749: out = 24'(72);
			22750: out = 24'(1620);
			22751: out = 24'(16072);
			22752: out = 24'(9328);
			22753: out = 24'(10520);
			22754: out = 24'(22072);
			22755: out = 24'(10064);
			22756: out = 24'(-7076);
			22757: out = 24'(-12428);
			22758: out = 24'(-1068);
			22759: out = 24'(-7496);
			22760: out = 24'(-11112);
			22761: out = 24'(-11040);
			22762: out = 24'(3724);
			22763: out = 24'(14328);
			22764: out = 24'(17756);
			22765: out = 24'(5928);
			22766: out = 24'(-4592);
			22767: out = 24'(-11320);
			22768: out = 24'(-19472);
			22769: out = 24'(-23968);
			22770: out = 24'(-14868);
			22771: out = 24'(-1296);
			22772: out = 24'(132);
			22773: out = 24'(-1976);
			22774: out = 24'(156);
			22775: out = 24'(-456);
			22776: out = 24'(18372);
			22777: out = 24'(-11164);
			22778: out = 24'(-15236);
			22779: out = 24'(2340);
			22780: out = 24'(-1424);
			22781: out = 24'(-9612);
			22782: out = 24'(-4988);
			22783: out = 24'(13340);
			22784: out = 24'(21944);
			22785: out = 24'(4248);
			22786: out = 24'(-8448);
			22787: out = 24'(-17856);
			22788: out = 24'(-27200);
			22789: out = 24'(-4292);
			22790: out = 24'(17140);
			22791: out = 24'(21108);
			22792: out = 24'(6572);
			22793: out = 24'(-14652);
			22794: out = 24'(-5016);
			22795: out = 24'(5268);
			22796: out = 24'(-2124);
			22797: out = 24'(-23476);
			22798: out = 24'(5540);
			22799: out = 24'(19912);
			22800: out = 24'(-1528);
			22801: out = 24'(-33780);
			22802: out = 24'(11220);
			22803: out = 24'(37116);
			22804: out = 24'(8040);
			22805: out = 24'(-40752);
			22806: out = 24'(-27388);
			22807: out = 24'(2684);
			22808: out = 24'(1604);
			22809: out = 24'(-25284);
			22810: out = 24'(-16848);
			22811: out = 24'(14856);
			22812: out = 24'(36476);
			22813: out = 24'(26920);
			22814: out = 24'(12224);
			22815: out = 24'(5780);
			22816: out = 24'(4696);
			22817: out = 24'(-5732);
			22818: out = 24'(-19108);
			22819: out = 24'(-30772);
			22820: out = 24'(-19844);
			22821: out = 24'(7920);
			22822: out = 24'(31068);
			22823: out = 24'(20172);
			22824: out = 24'(4904);
			22825: out = 24'(-1428);
			22826: out = 24'(1968);
			22827: out = 24'(-4300);
			22828: out = 24'(-6252);
			22829: out = 24'(652);
			22830: out = 24'(9644);
			22831: out = 24'(-368);
			22832: out = 24'(-4216);
			22833: out = 24'(-1052);
			22834: out = 24'(8500);
			22835: out = 24'(8244);
			22836: out = 24'(2572);
			22837: out = 24'(-12156);
			22838: out = 24'(-20888);
			22839: out = 24'(-14772);
			22840: out = 24'(2584);
			22841: out = 24'(12308);
			22842: out = 24'(13804);
			22843: out = 24'(16360);
			22844: out = 24'(6524);
			22845: out = 24'(2560);
			22846: out = 24'(-6112);
			22847: out = 24'(-12488);
			22848: out = 24'(-13640);
			22849: out = 24'(-3044);
			22850: out = 24'(-1960);
			22851: out = 24'(-2936);
			22852: out = 24'(5836);
			22853: out = 24'(8172);
			22854: out = 24'(-2776);
			22855: out = 24'(-14656);
			22856: out = 24'(-20008);
			22857: out = 24'(-580);
			22858: out = 24'(1312);
			22859: out = 24'(1392);
			22860: out = 24'(7368);
			22861: out = 24'(22616);
			22862: out = 24'(5780);
			22863: out = 24'(-5120);
			22864: out = 24'(2488);
			22865: out = 24'(568);
			22866: out = 24'(-30244);
			22867: out = 24'(-42804);
			22868: out = 24'(-13896);
			22869: out = 24'(11120);
			22870: out = 24'(6816);
			22871: out = 24'(-1320);
			22872: out = 24'(8464);
			22873: out = 24'(15420);
			22874: out = 24'(13852);
			22875: out = 24'(1372);
			22876: out = 24'(-5112);
			22877: out = 24'(-4344);
			22878: out = 24'(1952);
			22879: out = 24'(1600);
			22880: out = 24'(-668);
			22881: out = 24'(848);
			22882: out = 24'(11936);
			22883: out = 24'(11132);
			22884: out = 24'(-3928);
			22885: out = 24'(-20696);
			22886: out = 24'(-11764);
			22887: out = 24'(-3084);
			22888: out = 24'(176);
			22889: out = 24'(-6236);
			22890: out = 24'(-5984);
			22891: out = 24'(5092);
			22892: out = 24'(20280);
			22893: out = 24'(17696);
			22894: out = 24'(-244);
			22895: out = 24'(-5028);
			22896: out = 24'(2296);
			22897: out = 24'(6388);
			22898: out = 24'(1656);
			22899: out = 24'(-4508);
			22900: out = 24'(-1804);
			22901: out = 24'(-396);
			22902: out = 24'(236);
			22903: out = 24'(-1348);
			22904: out = 24'(8268);
			22905: out = 24'(5608);
			22906: out = 24'(-800);
			22907: out = 24'(-848);
			22908: out = 24'(29008);
			22909: out = 24'(28304);
			22910: out = 24'(-236);
			22911: out = 24'(-32208);
			22912: out = 24'(-17292);
			22913: out = 24'(-9628);
			22914: out = 24'(-5936);
			22915: out = 24'(3836);
			22916: out = 24'(21156);
			22917: out = 24'(10496);
			22918: out = 24'(-1268);
			22919: out = 24'(-424);
			22920: out = 24'(1960);
			22921: out = 24'(-11500);
			22922: out = 24'(-11428);
			22923: out = 24'(5032);
			22924: out = 24'(5424);
			22925: out = 24'(980);
			22926: out = 24'(5900);
			22927: out = 24'(17048);
			22928: out = 24'(6732);
			22929: out = 24'(-16812);
			22930: out = 24'(-27420);
			22931: out = 24'(-12000);
			22932: out = 24'(1016);
			22933: out = 24'(1988);
			22934: out = 24'(-4756);
			22935: out = 24'(-1944);
			22936: out = 24'(-2368);
			22937: out = 24'(-9256);
			22938: out = 24'(-15460);
			22939: out = 24'(3212);
			22940: out = 24'(23924);
			22941: out = 24'(17036);
			22942: out = 24'(-5204);
			22943: out = 24'(-9276);
			22944: out = 24'(1852);
			22945: out = 24'(-1336);
			22946: out = 24'(-3448);
			22947: out = 24'(-2796);
			22948: out = 24'(-1916);
			22949: out = 24'(-13248);
			22950: out = 24'(-18212);
			22951: out = 24'(-16000);
			22952: out = 24'(-7932);
			22953: out = 24'(-1920);
			22954: out = 24'(15580);
			22955: out = 24'(22776);
			22956: out = 24'(15600);
			22957: out = 24'(-5404);
			22958: out = 24'(-13568);
			22959: out = 24'(-20348);
			22960: out = 24'(-12824);
			22961: out = 24'(-1668);
			22962: out = 24'(592);
			22963: out = 24'(6388);
			22964: out = 24'(8284);
			22965: out = 24'(5940);
			22966: out = 24'(300);
			22967: out = 24'(6760);
			22968: out = 24'(8);
			22969: out = 24'(-11484);
			22970: out = 24'(-6948);
			22971: out = 24'(25956);
			22972: out = 24'(36520);
			22973: out = 24'(12536);
			22974: out = 24'(-23928);
			22975: out = 24'(-23164);
			22976: out = 24'(-16700);
			22977: out = 24'(-7196);
			22978: out = 24'(-3548);
			22979: out = 24'(1296);
			22980: out = 24'(12108);
			22981: out = 24'(22956);
			22982: out = 24'(14032);
			22983: out = 24'(-19852);
			22984: out = 24'(-4316);
			22985: out = 24'(5544);
			22986: out = 24'(4572);
			22987: out = 24'(-316);
			22988: out = 24'(5496);
			22989: out = 24'(7844);
			22990: out = 24'(3500);
			22991: out = 24'(988);
			22992: out = 24'(8360);
			22993: out = 24'(15704);
			22994: out = 24'(9512);
			22995: out = 24'(-2428);
			22996: out = 24'(-1512);
			22997: out = 24'(-9892);
			22998: out = 24'(-13056);
			22999: out = 24'(-4044);
			23000: out = 24'(6036);
			23001: out = 24'(39564);
			23002: out = 24'(27792);
			23003: out = 24'(-556);
			23004: out = 24'(-8624);
			23005: out = 24'(-3376);
			23006: out = 24'(-17092);
			23007: out = 24'(-42420);
			23008: out = 24'(-38148);
			23009: out = 24'(-816);
			23010: out = 24'(32120);
			23011: out = 24'(28180);
			23012: out = 24'(10008);
			23013: out = 24'(1648);
			23014: out = 24'(928);
			23015: out = 24'(-10424);
			23016: out = 24'(-19400);
			23017: out = 24'(-5084);
			23018: out = 24'(968);
			23019: out = 24'(3532);
			23020: out = 24'(11104);
			23021: out = 24'(20160);
			23022: out = 24'(4428);
			23023: out = 24'(-22648);
			23024: out = 24'(-25308);
			23025: out = 24'(1792);
			23026: out = 24'(6144);
			23027: out = 24'(-3164);
			23028: out = 24'(-4740);
			23029: out = 24'(7968);
			23030: out = 24'(6552);
			23031: out = 24'(-7260);
			23032: out = 24'(-5052);
			23033: out = 24'(11508);
			23034: out = 24'(-2264);
			23035: out = 24'(-25600);
			23036: out = 24'(-35832);
			23037: out = 24'(-13172);
			23038: out = 24'(1356);
			23039: out = 24'(25816);
			23040: out = 24'(15408);
			23041: out = 24'(6340);
			23042: out = 24'(5816);
			23043: out = 24'(2308);
			23044: out = 24'(-19680);
			23045: out = 24'(-32052);
			23046: out = 24'(-19188);
			23047: out = 24'(-1436);
			23048: out = 24'(1788);
			23049: out = 24'(3384);
			23050: out = 24'(14172);
			23051: out = 24'(15844);
			23052: out = 24'(7020);
			23053: out = 24'(-10028);
			23054: out = 24'(-23256);
			23055: out = 24'(-43788);
			23056: out = 24'(-17132);
			23057: out = 24'(-2172);
			23058: out = 24'(6020);
			23059: out = 24'(15836);
			23060: out = 24'(24244);
			23061: out = 24'(11784);
			23062: out = 24'(-2048);
			23063: out = 24'(2080);
			23064: out = 24'(-428);
			23065: out = 24'(2688);
			23066: out = 24'(-4084);
			23067: out = 24'(-8360);
			23068: out = 24'(10100);
			23069: out = 24'(7536);
			23070: out = 24'(-192);
			23071: out = 24'(5172);
			23072: out = 24'(22068);
			23073: out = 24'(25648);
			23074: out = 24'(5716);
			23075: out = 24'(-15296);
			23076: out = 24'(-9088);
			23077: out = 24'(16092);
			23078: out = 24'(26664);
			23079: out = 24'(13420);
			23080: out = 24'(-4824);
			23081: out = 24'(1020);
			23082: out = 24'(11908);
			23083: out = 24'(11776);
			23084: out = 24'(-4336);
			23085: out = 24'(-6676);
			23086: out = 24'(-9596);
			23087: out = 24'(7044);
			23088: out = 24'(23252);
			23089: out = 24'(24376);
			23090: out = 24'(8872);
			23091: out = 24'(5992);
			23092: out = 24'(2956);
			23093: out = 24'(-22028);
			23094: out = 24'(-20288);
			23095: out = 24'(-1444);
			23096: out = 24'(11780);
			23097: out = 24'(-4052);
			23098: out = 24'(-1076);
			23099: out = 24'(-3104);
			23100: out = 24'(-692);
			23101: out = 24'(-3424);
			23102: out = 24'(-11540);
			23103: out = 24'(-19616);
			23104: out = 24'(-18556);
			23105: out = 24'(-10072);
			23106: out = 24'(1216);
			23107: out = 24'(384);
			23108: out = 24'(440);
			23109: out = 24'(12812);
			23110: out = 24'(29172);
			23111: out = 24'(25952);
			23112: out = 24'(1112);
			23113: out = 24'(-26156);
			23114: out = 24'(-40652);
			23115: out = 24'(-11244);
			23116: out = 24'(-2652);
			23117: out = 24'(-7932);
			23118: out = 24'(-11668);
			23119: out = 24'(-1516);
			23120: out = 24'(-960);
			23121: out = 24'(6520);
			23122: out = 24'(15552);
			23123: out = 24'(-52);
			23124: out = 24'(-18724);
			23125: out = 24'(-15400);
			23126: out = 24'(6764);
			23127: out = 24'(-2464);
			23128: out = 24'(2456);
			23129: out = 24'(-6788);
			23130: out = 24'(-14520);
			23131: out = 24'(-27436);
			23132: out = 24'(-232);
			23133: out = 24'(4800);
			23134: out = 24'(7644);
			23135: out = 24'(13476);
			23136: out = 24'(3056);
			23137: out = 24'(-8648);
			23138: out = 24'(-5400);
			23139: out = 24'(9988);
			23140: out = 24'(16544);
			23141: out = 24'(-1752);
			23142: out = 24'(-18148);
			23143: out = 24'(-17344);
			23144: out = 24'(-11496);
			23145: out = 24'(3308);
			23146: out = 24'(17068);
			23147: out = 24'(23664);
			23148: out = 24'(15860);
			23149: out = 24'(3648);
			23150: out = 24'(-7492);
			23151: out = 24'(-13048);
			23152: out = 24'(-10060);
			23153: out = 24'(4424);
			23154: out = 24'(5108);
			23155: out = 24'(-7156);
			23156: out = 24'(-6488);
			23157: out = 24'(18644);
			23158: out = 24'(41420);
			23159: out = 24'(22048);
			23160: out = 24'(-12420);
			23161: out = 24'(-1016);
			23162: out = 24'(-244);
			23163: out = 24'(-11632);
			23164: out = 24'(-23568);
			23165: out = 24'(-2764);
			23166: out = 24'(17280);
			23167: out = 24'(17188);
			23168: out = 24'(-576);
			23169: out = 24'(-2100);
			23170: out = 24'(10684);
			23171: out = 24'(26444);
			23172: out = 24'(17956);
			23173: out = 24'(-5184);
			23174: out = 24'(-19548);
			23175: out = 24'(-17716);
			23176: out = 24'(-7620);
			23177: out = 24'(1484);
			23178: out = 24'(15220);
			23179: out = 24'(13728);
			23180: out = 24'(4388);
			23181: out = 24'(-9456);
			23182: out = 24'(-8188);
			23183: out = 24'(-14720);
			23184: out = 24'(-5824);
			23185: out = 24'(-1272);
			23186: out = 24'(524);
			23187: out = 24'(2816);
			23188: out = 24'(18568);
			23189: out = 24'(9824);
			23190: out = 24'(-24880);
			23191: out = 24'(-39328);
			23192: out = 24'(-23824);
			23193: out = 24'(-6044);
			23194: out = 24'(-2204);
			23195: out = 24'(16828);
			23196: out = 24'(26208);
			23197: out = 24'(20700);
			23198: out = 24'(1244);
			23199: out = 24'(-3920);
			23200: out = 24'(-17728);
			23201: out = 24'(-23408);
			23202: out = 24'(-17836);
			23203: out = 24'(9300);
			23204: out = 24'(14400);
			23205: out = 24'(14996);
			23206: out = 24'(4904);
			23207: out = 24'(860);
			23208: out = 24'(-2688);
			23209: out = 24'(20780);
			23210: out = 24'(27056);
			23211: out = 24'(620);
			23212: out = 24'(-31484);
			23213: out = 24'(-53340);
			23214: out = 24'(-38584);
			23215: out = 24'(-2860);
			23216: out = 24'(12356);
			23217: out = 24'(11084);
			23218: out = 24'(8112);
			23219: out = 24'(18956);
			23220: out = 24'(19348);
			23221: out = 24'(-1360);
			23222: out = 24'(-33628);
			23223: out = 24'(-27332);
			23224: out = 24'(8104);
			23225: out = 24'(19292);
			23226: out = 24'(-9372);
			23227: out = 24'(-15600);
			23228: out = 24'(14540);
			23229: out = 24'(16720);
			23230: out = 24'(-9904);
			23231: out = 24'(-19596);
			23232: out = 24'(9464);
			23233: out = 24'(28640);
			23234: out = 24'(15800);
			23235: out = 24'(-132);
			23236: out = 24'(420);
			23237: out = 24'(-6228);
			23238: out = 24'(-3900);
			23239: out = 24'(-3060);
			23240: out = 24'(84);
			23241: out = 24'(-4648);
			23242: out = 24'(14588);
			23243: out = 24'(12316);
			23244: out = 24'(-508);
			23245: out = 24'(-12620);
			23246: out = 24'(-12612);
			23247: out = 24'(248);
			23248: out = 24'(10060);
			23249: out = 24'(8020);
			23250: out = 24'(-3884);
			23251: out = 24'(2768);
			23252: out = 24'(6644);
			23253: out = 24'(-2780);
			23254: out = 24'(-18960);
			23255: out = 24'(-5856);
			23256: out = 24'(5784);
			23257: out = 24'(4560);
			23258: out = 24'(424);
			23259: out = 24'(-1260);
			23260: out = 24'(4516);
			23261: out = 24'(5012);
			23262: out = 24'(-3412);
			23263: out = 24'(-28448);
			23264: out = 24'(-24260);
			23265: out = 24'(-5128);
			23266: out = 24'(10020);
			23267: out = 24'(22604);
			23268: out = 24'(25648);
			23269: out = 24'(18804);
			23270: out = 24'(692);
			23271: out = 24'(-10500);
			23272: out = 24'(-20600);
			23273: out = 24'(-12400);
			23274: out = 24'(-3708);
			23275: out = 24'(-4392);
			23276: out = 24'(-17532);
			23277: out = 24'(-10252);
			23278: out = 24'(7348);
			23279: out = 24'(17136);
			23280: out = 24'(13940);
			23281: out = 24'(15988);
			23282: out = 24'(8436);
			23283: out = 24'(-16996);
			23284: out = 24'(-28768);
			23285: out = 24'(-21488);
			23286: out = 24'(-1636);
			23287: out = 24'(2388);
			23288: out = 24'(10184);
			23289: out = 24'(-936);
			23290: out = 24'(15232);
			23291: out = 24'(29092);
			23292: out = 24'(22120);
			23293: out = 24'(-15988);
			23294: out = 24'(-16196);
			23295: out = 24'(11352);
			23296: out = 24'(29836);
			23297: out = 24'(9588);
			23298: out = 24'(640);
			23299: out = 24'(-6072);
			23300: out = 24'(-12388);
			23301: out = 24'(-7160);
			23302: out = 24'(1608);
			23303: out = 24'(-4628);
			23304: out = 24'(-7664);
			23305: out = 24'(22376);
			23306: out = 24'(31284);
			23307: out = 24'(3484);
			23308: out = 24'(-27620);
			23309: out = 24'(-16540);
			23310: out = 24'(-5848);
			23311: out = 24'(-22628);
			23312: out = 24'(-38344);
			23313: out = 24'(-8060);
			23314: out = 24'(10036);
			23315: out = 24'(8168);
			23316: out = 24'(2208);
			23317: out = 24'(21472);
			23318: out = 24'(33636);
			23319: out = 24'(21084);
			23320: out = 24'(-12840);
			23321: out = 24'(-36360);
			23322: out = 24'(-20972);
			23323: out = 24'(-13992);
			23324: out = 24'(-6376);
			23325: out = 24'(5280);
			23326: out = 24'(26388);
			23327: out = 24'(18196);
			23328: out = 24'(17140);
			23329: out = 24'(11072);
			23330: out = 24'(-5796);
			23331: out = 24'(-36356);
			23332: out = 24'(-22240);
			23333: out = 24'(9736);
			23334: out = 24'(14088);
			23335: out = 24'(2696);
			23336: out = 24'(-5524);
			23337: out = 24'(-1472);
			23338: out = 24'(2500);
			23339: out = 24'(120);
			23340: out = 24'(84);
			23341: out = 24'(-4368);
			23342: out = 24'(-14584);
			23343: out = 24'(-22560);
			23344: out = 24'(-1108);
			23345: out = 24'(12876);
			23346: out = 24'(6472);
			23347: out = 24'(-2756);
			23348: out = 24'(4116);
			23349: out = 24'(4340);
			23350: out = 24'(-13128);
			23351: out = 24'(-24104);
			23352: out = 24'(-9628);
			23353: out = 24'(18448);
			23354: out = 24'(24540);
			23355: out = 24'(16684);
			23356: out = 24'(9512);
			23357: out = 24'(14680);
			23358: out = 24'(336);
			23359: out = 24'(-24752);
			23360: out = 24'(-44240);
			23361: out = 24'(-12332);
			23362: out = 24'(3616);
			23363: out = 24'(2968);
			23364: out = 24'(18628);
			23365: out = 24'(41056);
			23366: out = 24'(29736);
			23367: out = 24'(-1340);
			23368: out = 24'(-15644);
			23369: out = 24'(-20460);
			23370: out = 24'(-22648);
			23371: out = 24'(-17620);
			23372: out = 24'(4588);
			23373: out = 24'(20744);
			23374: out = 24'(20580);
			23375: out = 24'(15092);
			23376: out = 24'(16640);
			23377: out = 24'(12272);
			23378: out = 24'(3316);
			23379: out = 24'(-4408);
			23380: out = 24'(-6392);
			23381: out = 24'(-12980);
			23382: out = 24'(-4168);
			23383: out = 24'(3048);
			23384: out = 24'(8604);
			23385: out = 24'(16388);
			23386: out = 24'(9436);
			23387: out = 24'(11224);
			23388: out = 24'(11024);
			23389: out = 24'(7984);
			23390: out = 24'(-5716);
			23391: out = 24'(-5400);
			23392: out = 24'(-12016);
			23393: out = 24'(-21108);
			23394: out = 24'(-21984);
			23395: out = 24'(20212);
			23396: out = 24'(36400);
			23397: out = 24'(10132);
			23398: out = 24'(-22608);
			23399: out = 24'(-33812);
			23400: out = 24'(-27304);
			23401: out = 24'(-14088);
			23402: out = 24'(7648);
			23403: out = 24'(9276);
			23404: out = 24'(10192);
			23405: out = 24'(11108);
			23406: out = 24'(15572);
			23407: out = 24'(-64);
			23408: out = 24'(-8880);
			23409: out = 24'(-16496);
			23410: out = 24'(-19428);
			23411: out = 24'(-9316);
			23412: out = 24'(2040);
			23413: out = 24'(12224);
			23414: out = 24'(16472);
			23415: out = 24'(16452);
			23416: out = 24'(2312);
			23417: out = 24'(1548);
			23418: out = 24'(12748);
			23419: out = 24'(13424);
			23420: out = 24'(12);
			23421: out = 24'(-15044);
			23422: out = 24'(-12500);
			23423: out = 24'(-972);
			23424: out = 24'(9048);
			23425: out = 24'(2608);
			23426: out = 24'(-808);
			23427: out = 24'(1716);
			23428: out = 24'(6256);
			23429: out = 24'(-11696);
			23430: out = 24'(-24984);
			23431: out = 24'(-21628);
			23432: out = 24'(-5340);
			23433: out = 24'(-2484);
			23434: out = 24'(7024);
			23435: out = 24'(19160);
			23436: out = 24'(21464);
			23437: out = 24'(4476);
			23438: out = 24'(-11860);
			23439: out = 24'(-25424);
			23440: out = 24'(-30140);
			23441: out = 24'(-17116);
			23442: out = 24'(4548);
			23443: out = 24'(7760);
			23444: out = 24'(-712);
			23445: out = 24'(-12824);
			23446: out = 24'(18172);
			23447: out = 24'(27140);
			23448: out = 24'(-1272);
			23449: out = 24'(-28664);
			23450: out = 24'(-6876);
			23451: out = 24'(13256);
			23452: out = 24'(-2664);
			23453: out = 24'(-33008);
			23454: out = 24'(-14012);
			23455: out = 24'(7184);
			23456: out = 24'(3684);
			23457: out = 24'(-1356);
			23458: out = 24'(-1956);
			23459: out = 24'(12552);
			23460: out = 24'(13344);
			23461: out = 24'(-256);
			23462: out = 24'(-472);
			23463: out = 24'(6800);
			23464: out = 24'(10760);
			23465: out = 24'(6320);
			23466: out = 24'(10748);
			23467: out = 24'(2500);
			23468: out = 24'(-2252);
			23469: out = 24'(184);
			23470: out = 24'(1800);
			23471: out = 24'(6392);
			23472: out = 24'(6152);
			23473: out = 24'(7772);
			23474: out = 24'(8964);
			23475: out = 24'(10368);
			23476: out = 24'(4588);
			23477: out = 24'(1704);
			23478: out = 24'(404);
			23479: out = 24'(-100);
			23480: out = 24'(-10696);
			23481: out = 24'(-4076);
			23482: out = 24'(16880);
			23483: out = 24'(9308);
			23484: out = 24'(852);
			23485: out = 24'(4128);
			23486: out = 24'(14008);
			23487: out = 24'(-1936);
			23488: out = 24'(-15496);
			23489: out = 24'(-20632);
			23490: out = 24'(-15688);
			23491: out = 24'(-20240);
			23492: out = 24'(-13804);
			23493: out = 24'(1896);
			23494: out = 24'(22908);
			23495: out = 24'(26272);
			23496: out = 24'(-3484);
			23497: out = 24'(-27568);
			23498: out = 24'(-21476);
			23499: out = 24'(3948);
			23500: out = 24'(-3852);
			23501: out = 24'(-4548);
			23502: out = 24'(-636);
			23503: out = 24'(10788);
			23504: out = 24'(28252);
			23505: out = 24'(15656);
			23506: out = 24'(-9376);
			23507: out = 24'(-21052);
			23508: out = 24'(-1752);
			23509: out = 24'(968);
			23510: out = 24'(-9708);
			23511: out = 24'(-17296);
			23512: out = 24'(1284);
			23513: out = 24'(12552);
			23514: out = 24'(10208);
			23515: out = 24'(-8960);
			23516: out = 24'(-17252);
			23517: out = 24'(-25416);
			23518: out = 24'(-608);
			23519: out = 24'(9496);
			23520: out = 24'(-2264);
			23521: out = 24'(-17284);
			23522: out = 24'(368);
			23523: out = 24'(13972);
			23524: out = 24'(6892);
			23525: out = 24'(-2820);
			23526: out = 24'(756);
			23527: out = 24'(-4412);
			23528: out = 24'(-25552);
			23529: out = 24'(-34272);
			23530: out = 24'(-9784);
			23531: out = 24'(25440);
			23532: out = 24'(34616);
			23533: out = 24'(21656);
			23534: out = 24'(5200);
			23535: out = 24'(2628);
			23536: out = 24'(-1232);
			23537: out = 24'(-13572);
			23538: out = 24'(-31992);
			23539: out = 24'(-14296);
			23540: out = 24'(15808);
			23541: out = 24'(26836);
			23542: out = 24'(17724);
			23543: out = 24'(14476);
			23544: out = 24'(20688);
			23545: out = 24'(20104);
			23546: out = 24'(-1748);
			23547: out = 24'(-9692);
			23548: out = 24'(-19252);
			23549: out = 24'(-22628);
			23550: out = 24'(-9864);
			23551: out = 24'(5216);
			23552: out = 24'(15804);
			23553: out = 24'(11940);
			23554: out = 24'(6952);
			23555: out = 24'(10232);
			23556: out = 24'(19800);
			23557: out = 24'(13216);
			23558: out = 24'(-6304);
			23559: out = 24'(-30432);
			23560: out = 24'(-19924);
			23561: out = 24'(-5592);
			23562: out = 24'(-128);
			23563: out = 24'(-1460);
			23564: out = 24'(12408);
			23565: out = 24'(13764);
			23566: out = 24'(5424);
			23567: out = 24'(-5808);
			23568: out = 24'(-1536);
			23569: out = 24'(-2784);
			23570: out = 24'(6484);
			23571: out = 24'(20384);
			23572: out = 24'(17868);
			23573: out = 24'(-13500);
			23574: out = 24'(-22572);
			23575: out = 24'(6632);
			23576: out = 24'(9552);
			23577: out = 24'(-7332);
			23578: out = 24'(-29864);
			23579: out = 24'(-25916);
			23580: out = 24'(-6648);
			23581: out = 24'(8056);
			23582: out = 24'(11116);
			23583: out = 24'(12992);
			23584: out = 24'(7752);
			23585: out = 24'(-896);
			23586: out = 24'(-15276);
			23587: out = 24'(-16792);
			23588: out = 24'(-3168);
			23589: out = 24'(7888);
			23590: out = 24'(8452);
			23591: out = 24'(4136);
			23592: out = 24'(2704);
			23593: out = 24'(8500);
			23594: out = 24'(5024);
			23595: out = 24'(-4748);
			23596: out = 24'(-13436);
			23597: out = 24'(-11872);
			23598: out = 24'(-12340);
			23599: out = 24'(-11460);
			23600: out = 24'(-12412);
			23601: out = 24'(-13296);
			23602: out = 24'(18568);
			23603: out = 24'(38468);
			23604: out = 24'(27208);
			23605: out = 24'(-3908);
			23606: out = 24'(-27844);
			23607: out = 24'(-27964);
			23608: out = 24'(-22696);
			23609: out = 24'(-24832);
			23610: out = 24'(-1712);
			23611: out = 24'(6444);
			23612: out = 24'(4356);
			23613: out = 24'(-4036);
			23614: out = 24'(1760);
			23615: out = 24'(11752);
			23616: out = 24'(19820);
			23617: out = 24'(10208);
			23618: out = 24'(-10084);
			23619: out = 24'(-22076);
			23620: out = 24'(-11400);
			23621: out = 24'(6304);
			23622: out = 24'(12872);
			23623: out = 24'(3072);
			23624: out = 24'(-1036);
			23625: out = 24'(632);
			23626: out = 24'(16);
			23627: out = 24'(832);
			23628: out = 24'(-476);
			23629: out = 24'(2216);
			23630: out = 24'(8892);
			23631: out = 24'(15568);
			23632: out = 24'(26544);
			23633: out = 24'(29292);
			23634: out = 24'(17960);
			23635: out = 24'(-1552);
			23636: out = 24'(-11552);
			23637: out = 24'(-11468);
			23638: out = 24'(-8168);
			23639: out = 24'(-4532);
			23640: out = 24'(3540);
			23641: out = 24'(15384);
			23642: out = 24'(20920);
			23643: out = 24'(12008);
			23644: out = 24'(-5916);
			23645: out = 24'(-13844);
			23646: out = 24'(-8284);
			23647: out = 24'(-840);
			23648: out = 24'(-880);
			23649: out = 24'(2360);
			23650: out = 24'(13892);
			23651: out = 24'(22444);
			23652: out = 24'(7348);
			23653: out = 24'(1260);
			23654: out = 24'(-6828);
			23655: out = 24'(-10412);
			23656: out = 24'(-13960);
			23657: out = 24'(-18160);
			23658: out = 24'(-22212);
			23659: out = 24'(-12088);
			23660: out = 24'(7172);
			23661: out = 24'(15228);
			23662: out = 24'(3740);
			23663: out = 24'(-9524);
			23664: out = 24'(-12372);
			23665: out = 24'(-18936);
			23666: out = 24'(-15412);
			23667: out = 24'(144);
			23668: out = 24'(17544);
			23669: out = 24'(5656);
			23670: out = 24'(-5656);
			23671: out = 24'(-11836);
			23672: out = 24'(1172);
			23673: out = 24'(3768);
			23674: out = 24'(10860);
			23675: out = 24'(-19968);
			23676: out = 24'(-45352);
			23677: out = 24'(-29716);
			23678: out = 24'(9420);
			23679: out = 24'(21136);
			23680: out = 24'(13232);
			23681: out = 24'(12008);
			23682: out = 24'(15264);
			23683: out = 24'(7296);
			23684: out = 24'(-10092);
			23685: out = 24'(-17808);
			23686: out = 24'(-12060);
			23687: out = 24'(9324);
			23688: out = 24'(19824);
			23689: out = 24'(8156);
			23690: out = 24'(-28736);
			23691: out = 24'(-9008);
			23692: out = 24'(12176);
			23693: out = 24'(12492);
			23694: out = 24'(-3908);
			23695: out = 24'(-1628);
			23696: out = 24'(4432);
			23697: out = 24'(8004);
			23698: out = 24'(11204);
			23699: out = 24'(14560);
			23700: out = 24'(17652);
			23701: out = 24'(6844);
			23702: out = 24'(-10844);
			23703: out = 24'(-19088);
			23704: out = 24'(-7112);
			23705: out = 24'(-312);
			23706: out = 24'(-7696);
			23707: out = 24'(-17796);
			23708: out = 24'(-5636);
			23709: out = 24'(9684);
			23710: out = 24'(16780);
			23711: out = 24'(12596);
			23712: out = 24'(28004);
			23713: out = 24'(16664);
			23714: out = 24'(-10360);
			23715: out = 24'(-29252);
			23716: out = 24'(3540);
			23717: out = 24'(12668);
			23718: out = 24'(1260);
			23719: out = 24'(-12968);
			23720: out = 24'(-11952);
			23721: out = 24'(5516);
			23722: out = 24'(25076);
			23723: out = 24'(25052);
			23724: out = 24'(7692);
			23725: out = 24'(-2780);
			23726: out = 24'(8612);
			23727: out = 24'(13680);
			23728: out = 24'(-6276);
			23729: out = 24'(-35800);
			23730: out = 24'(-17512);
			23731: out = 24'(25340);
			23732: out = 24'(28876);
			23733: out = 24'(280);
			23734: out = 24'(-28556);
			23735: out = 24'(-22616);
			23736: out = 24'(-1148);
			23737: out = 24'(-14076);
			23738: out = 24'(-22636);
			23739: out = 24'(-15964);
			23740: out = 24'(1824);
			23741: out = 24'(1300);
			23742: out = 24'(8984);
			23743: out = 24'(8552);
			23744: out = 24'(5224);
			23745: out = 24'(-1080);
			23746: out = 24'(-8128);
			23747: out = 24'(-17636);
			23748: out = 24'(-14232);
			23749: out = 24'(296);
			23750: out = 24'(7384);
			23751: out = 24'(-8964);
			23752: out = 24'(-28020);
			23753: out = 24'(-26932);
			23754: out = 24'(-6924);
			23755: out = 24'(9492);
			23756: out = 24'(16780);
			23757: out = 24'(14636);
			23758: out = 24'(-1708);
			23759: out = 24'(-10032);
			23760: out = 24'(-5908);
			23761: out = 24'(1776);
			23762: out = 24'(1032);
			23763: out = 24'(-20);
			23764: out = 24'(2644);
			23765: out = 24'(-896);
			23766: out = 24'(-17880);
			23767: out = 24'(-19264);
			23768: out = 24'(192);
			23769: out = 24'(16816);
			23770: out = 24'(5036);
			23771: out = 24'(24);
			23772: out = 24'(2644);
			23773: out = 24'(20016);
			23774: out = 24'(20804);
			23775: out = 24'(1000);
			23776: out = 24'(-33556);
			23777: out = 24'(-29128);
			23778: out = 24'(10548);
			23779: out = 24'(22532);
			23780: out = 24'(17916);
			23781: out = 24'(392);
			23782: out = 24'(108);
			23783: out = 24'(9016);
			23784: out = 24'(17872);
			23785: out = 24'(-724);
			23786: out = 24'(-17104);
			23787: out = 24'(-8676);
			23788: out = 24'(12676);
			23789: out = 24'(13076);
			23790: out = 24'(1364);
			23791: out = 24'(-3384);
			23792: out = 24'(-884);
			23793: out = 24'(10484);
			23794: out = 24'(21072);
			23795: out = 24'(22060);
			23796: out = 24'(9804);
			23797: out = 24'(-6928);
			23798: out = 24'(-17156);
			23799: out = 24'(-20248);
			23800: out = 24'(-18336);
			23801: out = 24'(-6500);
			23802: out = 24'(17208);
			23803: out = 24'(30828);
			23804: out = 24'(18960);
			23805: out = 24'(-532);
			23806: out = 24'(-5852);
			23807: out = 24'(5412);
			23808: out = 24'(13504);
			23809: out = 24'(-3264);
			23810: out = 24'(-1140);
			23811: out = 24'(14528);
			23812: out = 24'(18352);
			23813: out = 24'(-18304);
			23814: out = 24'(-36452);
			23815: out = 24'(-34232);
			23816: out = 24'(-13044);
			23817: out = 24'(-1580);
			23818: out = 24'(28076);
			23819: out = 24'(25216);
			23820: out = 24'(4312);
			23821: out = 24'(-11064);
			23822: out = 24'(2428);
			23823: out = 24'(4628);
			23824: out = 24'(-7532);
			23825: out = 24'(-18400);
			23826: out = 24'(-2800);
			23827: out = 24'(-1072);
			23828: out = 24'(-8544);
			23829: out = 24'(-9680);
			23830: out = 24'(-1436);
			23831: out = 24'(8452);
			23832: out = 24'(4836);
			23833: out = 24'(-7064);
			23834: out = 24'(-10788);
			23835: out = 24'(-1404);
			23836: out = 24'(1888);
			23837: out = 24'(-9420);
			23838: out = 24'(-16516);
			23839: out = 24'(-9212);
			23840: out = 24'(16292);
			23841: out = 24'(27248);
			23842: out = 24'(13680);
			23843: out = 24'(-1676);
			23844: out = 24'(-9388);
			23845: out = 24'(-17740);
			23846: out = 24'(-31800);
			23847: out = 24'(-29488);
			23848: out = 24'(-10560);
			23849: out = 24'(14064);
			23850: out = 24'(21592);
			23851: out = 24'(11756);
			23852: out = 24'(1992);
			23853: out = 24'(5800);
			23854: out = 24'(15596);
			23855: out = 24'(14552);
			23856: out = 24'(-4568);
			23857: out = 24'(-19060);
			23858: out = 24'(-12960);
			23859: out = 24'(1120);
			23860: out = 24'(23588);
			23861: out = 24'(5668);
			23862: out = 24'(-22540);
			23863: out = 24'(-31064);
			23864: out = 24'(-2556);
			23865: out = 24'(2420);
			23866: out = 24'(5328);
			23867: out = 24'(21208);
			23868: out = 24'(22776);
			23869: out = 24'(27568);
			23870: out = 24'(10892);
			23871: out = 24'(-11024);
			23872: out = 24'(-30416);
			23873: out = 24'(-7572);
			23874: out = 24'(2284);
			23875: out = 24'(-1024);
			23876: out = 24'(212);
			23877: out = 24'(-1116);
			23878: out = 24'(3644);
			23879: out = 24'(11944);
			23880: out = 24'(23492);
			23881: out = 24'(28992);
			23882: out = 24'(13876);
			23883: out = 24'(-13836);
			23884: out = 24'(-29600);
			23885: out = 24'(-3212);
			23886: out = 24'(220);
			23887: out = 24'(920);
			23888: out = 24'(10164);
			23889: out = 24'(19904);
			23890: out = 24'(24948);
			23891: out = 24'(10616);
			23892: out = 24'(-7340);
			23893: out = 24'(-12456);
			23894: out = 24'(-7808);
			23895: out = 24'(-3156);
			23896: out = 24'(-2024);
			23897: out = 24'(-120);
			23898: out = 24'(12744);
			23899: out = 24'(20956);
			23900: out = 24'(18408);
			23901: out = 24'(-1548);
			23902: out = 24'(-20648);
			23903: out = 24'(-36496);
			23904: out = 24'(-21460);
			23905: out = 24'(1684);
			23906: out = 24'(-720);
			23907: out = 24'(5744);
			23908: out = 24'(15024);
			23909: out = 24'(3456);
			23910: out = 24'(-42540);
			23911: out = 24'(-21556);
			23912: out = 24'(15812);
			23913: out = 24'(21276);
			23914: out = 24'(-18392);
			23915: out = 24'(-18936);
			23916: out = 24'(-236);
			23917: out = 24'(13420);
			23918: out = 24'(-3740);
			23919: out = 24'(1824);
			23920: out = 24'(-12012);
			23921: out = 24'(-14000);
			23922: out = 24'(-9916);
			23923: out = 24'(-3768);
			23924: out = 24'(-292);
			23925: out = 24'(1120);
			23926: out = 24'(488);
			23927: out = 24'(132);
			23928: out = 24'(-2980);
			23929: out = 24'(-1928);
			23930: out = 24'(3208);
			23931: out = 24'(5736);
			23932: out = 24'(-12912);
			23933: out = 24'(-24020);
			23934: out = 24'(-11856);
			23935: out = 24'(8008);
			23936: out = 24'(3004);
			23937: out = 24'(-9756);
			23938: out = 24'(-9400);
			23939: out = 24'(3244);
			23940: out = 24'(7960);
			23941: out = 24'(-2520);
			23942: out = 24'(-1908);
			23943: out = 24'(10132);
			23944: out = 24'(6824);
			23945: out = 24'(2800);
			23946: out = 24'(-776);
			23947: out = 24'(900);
			23948: out = 24'(1044);
			23949: out = 24'(488);
			23950: out = 24'(9396);
			23951: out = 24'(20420);
			23952: out = 24'(20436);
			23953: out = 24'(-376);
			23954: out = 24'(-12344);
			23955: out = 24'(-14604);
			23956: out = 24'(-9332);
			23957: out = 24'(-5216);
			23958: out = 24'(11420);
			23959: out = 24'(14604);
			23960: out = 24'(4616);
			23961: out = 24'(1212);
			23962: out = 24'(6656);
			23963: out = 24'(13828);
			23964: out = 24'(15048);
			23965: out = 24'(8480);
			23966: out = 24'(2624);
			23967: out = 24'(-13284);
			23968: out = 24'(-23424);
			23969: out = 24'(-13324);
			23970: out = 24'(-2352);
			23971: out = 24'(3184);
			23972: out = 24'(4376);
			23973: out = 24'(8604);
			23974: out = 24'(23188);
			23975: out = 24'(15768);
			23976: out = 24'(5812);
			23977: out = 24'(7856);
			23978: out = 24'(13608);
			23979: out = 24'(9624);
			23980: out = 24'(-3720);
			23981: out = 24'(-14784);
			23982: out = 24'(-19740);
			23983: out = 24'(-3428);
			23984: out = 24'(4352);
			23985: out = 24'(620);
			23986: out = 24'(716);
			23987: out = 24'(11240);
			23988: out = 24'(17996);
			23989: out = 24'(3868);
			23990: out = 24'(-21740);
			23991: out = 24'(-24924);
			23992: out = 24'(-8272);
			23993: out = 24'(3560);
			23994: out = 24'(-5772);
			23995: out = 24'(-24488);
			23996: out = 24'(-7204);
			23997: out = 24'(19000);
			23998: out = 24'(11168);
			23999: out = 24'(-35852);
			24000: out = 24'(-37956);
			24001: out = 24'(-5032);
			24002: out = 24'(16792);
			24003: out = 24'(-880);
			24004: out = 24'(-9020);
			24005: out = 24'(-2072);
			24006: out = 24'(9432);
			24007: out = 24'(480);
			24008: out = 24'(-4556);
			24009: out = 24'(-5124);
			24010: out = 24'(8688);
			24011: out = 24'(13800);
			24012: out = 24'(-652);
			24013: out = 24'(-29320);
			24014: out = 24'(-32920);
			24015: out = 24'(-6092);
			24016: out = 24'(14768);
			24017: out = 24'(456);
			24018: out = 24'(-25348);
			24019: out = 24'(-26272);
			24020: out = 24'(4764);
			24021: out = 24'(16812);
			24022: out = 24'(15092);
			24023: out = 24'(11128);
			24024: out = 24'(11468);
			24025: out = 24'(17328);
			24026: out = 24'(-36);
			24027: out = 24'(-23228);
			24028: out = 24'(-24404);
			24029: out = 24'(12852);
			24030: out = 24'(11604);
			24031: out = 24'(-14208);
			24032: out = 24'(-23060);
			24033: out = 24'(15656);
			24034: out = 24'(32816);
			24035: out = 24'(27160);
			24036: out = 24'(13608);
			24037: out = 24'(7064);
			24038: out = 24'(7188);
			24039: out = 24'(2892);
			24040: out = 24'(-272);
			24041: out = 24'(-788);
			24042: out = 24'(-2660);
			24043: out = 24'(-6636);
			24044: out = 24'(4804);
			24045: out = 24'(21780);
			24046: out = 24'(11500);
			24047: out = 24'(-1724);
			24048: out = 24'(-16);
			24049: out = 24'(8764);
			24050: out = 24'(80);
			24051: out = 24'(-3504);
			24052: out = 24'(10600);
			24053: out = 24'(22816);
			24054: out = 24'(8344);
			24055: out = 24'(-12052);
			24056: out = 24'(-10496);
			24057: out = 24'(-92);
			24058: out = 24'(-5664);
			24059: out = 24'(-3528);
			24060: out = 24'(13884);
			24061: out = 24'(19552);
			24062: out = 24'(-6292);
			24063: out = 24'(-27340);
			24064: out = 24'(-27652);
			24065: out = 24'(-12388);
			24066: out = 24'(-2100);
			24067: out = 24'(18312);
			24068: out = 24'(21680);
			24069: out = 24'(12856);
			24070: out = 24'(-4128);
			24071: out = 24'(544);
			24072: out = 24'(-2812);
			24073: out = 24'(3424);
			24074: out = 24'(3284);
			24075: out = 24'(-5668);
			24076: out = 24'(-11696);
			24077: out = 24'(-13972);
			24078: out = 24'(-20220);
			24079: out = 24'(-30676);
			24080: out = 24'(-23768);
			24081: out = 24'(-4236);
			24082: out = 24'(14936);
			24083: out = 24'(13384);
			24084: out = 24'(-244);
			24085: out = 24'(-7076);
			24086: out = 24'(7100);
			24087: out = 24'(13536);
			24088: out = 24'(-5620);
			24089: out = 24'(-18196);
			24090: out = 24'(-5692);
			24091: out = 24'(8716);
			24092: out = 24'(2820);
			24093: out = 24'(-18092);
			24094: out = 24'(-11832);
			24095: out = 24'(3604);
			24096: out = 24'(996);
			24097: out = 24'(15304);
			24098: out = 24'(22444);
			24099: out = 24'(12656);
			24100: out = 24'(-14096);
			24101: out = 24'(-13720);
			24102: out = 24'(-816);
			24103: out = 24'(10228);
			24104: out = 24'(6432);
			24105: out = 24'(17836);
			24106: out = 24'(3236);
			24107: out = 24'(2044);
			24108: out = 24'(7652);
			24109: out = 24'(4912);
			24110: out = 24'(-12036);
			24111: out = 24'(-32640);
			24112: out = 24'(-31576);
			24113: out = 24'(-836);
			24114: out = 24'(13964);
			24115: out = 24'(18484);
			24116: out = 24'(14248);
			24117: out = 24'(10144);
			24118: out = 24'(10112);
			24119: out = 24'(3552);
			24120: out = 24'(-1344);
			24121: out = 24'(-380);
			24122: out = 24'(-1408);
			24123: out = 24'(288);
			24124: out = 24'(-3020);
			24125: out = 24'(-9392);
			24126: out = 24'(-10436);
			24127: out = 24'(-12168);
			24128: out = 24'(-2120);
			24129: out = 24'(12832);
			24130: out = 24'(24560);
			24131: out = 24'(9572);
			24132: out = 24'(6856);
			24133: out = 24'(12248);
			24134: out = 24'(14108);
			24135: out = 24'(-2756);
			24136: out = 24'(-3828);
			24137: out = 24'(2768);
			24138: out = 24'(4000);
			24139: out = 24'(-10884);
			24140: out = 24'(-20356);
			24141: out = 24'(-24600);
			24142: out = 24'(-18756);
			24143: out = 24'(-44);
			24144: out = 24'(19708);
			24145: out = 24'(27184);
			24146: out = 24'(19240);
			24147: out = 24'(1444);
			24148: out = 24'(-3604);
			24149: out = 24'(-9180);
			24150: out = 24'(-13512);
			24151: out = 24'(-13400);
			24152: out = 24'(17484);
			24153: out = 24'(23844);
			24154: out = 24'(13552);
			24155: out = 24'(-4108);
			24156: out = 24'(-12812);
			24157: out = 24'(-27276);
			24158: out = 24'(-19068);
			24159: out = 24'(9056);
			24160: out = 24'(21552);
			24161: out = 24'(19180);
			24162: out = 24'(7456);
			24163: out = 24'(104);
			24164: out = 24'(-5232);
			24165: out = 24'(6108);
			24166: out = 24'(9708);
			24167: out = 24'(5160);
			24168: out = 24'(-6404);
			24169: out = 24'(-10804);
			24170: out = 24'(-13144);
			24171: out = 24'(-8256);
			24172: out = 24'(-1072);
			24173: out = 24'(-452);
			24174: out = 24'(-3448);
			24175: out = 24'(-5060);
			24176: out = 24'(-4328);
			24177: out = 24'(-416);
			24178: out = 24'(-5908);
			24179: out = 24'(-7560);
			24180: out = 24'(-308);
			24181: out = 24'(15584);
			24182: out = 24'(15148);
			24183: out = 24'(12884);
			24184: out = 24'(3904);
			24185: out = 24'(-8380);
			24186: out = 24'(-15240);
			24187: out = 24'(-12348);
			24188: out = 24'(-15640);
			24189: out = 24'(-23916);
			24190: out = 24'(-3356);
			24191: out = 24'(17840);
			24192: out = 24'(17732);
			24193: out = 24'(-5528);
			24194: out = 24'(-12424);
			24195: out = 24'(-6452);
			24196: out = 24'(7284);
			24197: out = 24'(5144);
			24198: out = 24'(-12984);
			24199: out = 24'(-13784);
			24200: out = 24'(520);
			24201: out = 24'(10672);
			24202: out = 24'(6308);
			24203: out = 24'(6480);
			24204: out = 24'(6736);
			24205: out = 24'(3624);
			24206: out = 24'(-5956);
			24207: out = 24'(-19976);
			24208: out = 24'(-17016);
			24209: out = 24'(-3928);
			24210: out = 24'(4956);
			24211: out = 24'(16116);
			24212: out = 24'(4716);
			24213: out = 24'(1076);
			24214: out = 24'(16644);
			24215: out = 24'(38920);
			24216: out = 24'(13132);
			24217: out = 24'(-25208);
			24218: out = 24'(-37208);
			24219: out = 24'(-3948);
			24220: out = 24'(-824);
			24221: out = 24'(-3392);
			24222: out = 24'(848);
			24223: out = 24'(16524);
			24224: out = 24'(18432);
			24225: out = 24'(1340);
			24226: out = 24'(-15148);
			24227: out = 24'(-1596);
			24228: out = 24'(23592);
			24229: out = 24'(33300);
			24230: out = 24'(11848);
			24231: out = 24'(-10128);
			24232: out = 24'(-6416);
			24233: out = 24'(8112);
			24234: out = 24'(4992);
			24235: out = 24'(-10436);
			24236: out = 24'(-22968);
			24237: out = 24'(-3600);
			24238: out = 24'(-4);
			24239: out = 24'(-5988);
			24240: out = 24'(820);
			24241: out = 24'(23788);
			24242: out = 24'(23116);
			24243: out = 24'(5344);
			24244: out = 24'(-5436);
			24245: out = 24'(-6828);
			24246: out = 24'(-3016);
			24247: out = 24'(-2060);
			24248: out = 24'(-2152);
			24249: out = 24'(-12420);
			24250: out = 24'(-7564);
			24251: out = 24'(-3164);
			24252: out = 24'(1760);
			24253: out = 24'(14048);
			24254: out = 24'(3052);
			24255: out = 24'(-12572);
			24256: out = 24'(-27764);
			24257: out = 24'(-32352);
			24258: out = 24'(-16744);
			24259: out = 24'(6236);
			24260: out = 24'(17576);
			24261: out = 24'(13900);
			24262: out = 24'(1464);
			24263: out = 24'(-5032);
			24264: out = 24'(-13648);
			24265: out = 24'(-21236);
			24266: out = 24'(-4936);
			24267: out = 24'(10624);
			24268: out = 24'(12436);
			24269: out = 24'(-7920);
			24270: out = 24'(-29668);
			24271: out = 24'(-11744);
			24272: out = 24'(24416);
			24273: out = 24'(31808);
			24274: out = 24'(6040);
			24275: out = 24'(-9532);
			24276: out = 24'(2848);
			24277: out = 24'(17316);
			24278: out = 24'(5464);
			24279: out = 24'(-14076);
			24280: out = 24'(-17804);
			24281: out = 24'(-2952);
			24282: out = 24'(6040);
			24283: out = 24'(7404);
			24284: out = 24'(-1684);
			24285: out = 24'(-3612);
			24286: out = 24'(336);
			24287: out = 24'(6332);
			24288: out = 24'(1136);
			24289: out = 24'(1864);
			24290: out = 24'(7232);
			24291: out = 24'(4852);
			24292: out = 24'(1172);
			24293: out = 24'(-9880);
			24294: out = 24'(-13868);
			24295: out = 24'(-3288);
			24296: out = 24'(-2032);
			24297: out = 24'(1472);
			24298: out = 24'(3352);
			24299: out = 24'(8372);
			24300: out = 24'(19160);
			24301: out = 24'(15324);
			24302: out = 24'(-2660);
			24303: out = 24'(-12836);
			24304: out = 24'(7532);
			24305: out = 24'(17488);
			24306: out = 24'(3908);
			24307: out = 24'(-20320);
			24308: out = 24'(-16772);
			24309: out = 24'(-15408);
			24310: out = 24'(-576);
			24311: out = 24'(6820);
			24312: out = 24'(6636);
			24313: out = 24'(7596);
			24314: out = 24'(18280);
			24315: out = 24'(17688);
			24316: out = 24'(-5964);
			24317: out = 24'(-22264);
			24318: out = 24'(-30068);
			24319: out = 24'(-15592);
			24320: out = 24'(940);
			24321: out = 24'(10108);
			24322: out = 24'(1748);
			24323: out = 24'(2696);
			24324: out = 24'(5244);
			24325: out = 24'(180);
			24326: out = 24'(-15444);
			24327: out = 24'(-12712);
			24328: out = 24'(-1464);
			24329: out = 24'(200);
			24330: out = 24'(-552);
			24331: out = 24'(9540);
			24332: out = 24'(12920);
			24333: out = 24'(-2992);
			24334: out = 24'(-6444);
			24335: out = 24'(-2388);
			24336: out = 24'(5472);
			24337: out = 24'(6800);
			24338: out = 24'(15172);
			24339: out = 24'(7028);
			24340: out = 24'(-6440);
			24341: out = 24'(-14604);
			24342: out = 24'(-4356);
			24343: out = 24'(1680);
			24344: out = 24'(2008);
			24345: out = 24'(-548);
			24346: out = 24'(-636);
			24347: out = 24'(-8264);
			24348: out = 24'(-18604);
			24349: out = 24'(-16780);
			24350: out = 24'(3176);
			24351: out = 24'(19036);
			24352: out = 24'(14548);
			24353: out = 24'(-1520);
			24354: out = 24'(-12276);
			24355: out = 24'(-21836);
			24356: out = 24'(-14984);
			24357: out = 24'(-5116);
			24358: out = 24'(2152);
			24359: out = 24'(7364);
			24360: out = 24'(19772);
			24361: out = 24'(27072);
			24362: out = 24'(16580);
			24363: out = 24'(-7296);
			24364: out = 24'(-26160);
			24365: out = 24'(-24776);
			24366: out = 24'(-12208);
			24367: out = 24'(1620);
			24368: out = 24'(8168);
			24369: out = 24'(20476);
			24370: out = 24'(20752);
			24371: out = 24'(6804);
			24372: out = 24'(-15880);
			24373: out = 24'(-8028);
			24374: out = 24'(2352);
			24375: out = 24'(-1972);
			24376: out = 24'(-9572);
			24377: out = 24'(-3940);
			24378: out = 24'(1568);
			24379: out = 24'(-20);
			24380: out = 24'(1164);
			24381: out = 24'(12200);
			24382: out = 24'(17520);
			24383: out = 24'(12236);
			24384: out = 24'(2736);
			24385: out = 24'(3004);
			24386: out = 24'(-5336);
			24387: out = 24'(-11024);
			24388: out = 24'(-1852);
			24389: out = 24'(7340);
			24390: out = 24'(9176);
			24391: out = 24'(1632);
			24392: out = 24'(-3972);
			24393: out = 24'(-764);
			24394: out = 24'(-2296);
			24395: out = 24'(-5580);
			24396: out = 24'(-616);
			24397: out = 24'(14540);
			24398: out = 24'(11780);
			24399: out = 24'(5676);
			24400: out = 24'(10928);
			24401: out = 24'(26692);
			24402: out = 24'(-2640);
			24403: out = 24'(-32364);
			24404: out = 24'(-34944);
			24405: out = 24'(-2184);
			24406: out = 24'(-8076);
			24407: out = 24'(-5336);
			24408: out = 24'(-652);
			24409: out = 24'(8152);
			24410: out = 24'(11476);
			24411: out = 24'(5340);
			24412: out = 24'(-4240);
			24413: out = 24'(-1364);
			24414: out = 24'(3992);
			24415: out = 24'(1824);
			24416: out = 24'(-21188);
			24417: out = 24'(-34864);
			24418: out = 24'(-13528);
			24419: out = 24'(13576);
			24420: out = 24'(12388);
			24421: out = 24'(-3528);
			24422: out = 24'(-588);
			24423: out = 24'(16840);
			24424: out = 24'(18696);
			24425: out = 24'(-2368);
			24426: out = 24'(-20328);
			24427: out = 24'(-7152);
			24428: out = 24'(7412);
			24429: out = 24'(5412);
			24430: out = 24'(-4136);
			24431: out = 24'(136);
			24432: out = 24'(16696);
			24433: out = 24'(23696);
			24434: out = 24'(6740);
			24435: out = 24'(-19996);
			24436: out = 24'(-22576);
			24437: out = 24'(-4704);
			24438: out = 24'(8920);
			24439: out = 24'(13120);
			24440: out = 24'(6176);
			24441: out = 24'(13716);
			24442: out = 24'(13896);
			24443: out = 24'(-2628);
			24444: out = 24'(-20420);
			24445: out = 24'(-5396);
			24446: out = 24'(15928);
			24447: out = 24'(10144);
			24448: out = 24'(-7808);
			24449: out = 24'(-11136);
			24450: out = 24'(9020);
			24451: out = 24'(22492);
			24452: out = 24'(14980);
			24453: out = 24'(-8720);
			24454: out = 24'(-17088);
			24455: out = 24'(-9372);
			24456: out = 24'(-5936);
			24457: out = 24'(-4224);
			24458: out = 24'(-3852);
			24459: out = 24'(4308);
			24460: out = 24'(13936);
			24461: out = 24'(1992);
			24462: out = 24'(-13016);
			24463: out = 24'(-18992);
			24464: out = 24'(-8764);
			24465: out = 24'(6712);
			24466: out = 24'(4176);
			24467: out = 24'(-5688);
			24468: out = 24'(-412);
			24469: out = 24'(12408);
			24470: out = 24'(17888);
			24471: out = 24'(1180);
			24472: out = 24'(-13240);
			24473: out = 24'(-12712);
			24474: out = 24'(-1140);
			24475: out = 24'(-10700);
			24476: out = 24'(-13704);
			24477: out = 24'(10888);
			24478: out = 24'(15012);
			24479: out = 24'(5344);
			24480: out = 24'(1784);
			24481: out = 24'(16320);
			24482: out = 24'(14520);
			24483: out = 24'(-8636);
			24484: out = 24'(-28456);
			24485: out = 24'(-17520);
			24486: out = 24'(-3424);
			24487: out = 24'(3928);
			24488: out = 24'(1720);
			24489: out = 24'(12568);
			24490: out = 24'(28796);
			24491: out = 24'(17212);
			24492: out = 24'(-19236);
			24493: out = 24'(-44548);
			24494: out = 24'(-26268);
			24495: out = 24'(6928);
			24496: out = 24'(20592);
			24497: out = 24'(5360);
			24498: out = 24'(-10400);
			24499: out = 24'(-7036);
			24500: out = 24'(6456);
			24501: out = 24'(5780);
			24502: out = 24'(-912);
			24503: out = 24'(-1656);
			24504: out = 24'(18136);
			24505: out = 24'(12724);
			24506: out = 24'(-14860);
			24507: out = 24'(-20232);
			24508: out = 24'(-648);
			24509: out = 24'(15596);
			24510: out = 24'(5768);
			24511: out = 24'(-2356);
			24512: out = 24'(-4512);
			24513: out = 24'(14096);
			24514: out = 24'(15268);
			24515: out = 24'(-1476);
			24516: out = 24'(-2760);
			24517: out = 24'(9604);
			24518: out = 24'(9212);
			24519: out = 24'(-8984);
			24520: out = 24'(-21888);
			24521: out = 24'(-8952);
			24522: out = 24'(2136);
			24523: out = 24'(-2296);
			24524: out = 24'(488);
			24525: out = 24'(3244);
			24526: out = 24'(8360);
			24527: out = 24'(9256);
			24528: out = 24'(14776);
			24529: out = 24'(-2136);
			24530: out = 24'(-5352);
			24531: out = 24'(1772);
			24532: out = 24'(7532);
			24533: out = 24'(64);
			24534: out = 24'(-11644);
			24535: out = 24'(-13972);
			24536: out = 24'(-1604);
			24537: out = 24'(18160);
			24538: out = 24'(13960);
			24539: out = 24'(2256);
			24540: out = 24'(-364);
			24541: out = 24'(3728);
			24542: out = 24'(1520);
			24543: out = 24'(-12212);
			24544: out = 24'(-25496);
			24545: out = 24'(-21752);
			24546: out = 24'(-5952);
			24547: out = 24'(7216);
			24548: out = 24'(6708);
			24549: out = 24'(-92);
			24550: out = 24'(-1072);
			24551: out = 24'(3788);
			24552: out = 24'(6264);
			24553: out = 24'(5524);
			24554: out = 24'(-1056);
			24555: out = 24'(-9312);
			24556: out = 24'(-20372);
			24557: out = 24'(-18160);
			24558: out = 24'(-3484);
			24559: out = 24'(16572);
			24560: out = 24'(6360);
			24561: out = 24'(-12364);
			24562: out = 24'(-3064);
			24563: out = 24'(16088);
			24564: out = 24'(20252);
			24565: out = 24'(13624);
			24566: out = 24'(14312);
			24567: out = 24'(-4280);
			24568: out = 24'(-16896);
			24569: out = 24'(-13780);
			24570: out = 24'(-256);
			24571: out = 24'(276);
			24572: out = 24'(-20328);
			24573: out = 24'(-22120);
			24574: out = 24'(7832);
			24575: out = 24'(7000);
			24576: out = 24'(9284);
			24577: out = 24'(4336);
			24578: out = 24'(7760);
			24579: out = 24'(4444);
			24580: out = 24'(10180);
			24581: out = 24'(-896);
			24582: out = 24'(-15564);
			24583: out = 24'(-22036);
			24584: out = 24'(-19568);
			24585: out = 24'(-8828);
			24586: out = 24'(8492);
			24587: out = 24'(21140);
			24588: out = 24'(17432);
			24589: out = 24'(5108);
			24590: out = 24'(-1200);
			24591: out = 24'(-1204);
			24592: out = 24'(-10084);
			24593: out = 24'(-17176);
			24594: out = 24'(-11948);
			24595: out = 24'(3356);
			24596: out = 24'(5572);
			24597: out = 24'(10064);
			24598: out = 24'(5236);
			24599: out = 24'(-1808);
			24600: out = 24'(-3364);
			24601: out = 24'(3576);
			24602: out = 24'(9560);
			24603: out = 24'(6116);
			24604: out = 24'(-1296);
			24605: out = 24'(-14096);
			24606: out = 24'(-7124);
			24607: out = 24'(1364);
			24608: out = 24'(3160);
			24609: out = 24'(8504);
			24610: out = 24'(19420);
			24611: out = 24'(21696);
			24612: out = 24'(11392);
			24613: out = 24'(-196);
			24614: out = 24'(-18584);
			24615: out = 24'(-31976);
			24616: out = 24'(-20308);
			24617: out = 24'(13708);
			24618: out = 24'(23392);
			24619: out = 24'(-1112);
			24620: out = 24'(-23604);
			24621: out = 24'(-5192);
			24622: out = 24'(6052);
			24623: out = 24'(5820);
			24624: out = 24'(-2700);
			24625: out = 24'(2196);
			24626: out = 24'(12488);
			24627: out = 24'(11740);
			24628: out = 24'(-4472);
			24629: out = 24'(-20224);
			24630: out = 24'(-22144);
			24631: out = 24'(-8136);
			24632: out = 24'(9112);
			24633: out = 24'(12988);
			24634: out = 24'(396);
			24635: out = 24'(-4880);
			24636: out = 24'(2212);
			24637: out = 24'(9664);
			24638: out = 24'(5336);
			24639: out = 24'(-236);
			24640: out = 24'(-1180);
			24641: out = 24'(-1688);
			24642: out = 24'(-5700);
			24643: out = 24'(-21260);
			24644: out = 24'(-10520);
			24645: out = 24'(2452);
			24646: out = 24'(-3312);
			24647: out = 24'(-19284);
			24648: out = 24'(-3804);
			24649: out = 24'(28012);
			24650: out = 24'(37104);
			24651: out = 24'(6976);
			24652: out = 24'(-15884);
			24653: out = 24'(-24748);
			24654: out = 24'(-22360);
			24655: out = 24'(-29928);
			24656: out = 24'(-22284);
			24657: out = 24'(-10912);
			24658: out = 24'(12564);
			24659: out = 24'(29052);
			24660: out = 24'(26100);
			24661: out = 24'(-3324);
			24662: out = 24'(-17856);
			24663: out = 24'(-4532);
			24664: out = 24'(2060);
			24665: out = 24'(-5408);
			24666: out = 24'(-7388);
			24667: out = 24'(6184);
			24668: out = 24'(5988);
			24669: out = 24'(580);
			24670: out = 24'(-4252);
			24671: out = 24'(2120);
			24672: out = 24'(-724);
			24673: out = 24'(7388);
			24674: out = 24'(2960);
			24675: out = 24'(2156);
			24676: out = 24'(6408);
			24677: out = 24'(8080);
			24678: out = 24'(-7512);
			24679: out = 24'(-20024);
			24680: out = 24'(-10712);
			24681: out = 24'(3684);
			24682: out = 24'(10068);
			24683: out = 24'(-2584);
			24684: out = 24'(-17576);
			24685: out = 24'(-3584);
			24686: out = 24'(6260);
			24687: out = 24'(17580);
			24688: out = 24'(24372);
			24689: out = 24'(14312);
			24690: out = 24'(10272);
			24691: out = 24'(-11844);
			24692: out = 24'(-31500);
			24693: out = 24'(-14816);
			24694: out = 24'(-5016);
			24695: out = 24'(16568);
			24696: out = 24'(26444);
			24697: out = 24'(30332);
			24698: out = 24'(27112);
			24699: out = 24'(12728);
			24700: out = 24'(-37936);
			24701: out = 24'(-88608);
			24702: out = 24'(-24052);
			24703: out = 24'(25436);
			24704: out = 24'(33352);
			24705: out = 24'(10356);
			24706: out = 24'(2216);
			24707: out = 24'(6396);
			24708: out = 24'(7216);
			24709: out = 24'(-4464);
			24710: out = 24'(-9464);
			24711: out = 24'(-4044);
			24712: out = 24'(6612);
			24713: out = 24'(8308);
			24714: out = 24'(1572);
			24715: out = 24'(-3044);
			24716: out = 24'(-3288);
			24717: out = 24'(7064);
			24718: out = 24'(16008);
			24719: out = 24'(-12284);
			24720: out = 24'(-17636);
			24721: out = 24'(-5476);
			24722: out = 24'(6352);
			24723: out = 24'(-3604);
			24724: out = 24'(-2832);
			24725: out = 24'(7948);
			24726: out = 24'(14344);
			24727: out = 24'(1608);
			24728: out = 24'(-8908);
			24729: out = 24'(-8708);
			24730: out = 24'(-2948);
			24731: out = 24'(-4568);
			24732: out = 24'(-3828);
			24733: out = 24'(3408);
			24734: out = 24'(17540);
			24735: out = 24'(28504);
			24736: out = 24'(6964);
			24737: out = 24'(1776);
			24738: out = 24'(-10276);
			24739: out = 24'(-23856);
			24740: out = 24'(-22568);
			24741: out = 24'(-6552);
			24742: out = 24'(1412);
			24743: out = 24'(952);
			24744: out = 24'(6608);
			24745: out = 24'(10020);
			24746: out = 24'(-2060);
			24747: out = 24'(-17672);
			24748: out = 24'(-12640);
			24749: out = 24'(-6296);
			24750: out = 24'(-2124);
			24751: out = 24'(-3288);
			24752: out = 24'(2596);
			24753: out = 24'(5444);
			24754: out = 24'(10504);
			24755: out = 24'(6420);
			24756: out = 24'(-1528);
			24757: out = 24'(-13584);
			24758: out = 24'(-12268);
			24759: out = 24'(-5484);
			24760: out = 24'(2440);
			24761: out = 24'(84);
			24762: out = 24'(13996);
			24763: out = 24'(12776);
			24764: out = 24'(4408);
			24765: out = 24'(128);
			24766: out = 24'(8308);
			24767: out = 24'(7148);
			24768: out = 24'(448);
			24769: out = 24'(-3456);
			24770: out = 24'(8708);
			24771: out = 24'(-4084);
			24772: out = 24'(-19740);
			24773: out = 24'(-12584);
			24774: out = 24'(12332);
			24775: out = 24'(13416);
			24776: out = 24'(-7380);
			24777: out = 24'(-19932);
			24778: out = 24'(-4232);
			24779: out = 24'(19028);
			24780: out = 24'(19936);
			24781: out = 24'(4476);
			24782: out = 24'(-2976);
			24783: out = 24'(-1716);
			24784: out = 24'(-444);
			24785: out = 24'(-10668);
			24786: out = 24'(-24404);
			24787: out = 24'(-10252);
			24788: out = 24'(7964);
			24789: out = 24'(21132);
			24790: out = 24'(21728);
			24791: out = 24'(2088);
			24792: out = 24'(-4124);
			24793: out = 24'(-3784);
			24794: out = 24'(-6080);
			24795: out = 24'(-13612);
			24796: out = 24'(-13264);
			24797: out = 24'(-1708);
			24798: out = 24'(8244);
			24799: out = 24'(6468);
			24800: out = 24'(-1528);
			24801: out = 24'(408);
			24802: out = 24'(10984);
			24803: out = 24'(14484);
			24804: out = 24'(8772);
			24805: out = 24'(-1040);
			24806: out = 24'(-4764);
			24807: out = 24'(-5680);
			24808: out = 24'(-16768);
			24809: out = 24'(-14676);
			24810: out = 24'(-4756);
			24811: out = 24'(740);
			24812: out = 24'(1520);
			24813: out = 24'(6436);
			24814: out = 24'(16312);
			24815: out = 24'(15060);
			24816: out = 24'(540);
			24817: out = 24'(-1956);
			24818: out = 24'(9380);
			24819: out = 24'(13108);
			24820: out = 24'(1956);
			24821: out = 24'(-10408);
			24822: out = 24'(-6740);
			24823: out = 24'(-9180);
			24824: out = 24'(-19248);
			24825: out = 24'(5112);
			24826: out = 24'(29568);
			24827: out = 24'(24292);
			24828: out = 24'(-3236);
			24829: out = 24'(6180);
			24830: out = 24'(11924);
			24831: out = 24'(6680);
			24832: out = 24'(-12860);
			24833: out = 24'(-16408);
			24834: out = 24'(-9580);
			24835: out = 24'(4024);
			24836: out = 24'(7480);
			24837: out = 24'(-1112);
			24838: out = 24'(-292);
			24839: out = 24'(-4072);
			24840: out = 24'(-516);
			24841: out = 24'(8572);
			24842: out = 24'(7076);
			24843: out = 24'(-5388);
			24844: out = 24'(-10052);
			24845: out = 24'(-3692);
			24846: out = 24'(2780);
			24847: out = 24'(-21360);
			24848: out = 24'(-23568);
			24849: out = 24'(13100);
			24850: out = 24'(31204);
			24851: out = 24'(13664);
			24852: out = 24'(-19048);
			24853: out = 24'(-22132);
			24854: out = 24'(-2144);
			24855: out = 24'(928);
			24856: out = 24'(-22844);
			24857: out = 24'(-28372);
			24858: out = 24'(5644);
			24859: out = 24'(14508);
			24860: out = 24'(10644);
			24861: out = 24'(10572);
			24862: out = 24'(22948);
			24863: out = 24'(1672);
			24864: out = 24'(-4028);
			24865: out = 24'(3536);
			24866: out = 24'(17436);
			24867: out = 24'(-4568);
			24868: out = 24'(-8596);
			24869: out = 24'(-11944);
			24870: out = 24'(-10580);
			24871: out = 24'(-17704);
			24872: out = 24'(4120);
			24873: out = 24'(14236);
			24874: out = 24'(14068);
			24875: out = 24'(9064);
			24876: out = 24'(14144);
			24877: out = 24'(7496);
			24878: out = 24'(-8716);
			24879: out = 24'(-24240);
			24880: out = 24'(-12540);
			24881: out = 24'(-3008);
			24882: out = 24'(1100);
			24883: out = 24'(732);
			24884: out = 24'(9440);
			24885: out = 24'(3180);
			24886: out = 24'(-996);
			24887: out = 24'(2348);
			24888: out = 24'(14476);
			24889: out = 24'(3848);
			24890: out = 24'(-1908);
			24891: out = 24'(-1916);
			24892: out = 24'(-11960);
			24893: out = 24'(-7056);
			24894: out = 24'(-11772);
			24895: out = 24'(-11472);
			24896: out = 24'(708);
			24897: out = 24'(7856);
			24898: out = 24'(9908);
			24899: out = 24'(8688);
			24900: out = 24'(8220);
			24901: out = 24'(-3788);
			24902: out = 24'(1860);
			24903: out = 24'(7552);
			24904: out = 24'(720);
			24905: out = 24'(-26692);
			24906: out = 24'(-10680);
			24907: out = 24'(11752);
			24908: out = 24'(5772);
			24909: out = 24'(-30360);
			24910: out = 24'(-24188);
			24911: out = 24'(9192);
			24912: out = 24'(29392);
			24913: out = 24'(12256);
			24914: out = 24'(-348);
			24915: out = 24'(-4356);
			24916: out = 24'(840);
			24917: out = 24'(-3352);
			24918: out = 24'(-14968);
			24919: out = 24'(-9412);
			24920: out = 24'(11056);
			24921: out = 24'(19632);
			24922: out = 24'(16572);
			24923: out = 24'(1880);
			24924: out = 24'(5880);
			24925: out = 24'(14000);
			24926: out = 24'(4676);
			24927: out = 24'(-27356);
			24928: out = 24'(-31268);
			24929: out = 24'(-2288);
			24930: out = 24'(12628);
			24931: out = 24'(21064);
			24932: out = 24'(-6200);
			24933: out = 24'(-20584);
			24934: out = 24'(268);
			24935: out = 24'(18964);
			24936: out = 24'(15208);
			24937: out = 24'(-6268);
			24938: out = 24'(-15820);
			24939: out = 24'(-664);
			24940: out = 24'(548);
			24941: out = 24'(-16940);
			24942: out = 24'(-23392);
			24943: out = 24'(8768);
			24944: out = 24'(19708);
			24945: out = 24'(10940);
			24946: out = 24'(-3336);
			24947: out = 24'(-3060);
			24948: out = 24'(11560);
			24949: out = 24'(8280);
			24950: out = 24'(-5364);
			24951: out = 24'(-5764);
			24952: out = 24'(-2796);
			24953: out = 24'(10516);
			24954: out = 24'(11548);
			24955: out = 24'(-2312);
			24956: out = 24'(-22648);
			24957: out = 24'(-9008);
			24958: out = 24'(17748);
			24959: out = 24'(24452);
			24960: out = 24'(9996);
			24961: out = 24'(3468);
			24962: out = 24'(11464);
			24963: out = 24'(5816);
			24964: out = 24'(-21824);
			24965: out = 24'(-31244);
			24966: out = 24'(-5008);
			24967: out = 24'(16512);
			24968: out = 24'(3084);
			24969: out = 24'(696);
			24970: out = 24'(4092);
			24971: out = 24'(7740);
			24972: out = 24'(1392);
			24973: out = 24'(5016);
			24974: out = 24'(11352);
			24975: out = 24'(7928);
			24976: out = 24'(-11844);
			24977: out = 24'(-35532);
			24978: out = 24'(-27832);
			24979: out = 24'(-15072);
			24980: out = 24'(-8592);
			24981: out = 24'(1480);
			24982: out = 24'(18456);
			24983: out = 24'(24344);
			24984: out = 24'(13720);
			24985: out = 24'(-2692);
			24986: out = 24'(-15784);
			24987: out = 24'(-20024);
			24988: out = 24'(-11476);
			24989: out = 24'(4128);
			24990: out = 24'(8732);
			24991: out = 24'(3448);
			24992: out = 24'(-2644);
			24993: out = 24'(-5504);
			24994: out = 24'(-17060);
			24995: out = 24'(-5944);
			24996: out = 24'(6384);
			24997: out = 24'(8312);
			24998: out = 24'(3544);
			24999: out = 24'(-1168);
			25000: out = 24'(8168);
			25001: out = 24'(13796);
			25002: out = 24'(1544);
			25003: out = 24'(-8100);
			25004: out = 24'(-11712);
			25005: out = 24'(-9916);
			25006: out = 24'(-9076);
			25007: out = 24'(8032);
			25008: out = 24'(5348);
			25009: out = 24'(-6488);
			25010: out = 24'(-10380);
			25011: out = 24'(13324);
			25012: out = 24'(17616);
			25013: out = 24'(3728);
			25014: out = 24'(-11560);
			25015: out = 24'(-3100);
			25016: out = 24'(10732);
			25017: out = 24'(13136);
			25018: out = 24'(340);
			25019: out = 24'(-9200);
			25020: out = 24'(1640);
			25021: out = 24'(13468);
			25022: out = 24'(7812);
			25023: out = 24'(-12612);
			25024: out = 24'(-13632);
			25025: out = 24'(-12656);
			25026: out = 24'(-9732);
			25027: out = 24'(-9360);
			25028: out = 24'(6856);
			25029: out = 24'(1420);
			25030: out = 24'(7920);
			25031: out = 24'(23972);
			25032: out = 24'(26320);
			25033: out = 24'(7856);
			25034: out = 24'(-10424);
			25035: out = 24'(-13140);
			25036: out = 24'(-8904);
			25037: out = 24'(-17612);
			25038: out = 24'(-21000);
			25039: out = 24'(-532);
			25040: out = 24'(28672);
			25041: out = 24'(24712);
			25042: out = 24'(8004);
			25043: out = 24'(-2384);
			25044: out = 24'(-784);
			25045: out = 24'(-7124);
			25046: out = 24'(-8988);
			25047: out = 24'(856);
			25048: out = 24'(15704);
			25049: out = 24'(7912);
			25050: out = 24'(-2812);
			25051: out = 24'(-7960);
			25052: out = 24'(3844);
			25053: out = 24'(11872);
			25054: out = 24'(5184);
			25055: out = 24'(-19664);
			25056: out = 24'(-28964);
			25057: out = 24'(-1164);
			25058: out = 24'(18008);
			25059: out = 24'(18088);
			25060: out = 24'(-2412);
			25061: out = 24'(-16496);
			25062: out = 24'(-3912);
			25063: out = 24'(6392);
			25064: out = 24'(-3356);
			25065: out = 24'(-19472);
			25066: out = 24'(-21592);
			25067: out = 24'(128);
			25068: out = 24'(16852);
			25069: out = 24'(17776);
			25070: out = 24'(-1128);
			25071: out = 24'(936);
			25072: out = 24'(-15992);
			25073: out = 24'(-37064);
			25074: out = 24'(-41488);
			25075: out = 24'(-7360);
			25076: out = 24'(7680);
			25077: out = 24'(8036);
			25078: out = 24'(11892);
			25079: out = 24'(22732);
			25080: out = 24'(14392);
			25081: out = 24'(428);
			25082: out = 24'(-7744);
			25083: out = 24'(-9352);
			25084: out = 24'(-13536);
			25085: out = 24'(-7400);
			25086: out = 24'(1396);
			25087: out = 24'(-2308);
			25088: out = 24'(-1500);
			25089: out = 24'(13448);
			25090: out = 24'(20160);
			25091: out = 24'(-4808);
			25092: out = 24'(-17844);
			25093: out = 24'(-12976);
			25094: out = 24'(572);
			25095: out = 24'(484);
			25096: out = 24'(6600);
			25097: out = 24'(15868);
			25098: out = 24'(18804);
			25099: out = 24'(2064);
			25100: out = 24'(-10536);
			25101: out = 24'(-14280);
			25102: out = 24'(-1808);
			25103: out = 24'(6320);
			25104: out = 24'(1144);
			25105: out = 24'(1432);
			25106: out = 24'(5648);
			25107: out = 24'(4916);
			25108: out = 24'(940);
			25109: out = 24'(-1004);
			25110: out = 24'(5816);
			25111: out = 24'(7368);
			25112: out = 24'(-76);
			25113: out = 24'(-1456);
			25114: out = 24'(13176);
			25115: out = 24'(23252);
			25116: out = 24'(10644);
			25117: out = 24'(4860);
			25118: out = 24'(-19888);
			25119: out = 24'(-28424);
			25120: out = 24'(-10928);
			25121: out = 24'(17632);
			25122: out = 24'(8820);
			25123: out = 24'(-12112);
			25124: out = 24'(-9120);
			25125: out = 24'(26908);
			25126: out = 24'(26264);
			25127: out = 24'(6844);
			25128: out = 24'(-2160);
			25129: out = 24'(14108);
			25130: out = 24'(2124);
			25131: out = 24'(-16264);
			25132: out = 24'(-22284);
			25133: out = 24'(-1564);
			25134: out = 24'(856);
			25135: out = 24'(1664);
			25136: out = 24'(-3924);
			25137: out = 24'(-2668);
			25138: out = 24'(4528);
			25139: out = 24'(8780);
			25140: out = 24'(4704);
			25141: out = 24'(-1784);
			25142: out = 24'(-304);
			25143: out = 24'(-4340);
			25144: out = 24'(-2768);
			25145: out = 24'(-1092);
			25146: out = 24'(-4568);
			25147: out = 24'(-2032);
			25148: out = 24'(-2308);
			25149: out = 24'(-7072);
			25150: out = 24'(-9708);
			25151: out = 24'(-3412);
			25152: out = 24'(10496);
			25153: out = 24'(10632);
			25154: out = 24'(-3588);
			25155: out = 24'(-10116);
			25156: out = 24'(-6516);
			25157: out = 24'(-8204);
			25158: out = 24'(-18908);
			25159: out = 24'(-8536);
			25160: out = 24'(7036);
			25161: out = 24'(25576);
			25162: out = 24'(21552);
			25163: out = 24'(-1180);
			25164: out = 24'(-24584);
			25165: out = 24'(-26524);
			25166: out = 24'(-16852);
			25167: out = 24'(-5016);
			25168: out = 24'(6816);
			25169: out = 24'(20376);
			25170: out = 24'(16828);
			25171: out = 24'(-1560);
			25172: out = 24'(2828);
			25173: out = 24'(416);
			25174: out = 24'(-2620);
			25175: out = 24'(-3360);
			25176: out = 24'(-1504);
			25177: out = 24'(11972);
			25178: out = 24'(9392);
			25179: out = 24'(-4016);
			25180: out = 24'(-9832);
			25181: out = 24'(2220);
			25182: out = 24'(5044);
			25183: out = 24'(-4932);
			25184: out = 24'(-13100);
			25185: out = 24'(-2440);
			25186: out = 24'(1792);
			25187: out = 24'(-3464);
			25188: out = 24'(-9640);
			25189: out = 24'(-516);
			25190: out = 24'(10052);
			25191: out = 24'(17340);
			25192: out = 24'(13020);
			25193: out = 24'(16512);
			25194: out = 24'(-22204);
			25195: out = 24'(-39792);
			25196: out = 24'(-24588);
			25197: out = 24'(264);
			25198: out = 24'(7844);
			25199: out = 24'(21196);
			25200: out = 24'(30020);
			25201: out = 24'(11464);
			25202: out = 24'(-10856);
			25203: out = 24'(-22164);
			25204: out = 24'(-10160);
			25205: out = 24'(-908);
			25206: out = 24'(1816);
			25207: out = 24'(-9304);
			25208: out = 24'(1088);
			25209: out = 24'(27856);
			25210: out = 24'(39604);
			25211: out = 24'(13984);
			25212: out = 24'(-15872);
			25213: out = 24'(-22132);
			25214: out = 24'(-5688);
			25215: out = 24'(-3128);
			25216: out = 24'(-5428);
			25217: out = 24'(-988);
			25218: out = 24'(5844);
			25219: out = 24'(16660);
			25220: out = 24'(8352);
			25221: out = 24'(-3816);
			25222: out = 24'(-2876);
			25223: out = 24'(6452);
			25224: out = 24'(4948);
			25225: out = 24'(-6500);
			25226: out = 24'(-8284);
			25227: out = 24'(5852);
			25228: out = 24'(20620);
			25229: out = 24'(11148);
			25230: out = 24'(-13256);
			25231: out = 24'(-20460);
			25232: out = 24'(-7796);
			25233: out = 24'(4428);
			25234: out = 24'(-3980);
			25235: out = 24'(-23132);
			25236: out = 24'(-8200);
			25237: out = 24'(17656);
			25238: out = 24'(27464);
			25239: out = 24'(18092);
			25240: out = 24'(-1824);
			25241: out = 24'(-4324);
			25242: out = 24'(-3536);
			25243: out = 24'(-15028);
			25244: out = 24'(-33532);
			25245: out = 24'(-27412);
			25246: out = 24'(-4036);
			25247: out = 24'(11872);
			25248: out = 24'(23664);
			25249: out = 24'(10412);
			25250: out = 24'(1492);
			25251: out = 24'(-8616);
			25252: out = 24'(-20212);
			25253: out = 24'(-23344);
			25254: out = 24'(-4796);
			25255: out = 24'(14524);
			25256: out = 24'(16656);
			25257: out = 24'(-3048);
			25258: out = 24'(-4588);
			25259: out = 24'(3840);
			25260: out = 24'(5756);
			25261: out = 24'(3380);
			25262: out = 24'(1128);
			25263: out = 24'(-1448);
			25264: out = 24'(-2204);
			25265: out = 24'(8492);
			25266: out = 24'(14480);
			25267: out = 24'(8500);
			25268: out = 24'(-1564);
			25269: out = 24'(6252);
			25270: out = 24'(1268);
			25271: out = 24'(-8672);
			25272: out = 24'(-19428);
			25273: out = 24'(-12064);
			25274: out = 24'(-4084);
			25275: out = 24'(5392);
			25276: out = 24'(6468);
			25277: out = 24'(11188);
			25278: out = 24'(12484);
			25279: out = 24'(19316);
			25280: out = 24'(4112);
			25281: out = 24'(-24116);
			25282: out = 24'(-24116);
			25283: out = 24'(-8620);
			25284: out = 24'(8476);
			25285: out = 24'(17452);
			25286: out = 24'(27396);
			25287: out = 24'(14724);
			25288: out = 24'(-2356);
			25289: out = 24'(-10788);
			25290: out = 24'(-4692);
			25291: out = 24'(-216);
			25292: out = 24'(-7916);
			25293: out = 24'(-12808);
			25294: out = 24'(1448);
			25295: out = 24'(14104);
			25296: out = 24'(24772);
			25297: out = 24'(24128);
			25298: out = 24'(9324);
			25299: out = 24'(-11200);
			25300: out = 24'(-23324);
			25301: out = 24'(-14724);
			25302: out = 24'(-5300);
			25303: out = 24'(-5984);
			25304: out = 24'(-13288);
			25305: out = 24'(7332);
			25306: out = 24'(28360);
			25307: out = 24'(16060);
			25308: out = 24'(-16648);
			25309: out = 24'(-17076);
			25310: out = 24'(5268);
			25311: out = 24'(2664);
			25312: out = 24'(-9776);
			25313: out = 24'(-11972);
			25314: out = 24'(204);
			25315: out = 24'(-2492);
			25316: out = 24'(-1908);
			25317: out = 24'(-2672);
			25318: out = 24'(7484);
			25319: out = 24'(4552);
			25320: out = 24'(-10512);
			25321: out = 24'(-27928);
			25322: out = 24'(-10820);
			25323: out = 24'(21228);
			25324: out = 24'(28768);
			25325: out = 24'(3248);
			25326: out = 24'(-15128);
			25327: out = 24'(-9928);
			25328: out = 24'(-1848);
			25329: out = 24'(1564);
			25330: out = 24'(-6508);
			25331: out = 24'(-8668);
			25332: out = 24'(1492);
			25333: out = 24'(19992);
			25334: out = 24'(12404);
			25335: out = 24'(-14916);
			25336: out = 24'(-32956);
			25337: out = 24'(-4552);
			25338: out = 24'(13508);
			25339: out = 24'(6988);
			25340: out = 24'(-6740);
			25341: out = 24'(6092);
			25342: out = 24'(13484);
			25343: out = 24'(4788);
			25344: out = 24'(-15812);
			25345: out = 24'(-15276);
			25346: out = 24'(1192);
			25347: out = 24'(20480);
			25348: out = 24'(15656);
			25349: out = 24'(-5152);
			25350: out = 24'(-14228);
			25351: out = 24'(-8432);
			25352: out = 24'(-5472);
			25353: out = 24'(-9764);
			25354: out = 24'(7396);
			25355: out = 24'(19244);
			25356: out = 24'(18256);
			25357: out = 24'(2156);
			25358: out = 24'(1212);
			25359: out = 24'(-1264);
			25360: out = 24'(9848);
			25361: out = 24'(16576);
			25362: out = 24'(13960);
			25363: out = 24'(-1788);
			25364: out = 24'(-7868);
			25365: out = 24'(-10580);
			25366: out = 24'(-14768);
			25367: out = 24'(-13460);
			25368: out = 24'(3380);
			25369: out = 24'(18740);
			25370: out = 24'(21048);
			25371: out = 24'(14144);
			25372: out = 24'(6228);
			25373: out = 24'(-9280);
			25374: out = 24'(-22740);
			25375: out = 24'(-13524);
			25376: out = 24'(7108);
			25377: out = 24'(12184);
			25378: out = 24'(2096);
			25379: out = 24'(-1048);
			25380: out = 24'(-4272);
			25381: out = 24'(-12332);
			25382: out = 24'(-18900);
			25383: out = 24'(-10496);
			25384: out = 24'(-896);
			25385: out = 24'(4600);
			25386: out = 24'(8056);
			25387: out = 24'(13488);
			25388: out = 24'(860);
			25389: out = 24'(-3064);
			25390: out = 24'(1372);
			25391: out = 24'(4652);
			25392: out = 24'(9020);
			25393: out = 24'(-2688);
			25394: out = 24'(-1616);
			25395: out = 24'(5976);
			25396: out = 24'(14144);
			25397: out = 24'(-23004);
			25398: out = 24'(-28384);
			25399: out = 24'(-4244);
			25400: out = 24'(3216);
			25401: out = 24'(-15544);
			25402: out = 24'(-20108);
			25403: out = 24'(-2480);
			25404: out = 24'(7812);
			25405: out = 24'(4572);
			25406: out = 24'(-1308);
			25407: out = 24'(1980);
			25408: out = 24'(5288);
			25409: out = 24'(264);
			25410: out = 24'(-7104);
			25411: out = 24'(-16992);
			25412: out = 24'(-24136);
			25413: out = 24'(-13588);
			25414: out = 24'(-3144);
			25415: out = 24'(956);
			25416: out = 24'(-5684);
			25417: out = 24'(-3892);
			25418: out = 24'(19760);
			25419: out = 24'(38760);
			25420: out = 24'(18264);
			25421: out = 24'(-29072);
			25422: out = 24'(-24956);
			25423: out = 24'(2356);
			25424: out = 24'(12044);
			25425: out = 24'(-10552);
			25426: out = 24'(-11928);
			25427: out = 24'(-10112);
			25428: out = 24'(-7636);
			25429: out = 24'(-12496);
			25430: out = 24'(8104);
			25431: out = 24'(6692);
			25432: out = 24'(5276);
			25433: out = 24'(-2028);
			25434: out = 24'(1976);
			25435: out = 24'(96);
			25436: out = 24'(12480);
			25437: out = 24'(8760);
			25438: out = 24'(-13488);
			25439: out = 24'(-12540);
			25440: out = 24'(13620);
			25441: out = 24'(29196);
			25442: out = 24'(9156);
			25443: out = 24'(-18308);
			25444: out = 24'(-26640);
			25445: out = 24'(-8516);
			25446: out = 24'(8640);
			25447: out = 24'(15988);
			25448: out = 24'(4344);
			25449: out = 24'(2788);
			25450: out = 24'(12460);
			25451: out = 24'(16432);
			25452: out = 24'(2392);
			25453: out = 24'(-12280);
			25454: out = 24'(-9052);
			25455: out = 24'(6788);
			25456: out = 24'(27976);
			25457: out = 24'(18404);
			25458: out = 24'(-2296);
			25459: out = 24'(-10396);
			25460: out = 24'(-6252);
			25461: out = 24'(-3528);
			25462: out = 24'(-5204);
			25463: out = 24'(-3120);
			25464: out = 24'(-1240);
			25465: out = 24'(10868);
			25466: out = 24'(12436);
			25467: out = 24'(4940);
			25468: out = 24'(15164);
			25469: out = 24'(-836);
			25470: out = 24'(-8860);
			25471: out = 24'(-10780);
			25472: out = 24'(-716);
			25473: out = 24'(-28316);
			25474: out = 24'(-18140);
			25475: out = 24'(10404);
			25476: out = 24'(21488);
			25477: out = 24'(16464);
			25478: out = 24'(13144);
			25479: out = 24'(12536);
			25480: out = 24'(408);
			25481: out = 24'(-25236);
			25482: out = 24'(-27956);
			25483: out = 24'(-11092);
			25484: out = 24'(-144);
			25485: out = 24'(548);
			25486: out = 24'(2088);
			25487: out = 24'(18276);
			25488: out = 24'(23480);
			25489: out = 24'(-1824);
			25490: out = 24'(-32432);
			25491: out = 24'(-37204);
			25492: out = 24'(-15048);
			25493: out = 24'(-1972);
			25494: out = 24'(-3336);
			25495: out = 24'(-10604);
			25496: out = 24'(-720);
			25497: out = 24'(16416);
			25498: out = 24'(15616);
			25499: out = 24'(92);
			25500: out = 24'(-19256);
			25501: out = 24'(-29524);
			25502: out = 24'(-19136);
			25503: out = 24'(-692);
			25504: out = 24'(16984);
			25505: out = 24'(18384);
			25506: out = 24'(8164);
			25507: out = 24'(704);
			25508: out = 24'(3868);
			25509: out = 24'(-4604);
			25510: out = 24'(-29892);
			25511: out = 24'(-44312);
			25512: out = 24'(-18936);
			25513: out = 24'(15780);
			25514: out = 24'(20868);
			25515: out = 24'(29876);
			25516: out = 24'(20484);
			25517: out = 24'(9008);
			25518: out = 24'(-4580);
			25519: out = 24'(-1948);
			25520: out = 24'(-9768);
			25521: out = 24'(-13088);
			25522: out = 24'(-9700);
			25523: out = 24'(1804);
			25524: out = 24'(12204);
			25525: out = 24'(20708);
			25526: out = 24'(21752);
			25527: out = 24'(13936);
			25528: out = 24'(3588);
			25529: out = 24'(-9732);
			25530: out = 24'(-19180);
			25531: out = 24'(-17712);
			25532: out = 24'(5576);
			25533: out = 24'(19336);
			25534: out = 24'(22508);
			25535: out = 24'(18884);
			25536: out = 24'(17440);
			25537: out = 24'(-956);
			25538: out = 24'(-20460);
			25539: out = 24'(-24152);
			25540: out = 24'(-1500);
			25541: out = 24'(11500);
			25542: out = 24'(13180);
			25543: out = 24'(7084);
			25544: out = 24'(10152);
			25545: out = 24'(17320);
			25546: out = 24'(24456);
			25547: out = 24'(9696);
			25548: out = 24'(-19084);
			25549: out = 24'(-31664);
			25550: out = 24'(-13908);
			25551: out = 24'(4756);
			25552: out = 24'(4320);
			25553: out = 24'(556);
			25554: out = 24'(3340);
			25555: out = 24'(3340);
			25556: out = 24'(-7072);
			25557: out = 24'(-15984);
			25558: out = 24'(-6328);
			25559: out = 24'(2016);
			25560: out = 24'(-452);
			25561: out = 24'(7536);
			25562: out = 24'(1500);
			25563: out = 24'(9068);
			25564: out = 24'(13096);
			25565: out = 24'(3920);
			25566: out = 24'(-10424);
			25567: out = 24'(-19532);
			25568: out = 24'(-18128);
			25569: out = 24'(-7772);
			25570: out = 24'(6764);
			25571: out = 24'(18604);
			25572: out = 24'(20464);
			25573: out = 24'(10708);
			25574: out = 24'(208);
			25575: out = 24'(-9200);
			25576: out = 24'(-11144);
			25577: out = 24'(-10148);
			25578: out = 24'(-3728);
			25579: out = 24'(-12064);
			25580: out = 24'(-9964);
			25581: out = 24'(2940);
			25582: out = 24'(22552);
			25583: out = 24'(7980);
			25584: out = 24'(2180);
			25585: out = 24'(-2280);
			25586: out = 24'(-4832);
			25587: out = 24'(-29488);
			25588: out = 24'(-18804);
			25589: out = 24'(-4400);
			25590: out = 24'(2920);
			25591: out = 24'(13240);
			25592: out = 24'(27564);
			25593: out = 24'(18400);
			25594: out = 24'(-3852);
			25595: out = 24'(-2968);
			25596: out = 24'(-1348);
			25597: out = 24'(-4076);
			25598: out = 24'(-11824);
			25599: out = 24'(-9332);
			25600: out = 24'(-1528);
			25601: out = 24'(-1256);
			25602: out = 24'(-1076);
			25603: out = 24'(10940);
			25604: out = 24'(20384);
			25605: out = 24'(6812);
			25606: out = 24'(-19208);
			25607: out = 24'(-26964);
			25608: out = 24'(2524);
			25609: out = 24'(11108);
			25610: out = 24'(4304);
			25611: out = 24'(1768);
			25612: out = 24'(7792);
			25613: out = 24'(8396);
			25614: out = 24'(-3744);
			25615: out = 24'(-14824);
			25616: out = 24'(-12796);
			25617: out = 24'(2576);
			25618: out = 24'(4888);
			25619: out = 24'(-1528);
			25620: out = 24'(2240);
			25621: out = 24'(11376);
			25622: out = 24'(16848);
			25623: out = 24'(6604);
			25624: out = 24'(-9436);
			25625: out = 24'(-26316);
			25626: out = 24'(-10604);
			25627: out = 24'(6916);
			25628: out = 24'(6964);
			25629: out = 24'(1568);
			25630: out = 24'(4564);
			25631: out = 24'(15756);
			25632: out = 24'(15592);
			25633: out = 24'(-352);
			25634: out = 24'(-14668);
			25635: out = 24'(-14972);
			25636: out = 24'(-9452);
			25637: out = 24'(-10556);
			25638: out = 24'(-15796);
			25639: out = 24'(-3328);
			25640: out = 24'(18728);
			25641: out = 24'(24268);
			25642: out = 24'(4328);
			25643: out = 24'(-13380);
			25644: out = 24'(-12968);
			25645: out = 24'(-2140);
			25646: out = 24'(116);
			25647: out = 24'(-36);
			25648: out = 24'(3008);
			25649: out = 24'(5152);
			25650: out = 24'(-3840);
			25651: out = 24'(-18604);
			25652: out = 24'(-22480);
			25653: out = 24'(-10200);
			25654: out = 24'(956);
			25655: out = 24'(16648);
			25656: out = 24'(14012);
			25657: out = 24'(8588);
			25658: out = 24'(10260);
			25659: out = 24'(16404);
			25660: out = 24'(8144);
			25661: out = 24'(-9980);
			25662: out = 24'(-23300);
			25663: out = 24'(-13852);
			25664: out = 24'(-6128);
			25665: out = 24'(-680);
			25666: out = 24'(1584);
			25667: out = 24'(7052);
			25668: out = 24'(12532);
			25669: out = 24'(16308);
			25670: out = 24'(10620);
			25671: out = 24'(-32);
			25672: out = 24'(-14832);
			25673: out = 24'(-11288);
			25674: out = 24'(688);
			25675: out = 24'(5216);
			25676: out = 24'(-7704);
			25677: out = 24'(-5376);
			25678: out = 24'(5180);
			25679: out = 24'(7196);
			25680: out = 24'(-4700);
			25681: out = 24'(-14740);
			25682: out = 24'(-12436);
			25683: out = 24'(908);
			25684: out = 24'(13760);
			25685: out = 24'(10040);
			25686: out = 24'(180);
			25687: out = 24'(-1540);
			25688: out = 24'(5636);
			25689: out = 24'(7344);
			25690: out = 24'(-2852);
			25691: out = 24'(-9072);
			25692: out = 24'(1492);
			25693: out = 24'(4980);
			25694: out = 24'(1396);
			25695: out = 24'(-5668);
			25696: out = 24'(-1412);
			25697: out = 24'(4144);
			25698: out = 24'(13240);
			25699: out = 24'(10192);
			25700: out = 24'(532);
			25701: out = 24'(-564);
			25702: out = 24'(-8076);
			25703: out = 24'(-7768);
			25704: out = 24'(6776);
			25705: out = 24'(25204);
			25706: out = 24'(18956);
			25707: out = 24'(-3300);
			25708: out = 24'(-20584);
			25709: out = 24'(-19716);
			25710: out = 24'(-9388);
			25711: out = 24'(-2816);
			25712: out = 24'(2132);
			25713: out = 24'(5756);
			25714: out = 24'(1300);
			25715: out = 24'(2216);
			25716: out = 24'(13740);
			25717: out = 24'(17048);
			25718: out = 24'(-19952);
			25719: out = 24'(-27508);
			25720: out = 24'(-4696);
			25721: out = 24'(17712);
			25722: out = 24'(-456);
			25723: out = 24'(-12496);
			25724: out = 24'(-13704);
			25725: out = 24'(-3124);
			25726: out = 24'(32);
			25727: out = 24'(3556);
			25728: out = 24'(2300);
			25729: out = 24'(-288);
			25730: out = 24'(392);
			25731: out = 24'(-6780);
			25732: out = 24'(-2820);
			25733: out = 24'(-9192);
			25734: out = 24'(-16340);
			25735: out = 24'(6576);
			25736: out = 24'(25684);
			25737: out = 24'(13068);
			25738: out = 24'(-17516);
			25739: out = 24'(-21272);
			25740: out = 24'(-5692);
			25741: out = 24'(3160);
			25742: out = 24'(3304);
			25743: out = 24'(18636);
			25744: out = 24'(18540);
			25745: out = 24'(2764);
			25746: out = 24'(-17644);
			25747: out = 24'(-13284);
			25748: out = 24'(-3200);
			25749: out = 24'(8356);
			25750: out = 24'(7488);
			25751: out = 24'(2856);
			25752: out = 24'(708);
			25753: out = 24'(5768);
			25754: out = 24'(12548);
			25755: out = 24'(12408);
			25756: out = 24'(1336);
			25757: out = 24'(-6520);
			25758: out = 24'(1976);
			25759: out = 24'(15732);
			25760: out = 24'(7280);
			25761: out = 24'(1944);
			25762: out = 24'(-1708);
			25763: out = 24'(6124);
			25764: out = 24'(11880);
			25765: out = 24'(-4592);
			25766: out = 24'(-23456);
			25767: out = 24'(-18184);
			25768: out = 24'(10988);
			25769: out = 24'(8068);
			25770: out = 24'(3876);
			25771: out = 24'(-1908);
			25772: out = 24'(960);
			25773: out = 24'(-1624);
			25774: out = 24'(7176);
			25775: out = 24'(3656);
			25776: out = 24'(-4680);
			25777: out = 24'(-340);
			25778: out = 24'(-60);
			25779: out = 24'(-4980);
			25780: out = 24'(-10472);
			25781: out = 24'(-2516);
			25782: out = 24'(12328);
			25783: out = 24'(19264);
			25784: out = 24'(10880);
			25785: out = 24'(-484);
			25786: out = 24'(-1644);
			25787: out = 24'(284);
			25788: out = 24'(-8164);
			25789: out = 24'(-19828);
			25790: out = 24'(-224);
			25791: out = 24'(7556);
			25792: out = 24'(4956);
			25793: out = 24'(-424);
			25794: out = 24'(7956);
			25795: out = 24'(2092);
			25796: out = 24'(-5104);
			25797: out = 24'(-6824);
			25798: out = 24'(-916);
			25799: out = 24'(4332);
			25800: out = 24'(2108);
			25801: out = 24'(-2236);
			25802: out = 24'(-400);
			25803: out = 24'(-1448);
			25804: out = 24'(-3444);
			25805: out = 24'(-2180);
			25806: out = 24'(6936);
			25807: out = 24'(12148);
			25808: out = 24'(7296);
			25809: out = 24'(-6672);
			25810: out = 24'(-13200);
			25811: out = 24'(-2040);
			25812: out = 24'(4476);
			25813: out = 24'(2292);
			25814: out = 24'(-1232);
			25815: out = 24'(-1476);
			25816: out = 24'(-164);
			25817: out = 24'(-14600);
			25818: out = 24'(-28476);
			25819: out = 24'(-9880);
			25820: out = 24'(13772);
			25821: out = 24'(34936);
			25822: out = 24'(24468);
			25823: out = 24'(-3600);
			25824: out = 24'(-20216);
			25825: out = 24'(-11616);
			25826: out = 24'(-5560);
			25827: out = 24'(-16804);
			25828: out = 24'(-19088);
			25829: out = 24'(-8084);
			25830: out = 24'(9480);
			25831: out = 24'(11844);
			25832: out = 24'(1236);
			25833: out = 24'(2964);
			25834: out = 24'(9716);
			25835: out = 24'(428);
			25836: out = 24'(-26840);
			25837: out = 24'(-26264);
			25838: out = 24'(-4660);
			25839: out = 24'(12648);
			25840: out = 24'(7728);
			25841: out = 24'(7480);
			25842: out = 24'(5236);
			25843: out = 24'(7548);
			25844: out = 24'(7572);
			25845: out = 24'(472);
			25846: out = 24'(-11428);
			25847: out = 24'(-20940);
			25848: out = 24'(-15076);
			25849: out = 24'(8100);
			25850: out = 24'(17172);
			25851: out = 24'(10696);
			25852: out = 24'(-1308);
			25853: out = 24'(-10416);
			25854: out = 24'(-9708);
			25855: out = 24'(-9512);
			25856: out = 24'(1328);
			25857: out = 24'(20324);
			25858: out = 24'(16056);
			25859: out = 24'(2592);
			25860: out = 24'(-4032);
			25861: out = 24'(-584);
			25862: out = 24'(-9204);
			25863: out = 24'(-26808);
			25864: out = 24'(-32372);
			25865: out = 24'(-12036);
			25866: out = 24'(13296);
			25867: out = 24'(26572);
			25868: out = 24'(24760);
			25869: out = 24'(16968);
			25870: out = 24'(8884);
			25871: out = 24'(7980);
			25872: out = 24'(5128);
			25873: out = 24'(-9368);
			25874: out = 24'(-31636);
			25875: out = 24'(-35524);
			25876: out = 24'(-15180);
			25877: out = 24'(10172);
			25878: out = 24'(20812);
			25879: out = 24'(22480);
			25880: out = 24'(17936);
			25881: out = 24'(5668);
			25882: out = 24'(-8284);
			25883: out = 24'(-536);
			25884: out = 24'(-616);
			25885: out = 24'(-164);
			25886: out = 24'(752);
			25887: out = 24'(5652);
			25888: out = 24'(1308);
			25889: out = 24'(-2872);
			25890: out = 24'(-3120);
			25891: out = 24'(-332);
			25892: out = 24'(-2592);
			25893: out = 24'(-8264);
			25894: out = 24'(-7536);
			25895: out = 24'(1296);
			25896: out = 24'(2808);
			25897: out = 24'(6820);
			25898: out = 24'(10148);
			25899: out = 24'(4628);
			25900: out = 24'(-20812);
			25901: out = 24'(-23636);
			25902: out = 24'(-12356);
			25903: out = 24'(-8580);
			25904: out = 24'(-17344);
			25905: out = 24'(-9844);
			25906: out = 24'(20288);
			25907: out = 24'(36344);
			25908: out = 24'(20484);
			25909: out = 24'(-13220);
			25910: out = 24'(-16024);
			25911: out = 24'(-2988);
			25912: out = 24'(-5016);
			25913: out = 24'(-14276);
			25914: out = 24'(-9436);
			25915: out = 24'(1428);
			25916: out = 24'(5048);
			25917: out = 24'(14544);
			25918: out = 24'(16392);
			25919: out = 24'(6420);
			25920: out = 24'(-7328);
			25921: out = 24'(764);
			25922: out = 24'(892);
			25923: out = 24'(-4268);
			25924: out = 24'(-8512);
			25925: out = 24'(1240);
			25926: out = 24'(8032);
			25927: out = 24'(6380);
			25928: out = 24'(3556);
			25929: out = 24'(9860);
			25930: out = 24'(14004);
			25931: out = 24'(832);
			25932: out = 24'(-14876);
			25933: out = 24'(-9360);
			25934: out = 24'(11008);
			25935: out = 24'(13744);
			25936: out = 24'(748);
			25937: out = 24'(-5960);
			25938: out = 24'(-1424);
			25939: out = 24'(3460);
			25940: out = 24'(-7964);
			25941: out = 24'(-21344);
			25942: out = 24'(-11708);
			25943: out = 24'(3736);
			25944: out = 24'(15984);
			25945: out = 24'(14828);
			25946: out = 24'(8440);
			25947: out = 24'(-10884);
			25948: out = 24'(-7688);
			25949: out = 24'(1748);
			25950: out = 24'(-2072);
			25951: out = 24'(-10660);
			25952: out = 24'(-10312);
			25953: out = 24'(9980);
			25954: out = 24'(26768);
			25955: out = 24'(14920);
			25956: out = 24'(372);
			25957: out = 24'(-3916);
			25958: out = 24'(-1652);
			25959: out = 24'(-14404);
			25960: out = 24'(-24092);
			25961: out = 24'(-21512);
			25962: out = 24'(-2140);
			25963: out = 24'(7904);
			25964: out = 24'(16384);
			25965: out = 24'(3424);
			25966: out = 24'(-2076);
			25967: out = 24'(7328);
			25968: out = 24'(16188);
			25969: out = 24'(8424);
			25970: out = 24'(-1556);
			25971: out = 24'(-5008);
			25972: out = 24'(-12892);
			25973: out = 24'(-16924);
			25974: out = 24'(-8256);
			25975: out = 24'(10304);
			25976: out = 24'(13176);
			25977: out = 24'(15408);
			25978: out = 24'(11128);
			25979: out = 24'(5492);
			25980: out = 24'(-8492);
			25981: out = 24'(-9644);
			25982: out = 24'(-7012);
			25983: out = 24'(7580);
			25984: out = 24'(20384);
			25985: out = 24'(11340);
			25986: out = 24'(-10016);
			25987: out = 24'(-26432);
			25988: out = 24'(-29592);
			25989: out = 24'(-11280);
			25990: out = 24'(2268);
			25991: out = 24'(18952);
			25992: out = 24'(25096);
			25993: out = 24'(15640);
			25994: out = 24'(-3792);
			25995: out = 24'(1040);
			25996: out = 24'(14924);
			25997: out = 24'(6636);
			25998: out = 24'(-11992);
			25999: out = 24'(-18596);
			26000: out = 24'(-9628);
			26001: out = 24'(-336);
			26002: out = 24'(-476);
			26003: out = 24'(-1748);
			26004: out = 24'(-5796);
			26005: out = 24'(-620);
			26006: out = 24'(9896);
			26007: out = 24'(26776);
			26008: out = 24'(7888);
			26009: out = 24'(-29312);
			26010: out = 24'(-42352);
			26011: out = 24'(-2172);
			26012: out = 24'(17756);
			26013: out = 24'(4408);
			26014: out = 24'(1548);
			26015: out = 24'(12832);
			26016: out = 24'(9032);
			26017: out = 24'(-10048);
			26018: out = 24'(-11372);
			26019: out = 24'(4048);
			26020: out = 24'(4924);
			26021: out = 24'(-10264);
			26022: out = 24'(-8988);
			26023: out = 24'(16392);
			26024: out = 24'(26472);
			26025: out = 24'(6324);
			26026: out = 24'(-18520);
			26027: out = 24'(-11040);
			26028: out = 24'(-3212);
			26029: out = 24'(-3816);
			26030: out = 24'(-10304);
			26031: out = 24'(444);
			26032: out = 24'(-16244);
			26033: out = 24'(-12552);
			26034: out = 24'(9624);
			26035: out = 24'(24872);
			26036: out = 24'(-9008);
			26037: out = 24'(-32000);
			26038: out = 24'(-14936);
			26039: out = 24'(21020);
			26040: out = 24'(9424);
			26041: out = 24'(148);
			26042: out = 24'(6544);
			26043: out = 24'(15592);
			26044: out = 24'(-904);
			26045: out = 24'(-21776);
			26046: out = 24'(-17108);
			26047: out = 24'(6172);
			26048: out = 24'(-460);
			26049: out = 24'(1024);
			26050: out = 24'(3092);
			26051: out = 24'(5168);
			26052: out = 24'(-7076);
			26053: out = 24'(-564);
			26054: out = 24'(1128);
			26055: out = 24'(-908);
			26056: out = 24'(-1912);
			26057: out = 24'(6568);
			26058: out = 24'(19320);
			26059: out = 24'(14956);
			26060: out = 24'(-7108);
			26061: out = 24'(-18636);
			26062: out = 24'(-10888);
			26063: out = 24'(2588);
			26064: out = 24'(5536);
			26065: out = 24'(652);
			26066: out = 24'(500);
			26067: out = 24'(-2688);
			26068: out = 24'(-7052);
			26069: out = 24'(-6004);
			26070: out = 24'(10872);
			26071: out = 24'(12752);
			26072: out = 24'(152);
			26073: out = 24'(-12952);
			26074: out = 24'(-7936);
			26075: out = 24'(-836);
			26076: out = 24'(8116);
			26077: out = 24'(14648);
			26078: out = 24'(15340);
			26079: out = 24'(4412);
			26080: out = 24'(-1008);
			26081: out = 24'(-900);
			26082: out = 24'(-3080);
			26083: out = 24'(-14600);
			26084: out = 24'(-8280);
			26085: out = 24'(10648);
			26086: out = 24'(15920);
			26087: out = 24'(11284);
			26088: out = 24'(3636);
			26089: out = 24'(-4056);
			26090: out = 24'(-13272);
			26091: out = 24'(-3516);
			26092: out = 24'(6812);
			26093: out = 24'(3208);
			26094: out = 24'(-10416);
			26095: out = 24'(-5812);
			26096: out = 24'(8884);
			26097: out = 24'(10564);
			26098: out = 24'(-3648);
			26099: out = 24'(-19416);
			26100: out = 24'(-7832);
			26101: out = 24'(1800);
			26102: out = 24'(-704);
			26103: out = 24'(328);
			26104: out = 24'(11164);
			26105: out = 24'(11404);
			26106: out = 24'(4112);
			26107: out = 24'(5636);
			26108: out = 24'(976);
			26109: out = 24'(-11784);
			26110: out = 24'(-20044);
			26111: out = 24'(-4480);
			26112: out = 24'(-2988);
			26113: out = 24'(6516);
			26114: out = 24'(9256);
			26115: out = 24'(7424);
			26116: out = 24'(-6136);
			26117: out = 24'(-7940);
			26118: out = 24'(-3476);
			26119: out = 24'(3888);
			26120: out = 24'(5456);
			26121: out = 24'(3564);
			26122: out = 24'(3884);
			26123: out = 24'(12224);
			26124: out = 24'(17128);
			26125: out = 24'(-2824);
			26126: out = 24'(-27460);
			26127: out = 24'(-30236);
			26128: out = 24'(-9160);
			26129: out = 24'(-4156);
			26130: out = 24'(-5568);
			26131: out = 24'(-3852);
			26132: out = 24'(3680);
			26133: out = 24'(6568);
			26134: out = 24'(5664);
			26135: out = 24'(10116);
			26136: out = 24'(12228);
			26137: out = 24'(-2612);
			26138: out = 24'(-24468);
			26139: out = 24'(-24684);
			26140: out = 24'(-3056);
			26141: out = 24'(5084);
			26142: out = 24'(10704);
			26143: out = 24'(2764);
			26144: out = 24'(-5820);
			26145: out = 24'(-8316);
			26146: out = 24'(10740);
			26147: out = 24'(18840);
			26148: out = 24'(11268);
			26149: out = 24'(-736);
			26150: out = 24'(1960);
			26151: out = 24'(11156);
			26152: out = 24'(10180);
			26153: out = 24'(-4268);
			26154: out = 24'(-18896);
			26155: out = 24'(-12468);
			26156: out = 24'(-240);
			26157: out = 24'(1500);
			26158: out = 24'(-9220);
			26159: out = 24'(-2116);
			26160: out = 24'(5452);
			26161: out = 24'(12764);
			26162: out = 24'(21816);
			26163: out = 24'(11512);
			26164: out = 24'(-3740);
			26165: out = 24'(-18016);
			26166: out = 24'(-21084);
			26167: out = 24'(-11596);
			26168: out = 24'(-2008);
			26169: out = 24'(2744);
			26170: out = 24'(7896);
			26171: out = 24'(13152);
			26172: out = 24'(15204);
			26173: out = 24'(8128);
			26174: out = 24'(-3092);
			26175: out = 24'(-15444);
			26176: out = 24'(-3024);
			26177: out = 24'(6308);
			26178: out = 24'(2308);
			26179: out = 24'(-8624);
			26180: out = 24'(4132);
			26181: out = 24'(16072);
			26182: out = 24'(14276);
			26183: out = 24'(-1248);
			26184: out = 24'(4892);
			26185: out = 24'(3452);
			26186: out = 24'(1336);
			26187: out = 24'(-1552);
			26188: out = 24'(-2944);
			26189: out = 24'(-21440);
			26190: out = 24'(-26236);
			26191: out = 24'(-2196);
			26192: out = 24'(10240);
			26193: out = 24'(22964);
			26194: out = 24'(8632);
			26195: out = 24'(-5268);
			26196: out = 24'(-7904);
			26197: out = 24'(4712);
			26198: out = 24'(-4180);
			26199: out = 24'(-12124);
			26200: out = 24'(-3932);
			26201: out = 24'(-1704);
			26202: out = 24'(-17768);
			26203: out = 24'(-16092);
			26204: out = 24'(18152);
			26205: out = 24'(22608);
			26206: out = 24'(4116);
			26207: out = 24'(-11656);
			26208: out = 24'(5732);
			26209: out = 24'(17108);
			26210: out = 24'(16108);
			26211: out = 24'(-8716);
			26212: out = 24'(-27196);
			26213: out = 24'(-25788);
			26214: out = 24'(740);
			26215: out = 24'(12272);
			26216: out = 24'(3800);
			26217: out = 24'(-8228);
			26218: out = 24'(-3336);
			26219: out = 24'(8984);
			26220: out = 24'(13416);
			26221: out = 24'(7144);
			26222: out = 24'(-7464);
			26223: out = 24'(-7392);
			26224: out = 24'(-892);
			26225: out = 24'(-1956);
			26226: out = 24'(-20000);
			26227: out = 24'(-13612);
			26228: out = 24'(1748);
			26229: out = 24'(4236);
			26230: out = 24'(-4168);
			26231: out = 24'(2564);
			26232: out = 24'(22968);
			26233: out = 24'(28672);
			26234: out = 24'(4764);
			26235: out = 24'(-9704);
			26236: out = 24'(-14056);
			26237: out = 24'(-14040);
			26238: out = 24'(-19480);
			26239: out = 24'(-19644);
			26240: out = 24'(-4992);
			26241: out = 24'(14328);
			26242: out = 24'(20808);
			26243: out = 24'(18080);
			26244: out = 24'(5428);
			26245: out = 24'(-1900);
			26246: out = 24'(308);
			26247: out = 24'(-1092);
			26248: out = 24'(-888);
			26249: out = 24'(-12888);
			26250: out = 24'(-20556);
			26251: out = 24'(-2944);
			26252: out = 24'(5008);
			26253: out = 24'(2328);
			26254: out = 24'(-2528);
			26255: out = 24'(7520);
			26256: out = 24'(5516);
			26257: out = 24'(3496);
			26258: out = 24'(-3676);
			26259: out = 24'(-4540);
			26260: out = 24'(11264);
			26261: out = 24'(13060);
			26262: out = 24'(-1500);
			26263: out = 24'(-17372);
			26264: out = 24'(-16404);
			26265: out = 24'(-5032);
			26266: out = 24'(1512);
			26267: out = 24'(1828);
			26268: out = 24'(15052);
			26269: out = 24'(17396);
			26270: out = 24'(18060);
			26271: out = 24'(8128);
			26272: out = 24'(-3084);
			26273: out = 24'(-2876);
			26274: out = 24'(6232);
			26275: out = 24'(1212);
			26276: out = 24'(-16844);
			26277: out = 24'(-9016);
			26278: out = 24'(9860);
			26279: out = 24'(20928);
			26280: out = 24'(15688);
			26281: out = 24'(256);
			26282: out = 24'(-1088);
			26283: out = 24'(-5572);
			26284: out = 24'(-16872);
			26285: out = 24'(-25792);
			26286: out = 24'(-7324);
			26287: out = 24'(6496);
			26288: out = 24'(6940);
			26289: out = 24'(2292);
			26290: out = 24'(4856);
			26291: out = 24'(6808);
			26292: out = 24'(8732);
			26293: out = 24'(5988);
			26294: out = 24'(-3836);
			26295: out = 24'(-21324);
			26296: out = 24'(-20692);
			26297: out = 24'(-1816);
			26298: out = 24'(-1068);
			26299: out = 24'(-8708);
			26300: out = 24'(-11828);
			26301: out = 24'(-4136);
			26302: out = 24'(2452);
			26303: out = 24'(744);
			26304: out = 24'(8764);
			26305: out = 24'(20628);
			26306: out = 24'(11596);
			26307: out = 24'(-13904);
			26308: out = 24'(-25824);
			26309: out = 24'(-10872);
			26310: out = 24'(752);
			26311: out = 24'(-7800);
			26312: out = 24'(-17692);
			26313: out = 24'(-5380);
			26314: out = 24'(8720);
			26315: out = 24'(3988);
			26316: out = 24'(-12500);
			26317: out = 24'(-1448);
			26318: out = 24'(25488);
			26319: out = 24'(21120);
			26320: out = 24'(6148);
			26321: out = 24'(-1120);
			26322: out = 24'(1972);
			26323: out = 24'(-10100);
			26324: out = 24'(-4572);
			26325: out = 24'(3368);
			26326: out = 24'(9076);
			26327: out = 24'(2260);
			26328: out = 24'(12788);
			26329: out = 24'(10676);
			26330: out = 24'(-2140);
			26331: out = 24'(-14200);
			26332: out = 24'(13000);
			26333: out = 24'(17796);
			26334: out = 24'(48);
			26335: out = 24'(-19272);
			26336: out = 24'(1016);
			26337: out = 24'(11788);
			26338: out = 24'(6884);
			26339: out = 24'(-5764);
			26340: out = 24'(332);
			26341: out = 24'(9552);
			26342: out = 24'(15480);
			26343: out = 24'(7252);
			26344: out = 24'(-11284);
			26345: out = 24'(-15432);
			26346: out = 24'(-19412);
			26347: out = 24'(-15524);
			26348: out = 24'(-1184);
			26349: out = 24'(12136);
			26350: out = 24'(11912);
			26351: out = 24'(4460);
			26352: out = 24'(-1740);
			26353: out = 24'(-6304);
			26354: out = 24'(832);
			26355: out = 24'(12028);
			26356: out = 24'(12716);
			26357: out = 24'(-3028);
			26358: out = 24'(-12788);
			26359: out = 24'(-4456);
			26360: out = 24'(6232);
			26361: out = 24'(-1308);
			26362: out = 24'(-10428);
			26363: out = 24'(-7844);
			26364: out = 24'(6184);
			26365: out = 24'(12096);
			26366: out = 24'(-544);
			26367: out = 24'(-9168);
			26368: out = 24'(-6384);
			26369: out = 24'(1320);
			26370: out = 24'(7936);
			26371: out = 24'(3424);
			26372: out = 24'(-2672);
			26373: out = 24'(-2540);
			26374: out = 24'(-924);
			26375: out = 24'(5460);
			26376: out = 24'(-1172);
			26377: out = 24'(-10912);
			26378: out = 24'(-5808);
			26379: out = 24'(-1584);
			26380: out = 24'(812);
			26381: out = 24'(-1824);
			26382: out = 24'(-2992);
			26383: out = 24'(1132);
			26384: out = 24'(6752);
			26385: out = 24'(8248);
			26386: out = 24'(4620);
			26387: out = 24'(984);
			26388: out = 24'(-3272);
			26389: out = 24'(-1180);
			26390: out = 24'(2776);
			26391: out = 24'(120);
			26392: out = 24'(-9372);
			26393: out = 24'(-10580);
			26394: out = 24'(-744);
			26395: out = 24'(-1124);
			26396: out = 24'(1832);
			26397: out = 24'(-5708);
			26398: out = 24'(-6412);
			26399: out = 24'(7872);
			26400: out = 24'(30420);
			26401: out = 24'(29772);
			26402: out = 24'(7544);
			26403: out = 24'(-18380);
			26404: out = 24'(-20024);
			26405: out = 24'(-14464);
			26406: out = 24'(-5196);
			26407: out = 24'(-68);
			26408: out = 24'(-3148);
			26409: out = 24'(-6120);
			26410: out = 24'(-3996);
			26411: out = 24'(2388);
			26412: out = 24'(8360);
			26413: out = 24'(12680);
			26414: out = 24'(10872);
			26415: out = 24'(-916);
			26416: out = 24'(-19112);
			26417: out = 24'(-4492);
			26418: out = 24'(2780);
			26419: out = 24'(-6656);
			26420: out = 24'(-17076);
			26421: out = 24'(3540);
			26422: out = 24'(20408);
			26423: out = 24'(8884);
			26424: out = 24'(-18288);
			26425: out = 24'(-16380);
			26426: out = 24'(1064);
			26427: out = 24'(8040);
			26428: out = 24'(-2012);
			26429: out = 24'(1436);
			26430: out = 24'(-3136);
			26431: out = 24'(-2120);
			26432: out = 24'(4524);
			26433: out = 24'(20728);
			26434: out = 24'(-368);
			26435: out = 24'(-16556);
			26436: out = 24'(-12608);
			26437: out = 24'(9504);
			26438: out = 24'(1408);
			26439: out = 24'(-1180);
			26440: out = 24'(4356);
			26441: out = 24'(13996);
			26442: out = 24'(6296);
			26443: out = 24'(-1008);
			26444: out = 24'(-2648);
			26445: out = 24'(3712);
			26446: out = 24'(7788);
			26447: out = 24'(6004);
			26448: out = 24'(8192);
			26449: out = 24'(14256);
			26450: out = 24'(11772);
			26451: out = 24'(2604);
			26452: out = 24'(-8900);
			26453: out = 24'(-14808);
			26454: out = 24'(-13352);
			26455: out = 24'(-11384);
			26456: out = 24'(-4580);
			26457: out = 24'(2912);
			26458: out = 24'(9356);
			26459: out = 24'(19140);
			26460: out = 24'(17096);
			26461: out = 24'(3412);
			26462: out = 24'(-13160);
			26463: out = 24'(-16620);
			26464: out = 24'(-13132);
			26465: out = 24'(-7108);
			26466: out = 24'(-3120);
			26467: out = 24'(-140);
			26468: out = 24'(1372);
			26469: out = 24'(4952);
			26470: out = 24'(10136);
			26471: out = 24'(12640);
			26472: out = 24'(13860);
			26473: out = 24'(676);
			26474: out = 24'(-20252);
			26475: out = 24'(-36312);
			26476: out = 24'(-13196);
			26477: out = 24'(1008);
			26478: out = 24'(9904);
			26479: out = 24'(13704);
			26480: out = 24'(14076);
			26481: out = 24'(1060);
			26482: out = 24'(-4448);
			26483: out = 24'(1172);
			26484: out = 24'(780);
			26485: out = 24'(-1772);
			26486: out = 24'(-8184);
			26487: out = 24'(-8244);
			26488: out = 24'(384);
			26489: out = 24'(6468);
			26490: out = 24'(9464);
			26491: out = 24'(2312);
			26492: out = 24'(-14676);
			26493: out = 24'(-19144);
			26494: out = 24'(-6160);
			26495: out = 24'(14680);
			26496: out = 24'(17408);
			26497: out = 24'(-468);
			26498: out = 24'(-5308);
			26499: out = 24'(10700);
			26500: out = 24'(16120);
			26501: out = 24'(-4920);
			26502: out = 24'(-35136);
			26503: out = 24'(-24636);
			26504: out = 24'(11128);
			26505: out = 24'(16516);
			26506: out = 24'(10024);
			26507: out = 24'(500);
			26508: out = 24'(972);
			26509: out = 24'(1552);
			26510: out = 24'(-10888);
			26511: out = 24'(-7268);
			26512: out = 24'(4104);
			26513: out = 24'(4528);
			26514: out = 24'(9308);
			26515: out = 24'(1560);
			26516: out = 24'(-2692);
			26517: out = 24'(-2184);
			26518: out = 24'(16008);
			26519: out = 24'(1608);
			26520: out = 24'(-8996);
			26521: out = 24'(-7344);
			26522: out = 24'(8112);
			26523: out = 24'(1208);
			26524: out = 24'(-5304);
			26525: out = 24'(-13392);
			26526: out = 24'(-14360);
			26527: out = 24'(172);
			26528: out = 24'(21976);
			26529: out = 24'(20652);
			26530: out = 24'(-3216);
			26531: out = 24'(-9372);
			26532: out = 24'(-6836);
			26533: out = 24'(-5676);
			26534: out = 24'(-10052);
			26535: out = 24'(-4224);
			26536: out = 24'(10988);
			26537: out = 24'(11740);
			26538: out = 24'(-6512);
			26539: out = 24'(-20516);
			26540: out = 24'(-3080);
			26541: out = 24'(15024);
			26542: out = 24'(11288);
			26543: out = 24'(-268);
			26544: out = 24'(-5044);
			26545: out = 24'(1028);
			26546: out = 24'(-1724);
			26547: out = 24'(-13936);
			26548: out = 24'(-19448);
			26549: out = 24'(-2904);
			26550: out = 24'(16608);
			26551: out = 24'(17364);
			26552: out = 24'(-7112);
			26553: out = 24'(-12292);
			26554: out = 24'(-2700);
			26555: out = 24'(7496);
			26556: out = 24'(13488);
			26557: out = 24'(3012);
			26558: out = 24'(-1840);
			26559: out = 24'(1700);
			26560: out = 24'(7356);
			26561: out = 24'(-6388);
			26562: out = 24'(-13756);
			26563: out = 24'(-11028);
			26564: out = 24'(-6600);
			26565: out = 24'(-872);
			26566: out = 24'(2624);
			26567: out = 24'(11760);
			26568: out = 24'(22048);
			26569: out = 24'(27444);
			26570: out = 24'(3412);
			26571: out = 24'(-24140);
			26572: out = 24'(-29532);
			26573: out = 24'(-1648);
			26574: out = 24'(1320);
			26575: out = 24'(-1552);
			26576: out = 24'(2868);
			26577: out = 24'(13032);
			26578: out = 24'(14700);
			26579: out = 24'(2376);
			26580: out = 24'(-8792);
			26581: out = 24'(-3416);
			26582: out = 24'(-13040);
			26583: out = 24'(-8252);
			26584: out = 24'(824);
			26585: out = 24'(8408);
			26586: out = 24'(128);
			26587: out = 24'(3148);
			26588: out = 24'(7212);
			26589: out = 24'(5984);
			26590: out = 24'(-9476);
			26591: out = 24'(-3832);
			26592: out = 24'(1320);
			26593: out = 24'(-4316);
			26594: out = 24'(-18744);
			26595: out = 24'(-8648);
			26596: out = 24'(6928);
			26597: out = 24'(14788);
			26598: out = 24'(13000);
			26599: out = 24'(6696);
			26600: out = 24'(-1532);
			26601: out = 24'(-13240);
			26602: out = 24'(-22176);
			26603: out = 24'(-8708);
			26604: out = 24'(-968);
			26605: out = 24'(148);
			26606: out = 24'(2724);
			26607: out = 24'(15144);
			26608: out = 24'(12948);
			26609: out = 24'(-2980);
			26610: out = 24'(-15704);
			26611: out = 24'(-3200);
			26612: out = 24'(0);
			26613: out = 24'(-1244);
			26614: out = 24'(-1628);
			26615: out = 24'(6924);
			26616: out = 24'(14716);
			26617: out = 24'(13464);
			26618: out = 24'(2576);
			26619: out = 24'(-10612);
			26620: out = 24'(-12316);
			26621: out = 24'(-11852);
			26622: out = 24'(-2804);
			26623: out = 24'(9132);
			26624: out = 24'(708);
			26625: out = 24'(-400);
			26626: out = 24'(3732);
			26627: out = 24'(8108);
			26628: out = 24'(-16);
			26629: out = 24'(-648);
			26630: out = 24'(-544);
			26631: out = 24'(-2544);
			26632: out = 24'(-9224);
			26633: out = 24'(-2920);
			26634: out = 24'(12040);
			26635: out = 24'(21148);
			26636: out = 24'(10856);
			26637: out = 24'(-5808);
			26638: out = 24'(-11436);
			26639: out = 24'(-596);
			26640: out = 24'(7388);
			26641: out = 24'(9176);
			26642: out = 24'(-8284);
			26643: out = 24'(-19176);
			26644: out = 24'(-12440);
			26645: out = 24'(7012);
			26646: out = 24'(1288);
			26647: out = 24'(-7200);
			26648: out = 24'(-3372);
			26649: out = 24'(5004);
			26650: out = 24'(13232);
			26651: out = 24'(7464);
			26652: out = 24'(-4964);
			26653: out = 24'(-15428);
			26654: out = 24'(-3180);
			26655: out = 24'(6532);
			26656: out = 24'(3676);
			26657: out = 24'(-13676);
			26658: out = 24'(5216);
			26659: out = 24'(1996);
			26660: out = 24'(-2608);
			26661: out = 24'(-6204);
			26662: out = 24'(9240);
			26663: out = 24'(5020);
			26664: out = 24'(11308);
			26665: out = 24'(12908);
			26666: out = 24'(1380);
			26667: out = 24'(-24784);
			26668: out = 24'(-17876);
			26669: out = 24'(6280);
			26670: out = 24'(15576);
			26671: out = 24'(-8168);
			26672: out = 24'(-3680);
			26673: out = 24'(10828);
			26674: out = 24'(2712);
			26675: out = 24'(-18316);
			26676: out = 24'(-12140);
			26677: out = 24'(8940);
			26678: out = 24'(14900);
			26679: out = 24'(6796);
			26680: out = 24'(6936);
			26681: out = 24'(2724);
			26682: out = 24'(-15076);
			26683: out = 24'(-30880);
			26684: out = 24'(-11604);
			26685: out = 24'(14144);
			26686: out = 24'(18464);
			26687: out = 24'(5656);
			26688: out = 24'(-4420);
			26689: out = 24'(-12472);
			26690: out = 24'(-16012);
			26691: out = 24'(-8108);
			26692: out = 24'(5484);
			26693: out = 24'(6236);
			26694: out = 24'(-5928);
			26695: out = 24'(-9428);
			26696: out = 24'(12268);
			26697: out = 24'(23464);
			26698: out = 24'(6180);
			26699: out = 24'(-22576);
			26700: out = 24'(-18640);
			26701: out = 24'(-11048);
			26702: out = 24'(-1600);
			26703: out = 24'(472);
			26704: out = 24'(1064);
			26705: out = 24'(104);
			26706: out = 24'(4836);
			26707: out = 24'(10132);
			26708: out = 24'(7980);
			26709: out = 24'(4168);
			26710: out = 24'(1232);
			26711: out = 24'(2976);
			26712: out = 24'(-1712);
			26713: out = 24'(1592);
			26714: out = 24'(-16288);
			26715: out = 24'(-15932);
			26716: out = 24'(6720);
			26717: out = 24'(15312);
			26718: out = 24'(2180);
			26719: out = 24'(-13608);
			26720: out = 24'(-12724);
			26721: out = 24'(-232);
			26722: out = 24'(1420);
			26723: out = 24'(-268);
			26724: out = 24'(4956);
			26725: out = 24'(21676);
			26726: out = 24'(3448);
			26727: out = 24'(-2828);
			26728: out = 24'(-4720);
			26729: out = 24'(-6076);
			26730: out = 24'(-2116);
			26731: out = 24'(2880);
			26732: out = 24'(-3148);
			26733: out = 24'(-11768);
			26734: out = 24'(-1816);
			26735: out = 24'(25036);
			26736: out = 24'(34360);
			26737: out = 24'(12068);
			26738: out = 24'(-38148);
			26739: out = 24'(-23680);
			26740: out = 24'(-196);
			26741: out = 24'(4300);
			26742: out = 24'(-2696);
			26743: out = 24'(3780);
			26744: out = 24'(4748);
			26745: out = 24'(-6000);
			26746: out = 24'(-18072);
			26747: out = 24'(-252);
			26748: out = 24'(11692);
			26749: out = 24'(11404);
			26750: out = 24'(984);
			26751: out = 24'(-7824);
			26752: out = 24'(-7120);
			26753: out = 24'(3044);
			26754: out = 24'(8176);
			26755: out = 24'(4116);
			26756: out = 24'(-228);
			26757: out = 24'(3608);
			26758: out = 24'(4800);
			26759: out = 24'(3580);
			26760: out = 24'(-21356);
			26761: out = 24'(-16156);
			26762: out = 24'(1112);
			26763: out = 24'(-316);
			26764: out = 24'(1256);
			26765: out = 24'(8068);
			26766: out = 24'(16384);
			26767: out = 24'(11688);
			26768: out = 24'(2048);
			26769: out = 24'(-1368);
			26770: out = 24'(-2888);
			26771: out = 24'(-11592);
			26772: out = 24'(-8004);
			26773: out = 24'(-13444);
			26774: out = 24'(-3992);
			26775: out = 24'(9320);
			26776: out = 24'(13752);
			26777: out = 24'(10416);
			26778: out = 24'(4084);
			26779: out = 24'(-1040);
			26780: out = 24'(-588);
			26781: out = 24'(-11480);
			26782: out = 24'(-11584);
			26783: out = 24'(-6588);
			26784: out = 24'(2236);
			26785: out = 24'(6880);
			26786: out = 24'(18420);
			26787: out = 24'(16696);
			26788: out = 24'(1540);
			26789: out = 24'(-17912);
			26790: out = 24'(-13860);
			26791: out = 24'(-4188);
			26792: out = 24'(1028);
			26793: out = 24'(-268);
			26794: out = 24'(-1184);
			26795: out = 24'(-8856);
			26796: out = 24'(-9624);
			26797: out = 24'(1496);
			26798: out = 24'(25204);
			26799: out = 24'(16768);
			26800: out = 24'(-7612);
			26801: out = 24'(-20556);
			26802: out = 24'(-768);
			26803: out = 24'(7932);
			26804: out = 24'(11360);
			26805: out = 24'(16176);
			26806: out = 24'(6088);
			26807: out = 24'(1304);
			26808: out = 24'(-248);
			26809: out = 24'(-2520);
			26810: out = 24'(-15468);
			26811: out = 24'(-24356);
			26812: out = 24'(-16572);
			26813: out = 24'(2340);
			26814: out = 24'(8380);
			26815: out = 24'(14132);
			26816: out = 24'(15556);
			26817: out = 24'(13864);
			26818: out = 24'(512);
			26819: out = 24'(540);
			26820: out = 24'(-3648);
			26821: out = 24'(-4012);
			26822: out = 24'(-7212);
			26823: out = 24'(2860);
			26824: out = 24'(2856);
			26825: out = 24'(14076);
			26826: out = 24'(20200);
			26827: out = 24'(1136);
			26828: out = 24'(-21236);
			26829: out = 24'(-16140);
			26830: out = 24'(7844);
			26831: out = 24'(5780);
			26832: out = 24'(5708);
			26833: out = 24'(-2792);
			26834: out = 24'(-800);
			26835: out = 24'(7856);
			26836: out = 24'(12344);
			26837: out = 24'(5180);
			26838: out = 24'(-6632);
			26839: out = 24'(-12768);
			26840: out = 24'(-8180);
			26841: out = 24'(-4420);
			26842: out = 24'(-3500);
			26843: out = 24'(856);
			26844: out = 24'(6304);
			26845: out = 24'(3736);
			26846: out = 24'(-6964);
			26847: out = 24'(-4072);
			26848: out = 24'(17928);
			26849: out = 24'(22608);
			26850: out = 24'(-652);
			26851: out = 24'(-21680);
			26852: out = 24'(-11284);
			26853: out = 24'(10676);
			26854: out = 24'(6872);
			26855: out = 24'(-9328);
			26856: out = 24'(-7876);
			26857: out = 24'(-924);
			26858: out = 24'(-1604);
			26859: out = 24'(-11252);
			26860: out = 24'(-10408);
			26861: out = 24'(-2680);
			26862: out = 24'(14724);
			26863: out = 24'(21604);
			26864: out = 24'(15344);
			26865: out = 24'(-6648);
			26866: out = 24'(-5820);
			26867: out = 24'(-1984);
			26868: out = 24'(-1220);
			26869: out = 24'(-4304);
			26870: out = 24'(-9324);
			26871: out = 24'(-4184);
			26872: out = 24'(5032);
			26873: out = 24'(3208);
			26874: out = 24'(-1492);
			26875: out = 24'(-9796);
			26876: out = 24'(-4616);
			26877: out = 24'(5136);
			26878: out = 24'(5884);
			26879: out = 24'(-9768);
			26880: out = 24'(-12604);
			26881: out = 24'(4076);
			26882: out = 24'(10844);
			26883: out = 24'(5084);
			26884: out = 24'(-8508);
			26885: out = 24'(-10476);
			26886: out = 24'(-712);
			26887: out = 24'(4904);
			26888: out = 24'(2112);
			26889: out = 24'(-2200);
			26890: out = 24'(-3616);
			26891: out = 24'(-540);
			26892: out = 24'(4016);
			26893: out = 24'(11576);
			26894: out = 24'(13916);
			26895: out = 24'(6700);
			26896: out = 24'(-6020);
			26897: out = 24'(-8904);
			26898: out = 24'(-3340);
			26899: out = 24'(-1180);
			26900: out = 24'(-14128);
			26901: out = 24'(-16356);
			26902: out = 24'(-56);
			26903: out = 24'(14324);
			26904: out = 24'(20740);
			26905: out = 24'(8440);
			26906: out = 24'(-10352);
			26907: out = 24'(-18128);
			26908: out = 24'(-15460);
			26909: out = 24'(-2556);
			26910: out = 24'(3156);
			26911: out = 24'(2408);
			26912: out = 24'(1148);
			26913: out = 24'(14020);
			26914: out = 24'(21388);
			26915: out = 24'(17116);
			26916: out = 24'(-376);
			26917: out = 24'(-660);
			26918: out = 24'(-7340);
			26919: out = 24'(-18912);
			26920: out = 24'(-25348);
			26921: out = 24'(-4016);
			26922: out = 24'(3412);
			26923: out = 24'(-2732);
			26924: out = 24'(-2376);
			26925: out = 24'(16080);
			26926: out = 24'(13272);
			26927: out = 24'(-7140);
			26928: out = 24'(-21044);
			26929: out = 24'(-12292);
			26930: out = 24'(-636);
			26931: out = 24'(2704);
			26932: out = 24'(644);
			26933: out = 24'(13112);
			26934: out = 24'(9572);
			26935: out = 24'(5172);
			26936: out = 24'(-4492);
			26937: out = 24'(-17012);
			26938: out = 24'(-31004);
			26939: out = 24'(-17676);
			26940: out = 24'(7692);
			26941: out = 24'(20264);
			26942: out = 24'(4088);
			26943: out = 24'(5888);
			26944: out = 24'(14492);
			26945: out = 24'(4664);
			26946: out = 24'(-25276);
			26947: out = 24'(-27112);
			26948: out = 24'(344);
			26949: out = 24'(19312);
			26950: out = 24'(-272);
			26951: out = 24'(-5452);
			26952: out = 24'(4328);
			26953: out = 24'(13344);
			26954: out = 24'(5668);
			26955: out = 24'(-944);
			26956: out = 24'(-4664);
			26957: out = 24'(-1812);
			26958: out = 24'(2184);
			26959: out = 24'(-8388);
			26960: out = 24'(-12256);
			26961: out = 24'(2496);
			26962: out = 24'(19880);
			26963: out = 24'(24616);
			26964: out = 24'(-1504);
			26965: out = 24'(-25108);
			26966: out = 24'(-21776);
			26967: out = 24'(-2740);
			26968: out = 24'(-1556);
			26969: out = 24'(-7112);
			26970: out = 24'(556);
			26971: out = 24'(6868);
			26972: out = 24'(15872);
			26973: out = 24'(11680);
			26974: out = 24'(2408);
			26975: out = 24'(-12300);
			26976: out = 24'(3816);
			26977: out = 24'(9980);
			26978: out = 24'(5116);
			26979: out = 24'(-3632);
			26980: out = 24'(1952);
			26981: out = 24'(-216);
			26982: out = 24'(-5332);
			26983: out = 24'(-6212);
			26984: out = 24'(-6548);
			26985: out = 24'(836);
			26986: out = 24'(10096);
			26987: out = 24'(11500);
			26988: out = 24'(1528);
			26989: out = 24'(-2000);
			26990: out = 24'(6484);
			26991: out = 24'(11264);
			26992: out = 24'(8);
			26993: out = 24'(-15328);
			26994: out = 24'(-17184);
			26995: out = 24'(-11372);
			26996: out = 24'(-12276);
			26997: out = 24'(-15004);
			26998: out = 24'(-4028);
			26999: out = 24'(12816);
			27000: out = 24'(20004);
			27001: out = 24'(10100);
			27002: out = 24'(2688);
			27003: out = 24'(-3732);
			27004: out = 24'(-5240);
			27005: out = 24'(-1328);
			27006: out = 24'(7476);
			27007: out = 24'(268);
			27008: out = 24'(-12604);
			27009: out = 24'(-3144);
			27010: out = 24'(11924);
			27011: out = 24'(10560);
			27012: out = 24'(-4220);
			27013: out = 24'(-7748);
			27014: out = 24'(4020);
			27015: out = 24'(10416);
			27016: out = 24'(5396);
			27017: out = 24'(2980);
			27018: out = 24'(-304);
			27019: out = 24'(-2012);
			27020: out = 24'(-3016);
			27021: out = 24'(3612);
			27022: out = 24'(6748);
			27023: out = 24'(84);
			27024: out = 24'(-14208);
			27025: out = 24'(-15736);
			27026: out = 24'(-1856);
			27027: out = 24'(2608);
			27028: out = 24'(-8244);
			27029: out = 24'(-12700);
			27030: out = 24'(-388);
			27031: out = 24'(132);
			27032: out = 24'(-17328);
			27033: out = 24'(-21676);
			27034: out = 24'(8880);
			27035: out = 24'(8592);
			27036: out = 24'(4748);
			27037: out = 24'(2176);
			27038: out = 24'(9632);
			27039: out = 24'(3564);
			27040: out = 24'(-2412);
			27041: out = 24'(-4784);
			27042: out = 24'(2636);
			27043: out = 24'(5072);
			27044: out = 24'(2784);
			27045: out = 24'(-2760);
			27046: out = 24'(-1532);
			27047: out = 24'(2460);
			27048: out = 24'(17364);
			27049: out = 24'(18812);
			27050: out = 24'(8412);
			27051: out = 24'(-288);
			27052: out = 24'(-4356);
			27053: out = 24'(792);
			27054: out = 24'(-1780);
			27055: out = 24'(-13112);
			27056: out = 24'(-18120);
			27057: out = 24'(-3384);
			27058: out = 24'(11608);
			27059: out = 24'(11624);
			27060: out = 24'(1112);
			27061: out = 24'(4572);
			27062: out = 24'(12028);
			27063: out = 24'(9752);
			27064: out = 24'(-5760);
			27065: out = 24'(-632);
			27066: out = 24'(6556);
			27067: out = 24'(4816);
			27068: out = 24'(-6588);
			27069: out = 24'(-1984);
			27070: out = 24'(6904);
			27071: out = 24'(16568);
			27072: out = 24'(20620);
			27073: out = 24'(9548);
			27074: out = 24'(-2728);
			27075: out = 24'(-7952);
			27076: out = 24'(-3492);
			27077: out = 24'(-1696);
			27078: out = 24'(-2348);
			27079: out = 24'(-7692);
			27080: out = 24'(-7736);
			27081: out = 24'(6876);
			27082: out = 24'(7880);
			27083: out = 24'(5668);
			27084: out = 24'(4400);
			27085: out = 24'(4100);
			27086: out = 24'(6864);
			27087: out = 24'(104);
			27088: out = 24'(-13092);
			27089: out = 24'(-21252);
			27090: out = 24'(-3052);
			27091: out = 24'(2712);
			27092: out = 24'(-9060);
			27093: out = 24'(-21096);
			27094: out = 24'(-11588);
			27095: out = 24'(1612);
			27096: out = 24'(5116);
			27097: out = 24'(1448);
			27098: out = 24'(-3508);
			27099: out = 24'(10320);
			27100: out = 24'(16324);
			27101: out = 24'(9724);
			27102: out = 24'(-188);
			27103: out = 24'(-712);
			27104: out = 24'(-2228);
			27105: out = 24'(-3632);
			27106: out = 24'(-472);
			27107: out = 24'(-5480);
			27108: out = 24'(-8144);
			27109: out = 24'(-772);
			27110: out = 24'(13548);
			27111: out = 24'(12844);
			27112: out = 24'(3952);
			27113: out = 24'(-2788);
			27114: out = 24'(-44);
			27115: out = 24'(-1232);
			27116: out = 24'(-8628);
			27117: out = 24'(-14060);
			27118: out = 24'(-5640);
			27119: out = 24'(6284);
			27120: out = 24'(3080);
			27121: out = 24'(-7440);
			27122: out = 24'(-5544);
			27123: out = 24'(6920);
			27124: out = 24'(4868);
			27125: out = 24'(-12148);
			27126: out = 24'(-19300);
			27127: out = 24'(-748);
			27128: out = 24'(12688);
			27129: out = 24'(13092);
			27130: out = 24'(2580);
			27131: out = 24'(-3556);
			27132: out = 24'(-4624);
			27133: out = 24'(8712);
			27134: out = 24'(18952);
			27135: out = 24'(15908);
			27136: out = 24'(48);
			27137: out = 24'(-7208);
			27138: out = 24'(-6084);
			27139: out = 24'(-6972);
			27140: out = 24'(-15692);
			27141: out = 24'(-5820);
			27142: out = 24'(14996);
			27143: out = 24'(26584);
			27144: out = 24'(16180);
			27145: out = 24'(-15976);
			27146: out = 24'(-25504);
			27147: out = 24'(-12324);
			27148: out = 24'(-736);
			27149: out = 24'(2092);
			27150: out = 24'(-936);
			27151: out = 24'(3960);
			27152: out = 24'(13448);
			27153: out = 24'(11564);
			27154: out = 24'(3428);
			27155: out = 24'(-10384);
			27156: out = 24'(-14560);
			27157: out = 24'(1028);
			27158: out = 24'(6368);
			27159: out = 24'(3568);
			27160: out = 24'(-2928);
			27161: out = 24'(-4092);
			27162: out = 24'(-1928);
			27163: out = 24'(-492);
			27164: out = 24'(-2352);
			27165: out = 24'(-3176);
			27166: out = 24'(12644);
			27167: out = 24'(10048);
			27168: out = 24'(-3908);
			27169: out = 24'(-10688);
			27170: out = 24'(17016);
			27171: out = 24'(17656);
			27172: out = 24'(4256);
			27173: out = 24'(-10352);
			27174: out = 24'(-10320);
			27175: out = 24'(-2932);
			27176: out = 24'(2504);
			27177: out = 24'(-2228);
			27178: out = 24'(-6548);
			27179: out = 24'(-4092);
			27180: out = 24'(8956);
			27181: out = 24'(11184);
			27182: out = 24'(-3104);
			27183: out = 24'(-9572);
			27184: out = 24'(-5788);
			27185: out = 24'(236);
			27186: out = 24'(-2884);
			27187: out = 24'(-9220);
			27188: out = 24'(-6040);
			27189: out = 24'(3636);
			27190: out = 24'(5240);
			27191: out = 24'(-3836);
			27192: out = 24'(-12112);
			27193: out = 24'(-9780);
			27194: out = 24'(-2344);
			27195: out = 24'(-1160);
			27196: out = 24'(-5144);
			27197: out = 24'(-5628);
			27198: out = 24'(5588);
			27199: out = 24'(19676);
			27200: out = 24'(16036);
			27201: out = 24'(3392);
			27202: out = 24'(-11276);
			27203: out = 24'(-19052);
			27204: out = 24'(-5520);
			27205: out = 24'(-3780);
			27206: out = 24'(-2872);
			27207: out = 24'(120);
			27208: out = 24'(-760);
			27209: out = 24'(-4568);
			27210: out = 24'(-7896);
			27211: out = 24'(-4672);
			27212: out = 24'(-564);
			27213: out = 24'(732);
			27214: out = 24'(-2300);
			27215: out = 24'(-2824);
			27216: out = 24'(-756);
			27217: out = 24'(676);
			27218: out = 24'(-2592);
			27219: out = 24'(-1832);
			27220: out = 24'(2588);
			27221: out = 24'(5668);
			27222: out = 24'(3028);
			27223: out = 24'(1520);
			27224: out = 24'(-1040);
			27225: out = 24'(1048);
			27226: out = 24'(-10648);
			27227: out = 24'(-2352);
			27228: out = 24'(17424);
			27229: out = 24'(18340);
			27230: out = 24'(9360);
			27231: out = 24'(-2720);
			27232: out = 24'(-8348);
			27233: out = 24'(-9908);
			27234: out = 24'(-5180);
			27235: out = 24'(-1816);
			27236: out = 24'(-1128);
			27237: out = 24'(988);
			27238: out = 24'(5876);
			27239: out = 24'(17124);
			27240: out = 24'(13208);
			27241: out = 24'(-2492);
			27242: out = 24'(2208);
			27243: out = 24'(3800);
			27244: out = 24'(224);
			27245: out = 24'(-8156);
			27246: out = 24'(-568);
			27247: out = 24'(-1468);
			27248: out = 24'(-156);
			27249: out = 24'(-1248);
			27250: out = 24'(-100);
			27251: out = 24'(624);
			27252: out = 24'(1320);
			27253: out = 24'(-3928);
			27254: out = 24'(-9284);
			27255: out = 24'(-3060);
			27256: out = 24'(9932);
			27257: out = 24'(13424);
			27258: out = 24'(1652);
			27259: out = 24'(-5196);
			27260: out = 24'(-9332);
			27261: out = 24'(-140);
			27262: out = 24'(6752);
			27263: out = 24'(-444);
			27264: out = 24'(-10588);
			27265: out = 24'(-8680);
			27266: out = 24'(3868);
			27267: out = 24'(11924);
			27268: out = 24'(8856);
			27269: out = 24'(5232);
			27270: out = 24'(2808);
			27271: out = 24'(-6092);
			27272: out = 24'(-11208);
			27273: out = 24'(-18468);
			27274: out = 24'(-15644);
			27275: out = 24'(-5528);
			27276: out = 24'(-1096);
			27277: out = 24'(-916);
			27278: out = 24'(2408);
			27279: out = 24'(9864);
			27280: out = 24'(14616);
			27281: out = 24'(-1340);
			27282: out = 24'(-19688);
			27283: out = 24'(-22528);
			27284: out = 24'(-9348);
			27285: out = 24'(3252);
			27286: out = 24'(6612);
			27287: out = 24'(4272);
			27288: out = 24'(-1000);
			27289: out = 24'(-2444);
			27290: out = 24'(-5768);
			27291: out = 24'(-4116);
			27292: out = 24'(444);
			27293: out = 24'(912);
			27294: out = 24'(-7700);
			27295: out = 24'(-10492);
			27296: out = 24'(732);
			27297: out = 24'(12292);
			27298: out = 24'(14788);
			27299: out = 24'(10864);
			27300: out = 24'(5652);
			27301: out = 24'(-9580);
			27302: out = 24'(-2032);
			27303: out = 24'(2252);
			27304: out = 24'(256);
			27305: out = 24'(-12844);
			27306: out = 24'(-4096);
			27307: out = 24'(-1364);
			27308: out = 24'(2772);
			27309: out = 24'(5696);
			27310: out = 24'(13824);
			27311: out = 24'(4748);
			27312: out = 24'(-856);
			27313: out = 24'(1032);
			27314: out = 24'(15580);
			27315: out = 24'(1848);
			27316: out = 24'(-1980);
			27317: out = 24'(6732);
			27318: out = 24'(6964);
			27319: out = 24'(1276);
			27320: out = 24'(-880);
			27321: out = 24'(-4264);
			27322: out = 24'(-19248);
			27323: out = 24'(-18476);
			27324: out = 24'(56);
			27325: out = 24'(14628);
			27326: out = 24'(5972);
			27327: out = 24'(1020);
			27328: out = 24'(3476);
			27329: out = 24'(6928);
			27330: out = 24'(-4192);
			27331: out = 24'(-19368);
			27332: out = 24'(-20508);
			27333: out = 24'(-8496);
			27334: out = 24'(920);
			27335: out = 24'(8552);
			27336: out = 24'(11652);
			27337: out = 24'(12236);
			27338: out = 24'(4748);
			27339: out = 24'(724);
			27340: out = 24'(-14064);
			27341: out = 24'(-8600);
			27342: out = 24'(3100);
			27343: out = 24'(4600);
			27344: out = 24'(612);
			27345: out = 24'(-1032);
			27346: out = 24'(464);
			27347: out = 24'(-960);
			27348: out = 24'(-5524);
			27349: out = 24'(-3736);
			27350: out = 24'(3672);
			27351: out = 24'(8740);
			27352: out = 24'(13244);
			27353: out = 24'(-2580);
			27354: out = 24'(-13624);
			27355: out = 24'(-8480);
			27356: out = 24'(4712);
			27357: out = 24'(13012);
			27358: out = 24'(3888);
			27359: out = 24'(-9824);
			27360: out = 24'(-7420);
			27361: out = 24'(8220);
			27362: out = 24'(16096);
			27363: out = 24'(6336);
			27364: out = 24'(-3156);
			27365: out = 24'(-2536);
			27366: out = 24'(6700);
			27367: out = 24'(-544);
			27368: out = 24'(-17100);
			27369: out = 24'(-13228);
			27370: out = 24'(364);
			27371: out = 24'(4580);
			27372: out = 24'(-3540);
			27373: out = 24'(-11968);
			27374: out = 24'(6824);
			27375: out = 24'(12528);
			27376: out = 24'(-1676);
			27377: out = 24'(-17700);
			27378: out = 24'(-4556);
			27379: out = 24'(8896);
			27380: out = 24'(13836);
			27381: out = 24'(11196);
			27382: out = 24'(-6228);
			27383: out = 24'(-17672);
			27384: out = 24'(-13428);
			27385: out = 24'(868);
			27386: out = 24'(-76);
			27387: out = 24'(1360);
			27388: out = 24'(5140);
			27389: out = 24'(8272);
			27390: out = 24'(8352);
			27391: out = 24'(-5532);
			27392: out = 24'(-6692);
			27393: out = 24'(2572);
			27394: out = 24'(4188);
			27395: out = 24'(-15584);
			27396: out = 24'(-16248);
			27397: out = 24'(7764);
			27398: out = 24'(20320);
			27399: out = 24'(17516);
			27400: out = 24'(-9708);
			27401: out = 24'(-20684);
			27402: out = 24'(-7260);
			27403: out = 24'(-4056);
			27404: out = 24'(-8876);
			27405: out = 24'(-7236);
			27406: out = 24'(11064);
			27407: out = 24'(18156);
			27408: out = 24'(27688);
			27409: out = 24'(14940);
			27410: out = 24'(-7848);
			27411: out = 24'(-27748);
			27412: out = 24'(-7948);
			27413: out = 24'(9772);
			27414: out = 24'(9128);
			27415: out = 24'(-3992);
			27416: out = 24'(-1148);
			27417: out = 24'(3432);
			27418: out = 24'(3120);
			27419: out = 24'(-4576);
			27420: out = 24'(-36);
			27421: out = 24'(-764);
			27422: out = 24'(144);
			27423: out = 24'(-1216);
			27424: out = 24'(-3072);
			27425: out = 24'(-2368);
			27426: out = 24'(4496);
			27427: out = 24'(5760);
			27428: out = 24'(-3344);
			27429: out = 24'(-16792);
			27430: out = 24'(-10844);
			27431: out = 24'(3336);
			27432: out = 24'(1160);
			27433: out = 24'(-5896);
			27434: out = 24'(-13132);
			27435: out = 24'(-5940);
			27436: out = 24'(10356);
			27437: out = 24'(19224);
			27438: out = 24'(11252);
			27439: out = 24'(-7084);
			27440: out = 24'(-18416);
			27441: out = 24'(-16544);
			27442: out = 24'(372);
			27443: out = 24'(5360);
			27444: out = 24'(-1000);
			27445: out = 24'(-2576);
			27446: out = 24'(1112);
			27447: out = 24'(2972);
			27448: out = 24'(3648);
			27449: out = 24'(8340);
			27450: out = 24'(1808);
			27451: out = 24'(-7588);
			27452: out = 24'(-12100);
			27453: out = 24'(-7836);
			27454: out = 24'(1924);
			27455: out = 24'(6920);
			27456: out = 24'(8908);
			27457: out = 24'(3612);
			27458: out = 24'(-896);
			27459: out = 24'(-17524);
			27460: out = 24'(-13556);
			27461: out = 24'(2744);
			27462: out = 24'(620);
			27463: out = 24'(-356);
			27464: out = 24'(9712);
			27465: out = 24'(22928);
			27466: out = 24'(18860);
			27467: out = 24'(-5388);
			27468: out = 24'(-12888);
			27469: out = 24'(-1064);
			27470: out = 24'(4712);
			27471: out = 24'(6636);
			27472: out = 24'(1488);
			27473: out = 24'(-332);
			27474: out = 24'(568);
			27475: out = 24'(7252);
			27476: out = 24'(11612);
			27477: out = 24'(11440);
			27478: out = 24'(5672);
			27479: out = 24'(-232);
			27480: out = 24'(-5428);
			27481: out = 24'(-9180);
			27482: out = 24'(-8004);
			27483: out = 24'(1780);
			27484: out = 24'(7052);
			27485: out = 24'(4140);
			27486: out = 24'(-2456);
			27487: out = 24'(-3124);
			27488: out = 24'(-1416);
			27489: out = 24'(-896);
			27490: out = 24'(-9920);
			27491: out = 24'(-20788);
			27492: out = 24'(-3032);
			27493: out = 24'(13876);
			27494: out = 24'(20944);
			27495: out = 24'(11612);
			27496: out = 24'(1572);
			27497: out = 24'(-13084);
			27498: out = 24'(-14056);
			27499: out = 24'(-9212);
			27500: out = 24'(-8740);
			27501: out = 24'(-5504);
			27502: out = 24'(6136);
			27503: out = 24'(13600);
			27504: out = 24'(7604);
			27505: out = 24'(1148);
			27506: out = 24'(3900);
			27507: out = 24'(6588);
			27508: out = 24'(-2272);
			27509: out = 24'(-2596);
			27510: out = 24'(-2084);
			27511: out = 24'(756);
			27512: out = 24'(-952);
			27513: out = 24'(92);
			27514: out = 24'(-5252);
			27515: out = 24'(-3896);
			27516: out = 24'(308);
			27517: out = 24'(-3636);
			27518: out = 24'(-480);
			27519: out = 24'(124);
			27520: out = 24'(200);
			27521: out = 24'(-196);
			27522: out = 24'(2460);
			27523: out = 24'(-3580);
			27524: out = 24'(-8772);
			27525: out = 24'(-1552);
			27526: out = 24'(568);
			27527: out = 24'(7080);
			27528: out = 24'(5396);
			27529: out = 24'(-380);
			27530: out = 24'(-3148);
			27531: out = 24'(332);
			27532: out = 24'(1864);
			27533: out = 24'(16);
			27534: out = 24'(2156);
			27535: out = 24'(6152);
			27536: out = 24'(7216);
			27537: out = 24'(2892);
			27538: out = 24'(-3136);
			27539: out = 24'(-1988);
			27540: out = 24'(2548);
			27541: out = 24'(5384);
			27542: out = 24'(4360);
			27543: out = 24'(744);
			27544: out = 24'(-5540);
			27545: out = 24'(-10904);
			27546: out = 24'(-10848);
			27547: out = 24'(-1256);
			27548: out = 24'(876);
			27549: out = 24'(-528);
			27550: out = 24'(1320);
			27551: out = 24'(6804);
			27552: out = 24'(4804);
			27553: out = 24'(-2796);
			27554: out = 24'(-4440);
			27555: out = 24'(4492);
			27556: out = 24'(7972);
			27557: out = 24'(780);
			27558: out = 24'(-7312);
			27559: out = 24'(-2836);
			27560: out = 24'(444);
			27561: out = 24'(-112);
			27562: out = 24'(-6264);
			27563: out = 24'(-7360);
			27564: out = 24'(4896);
			27565: out = 24'(13836);
			27566: out = 24'(9076);
			27567: out = 24'(-6108);
			27568: out = 24'(-10860);
			27569: out = 24'(-11392);
			27570: out = 24'(-4564);
			27571: out = 24'(132);
			27572: out = 24'(12);
			27573: out = 24'(2920);
			27574: out = 24'(9828);
			27575: out = 24'(10400);
			27576: out = 24'(2092);
			27577: out = 24'(-1432);
			27578: out = 24'(3748);
			27579: out = 24'(6996);
			27580: out = 24'(3684);
			27581: out = 24'(-20716);
			27582: out = 24'(-13132);
			27583: out = 24'(5684);
			27584: out = 24'(3992);
			27585: out = 24'(-14180);
			27586: out = 24'(-21496);
			27587: out = 24'(-7272);
			27588: out = 24'(9924);
			27589: out = 24'(12348);
			27590: out = 24'(5432);
			27591: out = 24'(-1860);
			27592: out = 24'(-2200);
			27593: out = 24'(4800);
			27594: out = 24'(1316);
			27595: out = 24'(-6368);
			27596: out = 24'(-13632);
			27597: out = 24'(-10088);
			27598: out = 24'(3764);
			27599: out = 24'(14664);
			27600: out = 24'(9204);
			27601: out = 24'(-3692);
			27602: out = 24'(1272);
			27603: out = 24'(2040);
			27604: out = 24'(-9196);
			27605: out = 24'(-18456);
			27606: out = 24'(6184);
			27607: out = 24'(14856);
			27608: out = 24'(5344);
			27609: out = 24'(-12004);
			27610: out = 24'(-10924);
			27611: out = 24'(-3232);
			27612: out = 24'(240);
			27613: out = 24'(-4676);
			27614: out = 24'(-1608);
			27615: out = 24'(4964);
			27616: out = 24'(12772);
			27617: out = 24'(7132);
			27618: out = 24'(-7396);
			27619: out = 24'(-14456);
			27620: out = 24'(-4620);
			27621: out = 24'(7068);
			27622: out = 24'(5876);
			27623: out = 24'(-1460);
			27624: out = 24'(-5132);
			27625: out = 24'(2472);
			27626: out = 24'(6828);
			27627: out = 24'(580);
			27628: out = 24'(-5868);
			27629: out = 24'(472);
			27630: out = 24'(7956);
			27631: out = 24'(828);
			27632: out = 24'(-14288);
			27633: out = 24'(-10972);
			27634: out = 24'(9388);
			27635: out = 24'(20004);
			27636: out = 24'(10972);
			27637: out = 24'(-5784);
			27638: out = 24'(-13228);
			27639: out = 24'(-10624);
			27640: out = 24'(1456);
			27641: out = 24'(-1268);
			27642: out = 24'(-2544);
			27643: out = 24'(1848);
			27644: out = 24'(7576);
			27645: out = 24'(7956);
			27646: out = 24'(6852);
			27647: out = 24'(2080);
			27648: out = 24'(-9072);
			27649: out = 24'(-9728);
			27650: out = 24'(-3136);
			27651: out = 24'(2960);
			27652: out = 24'(-704);
			27653: out = 24'(672);
			27654: out = 24'(-2248);
			27655: out = 24'(-2652);
			27656: out = 24'(352);
			27657: out = 24'(7300);
			27658: out = 24'(-280);
			27659: out = 24'(-11736);
			27660: out = 24'(-11300);
			27661: out = 24'(6648);
			27662: out = 24'(7728);
			27663: out = 24'(236);
			27664: out = 24'(-1052);
			27665: out = 24'(7020);
			27666: out = 24'(3036);
			27667: out = 24'(-8212);
			27668: out = 24'(-5708);
			27669: out = 24'(15096);
			27670: out = 24'(2964);
			27671: out = 24'(-10768);
			27672: out = 24'(-7108);
			27673: out = 24'(18108);
			27674: out = 24'(19928);
			27675: out = 24'(8684);
			27676: out = 24'(-7248);
			27677: out = 24'(-7220);
			27678: out = 24'(-3016);
			27679: out = 24'(11872);
			27680: out = 24'(8772);
			27681: out = 24'(-3988);
			27682: out = 24'(-8644);
			27683: out = 24'(836);
			27684: out = 24'(4404);
			27685: out = 24'(-4824);
			27686: out = 24'(-6876);
			27687: out = 24'(84);
			27688: out = 24'(14672);
			27689: out = 24'(160);
			27690: out = 24'(-35480);
			27691: out = 24'(-32348);
			27692: out = 24'(1780);
			27693: out = 24'(23904);
			27694: out = 24'(9920);
			27695: out = 24'(-2796);
			27696: out = 24'(-4368);
			27697: out = 24'(6048);
			27698: out = 24'(2748);
			27699: out = 24'(-18960);
			27700: out = 24'(-20636);
			27701: out = 24'(-4048);
			27702: out = 24'(10764);
			27703: out = 24'(7240);
			27704: out = 24'(6784);
			27705: out = 24'(4728);
			27706: out = 24'(5612);
			27707: out = 24'(76);
			27708: out = 24'(-8424);
			27709: out = 24'(-21208);
			27710: out = 24'(-15808);
			27711: out = 24'(4320);
			27712: out = 24'(21192);
			27713: out = 24'(2596);
			27714: out = 24'(-10596);
			27715: out = 24'(3348);
			27716: out = 24'(17104);
			27717: out = 24'(10196);
			27718: out = 24'(-8616);
			27719: out = 24'(-11104);
			27720: out = 24'(-760);
			27721: out = 24'(8984);
			27722: out = 24'(-4424);
			27723: out = 24'(-12660);
			27724: out = 24'(2156);
			27725: out = 24'(7172);
			27726: out = 24'(2544);
			27727: out = 24'(-5352);
			27728: out = 24'(-4816);
			27729: out = 24'(-780);
			27730: out = 24'(-1844);
			27731: out = 24'(-360);
			27732: out = 24'(7844);
			27733: out = 24'(11996);
			27734: out = 24'(10180);
			27735: out = 24'(2556);
			27736: out = 24'(-5324);
			27737: out = 24'(-8132);
			27738: out = 24'(-5208);
			27739: out = 24'(892);
			27740: out = 24'(68);
			27741: out = 24'(-4676);
			27742: out = 24'(2432);
			27743: out = 24'(19240);
			27744: out = 24'(22140);
			27745: out = 24'(4772);
			27746: out = 24'(-4696);
			27747: out = 24'(-5492);
			27748: out = 24'(-4944);
			27749: out = 24'(-8756);
			27750: out = 24'(2444);
			27751: out = 24'(4676);
			27752: out = 24'(960);
			27753: out = 24'(-8648);
			27754: out = 24'(-10996);
			27755: out = 24'(-6020);
			27756: out = 24'(-292);
			27757: out = 24'(1156);
			27758: out = 24'(8932);
			27759: out = 24'(4688);
			27760: out = 24'(7604);
			27761: out = 24'(3064);
			27762: out = 24'(-9800);
			27763: out = 24'(-9292);
			27764: out = 24'(-444);
			27765: out = 24'(7920);
			27766: out = 24'(5584);
			27767: out = 24'(-4508);
			27768: out = 24'(-9508);
			27769: out = 24'(-4960);
			27770: out = 24'(700);
			27771: out = 24'(188);
			27772: out = 24'(5324);
			27773: out = 24'(12248);
			27774: out = 24'(12128);
			27775: out = 24'(-1528);
			27776: out = 24'(-16696);
			27777: out = 24'(-22172);
			27778: out = 24'(-9908);
			27779: out = 24'(9084);
			27780: out = 24'(12484);
			27781: out = 24'(12788);
			27782: out = 24'(11508);
			27783: out = 24'(3708);
			27784: out = 24'(-23588);
			27785: out = 24'(-32440);
			27786: out = 24'(-17392);
			27787: out = 24'(7220);
			27788: out = 24'(11996);
			27789: out = 24'(14324);
			27790: out = 24'(10184);
			27791: out = 24'(7944);
			27792: out = 24'(7164);
			27793: out = 24'(1808);
			27794: out = 24'(-7696);
			27795: out = 24'(-10004);
			27796: out = 24'(1084);
			27797: out = 24'(-544);
			27798: out = 24'(1956);
			27799: out = 24'(3316);
			27800: out = 24'(6488);
			27801: out = 24'(13516);
			27802: out = 24'(14252);
			27803: out = 24'(6652);
			27804: out = 24'(-1372);
			27805: out = 24'(-1396);
			27806: out = 24'(-516);
			27807: out = 24'(-1448);
			27808: out = 24'(508);
			27809: out = 24'(6572);
			27810: out = 24'(13524);
			27811: out = 24'(6764);
			27812: out = 24'(-3556);
			27813: out = 24'(-3976);
			27814: out = 24'(-2400);
			27815: out = 24'(-4620);
			27816: out = 24'(-5724);
			27817: out = 24'(3384);
			27818: out = 24'(2976);
			27819: out = 24'(6952);
			27820: out = 24'(3644);
			27821: out = 24'(-3092);
			27822: out = 24'(-9740);
			27823: out = 24'(-6284);
			27824: out = 24'(-4480);
			27825: out = 24'(-8592);
			27826: out = 24'(-11316);
			27827: out = 24'(1092);
			27828: out = 24'(20520);
			27829: out = 24'(26680);
			27830: out = 24'(9184);
			27831: out = 24'(-14972);
			27832: out = 24'(-30392);
			27833: out = 24'(-26132);
			27834: out = 24'(-10344);
			27835: out = 24'(3308);
			27836: out = 24'(7640);
			27837: out = 24'(6836);
			27838: out = 24'(4336);
			27839: out = 24'(176);
			27840: out = 24'(-4388);
			27841: out = 24'(-8248);
			27842: out = 24'(-7736);
			27843: out = 24'(-72);
			27844: out = 24'(5880);
			27845: out = 24'(7736);
			27846: out = 24'(2104);
			27847: out = 24'(-5776);
			27848: out = 24'(-7252);
			27849: out = 24'(472);
			27850: out = 24'(4968);
			27851: out = 24'(-1480);
			27852: out = 24'(-2740);
			27853: out = 24'(-1840);
			27854: out = 24'(1476);
			27855: out = 24'(1368);
			27856: out = 24'(-144);
			27857: out = 24'(-3180);
			27858: out = 24'(-1412);
			27859: out = 24'(2416);
			27860: out = 24'(1664);
			27861: out = 24'(-1748);
			27862: out = 24'(-4432);
			27863: out = 24'(-888);
			27864: out = 24'(7664);
			27865: out = 24'(5772);
			27866: out = 24'(5416);
			27867: out = 24'(9288);
			27868: out = 24'(10720);
			27869: out = 24'(2248);
			27870: out = 24'(-12632);
			27871: out = 24'(-16068);
			27872: out = 24'(-580);
			27873: out = 24'(12236);
			27874: out = 24'(11484);
			27875: out = 24'(1980);
			27876: out = 24'(-824);
			27877: out = 24'(-2780);
			27878: out = 24'(2464);
			27879: out = 24'(-5128);
			27880: out = 24'(-11616);
			27881: out = 24'(-1260);
			27882: out = 24'(6048);
			27883: out = 24'(3516);
			27884: out = 24'(-2100);
			27885: out = 24'(680);
			27886: out = 24'(17576);
			27887: out = 24'(13936);
			27888: out = 24'(-5764);
			27889: out = 24'(-20924);
			27890: out = 24'(-11648);
			27891: out = 24'(572);
			27892: out = 24'(4228);
			27893: out = 24'(-1704);
			27894: out = 24'(504);
			27895: out = 24'(3428);
			27896: out = 24'(12352);
			27897: out = 24'(10256);
			27898: out = 24'(-2872);
			27899: out = 24'(-19848);
			27900: out = 24'(-8424);
			27901: out = 24'(11256);
			27902: out = 24'(10084);
			27903: out = 24'(-12888);
			27904: out = 24'(-12436);
			27905: out = 24'(8620);
			27906: out = 24'(15892);
			27907: out = 24'(-2340);
			27908: out = 24'(-15400);
			27909: out = 24'(-9892);
			27910: out = 24'(-1048);
			27911: out = 24'(-11044);
			27912: out = 24'(-5920);
			27913: out = 24'(10500);
			27914: out = 24'(19824);
			27915: out = 24'(4584);
			27916: out = 24'(-10548);
			27917: out = 24'(-15152);
			27918: out = 24'(-5444);
			27919: out = 24'(-1664);
			27920: out = 24'(1880);
			27921: out = 24'(-10804);
			27922: out = 24'(-14928);
			27923: out = 24'(2036);
			27924: out = 24'(17040);
			27925: out = 24'(9900);
			27926: out = 24'(-7236);
			27927: out = 24'(-9444);
			27928: out = 24'(-2568);
			27929: out = 24'(10692);
			27930: out = 24'(7784);
			27931: out = 24'(-920);
			27932: out = 24'(-484);
			27933: out = 24'(4372);
			27934: out = 24'(36);
			27935: out = 24'(-7012);
			27936: out = 24'(-3400);
			27937: out = 24'(-216);
			27938: out = 24'(-7224);
			27939: out = 24'(-15648);
			27940: out = 24'(-6412);
			27941: out = 24'(4632);
			27942: out = 24'(13044);
			27943: out = 24'(9064);
			27944: out = 24'(1848);
			27945: out = 24'(-336);
			27946: out = 24'(-1080);
			27947: out = 24'(-11248);
			27948: out = 24'(-23736);
			27949: out = 24'(-8280);
			27950: out = 24'(2964);
			27951: out = 24'(14084);
			27952: out = 24'(11176);
			27953: out = 24'(-5000);
			27954: out = 24'(-9672);
			27955: out = 24'(100);
			27956: out = 24'(10524);
			27957: out = 24'(12480);
			27958: out = 24'(3952);
			27959: out = 24'(5460);
			27960: out = 24'(5536);
			27961: out = 24'(-5328);
			27962: out = 24'(-16008);
			27963: out = 24'(-7820);
			27964: out = 24'(5912);
			27965: out = 24'(6052);
			27966: out = 24'(1272);
			27967: out = 24'(-1620);
			27968: out = 24'(4612);
			27969: out = 24'(6548);
			27970: out = 24'(2952);
			27971: out = 24'(-7772);
			27972: out = 24'(-1188);
			27973: out = 24'(9080);
			27974: out = 24'(3788);
			27975: out = 24'(-8428);
			27976: out = 24'(-7904);
			27977: out = 24'(6708);
			27978: out = 24'(12800);
			27979: out = 24'(3420);
			27980: out = 24'(-8348);
			27981: out = 24'(-1000);
			27982: out = 24'(15264);
			27983: out = 24'(8032);
			27984: out = 24'(-9612);
			27985: out = 24'(-19320);
			27986: out = 24'(-6084);
			27987: out = 24'(10008);
			27988: out = 24'(11904);
			27989: out = 24'(-3484);
			27990: out = 24'(-7672);
			27991: out = 24'(14728);
			27992: out = 24'(15696);
			27993: out = 24'(2276);
			27994: out = 24'(-12288);
			27995: out = 24'(-7032);
			27996: out = 24'(8056);
			27997: out = 24'(12052);
			27998: out = 24'(-764);
			27999: out = 24'(-11388);
			28000: out = 24'(-2732);
			28001: out = 24'(4728);
			28002: out = 24'(-1672);
			28003: out = 24'(-13576);
			28004: out = 24'(-15048);
			28005: out = 24'(-2428);
			28006: out = 24'(4100);
			28007: out = 24'(928);
			28008: out = 24'(764);
			28009: out = 24'(14276);
			28010: out = 24'(16308);
			28011: out = 24'(-1120);
			28012: out = 24'(-16360);
			28013: out = 24'(-11060);
			28014: out = 24'(8112);
			28015: out = 24'(10484);
			28016: out = 24'(-5744);
			28017: out = 24'(-22056);
			28018: out = 24'(-10808);
			28019: out = 24'(8212);
			28020: out = 24'(13260);
			28021: out = 24'(3168);
			28022: out = 24'(-2744);
			28023: out = 24'(-2660);
			28024: out = 24'(-2168);
			28025: out = 24'(-15252);
			28026: out = 24'(-5876);
			28027: out = 24'(-1408);
			28028: out = 24'(3604);
			28029: out = 24'(14240);
			28030: out = 24'(4168);
			28031: out = 24'(-9792);
			28032: out = 24'(-12164);
			28033: out = 24'(-3696);
			28034: out = 24'(-8812);
			28035: out = 24'(-18996);
			28036: out = 24'(-8696);
			28037: out = 24'(18208);
			28038: out = 24'(22012);
			28039: out = 24'(-4868);
			28040: out = 24'(-24444);
			28041: out = 24'(-10940);
			28042: out = 24'(5664);
			28043: out = 24'(5332);
			28044: out = 24'(-4664);
			28045: out = 24'(-1080);
			28046: out = 24'(12144);
			28047: out = 24'(10928);
			28048: out = 24'(-1444);
			28049: out = 24'(-9196);
			28050: out = 24'(-5032);
			28051: out = 24'(-676);
			28052: out = 24'(5056);
			28053: out = 24'(10928);
			28054: out = 24'(15336);
			28055: out = 24'(14960);
			28056: out = 24'(8668);
			28057: out = 24'(1476);
			28058: out = 24'(-944);
			28059: out = 24'(-1084);
			28060: out = 24'(352);
			28061: out = 24'(-7912);
			28062: out = 24'(-20892);
			28063: out = 24'(-19292);
			28064: out = 24'(-6324);
			28065: out = 24'(13548);
			28066: out = 24'(21116);
			28067: out = 24'(13748);
			28068: out = 24'(-3132);
			28069: out = 24'(-6676);
			28070: out = 24'(-1612);
			28071: out = 24'(-652);
			28072: out = 24'(48);
			28073: out = 24'(-476);
			28074: out = 24'(36);
			28075: out = 24'(-288);
			28076: out = 24'(-212);
			28077: out = 24'(3560);
			28078: out = 24'(2708);
			28079: out = 24'(-6548);
			28080: out = 24'(-10608);
			28081: out = 24'(-13504);
			28082: out = 24'(-2828);
			28083: out = 24'(7804);
			28084: out = 24'(10044);
			28085: out = 24'(1764);
			28086: out = 24'(-1892);
			28087: out = 24'(-5936);
			28088: out = 24'(-12172);
			28089: out = 24'(-17516);
			28090: out = 24'(-6848);
			28091: out = 24'(5388);
			28092: out = 24'(7404);
			28093: out = 24'(740);
			28094: out = 24'(1192);
			28095: out = 24'(3380);
			28096: out = 24'(2400);
			28097: out = 24'(-172);
			28098: out = 24'(1584);
			28099: out = 24'(1460);
			28100: out = 24'(-2436);
			28101: out = 24'(-8504);
			28102: out = 24'(-4440);
			28103: out = 24'(6396);
			28104: out = 24'(20920);
			28105: out = 24'(23204);
			28106: out = 24'(9796);
			28107: out = 24'(-12232);
			28108: out = 24'(-11192);
			28109: out = 24'(9180);
			28110: out = 24'(7660);
			28111: out = 24'(-9860);
			28112: out = 24'(-14788);
			28113: out = 24'(5496);
			28114: out = 24'(12160);
			28115: out = 24'(11828);
			28116: out = 24'(36);
			28117: out = 24'(-2656);
			28118: out = 24'(-1684);
			28119: out = 24'(3272);
			28120: out = 24'(-6248);
			28121: out = 24'(-10252);
			28122: out = 24'(3204);
			28123: out = 24'(12768);
			28124: out = 24'(7372);
			28125: out = 24'(-8276);
			28126: out = 24'(-17796);
			28127: out = 24'(-10880);
			28128: out = 24'(-624);
			28129: out = 24'(2332);
			28130: out = 24'(-692);
			28131: out = 24'(204);
			28132: out = 24'(-2584);
			28133: out = 24'(-4796);
			28134: out = 24'(-6536);
			28135: out = 24'(-5652);
			28136: out = 24'(-1524);
			28137: out = 24'(2488);
			28138: out = 24'(1212);
			28139: out = 24'(-2812);
			28140: out = 24'(-4068);
			28141: out = 24'(6624);
			28142: out = 24'(12476);
			28143: out = 24'(3520);
			28144: out = 24'(840);
			28145: out = 24'(-1184);
			28146: out = 24'(976);
			28147: out = 24'(-968);
			28148: out = 24'(628);
			28149: out = 24'(-7604);
			28150: out = 24'(-4436);
			28151: out = 24'(3124);
			28152: out = 24'(104);
			28153: out = 24'(5996);
			28154: out = 24'(9152);
			28155: out = 24'(3588);
			28156: out = 24'(-9188);
			28157: out = 24'(-19308);
			28158: out = 24'(-13280);
			28159: out = 24'(-1960);
			28160: out = 24'(908);
			28161: out = 24'(12204);
			28162: out = 24'(9472);
			28163: out = 24'(-132);
			28164: out = 24'(-8192);
			28165: out = 24'(-328);
			28166: out = 24'(10828);
			28167: out = 24'(13996);
			28168: out = 24'(4664);
			28169: out = 24'(1076);
			28170: out = 24'(-12236);
			28171: out = 24'(-13352);
			28172: out = 24'(-4852);
			28173: out = 24'(8116);
			28174: out = 24'(1492);
			28175: out = 24'(872);
			28176: out = 24'(2052);
			28177: out = 24'(-272);
			28178: out = 24'(236);
			28179: out = 24'(-368);
			28180: out = 24'(-396);
			28181: out = 24'(728);
			28182: out = 24'(6628);
			28183: out = 24'(6428);
			28184: out = 24'(1444);
			28185: out = 24'(-4860);
			28186: out = 24'(-11132);
			28187: out = 24'(-7536);
			28188: out = 24'(-2720);
			28189: out = 24'(1324);
			28190: out = 24'(2352);
			28191: out = 24'(7216);
			28192: out = 24'(4804);
			28193: out = 24'(3260);
			28194: out = 24'(7508);
			28195: out = 24'(13468);
			28196: out = 24'(684);
			28197: out = 24'(-21208);
			28198: out = 24'(-29124);
			28199: out = 24'(-1584);
			28200: out = 24'(13168);
			28201: out = 24'(9376);
			28202: out = 24'(-120);
			28203: out = 24'(7528);
			28204: out = 24'(7332);
			28205: out = 24'(4644);
			28206: out = 24'(-3980);
			28207: out = 24'(-16152);
			28208: out = 24'(-11860);
			28209: out = 24'(996);
			28210: out = 24'(7484);
			28211: out = 24'(1648);
			28212: out = 24'(-2284);
			28213: out = 24'(-1404);
			28214: out = 24'(632);
			28215: out = 24'(-236);
			28216: out = 24'(-5064);
			28217: out = 24'(-2432);
			28218: out = 24'(-1904);
			28219: out = 24'(-10464);
			28220: out = 24'(-17592);
			28221: out = 24'(-9492);
			28222: out = 24'(6860);
			28223: out = 24'(10716);
			28224: out = 24'(1784);
			28225: out = 24'(-15048);
			28226: out = 24'(-13880);
			28227: out = 24'(-328);
			28228: out = 24'(5336);
			28229: out = 24'(2612);
			28230: out = 24'(156);
			28231: out = 24'(1736);
			28232: out = 24'(-516);
			28233: out = 24'(-13036);
			28234: out = 24'(-16660);
			28235: out = 24'(-2344);
			28236: out = 24'(17720);
			28237: out = 24'(19056);
			28238: out = 24'(10992);
			28239: out = 24'(2004);
			28240: out = 24'(1368);
			28241: out = 24'(-408);
			28242: out = 24'(-340);
			28243: out = 24'(-7672);
			28244: out = 24'(-7044);
			28245: out = 24'(8184);
			28246: out = 24'(14716);
			28247: out = 24'(7492);
			28248: out = 24'(-1124);
			28249: out = 24'(1148);
			28250: out = 24'(4596);
			28251: out = 24'(1040);
			28252: out = 24'(-3380);
			28253: out = 24'(2044);
			28254: out = 24'(6156);
			28255: out = 24'(5876);
			28256: out = 24'(-2748);
			28257: out = 24'(-7864);
			28258: out = 24'(-3604);
			28259: out = 24'(104);
			28260: out = 24'(-248);
			28261: out = 24'(552);
			28262: out = 24'(1704);
			28263: out = 24'(11052);
			28264: out = 24'(6608);
			28265: out = 24'(-2140);
			28266: out = 24'(-2272);
			28267: out = 24'(5372);
			28268: out = 24'(4544);
			28269: out = 24'(-5600);
			28270: out = 24'(-14264);
			28271: out = 24'(-14544);
			28272: out = 24'(-5256);
			28273: out = 24'(6624);
			28274: out = 24'(15656);
			28275: out = 24'(18024);
			28276: out = 24'(9492);
			28277: out = 24'(-2244);
			28278: out = 24'(-10436);
			28279: out = 24'(-14244);
			28280: out = 24'(-10212);
			28281: out = 24'(-5432);
			28282: out = 24'(-1844);
			28283: out = 24'(452);
			28284: out = 24'(204);
			28285: out = 24'(4340);
			28286: out = 24'(8196);
			28287: out = 24'(3320);
			28288: out = 24'(-5708);
			28289: out = 24'(-11892);
			28290: out = 24'(-6448);
			28291: out = 24'(1176);
			28292: out = 24'(8180);
			28293: out = 24'(1960);
			28294: out = 24'(3132);
			28295: out = 24'(7796);
			28296: out = 24'(7700);
			28297: out = 24'(-7212);
			28298: out = 24'(-7480);
			28299: out = 24'(1956);
			28300: out = 24'(-808);
			28301: out = 24'(16);
			28302: out = 24'(3292);
			28303: out = 24'(8680);
			28304: out = 24'(5848);
			28305: out = 24'(-1372);
			28306: out = 24'(-4744);
			28307: out = 24'(-1532);
			28308: out = 24'(-756);
			28309: out = 24'(-2544);
			28310: out = 24'(-4072);
			28311: out = 24'(-640);
			28312: out = 24'(3252);
			28313: out = 24'(7140);
			28314: out = 24'(-4152);
			28315: out = 24'(-10768);
			28316: out = 24'(-5884);
			28317: out = 24'(-744);
			28318: out = 24'(1040);
			28319: out = 24'(-5684);
			28320: out = 24'(-5948);
			28321: out = 24'(3356);
			28322: out = 24'(22512);
			28323: out = 24'(12060);
			28324: out = 24'(-8068);
			28325: out = 24'(-12192);
			28326: out = 24'(-2544);
			28327: out = 24'(296);
			28328: out = 24'(-10096);
			28329: out = 24'(-14644);
			28330: out = 24'(-1040);
			28331: out = 24'(19348);
			28332: out = 24'(21468);
			28333: out = 24'(6224);
			28334: out = 24'(-7644);
			28335: out = 24'(-8024);
			28336: out = 24'(-3732);
			28337: out = 24'(-3908);
			28338: out = 24'(-2172);
			28339: out = 24'(620);
			28340: out = 24'(9244);
			28341: out = 24'(8948);
			28342: out = 24'(-1384);
			28343: out = 24'(-5292);
			28344: out = 24'(-3140);
			28345: out = 24'(180);
			28346: out = 24'(-2292);
			28347: out = 24'(-10428);
			28348: out = 24'(-6604);
			28349: out = 24'(2640);
			28350: out = 24'(7064);
			28351: out = 24'(0);
			28352: out = 24'(3800);
			28353: out = 24'(4296);
			28354: out = 24'(-928);
			28355: out = 24'(-8628);
			28356: out = 24'(-8920);
			28357: out = 24'(-2760);
			28358: out = 24'(7196);
			28359: out = 24'(14008);
			28360: out = 24'(12608);
			28361: out = 24'(8168);
			28362: out = 24'(6980);
			28363: out = 24'(4864);
			28364: out = 24'(-5084);
			28365: out = 24'(-21016);
			28366: out = 24'(-23268);
			28367: out = 24'(-4400);
			28368: out = 24'(16584);
			28369: out = 24'(20144);
			28370: out = 24'(8904);
			28371: out = 24'(-4184);
			28372: out = 24'(-11404);
			28373: out = 24'(-5588);
			28374: out = 24'(-2420);
			28375: out = 24'(-6576);
			28376: out = 24'(-13780);
			28377: out = 24'(-1936);
			28378: out = 24'(5216);
			28379: out = 24'(9356);
			28380: out = 24'(11668);
			28381: out = 24'(4820);
			28382: out = 24'(1816);
			28383: out = 24'(-5316);
			28384: out = 24'(-10844);
			28385: out = 24'(-308);
			28386: out = 24'(-3820);
			28387: out = 24'(-9356);
			28388: out = 24'(-8096);
			28389: out = 24'(7892);
			28390: out = 24'(7652);
			28391: out = 24'(3864);
			28392: out = 24'(-1260);
			28393: out = 24'(536);
			28394: out = 24'(-3684);
			28395: out = 24'(-796);
			28396: out = 24'(-1068);
			28397: out = 24'(-2892);
			28398: out = 24'(-4056);
			28399: out = 24'(8508);
			28400: out = 24'(15100);
			28401: out = 24'(9268);
			28402: out = 24'(408);
			28403: out = 24'(2180);
			28404: out = 24'(4340);
			28405: out = 24'(-2040);
			28406: out = 24'(-10724);
			28407: out = 24'(-4196);
			28408: out = 24'(7440);
			28409: out = 24'(8736);
			28410: out = 24'(-4384);
			28411: out = 24'(-5808);
			28412: out = 24'(-5076);
			28413: out = 24'(-3008);
			28414: out = 24'(-3396);
			28415: out = 24'(-232);
			28416: out = 24'(4012);
			28417: out = 24'(8592);
			28418: out = 24'(4780);
			28419: out = 24'(-1680);
			28420: out = 24'(-5912);
			28421: out = 24'(7196);
			28422: out = 24'(20032);
			28423: out = 24'(10780);
			28424: out = 24'(-8528);
			28425: out = 24'(-15180);
			28426: out = 24'(-4868);
			28427: out = 24'(1004);
			28428: out = 24'(4992);
			28429: out = 24'(2292);
			28430: out = 24'(3320);
			28431: out = 24'(6464);
			28432: out = 24'(6912);
			28433: out = 24'(1796);
			28434: out = 24'(-1044);
			28435: out = 24'(1060);
			28436: out = 24'(-4196);
			28437: out = 24'(-7412);
			28438: out = 24'(-8444);
			28439: out = 24'(-1780);
			28440: out = 24'(-2044);
			28441: out = 24'(4868);
			28442: out = 24'(-2360);
			28443: out = 24'(-7784);
			28444: out = 24'(1300);
			28445: out = 24'(15640);
			28446: out = 24'(9084);
			28447: out = 24'(-3512);
			28448: out = 24'(-372);
			28449: out = 24'(3000);
			28450: out = 24'(-3972);
			28451: out = 24'(-16568);
			28452: out = 24'(-14520);
			28453: out = 24'(3336);
			28454: out = 24'(16060);
			28455: out = 24'(13900);
			28456: out = 24'(4408);
			28457: out = 24'(-3404);
			28458: out = 24'(-10088);
			28459: out = 24'(-12804);
			28460: out = 24'(-10960);
			28461: out = 24'(-9052);
			28462: out = 24'(-4536);
			28463: out = 24'(-1384);
			28464: out = 24'(304);
			28465: out = 24'(-172);
			28466: out = 24'(2068);
			28467: out = 24'(2380);
			28468: out = 24'(476);
			28469: out = 24'(-4220);
			28470: out = 24'(-10096);
			28471: out = 24'(-7780);
			28472: out = 24'(3748);
			28473: out = 24'(11108);
			28474: out = 24'(1240);
			28475: out = 24'(-4768);
			28476: out = 24'(-5688);
			28477: out = 24'(-5996);
			28478: out = 24'(-2096);
			28479: out = 24'(-6184);
			28480: out = 24'(244);
			28481: out = 24'(5148);
			28482: out = 24'(3148);
			28483: out = 24'(-7320);
			28484: out = 24'(2328);
			28485: out = 24'(14508);
			28486: out = 24'(10044);
			28487: out = 24'(-7792);
			28488: out = 24'(-9776);
			28489: out = 24'(-2628);
			28490: out = 24'(1016);
			28491: out = 24'(10844);
			28492: out = 24'(14336);
			28493: out = 24'(9332);
			28494: out = 24'(852);
			28495: out = 24'(-1480);
			28496: out = 24'(-536);
			28497: out = 24'(-6700);
			28498: out = 24'(-9268);
			28499: out = 24'(7284);
			28500: out = 24'(16264);
			28501: out = 24'(12720);
			28502: out = 24'(3524);
			28503: out = 24'(-1228);
			28504: out = 24'(1324);
			28505: out = 24'(-7448);
			28506: out = 24'(-9672);
			28507: out = 24'(4252);
			28508: out = 24'(15820);
			28509: out = 24'(7660);
			28510: out = 24'(-2492);
			28511: out = 24'(532);
			28512: out = 24'(4944);
			28513: out = 24'(1328);
			28514: out = 24'(-3000);
			28515: out = 24'(-1692);
			28516: out = 24'(-5248);
			28517: out = 24'(3972);
			28518: out = 24'(6892);
			28519: out = 24'(2248);
			28520: out = 24'(-10464);
			28521: out = 24'(-5536);
			28522: out = 24'(-1564);
			28523: out = 24'(1324);
			28524: out = 24'(1080);
			28525: out = 24'(824);
			28526: out = 24'(-908);
			28527: out = 24'(-3204);
			28528: out = 24'(-3512);
			28529: out = 24'(3220);
			28530: out = 24'(10848);
			28531: out = 24'(8468);
			28532: out = 24'(-6408);
			28533: out = 24'(-16600);
			28534: out = 24'(-18220);
			28535: out = 24'(-6560);
			28536: out = 24'(-1520);
			28537: out = 24'(-6040);
			28538: out = 24'(-9888);
			28539: out = 24'(3976);
			28540: out = 24'(16176);
			28541: out = 24'(11704);
			28542: out = 24'(552);
			28543: out = 24'(-1112);
			28544: out = 24'(1244);
			28545: out = 24'(-1560);
			28546: out = 24'(1424);
			28547: out = 24'(3900);
			28548: out = 24'(10136);
			28549: out = 24'(11116);
			28550: out = 24'(-2012);
			28551: out = 24'(-8064);
			28552: out = 24'(-9948);
			28553: out = 24'(-4448);
			28554: out = 24'(-224);
			28555: out = 24'(1124);
			28556: out = 24'(-11448);
			28557: out = 24'(-14308);
			28558: out = 24'(4132);
			28559: out = 24'(15700);
			28560: out = 24'(6516);
			28561: out = 24'(-12032);
			28562: out = 24'(-15984);
			28563: out = 24'(-8680);
			28564: out = 24'(-948);
			28565: out = 24'(-4840);
			28566: out = 24'(-6688);
			28567: out = 24'(6552);
			28568: out = 24'(9912);
			28569: out = 24'(3324);
			28570: out = 24'(-3172);
			28571: out = 24'(7680);
			28572: out = 24'(72);
			28573: out = 24'(-5420);
			28574: out = 24'(-9204);
			28575: out = 24'(-2260);
			28576: out = 24'(-7512);
			28577: out = 24'(5196);
			28578: out = 24'(13640);
			28579: out = 24'(12384);
			28580: out = 24'(-3164);
			28581: out = 24'(2840);
			28582: out = 24'(5272);
			28583: out = 24'(-5312);
			28584: out = 24'(-28332);
			28585: out = 24'(-10496);
			28586: out = 24'(8224);
			28587: out = 24'(10740);
			28588: out = 24'(7432);
			28589: out = 24'(6636);
			28590: out = 24'(3736);
			28591: out = 24'(-4196);
			28592: out = 24'(-11544);
			28593: out = 24'(-14472);
			28594: out = 24'(-6976);
			28595: out = 24'(3828);
			28596: out = 24'(6648);
			28597: out = 24'(8524);
			28598: out = 24'(-3808);
			28599: out = 24'(-6932);
			28600: out = 24'(1844);
			28601: out = 24'(6508);
			28602: out = 24'(2100);
			28603: out = 24'(-52);
			28604: out = 24'(1688);
			28605: out = 24'(-6360);
			28606: out = 24'(-1704);
			28607: out = 24'(3704);
			28608: out = 24'(6596);
			28609: out = 24'(576);
			28610: out = 24'(-7172);
			28611: out = 24'(-5676);
			28612: out = 24'(3560);
			28613: out = 24'(5596);
			28614: out = 24'(1544);
			28615: out = 24'(-2676);
			28616: out = 24'(7492);
			28617: out = 24'(19304);
			28618: out = 24'(7424);
			28619: out = 24'(-1628);
			28620: out = 24'(-3916);
			28621: out = 24'(-1284);
			28622: out = 24'(-840);
			28623: out = 24'(-9672);
			28624: out = 24'(-9584);
			28625: out = 24'(-1440);
			28626: out = 24'(684);
			28627: out = 24'(-328);
			28628: out = 24'(1084);
			28629: out = 24'(5692);
			28630: out = 24'(2780);
			28631: out = 24'(1240);
			28632: out = 24'(-14560);
			28633: out = 24'(-26768);
			28634: out = 24'(-21400);
			28635: out = 24'(10856);
			28636: out = 24'(19428);
			28637: out = 24'(13244);
			28638: out = 24'(6784);
			28639: out = 24'(8740);
			28640: out = 24'(2732);
			28641: out = 24'(-8084);
			28642: out = 24'(-15064);
			28643: out = 24'(-11352);
			28644: out = 24'(-2300);
			28645: out = 24'(-2052);
			28646: out = 24'(-6508);
			28647: out = 24'(-1864);
			28648: out = 24'(488);
			28649: out = 24'(-864);
			28650: out = 24'(-10264);
			28651: out = 24'(-11436);
			28652: out = 24'(-2596);
			28653: out = 24'(16320);
			28654: out = 24'(14396);
			28655: out = 24'(-4820);
			28656: out = 24'(-21044);
			28657: out = 24'(-2236);
			28658: out = 24'(13700);
			28659: out = 24'(8236);
			28660: out = 24'(-1856);
			28661: out = 24'(-12664);
			28662: out = 24'(-11428);
			28663: out = 24'(-5140);
			28664: out = 24'(4144);
			28665: out = 24'(12416);
			28666: out = 24'(18120);
			28667: out = 24'(15392);
			28668: out = 24'(4464);
			28669: out = 24'(-19152);
			28670: out = 24'(-23624);
			28671: out = 24'(-11024);
			28672: out = 24'(3872);
			28673: out = 24'(7660);
			28674: out = 24'(7228);
			28675: out = 24'(11980);
			28676: out = 24'(18816);
			28677: out = 24'(12812);
			28678: out = 24'(-2312);
			28679: out = 24'(-18588);
			28680: out = 24'(-20624);
			28681: out = 24'(-8260);
			28682: out = 24'(2980);
			28683: out = 24'(10308);
			28684: out = 24'(16652);
			28685: out = 24'(16124);
			28686: out = 24'(3204);
			28687: out = 24'(-14344);
			28688: out = 24'(-17688);
			28689: out = 24'(-7908);
			28690: out = 24'(-10856);
			28691: out = 24'(-10408);
			28692: out = 24'(2716);
			28693: out = 24'(20784);
			28694: out = 24'(13160);
			28695: out = 24'(364);
			28696: out = 24'(-8380);
			28697: out = 24'(2384);
			28698: out = 24'(12124);
			28699: out = 24'(16576);
			28700: out = 24'(-2236);
			28701: out = 24'(-15648);
			28702: out = 24'(-6984);
			28703: out = 24'(10884);
			28704: out = 24'(7372);
			28705: out = 24'(-5608);
			28706: out = 24'(-7592);
			28707: out = 24'(-4988);
			28708: out = 24'(-296);
			28709: out = 24'(-1024);
			28710: out = 24'(1924);
			28711: out = 24'(10356);
			28712: out = 24'(10068);
			28713: out = 24'(-4788);
			28714: out = 24'(-17028);
			28715: out = 24'(296);
			28716: out = 24'(8448);
			28717: out = 24'(9216);
			28718: out = 24'(-6784);
			28719: out = 24'(-21492);
			28720: out = 24'(-15812);
			28721: out = 24'(5952);
			28722: out = 24'(11552);
			28723: out = 24'(-968);
			28724: out = 24'(-552);
			28725: out = 24'(5664);
			28726: out = 24'(388);
			28727: out = 24'(-15696);
			28728: out = 24'(-8140);
			28729: out = 24'(7316);
			28730: out = 24'(16472);
			28731: out = 24'(7140);
			28732: out = 24'(-4592);
			28733: out = 24'(-14024);
			28734: out = 24'(-7524);
			28735: out = 24'(3168);
			28736: out = 24'(6892);
			28737: out = 24'(3456);
			28738: out = 24'(24);
			28739: out = 24'(444);
			28740: out = 24'(-1268);
			28741: out = 24'(-6648);
			28742: out = 24'(-7488);
			28743: out = 24'(4940);
			28744: out = 24'(13084);
			28745: out = 24'(9280);
			28746: out = 24'(-13304);
			28747: out = 24'(-13808);
			28748: out = 24'(2512);
			28749: out = 24'(-620);
			28750: out = 24'(-8236);
			28751: out = 24'(-7060);
			28752: out = 24'(2356);
			28753: out = 24'(-596);
			28754: out = 24'(736);
			28755: out = 24'(3712);
			28756: out = 24'(8368);
			28757: out = 24'(3736);
			28758: out = 24'(-1344);
			28759: out = 24'(-4704);
			28760: out = 24'(2828);
			28761: out = 24'(15344);
			28762: out = 24'(11044);
			28763: out = 24'(4764);
			28764: out = 24'(-7144);
			28765: out = 24'(-10468);
			28766: out = 24'(-10440);
			28767: out = 24'(14784);
			28768: out = 24'(13656);
			28769: out = 24'(-3996);
			28770: out = 24'(-17212);
			28771: out = 24'(-1484);
			28772: out = 24'(-5340);
			28773: out = 24'(-15872);
			28774: out = 24'(-9008);
			28775: out = 24'(11092);
			28776: out = 24'(7996);
			28777: out = 24'(-3384);
			28778: out = 24'(-1544);
			28779: out = 24'(-884);
			28780: out = 24'(3732);
			28781: out = 24'(6548);
			28782: out = 24'(5220);
			28783: out = 24'(-7272);
			28784: out = 24'(-14184);
			28785: out = 24'(-4448);
			28786: out = 24'(8460);
			28787: out = 24'(-508);
			28788: out = 24'(-4388);
			28789: out = 24'(356);
			28790: out = 24'(8648);
			28791: out = 24'(856);
			28792: out = 24'(-3328);
			28793: out = 24'(-4464);
			28794: out = 24'(6120);
			28795: out = 24'(13472);
			28796: out = 24'(8640);
			28797: out = 24'(1236);
			28798: out = 24'(-304);
			28799: out = 24'(-980);
			28800: out = 24'(328);
			28801: out = 24'(-10960);
			28802: out = 24'(-11452);
			28803: out = 24'(1244);
			28804: out = 24'(13336);
			28805: out = 24'(9592);
			28806: out = 24'(2596);
			28807: out = 24'(-756);
			28808: out = 24'(-344);
			28809: out = 24'(3688);
			28810: out = 24'(2556);
			28811: out = 24'(-3144);
			28812: out = 24'(-6180);
			28813: out = 24'(-14436);
			28814: out = 24'(-4520);
			28815: out = 24'(5352);
			28816: out = 24'(6776);
			28817: out = 24'(2072);
			28818: out = 24'(788);
			28819: out = 24'(-2940);
			28820: out = 24'(-5352);
			28821: out = 24'(-380);
			28822: out = 24'(6080);
			28823: out = 24'(3664);
			28824: out = 24'(-248);
			28825: out = 24'(7796);
			28826: out = 24'(15984);
			28827: out = 24'(9592);
			28828: out = 24'(-8284);
			28829: out = 24'(-15956);
			28830: out = 24'(-4180);
			28831: out = 24'(2212);
			28832: out = 24'(-8152);
			28833: out = 24'(-18440);
			28834: out = 24'(-2336);
			28835: out = 24'(6796);
			28836: out = 24'(2912);
			28837: out = 24'(-3028);
			28838: out = 24'(-504);
			28839: out = 24'(11560);
			28840: out = 24'(6440);
			28841: out = 24'(-10912);
			28842: out = 24'(-15568);
			28843: out = 24'(-4772);
			28844: out = 24'(6404);
			28845: out = 24'(4616);
			28846: out = 24'(-3424);
			28847: out = 24'(-9844);
			28848: out = 24'(-8100);
			28849: out = 24'(-1408);
			28850: out = 24'(5504);
			28851: out = 24'(296);
			28852: out = 24'(6184);
			28853: out = 24'(9900);
			28854: out = 24'(5180);
			28855: out = 24'(2900);
			28856: out = 24'(-1156);
			28857: out = 24'(5268);
			28858: out = 24'(10724);
			28859: out = 24'(6160);
			28860: out = 24'(-13852);
			28861: out = 24'(-19160);
			28862: out = 24'(-9124);
			28863: out = 24'(-1212);
			28864: out = 24'(-6216);
			28865: out = 24'(-3700);
			28866: out = 24'(7840);
			28867: out = 24'(12652);
			28868: out = 24'(8904);
			28869: out = 24'(-6572);
			28870: out = 24'(-14396);
			28871: out = 24'(-6712);
			28872: out = 24'(12256);
			28873: out = 24'(14844);
			28874: out = 24'(10264);
			28875: out = 24'(6004);
			28876: out = 24'(4260);
			28877: out = 24'(828);
			28878: out = 24'(-5300);
			28879: out = 24'(-15600);
			28880: out = 24'(-26940);
			28881: out = 24'(-14384);
			28882: out = 24'(932);
			28883: out = 24'(8860);
			28884: out = 24'(7196);
			28885: out = 24'(11504);
			28886: out = 24'(7848);
			28887: out = 24'(748);
			28888: out = 24'(-5908);
			28889: out = 24'(-3068);
			28890: out = 24'(-888);
			28891: out = 24'(460);
			28892: out = 24'(-196);
			28893: out = 24'(408);
			28894: out = 24'(4648);
			28895: out = 24'(10240);
			28896: out = 24'(8376);
			28897: out = 24'(-3872);
			28898: out = 24'(-20480);
			28899: out = 24'(-23900);
			28900: out = 24'(-11560);
			28901: out = 24'(3912);
			28902: out = 24'(16544);
			28903: out = 24'(16116);
			28904: out = 24'(11016);
			28905: out = 24'(5468);
			28906: out = 24'(-4420);
			28907: out = 24'(-11636);
			28908: out = 24'(-11308);
			28909: out = 24'(-4372);
			28910: out = 24'(-8420);
			28911: out = 24'(3764);
			28912: out = 24'(8456);
			28913: out = 24'(6628);
			28914: out = 24'(7228);
			28915: out = 24'(1384);
			28916: out = 24'(-4124);
			28917: out = 24'(-10220);
			28918: out = 24'(-12784);
			28919: out = 24'(-13640);
			28920: out = 24'(-3140);
			28921: out = 24'(13372);
			28922: out = 24'(24576);
			28923: out = 24'(6800);
			28924: out = 24'(-896);
			28925: out = 24'(-5096);
			28926: out = 24'(-9976);
			28927: out = 24'(-23104);
			28928: out = 24'(-14172);
			28929: out = 24'(3648);
			28930: out = 24'(14624);
			28931: out = 24'(7068);
			28932: out = 24'(7820);
			28933: out = 24'(6008);
			28934: out = 24'(4440);
			28935: out = 24'(2388);
			28936: out = 24'(8500);
			28937: out = 24'(4668);
			28938: out = 24'(-3444);
			28939: out = 24'(-7728);
			28940: out = 24'(-3988);
			28941: out = 24'(684);
			28942: out = 24'(2120);
			28943: out = 24'(-64);
			28944: out = 24'(7216);
			28945: out = 24'(-168);
			28946: out = 24'(-2200);
			28947: out = 24'(2916);
			28948: out = 24'(4056);
			28949: out = 24'(2440);
			28950: out = 24'(2944);
			28951: out = 24'(9784);
			28952: out = 24'(17876);
			28953: out = 24'(7460);
			28954: out = 24'(-6896);
			28955: out = 24'(-17372);
			28956: out = 24'(-18864);
			28957: out = 24'(-17796);
			28958: out = 24'(-6636);
			28959: out = 24'(3840);
			28960: out = 24'(6272);
			28961: out = 24'(676);
			28962: out = 24'(-360);
			28963: out = 24'(-840);
			28964: out = 24'(-3488);
			28965: out = 24'(-216);
			28966: out = 24'(784);
			28967: out = 24'(1548);
			28968: out = 24'(-1452);
			28969: out = 24'(948);
			28970: out = 24'(-9548);
			28971: out = 24'(-5836);
			28972: out = 24'(2356);
			28973: out = 24'(7308);
			28974: out = 24'(696);
			28975: out = 24'(-2080);
			28976: out = 24'(-12228);
			28977: out = 24'(-22880);
			28978: out = 24'(-5332);
			28979: out = 24'(10664);
			28980: out = 24'(9844);
			28981: out = 24'(-1048);
			28982: out = 24'(304);
			28983: out = 24'(6440);
			28984: out = 24'(-712);
			28985: out = 24'(-14292);
			28986: out = 24'(-3660);
			28987: out = 24'(4180);
			28988: out = 24'(8404);
			28989: out = 24'(1768);
			28990: out = 24'(-4664);
			28991: out = 24'(-5676);
			28992: out = 24'(-3352);
			28993: out = 24'(-312);
			28994: out = 24'(6408);
			28995: out = 24'(6824);
			28996: out = 24'(8040);
			28997: out = 24'(6072);
			28998: out = 24'(4804);
			28999: out = 24'(2284);
			29000: out = 24'(704);
			29001: out = 24'(-2236);
			29002: out = 24'(-2172);
			29003: out = 24'(-156);
			29004: out = 24'(5776);
			29005: out = 24'(7236);
			29006: out = 24'(6952);
			29007: out = 24'(6316);
			29008: out = 24'(3416);
			29009: out = 24'(-4276);
			29010: out = 24'(-8748);
			29011: out = 24'(-5432);
			29012: out = 24'(-5868);
			29013: out = 24'(-4532);
			29014: out = 24'(572);
			29015: out = 24'(8216);
			29016: out = 24'(10624);
			29017: out = 24'(11296);
			29018: out = 24'(9208);
			29019: out = 24'(4400);
			29020: out = 24'(-960);
			29021: out = 24'(-11904);
			29022: out = 24'(-10588);
			29023: out = 24'(-1168);
			29024: out = 24'(-1020);
			29025: out = 24'(5940);
			29026: out = 24'(6504);
			29027: out = 24'(5384);
			29028: out = 24'(684);
			29029: out = 24'(6396);
			29030: out = 24'(176);
			29031: out = 24'(-5796);
			29032: out = 24'(-5076);
			29033: out = 24'(5432);
			29034: out = 24'(2220);
			29035: out = 24'(-4168);
			29036: out = 24'(-4068);
			29037: out = 24'(10264);
			29038: out = 24'(10956);
			29039: out = 24'(4372);
			29040: out = 24'(-7844);
			29041: out = 24'(-10272);
			29042: out = 24'(-13648);
			29043: out = 24'(-740);
			29044: out = 24'(5652);
			29045: out = 24'(-1088);
			29046: out = 24'(-8372);
			29047: out = 24'(256);
			29048: out = 24'(6592);
			29049: out = 24'(-1372);
			29050: out = 24'(-20148);
			29051: out = 24'(-8048);
			29052: out = 24'(9884);
			29053: out = 24'(10008);
			29054: out = 24'(-7144);
			29055: out = 24'(-9348);
			29056: out = 24'(-7948);
			29057: out = 24'(-6680);
			29058: out = 24'(2904);
			29059: out = 24'(2344);
			29060: out = 24'(1212);
			29061: out = 24'(-872);
			29062: out = 24'(108);
			29063: out = 24'(-4792);
			29064: out = 24'(-4708);
			29065: out = 24'(-28);
			29066: out = 24'(4620);
			29067: out = 24'(856);
			29068: out = 24'(-5444);
			29069: out = 24'(-6880);
			29070: out = 24'(-2592);
			29071: out = 24'(-7788);
			29072: out = 24'(-11448);
			29073: out = 24'(-8624);
			29074: out = 24'(6260);
			29075: out = 24'(18228);
			29076: out = 24'(12456);
			29077: out = 24'(-3892);
			29078: out = 24'(-8076);
			29079: out = 24'(2888);
			29080: out = 24'(16256);
			29081: out = 24'(5876);
			29082: out = 24'(-11456);
			29083: out = 24'(-14032);
			29084: out = 24'(4064);
			29085: out = 24'(7784);
			29086: out = 24'(480);
			29087: out = 24'(-5312);
			29088: out = 24'(-3172);
			29089: out = 24'(-576);
			29090: out = 24'(2300);
			29091: out = 24'(5632);
			29092: out = 24'(7064);
			29093: out = 24'(1800);
			29094: out = 24'(204);
			29095: out = 24'(2144);
			29096: out = 24'(-616);
			29097: out = 24'(-2160);
			29098: out = 24'(-3860);
			29099: out = 24'(-1364);
			29100: out = 24'(2256);
			29101: out = 24'(-2316);
			29102: out = 24'(800);
			29103: out = 24'(8212);
			29104: out = 24'(9200);
			29105: out = 24'(-6236);
			29106: out = 24'(-9964);
			29107: out = 24'(-3952);
			29108: out = 24'(-1376);
			29109: out = 24'(-9532);
			29110: out = 24'(-4428);
			29111: out = 24'(10944);
			29112: out = 24'(17976);
			29113: out = 24'(6636);
			29114: out = 24'(-1796);
			29115: out = 24'(-1900);
			29116: out = 24'(-1936);
			29117: out = 24'(-8788);
			29118: out = 24'(-17980);
			29119: out = 24'(-7600);
			29120: out = 24'(6188);
			29121: out = 24'(6880);
			29122: out = 24'(13564);
			29123: out = 24'(13472);
			29124: out = 24'(8944);
			29125: out = 24'(-3592);
			29126: out = 24'(-9448);
			29127: out = 24'(-18144);
			29128: out = 24'(-11660);
			29129: out = 24'(5224);
			29130: out = 24'(16108);
			29131: out = 24'(12388);
			29132: out = 24'(2424);
			29133: out = 24'(1044);
			29134: out = 24'(2604);
			29135: out = 24'(-4512);
			29136: out = 24'(-22256);
			29137: out = 24'(-19448);
			29138: out = 24'(9832);
			29139: out = 24'(12524);
			29140: out = 24'(5320);
			29141: out = 24'(-2648);
			29142: out = 24'(1480);
			29143: out = 24'(5740);
			29144: out = 24'(-2624);
			29145: out = 24'(-11952);
			29146: out = 24'(-7792);
			29147: out = 24'(1288);
			29148: out = 24'(1828);
			29149: out = 24'(-2712);
			29150: out = 24'(-480);
			29151: out = 24'(6608);
			29152: out = 24'(9708);
			29153: out = 24'(-336);
			29154: out = 24'(-10476);
			29155: out = 24'(-6896);
			29156: out = 24'(-4640);
			29157: out = 24'(-3084);
			29158: out = 24'(-9344);
			29159: out = 24'(-11276);
			29160: out = 24'(-1392);
			29161: out = 24'(11364);
			29162: out = 24'(9420);
			29163: out = 24'(-3024);
			29164: out = 24'(-15164);
			29165: out = 24'(-4080);
			29166: out = 24'(1244);
			29167: out = 24'(-5132);
			29168: out = 24'(-8856);
			29169: out = 24'(3564);
			29170: out = 24'(12292);
			29171: out = 24'(8548);
			29172: out = 24'(400);
			29173: out = 24'(-160);
			29174: out = 24'(3628);
			29175: out = 24'(3196);
			29176: out = 24'(-3512);
			29177: out = 24'(200);
			29178: out = 24'(-2320);
			29179: out = 24'(-1464);
			29180: out = 24'(1248);
			29181: out = 24'(7404);
			29182: out = 24'(2008);
			29183: out = 24'(520);
			29184: out = 24'(1940);
			29185: out = 24'(340);
			29186: out = 24'(1420);
			29187: out = 24'(8220);
			29188: out = 24'(14468);
			29189: out = 24'(11992);
			29190: out = 24'(1840);
			29191: out = 24'(-4720);
			29192: out = 24'(-5652);
			29193: out = 24'(-3412);
			29194: out = 24'(-6148);
			29195: out = 24'(-3796);
			29196: out = 24'(-5132);
			29197: out = 24'(-6880);
			29198: out = 24'(4064);
			29199: out = 24'(11760);
			29200: out = 24'(8564);
			29201: out = 24'(-2812);
			29202: out = 24'(-2320);
			29203: out = 24'(-8176);
			29204: out = 24'(-8100);
			29205: out = 24'(-7760);
			29206: out = 24'(-1716);
			29207: out = 24'(2492);
			29208: out = 24'(11408);
			29209: out = 24'(9828);
			29210: out = 24'(-1596);
			29211: out = 24'(-9892);
			29212: out = 24'(-9688);
			29213: out = 24'(-6252);
			29214: out = 24'(-1744);
			29215: out = 24'(-656);
			29216: out = 24'(10652);
			29217: out = 24'(9308);
			29218: out = 24'(-3656);
			29219: out = 24'(-12592);
			29220: out = 24'(-4132);
			29221: out = 24'(136);
			29222: out = 24'(-4640);
			29223: out = 24'(-3892);
			29224: out = 24'(2336);
			29225: out = 24'(11304);
			29226: out = 24'(12788);
			29227: out = 24'(8492);
			29228: out = 24'(908);
			29229: out = 24'(-768);
			29230: out = 24'(36);
			29231: out = 24'(-972);
			29232: out = 24'(-5108);
			29233: out = 24'(-4952);
			29234: out = 24'(1300);
			29235: out = 24'(8328);
			29236: out = 24'(13136);
			29237: out = 24'(8184);
			29238: out = 24'(5884);
			29239: out = 24'(5064);
			29240: out = 24'(-1528);
			29241: out = 24'(-11376);
			29242: out = 24'(-14344);
			29243: out = 24'(-7540);
			29244: out = 24'(308);
			29245: out = 24'(9832);
			29246: out = 24'(14872);
			29247: out = 24'(15988);
			29248: out = 24'(7484);
			29249: out = 24'(-3816);
			29250: out = 24'(-17604);
			29251: out = 24'(-12204);
			29252: out = 24'(3480);
			29253: out = 24'(-1296);
			29254: out = 24'(-2332);
			29255: out = 24'(-2964);
			29256: out = 24'(1088);
			29257: out = 24'(3828);
			29258: out = 24'(6208);
			29259: out = 24'(6304);
			29260: out = 24'(5364);
			29261: out = 24'(548);
			29262: out = 24'(-4596);
			29263: out = 24'(-12056);
			29264: out = 24'(-10348);
			29265: out = 24'(3204);
			29266: out = 24'(2980);
			29267: out = 24'(3664);
			29268: out = 24'(-2732);
			29269: out = 24'(-4976);
			29270: out = 24'(-1692);
			29271: out = 24'(1392);
			29272: out = 24'(-9376);
			29273: out = 24'(-17148);
			29274: out = 24'(-452);
			29275: out = 24'(11356);
			29276: out = 24'(7552);
			29277: out = 24'(-2640);
			29278: out = 24'(620);
			29279: out = 24'(-544);
			29280: out = 24'(-6924);
			29281: out = 24'(-15860);
			29282: out = 24'(-10976);
			29283: out = 24'(-2344);
			29284: out = 24'(3820);
			29285: out = 24'(-176);
			29286: out = 24'(-1572);
			29287: out = 24'(-816);
			29288: out = 24'(6964);
			29289: out = 24'(-776);
			29290: out = 24'(-14952);
			29291: out = 24'(-12068);
			29292: out = 24'(-2920);
			29293: out = 24'(2404);
			29294: out = 24'(-184);
			29295: out = 24'(1612);
			29296: out = 24'(-2440);
			29297: out = 24'(-104);
			29298: out = 24'(768);
			29299: out = 24'(1260);
			29300: out = 24'(64);
			29301: out = 24'(8132);
			29302: out = 24'(11164);
			29303: out = 24'(3028);
			29304: out = 24'(-1352);
			29305: out = 24'(-8800);
			29306: out = 24'(-9612);
			29307: out = 24'(-7628);
			29308: out = 24'(-9692);
			29309: out = 24'(-2956);
			29310: out = 24'(7968);
			29311: out = 24'(15544);
			29312: out = 24'(13376);
			29313: out = 24'(3212);
			29314: out = 24'(-3080);
			29315: out = 24'(-1112);
			29316: out = 24'(-100);
			29317: out = 24'(1148);
			29318: out = 24'(-484);
			29319: out = 24'(1864);
			29320: out = 24'(960);
			29321: out = 24'(-1040);
			29322: out = 24'(180);
			29323: out = 24'(15504);
			29324: out = 24'(21564);
			29325: out = 24'(2052);
			29326: out = 24'(-26816);
			29327: out = 24'(-20932);
			29328: out = 24'(9944);
			29329: out = 24'(15496);
			29330: out = 24'(10816);
			29331: out = 24'(5104);
			29332: out = 24'(6676);
			29333: out = 24'(-2164);
			29334: out = 24'(-1256);
			29335: out = 24'(-9312);
			29336: out = 24'(-7376);
			29337: out = 24'(2212);
			29338: out = 24'(160);
			29339: out = 24'(784);
			29340: out = 24'(6700);
			29341: out = 24'(12628);
			29342: out = 24'(-296);
			29343: out = 24'(-7532);
			29344: out = 24'(-11960);
			29345: out = 24'(-4396);
			29346: out = 24'(2828);
			29347: out = 24'(5308);
			29348: out = 24'(-7692);
			29349: out = 24'(-7900);
			29350: out = 24'(13640);
			29351: out = 24'(20092);
			29352: out = 24'(-2952);
			29353: out = 24'(-28372);
			29354: out = 24'(-23996);
			29355: out = 24'(-1940);
			29356: out = 24'(3988);
			29357: out = 24'(-1752);
			29358: out = 24'(2648);
			29359: out = 24'(3256);
			29360: out = 24'(8608);
			29361: out = 24'(492);
			29362: out = 24'(-8424);
			29363: out = 24'(-7784);
			29364: out = 24'(4104);
			29365: out = 24'(6528);
			29366: out = 24'(-784);
			29367: out = 24'(-6824);
			29368: out = 24'(4024);
			29369: out = 24'(10360);
			29370: out = 24'(6316);
			29371: out = 24'(4);
			29372: out = 24'(-7528);
			29373: out = 24'(-2308);
			29374: out = 24'(4132);
			29375: out = 24'(4148);
			29376: out = 24'(628);
			29377: out = 24'(-3420);
			29378: out = 24'(-8928);
			29379: out = 24'(-12092);
			29380: out = 24'(344);
			29381: out = 24'(336);
			29382: out = 24'(548);
			29383: out = 24'(112);
			29384: out = 24'(428);
			29385: out = 24'(-6188);
			29386: out = 24'(-4604);
			29387: out = 24'(5048);
			29388: out = 24'(12996);
			29389: out = 24'(2864);
			29390: out = 24'(-10596);
			29391: out = 24'(-13388);
			29392: out = 24'(-376);
			29393: out = 24'(-700);
			29394: out = 24'(6140);
			29395: out = 24'(6860);
			29396: out = 24'(4520);
			29397: out = 24'(-2864);
			29398: out = 24'(-2140);
			29399: out = 24'(-4500);
			29400: out = 24'(-3612);
			29401: out = 24'(-352);
			29402: out = 24'(7512);
			29403: out = 24'(-1296);
			29404: out = 24'(-10352);
			29405: out = 24'(-1080);
			29406: out = 24'(14888);
			29407: out = 24'(12456);
			29408: out = 24'(1156);
			29409: out = 24'(1404);
			29410: out = 24'(5500);
			29411: out = 24'(2144);
			29412: out = 24'(-7936);
			29413: out = 24'(-9400);
			29414: out = 24'(-4400);
			29415: out = 24'(5116);
			29416: out = 24'(6524);
			29417: out = 24'(3900);
			29418: out = 24'(-204);
			29419: out = 24'(5468);
			29420: out = 24'(4400);
			29421: out = 24'(-3036);
			29422: out = 24'(-7488);
			29423: out = 24'(-4848);
			29424: out = 24'(3068);
			29425: out = 24'(9288);
			29426: out = 24'(13252);
			29427: out = 24'(4984);
			29428: out = 24'(4336);
			29429: out = 24'(1752);
			29430: out = 24'(-4920);
			29431: out = 24'(-10904);
			29432: out = 24'(-4208);
			29433: out = 24'(1032);
			29434: out = 24'(-1200);
			29435: out = 24'(500);
			29436: out = 24'(3988);
			29437: out = 24'(10132);
			29438: out = 24'(7728);
			29439: out = 24'(-3692);
			29440: out = 24'(-12788);
			29441: out = 24'(-9164);
			29442: out = 24'(-1148);
			29443: out = 24'(-616);
			29444: out = 24'(2148);
			29445: out = 24'(4536);
			29446: out = 24'(7084);
			29447: out = 24'(2372);
			29448: out = 24'(-1672);
			29449: out = 24'(-15556);
			29450: out = 24'(-12924);
			29451: out = 24'(5220);
			29452: out = 24'(5172);
			29453: out = 24'(3016);
			29454: out = 24'(-6472);
			29455: out = 24'(-4768);
			29456: out = 24'(5808);
			29457: out = 24'(8848);
			29458: out = 24'(-7160);
			29459: out = 24'(-20148);
			29460: out = 24'(-11776);
			29461: out = 24'(-1812);
			29462: out = 24'(-308);
			29463: out = 24'(-2672);
			29464: out = 24'(1968);
			29465: out = 24'(6440);
			29466: out = 24'(3676);
			29467: out = 24'(-1188);
			29468: out = 24'(2252);
			29469: out = 24'(6040);
			29470: out = 24'(12);
			29471: out = 24'(-13372);
			29472: out = 24'(-15016);
			29473: out = 24'(220);
			29474: out = 24'(7396);
			29475: out = 24'(2584);
			29476: out = 24'(-2588);
			29477: out = 24'(1404);
			29478: out = 24'(12336);
			29479: out = 24'(4760);
			29480: out = 24'(-12600);
			29481: out = 24'(-20212);
			29482: out = 24'(-17084);
			29483: out = 24'(-4300);
			29484: out = 24'(4728);
			29485: out = 24'(8400);
			29486: out = 24'(7708);
			29487: out = 24'(8180);
			29488: out = 24'(3876);
			29489: out = 24'(-5804);
			29490: out = 24'(-14568);
			29491: out = 24'(-6732);
			29492: out = 24'(7904);
			29493: out = 24'(12532);
			29494: out = 24'(-68);
			29495: out = 24'(232);
			29496: out = 24'(3812);
			29497: out = 24'(9020);
			29498: out = 24'(5196);
			29499: out = 24'(-9584);
			29500: out = 24'(-15688);
			29501: out = 24'(-2932);
			29502: out = 24'(12740);
			29503: out = 24'(5832);
			29504: out = 24'(-348);
			29505: out = 24'(-1532);
			29506: out = 24'(652);
			29507: out = 24'(-2344);
			29508: out = 24'(-6500);
			29509: out = 24'(-4200);
			29510: out = 24'(1288);
			29511: out = 24'(-160);
			29512: out = 24'(1096);
			29513: out = 24'(3836);
			29514: out = 24'(11932);
			29515: out = 24'(19120);
			29516: out = 24'(6940);
			29517: out = 24'(-3132);
			29518: out = 24'(-10992);
			29519: out = 24'(-14576);
			29520: out = 24'(-10172);
			29521: out = 24'(-4428);
			29522: out = 24'(1012);
			29523: out = 24'(7028);
			29524: out = 24'(10484);
			29525: out = 24'(5024);
			29526: out = 24'(-10384);
			29527: out = 24'(-19216);
			29528: out = 24'(-9008);
			29529: out = 24'(-3048);
			29530: out = 24'(-624);
			29531: out = 24'(6092);
			29532: out = 24'(19036);
			29533: out = 24'(9884);
			29534: out = 24'(-6428);
			29535: out = 24'(-13924);
			29536: out = 24'(-1864);
			29537: out = 24'(5804);
			29538: out = 24'(4408);
			29539: out = 24'(-1024);
			29540: out = 24'(3248);
			29541: out = 24'(9876);
			29542: out = 24'(12900);
			29543: out = 24'(3760);
			29544: out = 24'(-7796);
			29545: out = 24'(-14692);
			29546: out = 24'(-9052);
			29547: out = 24'(-2880);
			29548: out = 24'(3536);
			29549: out = 24'(9456);
			29550: out = 24'(13420);
			29551: out = 24'(4936);
			29552: out = 24'(-6548);
			29553: out = 24'(-8016);
			29554: out = 24'(4860);
			29555: out = 24'(6220);
			29556: out = 24'(-3764);
			29557: out = 24'(-11832);
			29558: out = 24'(-5384);
			29559: out = 24'(4096);
			29560: out = 24'(8940);
			29561: out = 24'(7864);
			29562: out = 24'(288);
			29563: out = 24'(3776);
			29564: out = 24'(3100);
			29565: out = 24'(-2344);
			29566: out = 24'(-9692);
			29567: out = 24'(-212);
			29568: out = 24'(4488);
			29569: out = 24'(3652);
			29570: out = 24'(-56);
			29571: out = 24'(2596);
			29572: out = 24'(640);
			29573: out = 24'(1012);
			29574: out = 24'(76);
			29575: out = 24'(-13304);
			29576: out = 24'(-17164);
			29577: out = 24'(-3924);
			29578: out = 24'(13856);
			29579: out = 24'(12464);
			29580: out = 24'(2088);
			29581: out = 24'(-4564);
			29582: out = 24'(-1012);
			29583: out = 24'(-752);
			29584: out = 24'(-7004);
			29585: out = 24'(-10700);
			29586: out = 24'(-1644);
			29587: out = 24'(8808);
			29588: out = 24'(8504);
			29589: out = 24'(-872);
			29590: out = 24'(-4936);
			29591: out = 24'(-1724);
			29592: out = 24'(6860);
			29593: out = 24'(-3860);
			29594: out = 24'(-10064);
			29595: out = 24'(-1948);
			29596: out = 24'(3692);
			29597: out = 24'(4444);
			29598: out = 24'(636);
			29599: out = 24'(2152);
			29600: out = 24'(6360);
			29601: out = 24'(7912);
			29602: out = 24'(-348);
			29603: out = 24'(-10160);
			29604: out = 24'(-11680);
			29605: out = 24'(-6428);
			29606: out = 24'(-224);
			29607: out = 24'(4708);
			29608: out = 24'(9724);
			29609: out = 24'(6624);
			29610: out = 24'(7392);
			29611: out = 24'(4176);
			29612: out = 24'(-1072);
			29613: out = 24'(-7524);
			29614: out = 24'(-7368);
			29615: out = 24'(-8808);
			29616: out = 24'(-7956);
			29617: out = 24'(440);
			29618: out = 24'(9356);
			29619: out = 24'(7140);
			29620: out = 24'(-3568);
			29621: out = 24'(-9164);
			29622: out = 24'(-12724);
			29623: out = 24'(-5336);
			29624: out = 24'(5584);
			29625: out = 24'(13708);
			29626: out = 24'(13452);
			29627: out = 24'(6616);
			29628: out = 24'(-2560);
			29629: out = 24'(-6880);
			29630: out = 24'(1336);
			29631: out = 24'(1140);
			29632: out = 24'(-428);
			29633: out = 24'(192);
			29634: out = 24'(1776);
			29635: out = 24'(5708);
			29636: out = 24'(7096);
			29637: out = 24'(5132);
			29638: out = 24'(-328);
			29639: out = 24'(1692);
			29640: out = 24'(-68);
			29641: out = 24'(-6972);
			29642: out = 24'(-15640);
			29643: out = 24'(-13132);
			29644: out = 24'(-3844);
			29645: out = 24'(8016);
			29646: out = 24'(12280);
			29647: out = 24'(7832);
			29648: out = 24'(-208);
			29649: out = 24'(-6652);
			29650: out = 24'(-15164);
			29651: out = 24'(-18576);
			29652: out = 24'(-24160);
			29653: out = 24'(-7676);
			29654: out = 24'(15172);
			29655: out = 24'(20164);
			29656: out = 24'(13968);
			29657: out = 24'(7448);
			29658: out = 24'(1620);
			29659: out = 24'(-7892);
			29660: out = 24'(-7488);
			29661: out = 24'(-1456);
			29662: out = 24'(5140);
			29663: out = 24'(7056);
			29664: out = 24'(6828);
			29665: out = 24'(6152);
			29666: out = 24'(-952);
			29667: out = 24'(-11184);
			29668: out = 24'(-9696);
			29669: out = 24'(-960);
			29670: out = 24'(3064);
			29671: out = 24'(-620);
			29672: out = 24'(1344);
			29673: out = 24'(7868);
			29674: out = 24'(13908);
			29675: out = 24'(8524);
			29676: out = 24'(-2856);
			29677: out = 24'(724);
			29678: out = 24'(3124);
			29679: out = 24'(-3404);
			29680: out = 24'(-12296);
			29681: out = 24'(-100);
			29682: out = 24'(8564);
			29683: out = 24'(9740);
			29684: out = 24'(4740);
			29685: out = 24'(-5040);
			29686: out = 24'(804);
			29687: out = 24'(5620);
			29688: out = 24'(204);
			29689: out = 24'(-17656);
			29690: out = 24'(-10744);
			29691: out = 24'(-4228);
			29692: out = 24'(-2076);
			29693: out = 24'(1428);
			29694: out = 24'(15160);
			29695: out = 24'(17752);
			29696: out = 24'(4756);
			29697: out = 24'(-11824);
			29698: out = 24'(-30392);
			29699: out = 24'(-14496);
			29700: out = 24'(10932);
			29701: out = 24'(16548);
			29702: out = 24'(9048);
			29703: out = 24'(1160);
			29704: out = 24'(9812);
			29705: out = 24'(16448);
			29706: out = 24'(4208);
			29707: out = 24'(-19560);
			29708: out = 24'(-24692);
			29709: out = 24'(-9948);
			29710: out = 24'(-1500);
			29711: out = 24'(-900);
			29712: out = 24'(-5168);
			29713: out = 24'(-1372);
			29714: out = 24'(7596);
			29715: out = 24'(6932);
			29716: out = 24'(3392);
			29717: out = 24'(-3056);
			29718: out = 24'(-7524);
			29719: out = 24'(-10092);
			29720: out = 24'(-1680);
			29721: out = 24'(4996);
			29722: out = 24'(8908);
			29723: out = 24'(18052);
			29724: out = 24'(10828);
			29725: out = 24'(-2608);
			29726: out = 24'(-10388);
			29727: out = 24'(-5200);
			29728: out = 24'(776);
			29729: out = 24'(-2672);
			29730: out = 24'(-7824);
			29731: out = 24'(-776);
			29732: out = 24'(10196);
			29733: out = 24'(13748);
			29734: out = 24'(3528);
			29735: out = 24'(-11056);
			29736: out = 24'(-5496);
			29737: out = 24'(-3832);
			29738: out = 24'(-1692);
			29739: out = 24'(276);
			29740: out = 24'(6892);
			29741: out = 24'(4836);
			29742: out = 24'(3064);
			29743: out = 24'(-3412);
			29744: out = 24'(-11796);
			29745: out = 24'(-16348);
			29746: out = 24'(-6848);
			29747: out = 24'(-336);
			29748: out = 24'(-4088);
			29749: out = 24'(548);
			29750: out = 24'(14724);
			29751: out = 24'(16188);
			29752: out = 24'(-2120);
			29753: out = 24'(-4360);
			29754: out = 24'(-1052);
			29755: out = 24'(-1008);
			29756: out = 24'(-12944);
			29757: out = 24'(-18688);
			29758: out = 24'(-7120);
			29759: out = 24'(8400);
			29760: out = 24'(9128);
			29761: out = 24'(1604);
			29762: out = 24'(-496);
			29763: out = 24'(2700);
			29764: out = 24'(1096);
			29765: out = 24'(-1608);
			29766: out = 24'(-5592);
			29767: out = 24'(5688);
			29768: out = 24'(15100);
			29769: out = 24'(10936);
			29770: out = 24'(-4712);
			29771: out = 24'(-6556);
			29772: out = 24'(2124);
			29773: out = 24'(5260);
			29774: out = 24'(-6112);
			29775: out = 24'(-7316);
			29776: out = 24'(716);
			29777: out = 24'(6824);
			29778: out = 24'(2568);
			29779: out = 24'(5052);
			29780: out = 24'(10316);
			29781: out = 24'(10768);
			29782: out = 24'(760);
			29783: out = 24'(-22760);
			29784: out = 24'(-28788);
			29785: out = 24'(-7956);
			29786: out = 24'(17652);
			29787: out = 24'(22656);
			29788: out = 24'(9096);
			29789: out = 24'(-6316);
			29790: out = 24'(-11884);
			29791: out = 24'(-848);
			29792: out = 24'(-1460);
			29793: out = 24'(-1724);
			29794: out = 24'(3096);
			29795: out = 24'(4056);
			29796: out = 24'(1660);
			29797: out = 24'(-976);
			29798: out = 24'(1356);
			29799: out = 24'(3980);
			29800: out = 24'(10044);
			29801: out = 24'(5520);
			29802: out = 24'(-4544);
			29803: out = 24'(-12284);
			29804: out = 24'(-2584);
			29805: out = 24'(4864);
			29806: out = 24'(4148);
			29807: out = 24'(-4000);
			29808: out = 24'(-2668);
			29809: out = 24'(-1584);
			29810: out = 24'(520);
			29811: out = 24'(-204);
			29812: out = 24'(6960);
			29813: out = 24'(1000);
			29814: out = 24'(-208);
			29815: out = 24'(-948);
			29816: out = 24'(648);
			29817: out = 24'(1412);
			29818: out = 24'(10368);
			29819: out = 24'(5824);
			29820: out = 24'(-15804);
			29821: out = 24'(-24288);
			29822: out = 24'(-6460);
			29823: out = 24'(8028);
			29824: out = 24'(-2516);
			29825: out = 24'(-17584);
			29826: out = 24'(-9656);
			29827: out = 24'(5112);
			29828: out = 24'(3200);
			29829: out = 24'(1844);
			29830: out = 24'(-496);
			29831: out = 24'(1256);
			29832: out = 24'(-832);
			29833: out = 24'(-4316);
			29834: out = 24'(-1688);
			29835: out = 24'(-124);
			29836: out = 24'(-4056);
			29837: out = 24'(-6244);
			29838: out = 24'(-1220);
			29839: out = 24'(1872);
			29840: out = 24'(-2936);
			29841: out = 24'(-8636);
			29842: out = 24'(-3660);
			29843: out = 24'(5900);
			29844: out = 24'(9224);
			29845: out = 24'(3904);
			29846: out = 24'(1280);
			29847: out = 24'(-3464);
			29848: out = 24'(-3604);
			29849: out = 24'(2248);
			29850: out = 24'(10548);
			29851: out = 24'(9188);
			29852: out = 24'(-24);
			29853: out = 24'(-8364);
			29854: out = 24'(-4468);
			29855: out = 24'(-880);
			29856: out = 24'(-1292);
			29857: out = 24'(-6468);
			29858: out = 24'(-2892);
			29859: out = 24'(4024);
			29860: out = 24'(16120);
			29861: out = 24'(15120);
			29862: out = 24'(6404);
			29863: out = 24'(7656);
			29864: out = 24'(12292);
			29865: out = 24'(6336);
			29866: out = 24'(-4268);
			29867: out = 24'(-992);
			29868: out = 24'(9312);
			29869: out = 24'(5688);
			29870: out = 24'(-10776);
			29871: out = 24'(-16760);
			29872: out = 24'(4256);
			29873: out = 24'(19184);
			29874: out = 24'(9896);
			29875: out = 24'(-11044);
			29876: out = 24'(-5772);
			29877: out = 24'(-732);
			29878: out = 24'(-4084);
			29879: out = 24'(-10696);
			29880: out = 24'(-4528);
			29881: out = 24'(3376);
			29882: out = 24'(4968);
			29883: out = 24'(-3544);
			29884: out = 24'(-14024);
			29885: out = 24'(-7076);
			29886: out = 24'(10700);
			29887: out = 24'(14424);
			29888: out = 24'(-4956);
			29889: out = 24'(-17164);
			29890: out = 24'(-6620);
			29891: out = 24'(8588);
			29892: out = 24'(488);
			29893: out = 24'(556);
			29894: out = 24'(5264);
			29895: out = 24'(15444);
			29896: out = 24'(9016);
			29897: out = 24'(4692);
			29898: out = 24'(-13944);
			29899: out = 24'(-15540);
			29900: out = 24'(-7424);
			29901: out = 24'(524);
			29902: out = 24'(-12024);
			29903: out = 24'(-10348);
			29904: out = 24'(2232);
			29905: out = 24'(8892);
			29906: out = 24'(-10020);
			29907: out = 24'(-9164);
			29908: out = 24'(8004);
			29909: out = 24'(13572);
			29910: out = 24'(-1156);
			29911: out = 24'(-4592);
			29912: out = 24'(592);
			29913: out = 24'(-3948);
			29914: out = 24'(712);
			29915: out = 24'(-1868);
			29916: out = 24'(-3696);
			29917: out = 24'(-4108);
			29918: out = 24'(6044);
			29919: out = 24'(3484);
			29920: out = 24'(-7920);
			29921: out = 24'(-16712);
			29922: out = 24'(-2452);
			29923: out = 24'(9760);
			29924: out = 24'(11004);
			29925: out = 24'(2212);
			29926: out = 24'(3080);
			29927: out = 24'(1196);
			29928: out = 24'(1160);
			29929: out = 24'(-7752);
			29930: out = 24'(-13752);
			29931: out = 24'(-5868);
			29932: out = 24'(11348);
			29933: out = 24'(14836);
			29934: out = 24'(5232);
			29935: out = 24'(-2260);
			29936: out = 24'(352);
			29937: out = 24'(-2060);
			29938: out = 24'(-12296);
			29939: out = 24'(-16736);
			29940: out = 24'(-116);
			29941: out = 24'(12040);
			29942: out = 24'(8104);
			29943: out = 24'(744);
			29944: out = 24'(7992);
			29945: out = 24'(10900);
			29946: out = 24'(1492);
			29947: out = 24'(-7512);
			29948: out = 24'(-22340);
			29949: out = 24'(-11800);
			29950: out = 24'(2848);
			29951: out = 24'(7156);
			29952: out = 24'(7128);
			29953: out = 24'(10884);
			29954: out = 24'(11708);
			29955: out = 24'(4116);
			29956: out = 24'(-1700);
			29957: out = 24'(-2976);
			29958: out = 24'(5948);
			29959: out = 24'(12380);
			29960: out = 24'(5716);
			29961: out = 24'(1084);
			29962: out = 24'(-1424);
			29963: out = 24'(308);
			29964: out = 24'(628);
			29965: out = 24'(-2408);
			29966: out = 24'(-2100);
			29967: out = 24'(5568);
			29968: out = 24'(11492);
			29969: out = 24'(7212);
			29970: out = 24'(-1428);
			29971: out = 24'(-940);
			29972: out = 24'(5784);
			29973: out = 24'(-880);
			29974: out = 24'(-4964);
			29975: out = 24'(-4500);
			29976: out = 24'(-564);
			29977: out = 24'(-3868);
			29978: out = 24'(-1740);
			29979: out = 24'(5320);
			29980: out = 24'(13576);
			29981: out = 24'(10284);
			29982: out = 24'(3672);
			29983: out = 24'(-7412);
			29984: out = 24'(-11156);
			29985: out = 24'(-8396);
			29986: out = 24'(-4040);
			29987: out = 24'(-2292);
			29988: out = 24'(3708);
			29989: out = 24'(13796);
			29990: out = 24'(21672);
			29991: out = 24'(12172);
			29992: out = 24'(-6216);
			29993: out = 24'(-19888);
			29994: out = 24'(-10928);
			29995: out = 24'(-8260);
			29996: out = 24'(-2640);
			29997: out = 24'(-1508);
			29998: out = 24'(-2956);
			29999: out = 24'(-2328);
			30000: out = 24'(4040);
			30001: out = 24'(2844);
			30002: out = 24'(-5812);
			30003: out = 24'(-5024);
			30004: out = 24'(2468);
			30005: out = 24'(-2732);
			30006: out = 24'(-19032);
			30007: out = 24'(-13856);
			30008: out = 24'(1956);
			30009: out = 24'(7584);
			30010: out = 24'(-3124);
			30011: out = 24'(-9052);
			30012: out = 24'(-2360);
			30013: out = 24'(1800);
			30014: out = 24'(-6680);
			30015: out = 24'(-13816);
			30016: out = 24'(-4176);
			30017: out = 24'(6904);
			30018: out = 24'(8224);
			30019: out = 24'(6792);
			30020: out = 24'(-8040);
			30021: out = 24'(-7968);
			30022: out = 24'(-3508);
			30023: out = 24'(-2668);
			30024: out = 24'(-2220);
			30025: out = 24'(-1112);
			30026: out = 24'(572);
			30027: out = 24'(1228);
			30028: out = 24'(9168);
			30029: out = 24'(7316);
			30030: out = 24'(8664);
			30031: out = 24'(10084);
			30032: out = 24'(3748);
			30033: out = 24'(-10324);
			30034: out = 24'(-20436);
			30035: out = 24'(-15512);
			30036: out = 24'(1260);
			30037: out = 24'(11248);
			30038: out = 24'(14088);
			30039: out = 24'(10924);
			30040: out = 24'(5888);
			30041: out = 24'(460);
			30042: out = 24'(-3612);
			30043: out = 24'(-6920);
			30044: out = 24'(-6960);
			30045: out = 24'(-592);
			30046: out = 24'(416);
			30047: out = 24'(-552);
			30048: out = 24'(2204);
			30049: out = 24'(12280);
			30050: out = 24'(11724);
			30051: out = 24'(5092);
			30052: out = 24'(-2160);
			30053: out = 24'(-2608);
			30054: out = 24'(3788);
			30055: out = 24'(10596);
			30056: out = 24'(9136);
			30057: out = 24'(-1836);
			30058: out = 24'(1452);
			30059: out = 24'(-5012);
			30060: out = 24'(-9520);
			30061: out = 24'(-7468);
			30062: out = 24'(-4072);
			30063: out = 24'(3188);
			30064: out = 24'(9392);
			30065: out = 24'(11700);
			30066: out = 24'(7736);
			30067: out = 24'(1520);
			30068: out = 24'(-5232);
			30069: out = 24'(-8368);
			30070: out = 24'(-3408);
			30071: out = 24'(-1656);
			30072: out = 24'(-184);
			30073: out = 24'(-1416);
			30074: out = 24'(-292);
			30075: out = 24'(-4160);
			30076: out = 24'(2444);
			30077: out = 24'(5892);
			30078: out = 24'(2448);
			30079: out = 24'(-7832);
			30080: out = 24'(404);
			30081: out = 24'(7656);
			30082: out = 24'(3660);
			30083: out = 24'(-2792);
			30084: out = 24'(-2732);
			30085: out = 24'(2712);
			30086: out = 24'(4868);
			30087: out = 24'(-1368);
			30088: out = 24'(-1020);
			30089: out = 24'(-5240);
			30090: out = 24'(-9408);
			30091: out = 24'(-8196);
			30092: out = 24'(-6360);
			30093: out = 24'(-4368);
			30094: out = 24'(-2168);
			30095: out = 24'(-380);
			30096: out = 24'(-268);
			30097: out = 24'(564);
			30098: out = 24'(1536);
			30099: out = 24'(-2456);
			30100: out = 24'(-8828);
			30101: out = 24'(-12768);
			30102: out = 24'(3208);
			30103: out = 24'(22376);
			30104: out = 24'(16504);
			30105: out = 24'(-5076);
			30106: out = 24'(-19540);
			30107: out = 24'(-13604);
			30108: out = 24'(-3832);
			30109: out = 24'(-1708);
			30110: out = 24'(-6460);
			30111: out = 24'(-5312);
			30112: out = 24'(1264);
			30113: out = 24'(12140);
			30114: out = 24'(7016);
			30115: out = 24'(-44);
			30116: out = 24'(1416);
			30117: out = 24'(7476);
			30118: out = 24'(3944);
			30119: out = 24'(-7944);
			30120: out = 24'(-14228);
			30121: out = 24'(-688);
			30122: out = 24'(6744);
			30123: out = 24'(8568);
			30124: out = 24'(4860);
			30125: out = 24'(2188);
			30126: out = 24'(-440);
			30127: out = 24'(16);
			30128: out = 24'(-2500);
			30129: out = 24'(-8080);
			30130: out = 24'(-6152);
			30131: out = 24'(2024);
			30132: out = 24'(5984);
			30133: out = 24'(-1960);
			30134: out = 24'(1088);
			30135: out = 24'(-272);
			30136: out = 24'(5372);
			30137: out = 24'(3212);
			30138: out = 24'(-6156);
			30139: out = 24'(-21796);
			30140: out = 24'(-13344);
			30141: out = 24'(3616);
			30142: out = 24'(6464);
			30143: out = 24'(-3100);
			30144: out = 24'(604);
			30145: out = 24'(6972);
			30146: out = 24'(-1468);
			30147: out = 24'(-10464);
			30148: out = 24'(-5404);
			30149: out = 24'(8540);
			30150: out = 24'(10692);
			30151: out = 24'(-7452);
			30152: out = 24'(-10268);
			30153: out = 24'(-2640);
			30154: out = 24'(616);
			30155: out = 24'(-11768);
			30156: out = 24'(-4228);
			30157: out = 24'(3996);
			30158: out = 24'(3604);
			30159: out = 24'(-1968);
			30160: out = 24'(848);
			30161: out = 24'(4356);
			30162: out = 24'(5348);
			30163: out = 24'(7016);
			30164: out = 24'(1084);
			30165: out = 24'(-1388);
			30166: out = 24'(-4336);
			30167: out = 24'(-7128);
			30168: out = 24'(-2964);
			30169: out = 24'(4904);
			30170: out = 24'(12084);
			30171: out = 24'(11252);
			30172: out = 24'(3480);
			30173: out = 24'(-2504);
			30174: out = 24'(1228);
			30175: out = 24'(6364);
			30176: out = 24'(-544);
			30177: out = 24'(-7824);
			30178: out = 24'(-7360);
			30179: out = 24'(4940);
			30180: out = 24'(13628);
			30181: out = 24'(9088);
			30182: out = 24'(-2808);
			30183: out = 24'(-8764);
			30184: out = 24'(-8272);
			30185: out = 24'(-9532);
			30186: out = 24'(-11220);
			30187: out = 24'(-2860);
			30188: out = 24'(9284);
			30189: out = 24'(4528);
			30190: out = 24'(-3424);
			30191: out = 24'(-7604);
			30192: out = 24'(-2704);
			30193: out = 24'(1864);
			30194: out = 24'(4576);
			30195: out = 24'(2432);
			30196: out = 24'(-412);
			30197: out = 24'(480);
			30198: out = 24'(-412);
			30199: out = 24'(944);
			30200: out = 24'(-5040);
			30201: out = 24'(-16824);
			30202: out = 24'(-14924);
			30203: out = 24'(-920);
			30204: out = 24'(8944);
			30205: out = 24'(2900);
			30206: out = 24'(-328);
			30207: out = 24'(-1748);
			30208: out = 24'(5260);
			30209: out = 24'(7580);
			30210: out = 24'(1364);
			30211: out = 24'(-2308);
			30212: out = 24'(-200);
			30213: out = 24'(-1060);
			30214: out = 24'(-5988);
			30215: out = 24'(-9780);
			30216: out = 24'(1860);
			30217: out = 24'(12052);
			30218: out = 24'(5160);
			30219: out = 24'(-4256);
			30220: out = 24'(-4068);
			30221: out = 24'(4340);
			30222: out = 24'(5116);
			30223: out = 24'(-2500);
			30224: out = 24'(-4748);
			30225: out = 24'(2580);
			30226: out = 24'(5780);
			30227: out = 24'(3652);
			30228: out = 24'(-10528);
			30229: out = 24'(-8612);
			30230: out = 24'(6388);
			30231: out = 24'(11212);
			30232: out = 24'(3960);
			30233: out = 24'(-7836);
			30234: out = 24'(-9420);
			30235: out = 24'(328);
			30236: out = 24'(-1884);
			30237: out = 24'(-1016);
			30238: out = 24'(3316);
			30239: out = 24'(8748);
			30240: out = 24'(3008);
			30241: out = 24'(1000);
			30242: out = 24'(0);
			30243: out = 24'(1056);
			30244: out = 24'(3964);
			30245: out = 24'(3652);
			30246: out = 24'(-3964);
			30247: out = 24'(-13820);
			30248: out = 24'(-18012);
			30249: out = 24'(-6572);
			30250: out = 24'(4436);
			30251: out = 24'(5996);
			30252: out = 24'(1092);
			30253: out = 24'(5604);
			30254: out = 24'(8836);
			30255: out = 24'(5920);
			30256: out = 24'(-3212);
			30257: out = 24'(-5916);
			30258: out = 24'(-5004);
			30259: out = 24'(1912);
			30260: out = 24'(6332);
			30261: out = 24'(3056);
			30262: out = 24'(-3592);
			30263: out = 24'(1720);
			30264: out = 24'(13880);
			30265: out = 24'(7340);
			30266: out = 24'(6056);
			30267: out = 24'(1904);
			30268: out = 24'(2212);
			30269: out = 24'(1036);
			30270: out = 24'(-944);
			30271: out = 24'(-6732);
			30272: out = 24'(-4084);
			30273: out = 24'(4172);
			30274: out = 24'(6568);
			30275: out = 24'(1584);
			30276: out = 24'(-256);
			30277: out = 24'(864);
			30278: out = 24'(268);
			30279: out = 24'(-10848);
			30280: out = 24'(-10664);
			30281: out = 24'(2296);
			30282: out = 24'(7612);
			30283: out = 24'(2580);
			30284: out = 24'(1536);
			30285: out = 24'(7420);
			30286: out = 24'(5124);
			30287: out = 24'(-380);
			30288: out = 24'(-4432);
			30289: out = 24'(-548);
			30290: out = 24'(3344);
			30291: out = 24'(-3320);
			30292: out = 24'(-3152);
			30293: out = 24'(7464);
			30294: out = 24'(15704);
			30295: out = 24'(1656);
			30296: out = 24'(-9516);
			30297: out = 24'(-11804);
			30298: out = 24'(-7112);
			30299: out = 24'(-7856);
			30300: out = 24'(-1508);
			30301: out = 24'(6584);
			30302: out = 24'(12340);
			30303: out = 24'(9200);
			30304: out = 24'(5424);
			30305: out = 24'(632);
			30306: out = 24'(-1596);
			30307: out = 24'(-6252);
			30308: out = 24'(436);
			30309: out = 24'(-36);
			30310: out = 24'(-432);
			30311: out = 24'(-1444);
			30312: out = 24'(540);
			30313: out = 24'(-11592);
			30314: out = 24'(-16000);
			30315: out = 24'(-3592);
			30316: out = 24'(15440);
			30317: out = 24'(11004);
			30318: out = 24'(-1876);
			30319: out = 24'(-10692);
			30320: out = 24'(-6940);
			30321: out = 24'(-2920);
			30322: out = 24'(4416);
			30323: out = 24'(2596);
			30324: out = 24'(-9320);
			30325: out = 24'(-13164);
			30326: out = 24'(-1212);
			30327: out = 24'(5528);
			30328: out = 24'(-3544);
			30329: out = 24'(-11380);
			30330: out = 24'(2696);
			30331: out = 24'(13008);
			30332: out = 24'(1136);
			30333: out = 24'(-2872);
			30334: out = 24'(-3184);
			30335: out = 24'(1848);
			30336: out = 24'(-2468);
			30337: out = 24'(-5624);
			30338: out = 24'(-9052);
			30339: out = 24'(236);
			30340: out = 24'(5948);
			30341: out = 24'(56);
			30342: out = 24'(-9800);
			30343: out = 24'(-7996);
			30344: out = 24'(1560);
			30345: out = 24'(6212);
			30346: out = 24'(-704);
			30347: out = 24'(-2164);
			30348: out = 24'(2924);
			30349: out = 24'(6308);
			30350: out = 24'(3124);
			30351: out = 24'(4252);
			30352: out = 24'(9624);
			30353: out = 24'(10380);
			30354: out = 24'(528);
			30355: out = 24'(-7812);
			30356: out = 24'(-8468);
			30357: out = 24'(-4000);
			30358: out = 24'(-2816);
			30359: out = 24'(764);
			30360: out = 24'(4564);
			30361: out = 24'(5328);
			30362: out = 24'(-1012);
			30363: out = 24'(-7840);
			30364: out = 24'(-7048);
			30365: out = 24'(2296);
			30366: out = 24'(8116);
			30367: out = 24'(9012);
			30368: out = 24'(3276);
			30369: out = 24'(1560);
			30370: out = 24'(1516);
			30371: out = 24'(2376);
			30372: out = 24'(-7112);
			30373: out = 24'(-7776);
			30374: out = 24'(-1936);
			30375: out = 24'(-3124);
			30376: out = 24'(-7992);
			30377: out = 24'(-5720);
			30378: out = 24'(3720);
			30379: out = 24'(7704);
			30380: out = 24'(7488);
			30381: out = 24'(2184);
			30382: out = 24'(-452);
			30383: out = 24'(116);
			30384: out = 24'(1404);
			30385: out = 24'(760);
			30386: out = 24'(-540);
			30387: out = 24'(816);
			30388: out = 24'(5472);
			30389: out = 24'(6800);
			30390: out = 24'(1296);
			30391: out = 24'(-7028);
			30392: out = 24'(-9320);
			30393: out = 24'(284);
			30394: out = 24'(6148);
			30395: out = 24'(-516);
			30396: out = 24'(-13880);
			30397: out = 24'(-5736);
			30398: out = 24'(3936);
			30399: out = 24'(4864);
			30400: out = 24'(320);
			30401: out = 24'(5116);
			30402: out = 24'(7376);
			30403: out = 24'(12);
			30404: out = 24'(-14024);
			30405: out = 24'(-18432);
			30406: out = 24'(-7400);
			30407: out = 24'(5612);
			30408: out = 24'(2892);
			30409: out = 24'(-12220);
			30410: out = 24'(-12688);
			30411: out = 24'(4176);
			30412: out = 24'(17388);
			30413: out = 24'(11236);
			30414: out = 24'(-8444);
			30415: out = 24'(-14724);
			30416: out = 24'(-2904);
			30417: out = 24'(5680);
			30418: out = 24'(3064);
			30419: out = 24'(-9440);
			30420: out = 24'(-10212);
			30421: out = 24'(2328);
			30422: out = 24'(436);
			30423: out = 24'(5976);
			30424: out = 24'(14036);
			30425: out = 24'(18584);
			30426: out = 24'(6664);
			30427: out = 24'(-4752);
			30428: out = 24'(-11464);
			30429: out = 24'(-5408);
			30430: out = 24'(6084);
			30431: out = 24'(12224);
			30432: out = 24'(6248);
			30433: out = 24'(-1500);
			30434: out = 24'(-60);
			30435: out = 24'(-8656);
			30436: out = 24'(-7316);
			30437: out = 24'(-2676);
			30438: out = 24'(708);
			30439: out = 24'(2160);
			30440: out = 24'(2672);
			30441: out = 24'(-684);
			30442: out = 24'(-3948);
			30443: out = 24'(6248);
			30444: out = 24'(5268);
			30445: out = 24'(2320);
			30446: out = 24'(-292);
			30447: out = 24'(208);
			30448: out = 24'(-3896);
			30449: out = 24'(-4272);
			30450: out = 24'(-1316);
			30451: out = 24'(-28);
			30452: out = 24'(708);
			30453: out = 24'(-1296);
			30454: out = 24'(-3060);
			30455: out = 24'(-4736);
			30456: out = 24'(-2408);
			30457: out = 24'(2888);
			30458: out = 24'(8344);
			30459: out = 24'(4748);
			30460: out = 24'(4164);
			30461: out = 24'(-1488);
			30462: out = 24'(8220);
			30463: out = 24'(16156);
			30464: out = 24'(8692);
			30465: out = 24'(-17792);
			30466: out = 24'(-19904);
			30467: out = 24'(-1344);
			30468: out = 24'(7072);
			30469: out = 24'(-5424);
			30470: out = 24'(-8940);
			30471: out = 24'(-2044);
			30472: out = 24'(-52);
			30473: out = 24'(404);
			30474: out = 24'(5108);
			30475: out = 24'(7124);
			30476: out = 24'(-1400);
			30477: out = 24'(964);
			30478: out = 24'(-2400);
			30479: out = 24'(-1156);
			30480: out = 24'(3148);
			30481: out = 24'(9532);
			30482: out = 24'(3460);
			30483: out = 24'(-7040);
			30484: out = 24'(-10352);
			30485: out = 24'(1832);
			30486: out = 24'(8920);
			30487: out = 24'(6528);
			30488: out = 24'(252);
			30489: out = 24'(104);
			30490: out = 24'(-352);
			30491: out = 24'(-3916);
			30492: out = 24'(-9348);
			30493: out = 24'(-7952);
			30494: out = 24'(2632);
			30495: out = 24'(6784);
			30496: out = 24'(3760);
			30497: out = 24'(-1180);
			30498: out = 24'(-6836);
			30499: out = 24'(-10788);
			30500: out = 24'(-9880);
			30501: out = 24'(-1332);
			30502: out = 24'(5712);
			30503: out = 24'(9336);
			30504: out = 24'(2476);
			30505: out = 24'(-2560);
			30506: out = 24'(2168);
			30507: out = 24'(5844);
			30508: out = 24'(2648);
			30509: out = 24'(-1228);
			30510: out = 24'(336);
			30511: out = 24'(-356);
			30512: out = 24'(-264);
			30513: out = 24'(1872);
			30514: out = 24'(5832);
			30515: out = 24'(-2792);
			30516: out = 24'(-3160);
			30517: out = 24'(-1112);
			30518: out = 24'(3220);
			30519: out = 24'(5544);
			30520: out = 24'(5076);
			30521: out = 24'(-860);
			30522: out = 24'(-5348);
			30523: out = 24'(636);
			30524: out = 24'(3916);
			30525: out = 24'(10276);
			30526: out = 24'(8948);
			30527: out = 24'(684);
			30528: out = 24'(-3096);
			30529: out = 24'(-1580);
			30530: out = 24'(-2592);
			30531: out = 24'(-8864);
			30532: out = 24'(-9736);
			30533: out = 24'(-1172);
			30534: out = 24'(6796);
			30535: out = 24'(2772);
			30536: out = 24'(-8820);
			30537: out = 24'(-13084);
			30538: out = 24'(-6304);
			30539: out = 24'(1224);
			30540: out = 24'(1916);
			30541: out = 24'(-5596);
			30542: out = 24'(-3536);
			30543: out = 24'(3212);
			30544: out = 24'(-1604);
			30545: out = 24'(-2832);
			30546: out = 24'(-8228);
			30547: out = 24'(-1892);
			30548: out = 24'(6328);
			30549: out = 24'(7568);
			30550: out = 24'(-6800);
			30551: out = 24'(-9004);
			30552: out = 24'(3300);
			30553: out = 24'(11424);
			30554: out = 24'(3988);
			30555: out = 24'(-2544);
			30556: out = 24'(-1720);
			30557: out = 24'(1656);
			30558: out = 24'(1364);
			30559: out = 24'(4308);
			30560: out = 24'(5012);
			30561: out = 24'(-760);
			30562: out = 24'(-10788);
			30563: out = 24'(-5848);
			30564: out = 24'(1136);
			30565: out = 24'(-4276);
			30566: out = 24'(-8276);
			30567: out = 24'(-6280);
			30568: out = 24'(1404);
			30569: out = 24'(5824);
			30570: out = 24'(17552);
			30571: out = 24'(13528);
			30572: out = 24'(9344);
			30573: out = 24'(3536);
			30574: out = 24'(-3012);
			30575: out = 24'(-16344);
			30576: out = 24'(-20012);
			30577: out = 24'(-12216);
			30578: out = 24'(1156);
			30579: out = 24'(10424);
			30580: out = 24'(13476);
			30581: out = 24'(8288);
			30582: out = 24'(-996);
			30583: out = 24'(-2356);
			30584: out = 24'(-8540);
			30585: out = 24'(-14268);
			30586: out = 24'(-12012);
			30587: out = 24'(572);
			30588: out = 24'(6668);
			30589: out = 24'(4456);
			30590: out = 24'(3264);
			30591: out = 24'(5604);
			30592: out = 24'(6144);
			30593: out = 24'(-5508);
			30594: out = 24'(-13704);
			30595: out = 24'(-1476);
			30596: out = 24'(4928);
			30597: out = 24'(3848);
			30598: out = 24'(-576);
			30599: out = 24'(3024);
			30600: out = 24'(-352);
			30601: out = 24'(1560);
			30602: out = 24'(-436);
			30603: out = 24'(-5828);
			30604: out = 24'(-6656);
			30605: out = 24'(-7708);
			30606: out = 24'(-3720);
			30607: out = 24'(1604);
			30608: out = 24'(6816);
			30609: out = 24'(6140);
			30610: out = 24'(8272);
			30611: out = 24'(4216);
			30612: out = 24'(-12004);
			30613: out = 24'(-16712);
			30614: out = 24'(-4752);
			30615: out = 24'(11128);
			30616: out = 24'(10668);
			30617: out = 24'(2752);
			30618: out = 24'(720);
			30619: out = 24'(8028);
			30620: out = 24'(8324);
			30621: out = 24'(3564);
			30622: out = 24'(-10704);
			30623: out = 24'(-12836);
			30624: out = 24'(-5448);
			30625: out = 24'(2348);
			30626: out = 24'(-13276);
			30627: out = 24'(-16524);
			30628: out = 24'(-60);
			30629: out = 24'(13256);
			30630: out = 24'(11488);
			30631: out = 24'(3792);
			30632: out = 24'(2068);
			30633: out = 24'(-1308);
			30634: out = 24'(-6412);
			30635: out = 24'(-16996);
			30636: out = 24'(-13196);
			30637: out = 24'(2680);
			30638: out = 24'(12284);
			30639: out = 24'(5008);
			30640: out = 24'(1312);
			30641: out = 24'(8736);
			30642: out = 24'(11596);
			30643: out = 24'(5828);
			30644: out = 24'(-1144);
			30645: out = 24'(-2520);
			30646: out = 24'(-2920);
			30647: out = 24'(-4296);
			30648: out = 24'(-2812);
			30649: out = 24'(2448);
			30650: out = 24'(5912);
			30651: out = 24'(1496);
			30652: out = 24'(-2168);
			30653: out = 24'(-1440);
			30654: out = 24'(2348);
			30655: out = 24'(5728);
			30656: out = 24'(4432);
			30657: out = 24'(-3456);
			30658: out = 24'(-11680);
			30659: out = 24'(4);
			30660: out = 24'(4468);
			30661: out = 24'(8064);
			30662: out = 24'(6848);
			30663: out = 24'(2372);
			30664: out = 24'(-3904);
			30665: out = 24'(-2372);
			30666: out = 24'(4412);
			30667: out = 24'(6688);
			30668: out = 24'(-9476);
			30669: out = 24'(-22896);
			30670: out = 24'(-18004);
			30671: out = 24'(2396);
			30672: out = 24'(7588);
			30673: out = 24'(4472);
			30674: out = 24'(-3200);
			30675: out = 24'(-3160);
			30676: out = 24'(-740);
			30677: out = 24'(5836);
			30678: out = 24'(3952);
			30679: out = 24'(1764);
			30680: out = 24'(11704);
			30681: out = 24'(9084);
			30682: out = 24'(-2916);
			30683: out = 24'(-11844);
			30684: out = 24'(-1904);
			30685: out = 24'(-848);
			30686: out = 24'(-2380);
			30687: out = 24'(-3760);
			30688: out = 24'(4032);
			30689: out = 24'(10212);
			30690: out = 24'(10600);
			30691: out = 24'(-128);
			30692: out = 24'(-9040);
			30693: out = 24'(-6276);
			30694: out = 24'(8520);
			30695: out = 24'(12904);
			30696: out = 24'(3140);
			30697: out = 24'(-3816);
			30698: out = 24'(-6460);
			30699: out = 24'(288);
			30700: out = 24'(7028);
			30701: out = 24'(5284);
			30702: out = 24'(-348);
			30703: out = 24'(-6716);
			30704: out = 24'(-5276);
			30705: out = 24'(1672);
			30706: out = 24'(5932);
			30707: out = 24'(2384);
			30708: out = 24'(-840);
			30709: out = 24'(36);
			30710: out = 24'(3676);
			30711: out = 24'(1224);
			30712: out = 24'(-788);
			30713: out = 24'(-324);
			30714: out = 24'(1956);
			30715: out = 24'(-8320);
			30716: out = 24'(-10188);
			30717: out = 24'(-400);
			30718: out = 24'(-1372);
			30719: out = 24'(2768);
			30720: out = 24'(-900);
			30721: out = 24'(-1872);
			30722: out = 24'(1516);
			30723: out = 24'(3988);
			30724: out = 24'(4908);
			30725: out = 24'(6680);
			30726: out = 24'(5024);
			30727: out = 24'(6632);
			30728: out = 24'(860);
			30729: out = 24'(192);
			30730: out = 24'(668);
			30731: out = 24'(340);
			30732: out = 24'(-12840);
			30733: out = 24'(-15588);
			30734: out = 24'(-8048);
			30735: out = 24'(-2688);
			30736: out = 24'(132);
			30737: out = 24'(10888);
			30738: out = 24'(18744);
			30739: out = 24'(10628);
			30740: out = 24'(-10140);
			30741: out = 24'(-12328);
			30742: out = 24'(-1980);
			30743: out = 24'(-1180);
			30744: out = 24'(2096);
			30745: out = 24'(2668);
			30746: out = 24'(3644);
			30747: out = 24'(100);
			30748: out = 24'(-4824);
			30749: out = 24'(-5684);
			30750: out = 24'(-6084);
			30751: out = 24'(-6624);
			30752: out = 24'(1896);
			30753: out = 24'(2372);
			30754: out = 24'(-1168);
			30755: out = 24'(-5608);
			30756: out = 24'(-2316);
			30757: out = 24'(4124);
			30758: out = 24'(7200);
			30759: out = 24'(4024);
			30760: out = 24'(-1304);
			30761: out = 24'(-8460);
			30762: out = 24'(-13288);
			30763: out = 24'(-11644);
			30764: out = 24'(-180);
			30765: out = 24'(6800);
			30766: out = 24'(12372);
			30767: out = 24'(8320);
			30768: out = 24'(60);
			30769: out = 24'(-4752);
			30770: out = 24'(-6672);
			30771: out = 24'(-7788);
			30772: out = 24'(-4196);
			30773: out = 24'(8516);
			30774: out = 24'(8808);
			30775: out = 24'(3916);
			30776: out = 24'(160);
			30777: out = 24'(6388);
			30778: out = 24'(-7924);
			30779: out = 24'(-9420);
			30780: out = 24'(-5548);
			30781: out = 24'(-2764);
			30782: out = 24'(-4572);
			30783: out = 24'(-1920);
			30784: out = 24'(3112);
			30785: out = 24'(6944);
			30786: out = 24'(8380);
			30787: out = 24'(6712);
			30788: out = 24'(5984);
			30789: out = 24'(5056);
			30790: out = 24'(-672);
			30791: out = 24'(-2204);
			30792: out = 24'(-6732);
			30793: out = 24'(-10184);
			30794: out = 24'(-6048);
			30795: out = 24'(8292);
			30796: out = 24'(14616);
			30797: out = 24'(3596);
			30798: out = 24'(-15388);
			30799: out = 24'(-10804);
			30800: out = 24'(604);
			30801: out = 24'(7948);
			30802: out = 24'(4932);
			30803: out = 24'(2320);
			30804: out = 24'(700);
			30805: out = 24'(2076);
			30806: out = 24'(1344);
			30807: out = 24'(1804);
			30808: out = 24'(3928);
			30809: out = 24'(10552);
			30810: out = 24'(10780);
			30811: out = 24'(-1928);
			30812: out = 24'(-16476);
			30813: out = 24'(-18396);
			30814: out = 24'(-7116);
			30815: out = 24'(-1280);
			30816: out = 24'(-5256);
			30817: out = 24'(-5240);
			30818: out = 24'(8460);
			30819: out = 24'(14048);
			30820: out = 24'(-6068);
			30821: out = 24'(-23772);
			30822: out = 24'(-9644);
			30823: out = 24'(18916);
			30824: out = 24'(21204);
			30825: out = 24'(2556);
			30826: out = 24'(-9308);
			30827: out = 24'(-5420);
			30828: out = 24'(-3632);
			30829: out = 24'(-6292);
			30830: out = 24'(-2136);
			30831: out = 24'(8152);
			30832: out = 24'(10808);
			30833: out = 24'(1724);
			30834: out = 24'(-1672);
			30835: out = 24'(-84);
			30836: out = 24'(-512);
			30837: out = 24'(1412);
			30838: out = 24'(140);
			30839: out = 24'(-696);
			30840: out = 24'(-556);
			30841: out = 24'(-584);
			30842: out = 24'(-1684);
			30843: out = 24'(-6764);
			30844: out = 24'(-7908);
			30845: out = 24'(1916);
			30846: out = 24'(7448);
			30847: out = 24'(4428);
			30848: out = 24'(-1744);
			30849: out = 24'(-2084);
			30850: out = 24'(4888);
			30851: out = 24'(3112);
			30852: out = 24'(-1412);
			30853: out = 24'(540);
			30854: out = 24'(-832);
			30855: out = 24'(236);
			30856: out = 24'(-764);
			30857: out = 24'(-516);
			30858: out = 24'(-3140);
			30859: out = 24'(3620);
			30860: out = 24'(6316);
			30861: out = 24'(4372);
			30862: out = 24'(-540);
			30863: out = 24'(-3796);
			30864: out = 24'(-7700);
			30865: out = 24'(-8880);
			30866: out = 24'(-6168);
			30867: out = 24'(5600);
			30868: out = 24'(7792);
			30869: out = 24'(3396);
			30870: out = 24'(148);
			30871: out = 24'(4848);
			30872: out = 24'(2820);
			30873: out = 24'(-5868);
			30874: out = 24'(-13508);
			30875: out = 24'(-2940);
			30876: out = 24'(-580);
			30877: out = 24'(-504);
			30878: out = 24'(-3464);
			30879: out = 24'(-3724);
			30880: out = 24'(2356);
			30881: out = 24'(13596);
			30882: out = 24'(14516);
			30883: out = 24'(-1344);
			30884: out = 24'(-13364);
			30885: out = 24'(-15100);
			30886: out = 24'(-8060);
			30887: out = 24'(-2088);
			30888: out = 24'(1772);
			30889: out = 24'(4992);
			30890: out = 24'(3932);
			30891: out = 24'(-3704);
			30892: out = 24'(-3660);
			30893: out = 24'(-2228);
			30894: out = 24'(4416);
			30895: out = 24'(6912);
			30896: out = 24'(540);
			30897: out = 24'(-2404);
			30898: out = 24'(1504);
			30899: out = 24'(5828);
			30900: out = 24'(-820);
			30901: out = 24'(-1448);
			30902: out = 24'(-2304);
			30903: out = 24'(3884);
			30904: out = 24'(10016);
			30905: out = 24'(-3316);
			30906: out = 24'(-17032);
			30907: out = 24'(-15944);
			30908: out = 24'(572);
			30909: out = 24'(10168);
			30910: out = 24'(9196);
			30911: out = 24'(1808);
			30912: out = 24'(-2204);
			30913: out = 24'(1404);
			30914: out = 24'(3300);
			30915: out = 24'(4968);
			30916: out = 24'(5704);
			30917: out = 24'(5568);
			30918: out = 24'(740);
			30919: out = 24'(-724);
			30920: out = 24'(-368);
			30921: out = 24'(-380);
			30922: out = 24'(-2640);
			30923: out = 24'(-1352);
			30924: out = 24'(-176);
			30925: out = 24'(-92);
			30926: out = 24'(1220);
			30927: out = 24'(1156);
			30928: out = 24'(-3512);
			30929: out = 24'(-6304);
			30930: out = 24'(-1180);
			30931: out = 24'(10028);
			30932: out = 24'(8372);
			30933: out = 24'(-3468);
			30934: out = 24'(-6320);
			30935: out = 24'(-1284);
			30936: out = 24'(4916);
			30937: out = 24'(3436);
			30938: out = 24'(-3164);
			30939: out = 24'(-5056);
			30940: out = 24'(-2796);
			30941: out = 24'(1996);
			30942: out = 24'(4900);
			30943: out = 24'(392);
			30944: out = 24'(-5952);
			30945: out = 24'(-3304);
			30946: out = 24'(6744);
			30947: out = 24'(5112);
			30948: out = 24'(-4108);
			30949: out = 24'(-11988);
			30950: out = 24'(-5460);
			30951: out = 24'(4220);
			30952: out = 24'(7760);
			30953: out = 24'(-4296);
			30954: out = 24'(-13644);
			30955: out = 24'(-3796);
			30956: out = 24'(3920);
			30957: out = 24'(3936);
			30958: out = 24'(-2652);
			30959: out = 24'(-3684);
			30960: out = 24'(-1376);
			30961: out = 24'(1280);
			30962: out = 24'(-4204);
			30963: out = 24'(-11252);
			30964: out = 24'(-11600);
			30965: out = 24'(2068);
			30966: out = 24'(10340);
			30967: out = 24'(5192);
			30968: out = 24'(-5552);
			30969: out = 24'(-7316);
			30970: out = 24'(-6612);
			30971: out = 24'(-10904);
			30972: out = 24'(-16080);
			30973: out = 24'(5168);
			30974: out = 24'(21820);
			30975: out = 24'(16996);
			30976: out = 24'(56);
			30977: out = 24'(-900);
			30978: out = 24'(5992);
			30979: out = 24'(1876);
			30980: out = 24'(-14320);
			30981: out = 24'(-2956);
			30982: out = 24'(3604);
			30983: out = 24'(5064);
			30984: out = 24'(-1284);
			30985: out = 24'(-1380);
			30986: out = 24'(-1512);
			30987: out = 24'(4304);
			30988: out = 24'(7900);
			30989: out = 24'(5728);
			30990: out = 24'(2624);
			30991: out = 24'(-3080);
			30992: out = 24'(-7176);
			30993: out = 24'(-1116);
			30994: out = 24'(5088);
			30995: out = 24'(14088);
			30996: out = 24'(13740);
			30997: out = 24'(5740);
			30998: out = 24'(-8288);
			30999: out = 24'(-7232);
			31000: out = 24'(-5660);
			31001: out = 24'(-11620);
			31002: out = 24'(-24636);
			31003: out = 24'(-4772);
			31004: out = 24'(15852);
			31005: out = 24'(14192);
			31006: out = 24'(1520);
			31007: out = 24'(-6816);
			31008: out = 24'(-2664);
			31009: out = 24'(-1328);
			31010: out = 24'(-6288);
			31011: out = 24'(-9516);
			31012: out = 24'(-1748);
			31013: out = 24'(1768);
			31014: out = 24'(-1964);
			31015: out = 24'(-596);
			31016: out = 24'(12368);
			31017: out = 24'(16156);
			31018: out = 24'(1632);
			31019: out = 24'(-15792);
			31020: out = 24'(-18348);
			31021: out = 24'(-9424);
			31022: out = 24'(-296);
			31023: out = 24'(2168);
			31024: out = 24'(6168);
			31025: out = 24'(4204);
			31026: out = 24'(4160);
			31027: out = 24'(11116);
			31028: out = 24'(3480);
			31029: out = 24'(-14752);
			31030: out = 24'(-24668);
			31031: out = 24'(-7260);
			31032: out = 24'(8276);
			31033: out = 24'(9424);
			31034: out = 24'(-5272);
			31035: out = 24'(-9784);
			31036: out = 24'(8912);
			31037: out = 24'(18464);
			31038: out = 24'(5432);
			31039: out = 24'(-13424);
			31040: out = 24'(-14784);
			31041: out = 24'(-3736);
			31042: out = 24'(3976);
			31043: out = 24'(4924);
			31044: out = 24'(6664);
			31045: out = 24'(6920);
			31046: out = 24'(124);
			31047: out = 24'(-8084);
			31048: out = 24'(-4676);
			31049: out = 24'(4100);
			31050: out = 24'(7192);
			31051: out = 24'(24);
			31052: out = 24'(-6048);
			31053: out = 24'(-5064);
			31054: out = 24'(-36);
			31055: out = 24'(-2472);
			31056: out = 24'(-9788);
			31057: out = 24'(-14412);
			31058: out = 24'(1404);
			31059: out = 24'(16084);
			31060: out = 24'(15720);
			31061: out = 24'(2468);
			31062: out = 24'(3312);
			31063: out = 24'(5392);
			31064: out = 24'(36);
			31065: out = 24'(-13564);
			31066: out = 24'(-7732);
			31067: out = 24'(-1300);
			31068: out = 24'(4712);
			31069: out = 24'(8332);
			31070: out = 24'(6452);
			31071: out = 24'(3772);
			31072: out = 24'(1688);
			31073: out = 24'(2380);
			31074: out = 24'(-412);
			31075: out = 24'(-572);
			31076: out = 24'(-8688);
			31077: out = 24'(-14340);
			31078: out = 24'(-1464);
			31079: out = 24'(8704);
			31080: out = 24'(13380);
			31081: out = 24'(8524);
			31082: out = 24'(156);
			31083: out = 24'(-132);
			31084: out = 24'(-1924);
			31085: out = 24'(-6816);
			31086: out = 24'(-7668);
			31087: out = 24'(368);
			31088: out = 24'(10336);
			31089: out = 24'(11708);
			31090: out = 24'(3864);
			31091: out = 24'(-1668);
			31092: out = 24'(-7704);
			31093: out = 24'(-9392);
			31094: out = 24'(-8876);
			31095: out = 24'(-8740);
			31096: out = 24'(-7116);
			31097: out = 24'(-2664);
			31098: out = 24'(5136);
			31099: out = 24'(11456);
			31100: out = 24'(12408);
			31101: out = 24'(5256);
			31102: out = 24'(-2836);
			31103: out = 24'(-7024);
			31104: out = 24'(-10780);
			31105: out = 24'(-10472);
			31106: out = 24'(-3576);
			31107: out = 24'(9244);
			31108: out = 24'(21524);
			31109: out = 24'(19748);
			31110: out = 24'(9700);
			31111: out = 24'(-552);
			31112: out = 24'(-9116);
			31113: out = 24'(-11120);
			31114: out = 24'(-11748);
			31115: out = 24'(-9608);
			31116: out = 24'(-1988);
			31117: out = 24'(4448);
			31118: out = 24'(7048);
			31119: out = 24'(4208);
			31120: out = 24'(644);
			31121: out = 24'(9368);
			31122: out = 24'(10892);
			31123: out = 24'(-328);
			31124: out = 24'(-16764);
			31125: out = 24'(-11704);
			31126: out = 24'(-8016);
			31127: out = 24'(-6892);
			31128: out = 24'(-6948);
			31129: out = 24'(8132);
			31130: out = 24'(8160);
			31131: out = 24'(8412);
			31132: out = 24'(6444);
			31133: out = 24'(132);
			31134: out = 24'(-6904);
			31135: out = 24'(-9780);
			31136: out = 24'(-6224);
			31137: out = 24'(2096);
			31138: out = 24'(-3532);
			31139: out = 24'(-2004);
			31140: out = 24'(1856);
			31141: out = 24'(1392);
			31142: out = 24'(-6988);
			31143: out = 24'(-5976);
			31144: out = 24'(4300);
			31145: out = 24'(11824);
			31146: out = 24'(8620);
			31147: out = 24'(-3584);
			31148: out = 24'(-9808);
			31149: out = 24'(-3264);
			31150: out = 24'(5364);
			31151: out = 24'(7232);
			31152: out = 24'(3480);
			31153: out = 24'(1788);
			31154: out = 24'(-416);
			31155: out = 24'(7448);
			31156: out = 24'(1216);
			31157: out = 24'(-4876);
			31158: out = 24'(1408);
			31159: out = 24'(6332);
			31160: out = 24'(2896);
			31161: out = 24'(-6820);
			31162: out = 24'(-6688);
			31163: out = 24'(3908);
			31164: out = 24'(11432);
			31165: out = 24'(6432);
			31166: out = 24'(-724);
			31167: out = 24'(-540);
			31168: out = 24'(6056);
			31169: out = 24'(3452);
			31170: out = 24'(-4672);
			31171: out = 24'(-4012);
			31172: out = 24'(7316);
			31173: out = 24'(12968);
			31174: out = 24'(5980);
			31175: out = 24'(-5296);
			31176: out = 24'(-5856);
			31177: out = 24'(-2008);
			31178: out = 24'(-1496);
			31179: out = 24'(-5264);
			31180: out = 24'(-964);
			31181: out = 24'(676);
			31182: out = 24'(3524);
			31183: out = 24'(4612);
			31184: out = 24'(-2556);
			31185: out = 24'(-1732);
			31186: out = 24'(2608);
			31187: out = 24'(4452);
			31188: out = 24'(-3288);
			31189: out = 24'(-3268);
			31190: out = 24'(-2192);
			31191: out = 24'(-884);
			31192: out = 24'(-1004);
			31193: out = 24'(4372);
			31194: out = 24'(5728);
			31195: out = 24'(3344);
			31196: out = 24'(-920);
			31197: out = 24'(4804);
			31198: out = 24'(-1116);
			31199: out = 24'(-8632);
			31200: out = 24'(-8068);
			31201: out = 24'(252);
			31202: out = 24'(5148);
			31203: out = 24'(2676);
			31204: out = 24'(-1036);
			31205: out = 24'(-832);
			31206: out = 24'(1064);
			31207: out = 24'(-3008);
			31208: out = 24'(-9284);
			31209: out = 24'(-11228);
			31210: out = 24'(-736);
			31211: out = 24'(2968);
			31212: out = 24'(-464);
			31213: out = 24'(-5136);
			31214: out = 24'(-5072);
			31215: out = 24'(1212);
			31216: out = 24'(9840);
			31217: out = 24'(10896);
			31218: out = 24'(1164);
			31219: out = 24'(-15608);
			31220: out = 24'(-20984);
			31221: out = 24'(-14140);
			31222: out = 24'(-11504);
			31223: out = 24'(-7660);
			31224: out = 24'(608);
			31225: out = 24'(10852);
			31226: out = 24'(10608);
			31227: out = 24'(3424);
			31228: out = 24'(-5036);
			31229: out = 24'(-4328);
			31230: out = 24'(1756);
			31231: out = 24'(516);
			31232: out = 24'(-5664);
			31233: out = 24'(-7248);
			31234: out = 24'(3092);
			31235: out = 24'(14728);
			31236: out = 24'(18684);
			31237: out = 24'(7564);
			31238: out = 24'(-6860);
			31239: out = 24'(-8808);
			31240: out = 24'(-5820);
			31241: out = 24'(-6120);
			31242: out = 24'(-8388);
			31243: out = 24'(-1088);
			31244: out = 24'(12492);
			31245: out = 24'(18960);
			31246: out = 24'(10960);
			31247: out = 24'(-580);
			31248: out = 24'(-8984);
			31249: out = 24'(-4136);
			31250: out = 24'(584);
			31251: out = 24'(-1080);
			31252: out = 24'(-8580);
			31253: out = 24'(3132);
			31254: out = 24'(17880);
			31255: out = 24'(17268);
			31256: out = 24'(700);
			31257: out = 24'(-10368);
			31258: out = 24'(-9000);
			31259: out = 24'(-1216);
			31260: out = 24'(1036);
			31261: out = 24'(1432);
			31262: out = 24'(-16);
			31263: out = 24'(-624);
			31264: out = 24'(-292);
			31265: out = 24'(4280);
			31266: out = 24'(9792);
			31267: out = 24'(11412);
			31268: out = 24'(2340);
			31269: out = 24'(-7376);
			31270: out = 24'(-17988);
			31271: out = 24'(-13580);
			31272: out = 24'(-1012);
			31273: out = 24'(5296);
			31274: out = 24'(1000);
			31275: out = 24'(2416);
			31276: out = 24'(7056);
			31277: out = 24'(-1056);
			31278: out = 24'(668);
			31279: out = 24'(3276);
			31280: out = 24'(4100);
			31281: out = 24'(-3888);
			31282: out = 24'(312);
			31283: out = 24'(592);
			31284: out = 24'(-5128);
			31285: out = 24'(-16716);
			31286: out = 24'(-4020);
			31287: out = 24'(2484);
			31288: out = 24'(7016);
			31289: out = 24'(2800);
			31290: out = 24'(-9724);
			31291: out = 24'(-13944);
			31292: out = 24'(-1036);
			31293: out = 24'(12236);
			31294: out = 24'(5108);
			31295: out = 24'(-8724);
			31296: out = 24'(-14092);
			31297: out = 24'(-4772);
			31298: out = 24'(1188);
			31299: out = 24'(-428);
			31300: out = 24'(92);
			31301: out = 24'(12840);
			31302: out = 24'(18256);
			31303: out = 24'(4820);
			31304: out = 24'(-24568);
			31305: out = 24'(-32152);
			31306: out = 24'(-11532);
			31307: out = 24'(-732);
			31308: out = 24'(-328);
			31309: out = 24'(1492);
			31310: out = 24'(11428);
			31311: out = 24'(17700);
			31312: out = 24'(11476);
			31313: out = 24'(2504);
			31314: out = 24'(-5672);
			31315: out = 24'(-15264);
			31316: out = 24'(-16312);
			31317: out = 24'(-6828);
			31318: out = 24'(3644);
			31319: out = 24'(6428);
			31320: out = 24'(4592);
			31321: out = 24'(8992);
			31322: out = 24'(10772);
			31323: out = 24'(4464);
			31324: out = 24'(-5728);
			31325: out = 24'(-1732);
			31326: out = 24'(1368);
			31327: out = 24'(-3716);
			31328: out = 24'(-3772);
			31329: out = 24'(7568);
			31330: out = 24'(17792);
			31331: out = 24'(13888);
			31332: out = 24'(-176);
			31333: out = 24'(-6268);
			31334: out = 24'(-8612);
			31335: out = 24'(-9168);
			31336: out = 24'(-6208);
			31337: out = 24'(-1492);
			31338: out = 24'(7892);
			31339: out = 24'(15872);
			31340: out = 24'(16408);
			31341: out = 24'(8752);
			31342: out = 24'(-332);
			31343: out = 24'(-3940);
			31344: out = 24'(-3428);
			31345: out = 24'(-3092);
			31346: out = 24'(-6612);
			31347: out = 24'(-4476);
			31348: out = 24'(3588);
			31349: out = 24'(10388);
			31350: out = 24'(6672);
			31351: out = 24'(5260);
			31352: out = 24'(7104);
			31353: out = 24'(3056);
			31354: out = 24'(-20084);
			31355: out = 24'(-33424);
			31356: out = 24'(-21764);
			31357: out = 24'(4628);
			31358: out = 24'(20620);
			31359: out = 24'(19656);
			31360: out = 24'(11424);
			31361: out = 24'(3544);
			31362: out = 24'(-4660);
			31363: out = 24'(-13460);
			31364: out = 24'(-16760);
			31365: out = 24'(-12288);
			31366: out = 24'(-7424);
			31367: out = 24'(-16);
			31368: out = 24'(2248);
			31369: out = 24'(620);
			31370: out = 24'(-2088);
			31371: out = 24'(5752);
			31372: out = 24'(8208);
			31373: out = 24'(1272);
			31374: out = 24'(-9200);
			31375: out = 24'(-9692);
			31376: out = 24'(-2240);
			31377: out = 24'(1400);
			31378: out = 24'(-3408);
			31379: out = 24'(-3988);
			31380: out = 24'(-1728);
			31381: out = 24'(1260);
			31382: out = 24'(-1608);
			31383: out = 24'(-7708);
			31384: out = 24'(-5348);
			31385: out = 24'(5568);
			31386: out = 24'(10516);
			31387: out = 24'(-128);
			31388: out = 24'(-3500);
			31389: out = 24'(-2536);
			31390: out = 24'(1288);
			31391: out = 24'(-508);
			31392: out = 24'(-3020);
			31393: out = 24'(-3004);
			31394: out = 24'(5252);
			31395: out = 24'(10984);
			31396: out = 24'(9316);
			31397: out = 24'(-3876);
			31398: out = 24'(-9488);
			31399: out = 24'(-5564);
			31400: out = 24'(-228);
			31401: out = 24'(-2260);
			31402: out = 24'(3676);
			31403: out = 24'(12648);
			31404: out = 24'(7016);
			31405: out = 24'(36);
			31406: out = 24'(-1720);
			31407: out = 24'(3892);
			31408: out = 24'(2804);
			31409: out = 24'(4804);
			31410: out = 24'(696);
			31411: out = 24'(-28);
			31412: out = 24'(-1028);
			31413: out = 24'(-1808);
			31414: out = 24'(-6388);
			31415: out = 24'(-4552);
			31416: out = 24'(716);
			31417: out = 24'(5828);
			31418: out = 24'(1436);
			31419: out = 24'(-368);
			31420: out = 24'(-1680);
			31421: out = 24'(-8448);
			31422: out = 24'(-388);
			31423: out = 24'(12092);
			31424: out = 24'(12776);
			31425: out = 24'(-688);
			31426: out = 24'(-12620);
			31427: out = 24'(-5940);
			31428: out = 24'(3324);
			31429: out = 24'(-1120);
			31430: out = 24'(180);
			31431: out = 24'(-1544);
			31432: out = 24'(-6052);
			31433: out = 24'(-10124);
			31434: out = 24'(4808);
			31435: out = 24'(10736);
			31436: out = 24'(6816);
			31437: out = 24'(-968);
			31438: out = 24'(1296);
			31439: out = 24'(392);
			31440: out = 24'(-8120);
			31441: out = 24'(-15916);
			31442: out = 24'(-5400);
			31443: out = 24'(7836);
			31444: out = 24'(10584);
			31445: out = 24'(1948);
			31446: out = 24'(-1928);
			31447: out = 24'(-3724);
			31448: out = 24'(-232);
			31449: out = 24'(-1136);
			31450: out = 24'(-3352);
			31451: out = 24'(-17740);
			31452: out = 24'(-5392);
			31453: out = 24'(6040);
			31454: out = 24'(4360);
			31455: out = 24'(-3312);
			31456: out = 24'(2528);
			31457: out = 24'(8464);
			31458: out = 24'(1360);
			31459: out = 24'(-12552);
			31460: out = 24'(-22328);
			31461: out = 24'(-12592);
			31462: out = 24'(2800);
			31463: out = 24'(6324);
			31464: out = 24'(7008);
			31465: out = 24'(9544);
			31466: out = 24'(11452);
			31467: out = 24'(3900);
			31468: out = 24'(-4396);
			31469: out = 24'(-7184);
			31470: out = 24'(1056);
			31471: out = 24'(5144);
			31472: out = 24'(1088);
			31473: out = 24'(-7988);
			31474: out = 24'(-2140);
			31475: out = 24'(7096);
			31476: out = 24'(3952);
			31477: out = 24'(-13236);
			31478: out = 24'(-14556);
			31479: out = 24'(-972);
			31480: out = 24'(5736);
			31481: out = 24'(2436);
			31482: out = 24'(-2888);
			31483: out = 24'(-3464);
			31484: out = 24'(-964);
			31485: out = 24'(5572);
			31486: out = 24'(10868);
			31487: out = 24'(8436);
			31488: out = 24'(-992);
			31489: out = 24'(1028);
			31490: out = 24'(-228);
			31491: out = 24'(-36);
			31492: out = 24'(-4020);
			31493: out = 24'(-7780);
			31494: out = 24'(-2616);
			31495: out = 24'(7480);
			31496: out = 24'(10652);
			31497: out = 24'(4252);
			31498: out = 24'(5396);
			31499: out = 24'(6852);
			31500: out = 24'(448);
			31501: out = 24'(-14804);
			31502: out = 24'(-15340);
			31503: out = 24'(-5696);
			31504: out = 24'(7800);
			31505: out = 24'(11296);
			31506: out = 24'(14268);
			31507: out = 24'(7212);
			31508: out = 24'(6676);
			31509: out = 24'(5640);
			31510: out = 24'(-2488);
			31511: out = 24'(-15548);
			31512: out = 24'(-14716);
			31513: out = 24'(-2428);
			31514: out = 24'(5524);
			31515: out = 24'(6584);
			31516: out = 24'(2556);
			31517: out = 24'(-1316);
			31518: out = 24'(-1840);
			31519: out = 24'(4276);
			31520: out = 24'(8336);
			31521: out = 24'(1376);
			31522: out = 24'(-12968);
			31523: out = 24'(-11096);
			31524: out = 24'(-7108);
			31525: out = 24'(-3564);
			31526: out = 24'(-4352);
			31527: out = 24'(896);
			31528: out = 24'(4032);
			31529: out = 24'(7084);
			31530: out = 24'(3872);
			31531: out = 24'(744);
			31532: out = 24'(-7416);
			31533: out = 24'(-6036);
			31534: out = 24'(-4688);
			31535: out = 24'(-7924);
			31536: out = 24'(-10176);
			31537: out = 24'(-488);
			31538: out = 24'(9872);
			31539: out = 24'(10476);
			31540: out = 24'(8480);
			31541: out = 24'(88);
			31542: out = 24'(-8296);
			31543: out = 24'(-12308);
			31544: out = 24'(-10348);
			31545: out = 24'(-1780);
			31546: out = 24'(712);
			31547: out = 24'(-1908);
			31548: out = 24'(968);
			31549: out = 24'(1924);
			31550: out = 24'(4024);
			31551: out = 24'(3600);
			31552: out = 24'(248);
			31553: out = 24'(-2844);
			31554: out = 24'(-5620);
			31555: out = 24'(-3316);
			31556: out = 24'(3816);
			31557: out = 24'(10452);
			31558: out = 24'(8600);
			31559: out = 24'(3064);
			31560: out = 24'(432);
			31561: out = 24'(1916);
			31562: out = 24'(-440);
			31563: out = 24'(-5428);
			31564: out = 24'(-7060);
			31565: out = 24'(956);
			31566: out = 24'(8492);
			31567: out = 24'(11016);
			31568: out = 24'(3104);
			31569: out = 24'(-5164);
			31570: out = 24'(-2424);
			31571: out = 24'(8860);
			31572: out = 24'(7736);
			31573: out = 24'(-7420);
			31574: out = 24'(-8580);
			31575: out = 24'(3524);
			31576: out = 24'(11984);
			31577: out = 24'(4364);
			31578: out = 24'(-4628);
			31579: out = 24'(72);
			31580: out = 24'(10744);
			31581: out = 24'(8732);
			31582: out = 24'(-3384);
			31583: out = 24'(-12592);
			31584: out = 24'(-6428);
			31585: out = 24'(3696);
			31586: out = 24'(5004);
			31587: out = 24'(1052);
			31588: out = 24'(1148);
			31589: out = 24'(4872);
			31590: out = 24'(4436);
			31591: out = 24'(-1136);
			31592: out = 24'(-3740);
			31593: out = 24'(-1140);
			31594: out = 24'(-864);
			31595: out = 24'(-1684);
			31596: out = 24'(-2508);
			31597: out = 24'(4500);
			31598: out = 24'(10644);
			31599: out = 24'(12188);
			31600: out = 24'(-9852);
			31601: out = 24'(-17208);
			31602: out = 24'(-2492);
			31603: out = 24'(10400);
			31604: out = 24'(4040);
			31605: out = 24'(-10868);
			31606: out = 24'(-17136);
			31607: out = 24'(-11568);
			31608: out = 24'(4632);
			31609: out = 24'(5104);
			31610: out = 24'(-6340);
			31611: out = 24'(-15560);
			31612: out = 24'(276);
			31613: out = 24'(6148);
			31614: out = 24'(1652);
			31615: out = 24'(-6332);
			31616: out = 24'(144);
			31617: out = 24'(-5508);
			31618: out = 24'(-9684);
			31619: out = 24'(-7944);
			31620: out = 24'(984);
			31621: out = 24'(5008);
			31622: out = 24'(9320);
			31623: out = 24'(10992);
			31624: out = 24'(6704);
			31625: out = 24'(-4732);
			31626: out = 24'(-13260);
			31627: out = 24'(-10772);
			31628: out = 24'(-1236);
			31629: out = 24'(-5148);
			31630: out = 24'(-2396);
			31631: out = 24'(3688);
			31632: out = 24'(5536);
			31633: out = 24'(1868);
			31634: out = 24'(-4564);
			31635: out = 24'(-304);
			31636: out = 24'(9268);
			31637: out = 24'(5508);
			31638: out = 24'(3620);
			31639: out = 24'(-404);
			31640: out = 24'(-2276);
			31641: out = 24'(-3828);
			31642: out = 24'(-188);
			31643: out = 24'(984);
			31644: out = 24'(-200);
			31645: out = 24'(-1204);
			31646: out = 24'(4960);
			31647: out = 24'(3980);
			31648: out = 24'(-5396);
			31649: out = 24'(-13452);
			31650: out = 24'(-3376);
			31651: out = 24'(9356);
			31652: out = 24'(9460);
			31653: out = 24'(-2204);
			31654: out = 24'(-4796);
			31655: out = 24'(3100);
			31656: out = 24'(10196);
			31657: out = 24'(3952);
			31658: out = 24'(-752);
			31659: out = 24'(-10908);
			31660: out = 24'(1088);
			31661: out = 24'(13256);
			31662: out = 24'(11276);
			31663: out = 24'(-3996);
			31664: out = 24'(-72);
			31665: out = 24'(12128);
			31666: out = 24'(12812);
			31667: out = 24'(-456);
			31668: out = 24'(-11176);
			31669: out = 24'(-9364);
			31670: out = 24'(3056);
			31671: out = 24'(8888);
			31672: out = 24'(16532);
			31673: out = 24'(9392);
			31674: out = 24'(-1556);
			31675: out = 24'(-5260);
			31676: out = 24'(-3168);
			31677: out = 24'(-6588);
			31678: out = 24'(-7152);
			31679: out = 24'(2028);
			31680: out = 24'(6468);
			31681: out = 24'(92);
			31682: out = 24'(-4740);
			31683: out = 24'(2544);
			31684: out = 24'(9012);
			31685: out = 24'(3924);
			31686: out = 24'(-2832);
			31687: out = 24'(496);
			31688: out = 24'(3512);
			31689: out = 24'(1936);
			31690: out = 24'(-9384);
			31691: out = 24'(-18736);
			31692: out = 24'(-14484);
			31693: out = 24'(-48);
			31694: out = 24'(11552);
			31695: out = 24'(6548);
			31696: out = 24'(-11268);
			31697: out = 24'(-17304);
			31698: out = 24'(-7132);
			31699: out = 24'(3972);
			31700: out = 24'(268);
			31701: out = 24'(1308);
			31702: out = 24'(-2316);
			31703: out = 24'(-592);
			31704: out = 24'(1428);
			31705: out = 24'(568);
			31706: out = 24'(-2040);
			31707: out = 24'(-456);
			31708: out = 24'(2116);
			31709: out = 24'(-164);
			31710: out = 24'(-10600);
			31711: out = 24'(-17476);
			31712: out = 24'(-13612);
			31713: out = 24'(-5548);
			31714: out = 24'(1992);
			31715: out = 24'(4600);
			31716: out = 24'(9008);
			31717: out = 24'(12028);
			31718: out = 24'(2836);
			31719: out = 24'(-11012);
			31720: out = 24'(-15920);
			31721: out = 24'(-7440);
			31722: out = 24'(1232);
			31723: out = 24'(7008);
			31724: out = 24'(9748);
			31725: out = 24'(10996);
			31726: out = 24'(5908);
			31727: out = 24'(3288);
			31728: out = 24'(128);
			31729: out = 24'(-3708);
			31730: out = 24'(-7748);
			31731: out = 24'(-1724);
			31732: out = 24'(7832);
			31733: out = 24'(12568);
			31734: out = 24'(6308);
			31735: out = 24'(3084);
			31736: out = 24'(3068);
			31737: out = 24'(7288);
			31738: out = 24'(4444);
			31739: out = 24'(-10520);
			31740: out = 24'(-16604);
			31741: out = 24'(-6148);
			31742: out = 24'(7748);
			31743: out = 24'(10616);
			31744: out = 24'(4112);
			31745: out = 24'(2708);
			31746: out = 24'(5768);
			31747: out = 24'(3080);
			31748: out = 24'(1824);
			31749: out = 24'(120);
			31750: out = 24'(804);
			31751: out = 24'(5660);
			31752: out = 24'(-368);
			31753: out = 24'(4204);
			31754: out = 24'(5272);
			31755: out = 24'(-1196);
			31756: out = 24'(-472);
			31757: out = 24'(4128);
			31758: out = 24'(6772);
			31759: out = 24'(4228);
			31760: out = 24'(4740);
			31761: out = 24'(-616);
			31762: out = 24'(-7896);
			31763: out = 24'(-10000);
			31764: out = 24'(-568);
			31765: out = 24'(4020);
			31766: out = 24'(3176);
			31767: out = 24'(792);
			31768: out = 24'(972);
			31769: out = 24'(-28);
			31770: out = 24'(-6024);
			31771: out = 24'(-8208);
			31772: out = 24'(-2536);
			31773: out = 24'(-4660);
			31774: out = 24'(-10144);
			31775: out = 24'(-13352);
			31776: out = 24'(-9132);
			31777: out = 24'(-4900);
			31778: out = 24'(528);
			31779: out = 24'(4320);
			31780: out = 24'(4372);
			31781: out = 24'(-4024);
			31782: out = 24'(-9232);
			31783: out = 24'(-6980);
			31784: out = 24'(-204);
			31785: out = 24'(-924);
			31786: out = 24'(-7460);
			31787: out = 24'(-7564);
			31788: out = 24'(5352);
			31789: out = 24'(14464);
			31790: out = 24'(5544);
			31791: out = 24'(-11052);
			31792: out = 24'(-13076);
			31793: out = 24'(1024);
			31794: out = 24'(10160);
			31795: out = 24'(4936);
			31796: out = 24'(-3392);
			31797: out = 24'(-5032);
			31798: out = 24'(68);
			31799: out = 24'(424);
			31800: out = 24'(3068);
			31801: out = 24'(6564);
			31802: out = 24'(5568);
			31803: out = 24'(-2064);
			31804: out = 24'(-3144);
			31805: out = 24'(2364);
			31806: out = 24'(5368);
			31807: out = 24'(1260);
			31808: out = 24'(-1820);
			31809: out = 24'(24);
			31810: out = 24'(6808);
			31811: out = 24'(6496);
			31812: out = 24'(7244);
			31813: out = 24'(-464);
			31814: out = 24'(-9404);
			31815: out = 24'(-10692);
			31816: out = 24'(6316);
			31817: out = 24'(13896);
			31818: out = 24'(7364);
			31819: out = 24'(324);
			31820: out = 24'(3420);
			31821: out = 24'(4496);
			31822: out = 24'(-2412);
			31823: out = 24'(-10568);
			31824: out = 24'(-6432);
			31825: out = 24'(4240);
			31826: out = 24'(13816);
			31827: out = 24'(14968);
			31828: out = 24'(6448);
			31829: out = 24'(-1484);
			31830: out = 24'(-2480);
			31831: out = 24'(-1188);
			31832: out = 24'(-2620);
			31833: out = 24'(-7012);
			31834: out = 24'(-1484);
			31835: out = 24'(7784);
			31836: out = 24'(5764);
			31837: out = 24'(-6992);
			31838: out = 24'(-12624);
			31839: out = 24'(-6044);
			31840: out = 24'(-908);
			31841: out = 24'(6248);
			31842: out = 24'(3960);
			31843: out = 24'(-2420);
			31844: out = 24'(-9072);
			31845: out = 24'(-1116);
			31846: out = 24'(-3672);
			31847: out = 24'(-9320);
			31848: out = 24'(-8292);
			31849: out = 24'(8932);
			31850: out = 24'(13040);
			31851: out = 24'(6636);
			31852: out = 24'(-1752);
			31853: out = 24'(-2608);
			31854: out = 24'(-4368);
			31855: out = 24'(-7776);
			31856: out = 24'(-10436);
			31857: out = 24'(-3668);
			31858: out = 24'(-1448);
			31859: out = 24'(3664);
			31860: out = 24'(4740);
			31861: out = 24'(1524);
			31862: out = 24'(-96);
			31863: out = 24'(924);
			31864: out = 24'(172);
			31865: out = 24'(-6108);
			31866: out = 24'(-11704);
			31867: out = 24'(-12556);
			31868: out = 24'(-4884);
			31869: out = 24'(3048);
			31870: out = 24'(1764);
			31871: out = 24'(-1456);
			31872: out = 24'(3152);
			31873: out = 24'(13356);
			31874: out = 24'(10384);
			31875: out = 24'(2552);
			31876: out = 24'(-16056);
			31877: out = 24'(-22560);
			31878: out = 24'(-11504);
			31879: out = 24'(-4548);
			31880: out = 24'(-2860);
			31881: out = 24'(4308);
			31882: out = 24'(16728);
			31883: out = 24'(11720);
			31884: out = 24'(28);
			31885: out = 24'(-8016);
			31886: out = 24'(-4228);
			31887: out = 24'(-248);
			31888: out = 24'(972);
			31889: out = 24'(2216);
			31890: out = 24'(8172);
			31891: out = 24'(11676);
			31892: out = 24'(6704);
			31893: out = 24'(-3616);
			31894: out = 24'(-7796);
			31895: out = 24'(-1692);
			31896: out = 24'(996);
			31897: out = 24'(-72);
			31898: out = 24'(-2432);
			31899: out = 24'(2044);
			31900: out = 24'(8816);
			31901: out = 24'(15432);
			31902: out = 24'(8824);
			31903: out = 24'(-6196);
			31904: out = 24'(-23268);
			31905: out = 24'(-10196);
			31906: out = 24'(4564);
			31907: out = 24'(6264);
			31908: out = 24'(2508);
			31909: out = 24'(5524);
			31910: out = 24'(8072);
			31911: out = 24'(5976);
			31912: out = 24'(5528);
			31913: out = 24'(-64);
			31914: out = 24'(-1360);
			31915: out = 24'(-5744);
			31916: out = 24'(-10452);
			31917: out = 24'(-4108);
			31918: out = 24'(3248);
			31919: out = 24'(4436);
			31920: out = 24'(1620);
			31921: out = 24'(4904);
			31922: out = 24'(3304);
			31923: out = 24'(-2448);
			31924: out = 24'(-6904);
			31925: out = 24'(-4796);
			31926: out = 24'(516);
			31927: out = 24'(304);
			31928: out = 24'(-4592);
			31929: out = 24'(-10304);
			31930: out = 24'(4188);
			31931: out = 24'(7712);
			31932: out = 24'(2812);
			31933: out = 24'(-2484);
			31934: out = 24'(1500);
			31935: out = 24'(428);
			31936: out = 24'(304);
			31937: out = 24'(1120);
			31938: out = 24'(284);
			31939: out = 24'(-892);
			31940: out = 24'(860);
			31941: out = 24'(-3976);
			31942: out = 24'(-19788);
			31943: out = 24'(-24480);
			31944: out = 24'(-4784);
			31945: out = 24'(16232);
			31946: out = 24'(14760);
			31947: out = 24'(-3472);
			31948: out = 24'(-6884);
			31949: out = 24'(-960);
			31950: out = 24'(-5276);
			31951: out = 24'(-14828);
			31952: out = 24'(-7072);
			31953: out = 24'(7084);
			31954: out = 24'(6096);
			31955: out = 24'(2400);
			31956: out = 24'(-908);
			31957: out = 24'(3640);
			31958: out = 24'(4868);
			31959: out = 24'(-1272);
			31960: out = 24'(-8352);
			31961: out = 24'(-9096);
			31962: out = 24'(-2772);
			31963: out = 24'(6024);
			31964: out = 24'(8172);
			31965: out = 24'(3972);
			31966: out = 24'(-652);
			31967: out = 24'(1244);
			31968: out = 24'(4740);
			31969: out = 24'(3912);
			31970: out = 24'(-4356);
			31971: out = 24'(-12396);
			31972: out = 24'(-12776);
			31973: out = 24'(-504);
			31974: out = 24'(10784);
			31975: out = 24'(11628);
			31976: out = 24'(6800);
			31977: out = 24'(1220);
			31978: out = 24'(212);
			31979: out = 24'(-388);
			31980: out = 24'(-1808);
			31981: out = 24'(-5936);
			31982: out = 24'(-2264);
			31983: out = 24'(3888);
			31984: out = 24'(5508);
			31985: out = 24'(2636);
			31986: out = 24'(3784);
			31987: out = 24'(4900);
			31988: out = 24'(-1668);
			31989: out = 24'(-8648);
			31990: out = 24'(-10888);
			31991: out = 24'(-2424);
			31992: out = 24'(6280);
			31993: out = 24'(6112);
			31994: out = 24'(1076);
			31995: out = 24'(3944);
			31996: out = 24'(15484);
			31997: out = 24'(19444);
			31998: out = 24'(6272);
			31999: out = 24'(-10780);
			32000: out = 24'(-12248);
			32001: out = 24'(-680);
			32002: out = 24'(9700);
			32003: out = 24'(1212);
			32004: out = 24'(-7996);
			32005: out = 24'(-968);
			32006: out = 24'(8192);
			32007: out = 24'(5588);
			32008: out = 24'(-7320);
			32009: out = 24'(-14072);
			32010: out = 24'(-4136);
			32011: out = 24'(260);
			32012: out = 24'(-1640);
			32013: out = 24'(-1860);
			32014: out = 24'(-636);
			32015: out = 24'(3288);
			32016: out = 24'(1696);
			32017: out = 24'(-740);
			32018: out = 24'(-2800);
			32019: out = 24'(5788);
			32020: out = 24'(3692);
			32021: out = 24'(-1772);
			32022: out = 24'(-2780);
			32023: out = 24'(-7748);
			32024: out = 24'(-10532);
			32025: out = 24'(-8080);
			32026: out = 24'(-1244);
			32027: out = 24'(1912);
			32028: out = 24'(900);
			32029: out = 24'(888);
			32030: out = 24'(1948);
			32031: out = 24'(428);
			32032: out = 24'(-4632);
			32033: out = 24'(-6264);
			32034: out = 24'(-7144);
			32035: out = 24'(-11852);
			32036: out = 24'(-12960);
			32037: out = 24'(-2440);
			32038: out = 24'(8988);
			32039: out = 24'(6772);
			32040: out = 24'(-6376);
			32041: out = 24'(-5940);
			32042: out = 24'(6680);
			32043: out = 24'(8972);
			32044: out = 24'(-4000);
			32045: out = 24'(-18624);
			32046: out = 24'(-13500);
			32047: out = 24'(3692);
			32048: out = 24'(6056);
			32049: out = 24'(4376);
			32050: out = 24'(2096);
			32051: out = 24'(3140);
			32052: out = 24'(636);
			32053: out = 24'(2696);
			32054: out = 24'(940);
			32055: out = 24'(-2852);
			32056: out = 24'(-4756);
			32057: out = 24'(5480);
			32058: out = 24'(11528);
			32059: out = 24'(8128);
			32060: out = 24'(396);
			32061: out = 24'(120);
			32062: out = 24'(5196);
			32063: out = 24'(7724);
			32064: out = 24'(4868);
			32065: out = 24'(624);
			32066: out = 24'(-2804);
			32067: out = 24'(-4980);
			32068: out = 24'(-2136);
			32069: out = 24'(5192);
			32070: out = 24'(6680);
			32071: out = 24'(1460);
			32072: out = 24'(-1880);
			32073: out = 24'(-208);
			32074: out = 24'(1096);
			32075: out = 24'(-6148);
			32076: out = 24'(-8180);
			32077: out = 24'(2920);
			32078: out = 24'(9840);
			32079: out = 24'(8112);
			32080: out = 24'(4932);
			32081: out = 24'(5188);
			32082: out = 24'(5952);
			32083: out = 24'(-9664);
			32084: out = 24'(-16904);
			32085: out = 24'(-3716);
			32086: out = 24'(8940);
			32087: out = 24'(9896);
			32088: out = 24'(2368);
			32089: out = 24'(512);
			32090: out = 24'(5032);
			32091: out = 24'(9760);
			32092: out = 24'(5468);
			32093: out = 24'(-4464);
			32094: out = 24'(-10368);
			32095: out = 24'(-6724);
			32096: out = 24'(56);
			32097: out = 24'(-2236);
			32098: out = 24'(-10400);
			32099: out = 24'(-1392);
			32100: out = 24'(5432);
			32101: out = 24'(5560);
			32102: out = 24'(404);
			32103: out = 24'(-2448);
			32104: out = 24'(-480);
			32105: out = 24'(-4340);
			32106: out = 24'(-11896);
			32107: out = 24'(-9948);
			32108: out = 24'(-2696);
			32109: out = 24'(3124);
			32110: out = 24'(4144);
			32111: out = 24'(5832);
			32112: out = 24'(824);
			32113: out = 24'(-1388);
			32114: out = 24'(-2988);
			32115: out = 24'(-4976);
			32116: out = 24'(-9424);
			32117: out = 24'(-13616);
			32118: out = 24'(-11284);
			32119: out = 24'(-972);
			32120: out = 24'(10264);
			32121: out = 24'(8996);
			32122: out = 24'(1244);
			32123: out = 24'(-3704);
			32124: out = 24'(908);
			32125: out = 24'(5824);
			32126: out = 24'(8192);
			32127: out = 24'(2544);
			32128: out = 24'(-5692);
			32129: out = 24'(-14032);
			32130: out = 24'(-6756);
			32131: out = 24'(4292);
			32132: out = 24'(7256);
			32133: out = 24'(-660);
			32134: out = 24'(292);
			32135: out = 24'(2680);
			32136: out = 24'(-700);
			32137: out = 24'(-5048);
			32138: out = 24'(-2404);
			32139: out = 24'(4628);
			32140: out = 24'(6320);
			32141: out = 24'(-3468);
			32142: out = 24'(4144);
			32143: out = 24'(10852);
			32144: out = 24'(7536);
			32145: out = 24'(-4240);
			32146: out = 24'(-6672);
			32147: out = 24'(-136);
			32148: out = 24'(7724);
			32149: out = 24'(6104);
			32150: out = 24'(6892);
			32151: out = 24'(-3660);
			32152: out = 24'(-8688);
			32153: out = 24'(-2868);
			32154: out = 24'(4636);
			32155: out = 24'(6832);
			32156: out = 24'(9096);
			32157: out = 24'(11656);
			32158: out = 24'(4784);
			32159: out = 24'(-3292);
			32160: out = 24'(-9564);
			32161: out = 24'(-6680);
			32162: out = 24'(-744);
			32163: out = 24'(6252);
			32164: out = 24'(3416);
			32165: out = 24'(-1288);
			32166: out = 24'(-80);
			32167: out = 24'(-772);
			32168: out = 24'(888);
			32169: out = 24'(-1116);
			32170: out = 24'(-7100);
			32171: out = 24'(1140);
			32172: out = 24'(-2856);
			32173: out = 24'(-3568);
			32174: out = 24'(1696);
			32175: out = 24'(9812);
			32176: out = 24'(7052);
			32177: out = 24'(2284);
			32178: out = 24'(-2444);
			32179: out = 24'(-8868);
			32180: out = 24'(-18056);
			32181: out = 24'(-12580);
			32182: out = 24'(2524);
			32183: out = 24'(4336);
			32184: out = 24'(8856);
			32185: out = 24'(1544);
			32186: out = 24'(3732);
			32187: out = 24'(11736);
			32188: out = 24'(6616);
			32189: out = 24'(-6164);
			32190: out = 24'(-9392);
			32191: out = 24'(-2252);
			32192: out = 24'(-8728);
			32193: out = 24'(-10528);
			32194: out = 24'(-4300);
			32195: out = 24'(8740);
			32196: out = 24'(9220);
			32197: out = 24'(3820);
			32198: out = 24'(-6896);
			32199: out = 24'(-8988);
			32200: out = 24'(-4504);
			32201: out = 24'(-3364);
			32202: out = 24'(-8012);
			32203: out = 24'(-6984);
			32204: out = 24'(4216);
			32205: out = 24'(14932);
			32206: out = 24'(11284);
			32207: out = 24'(-1676);
			32208: out = 24'(-9160);
			32209: out = 24'(1048);
			32210: out = 24'(-2092);
			32211: out = 24'(-10952);
			32212: out = 24'(-11028);
			32213: out = 24'(1612);
			32214: out = 24'(7700);
			32215: out = 24'(1884);
			32216: out = 24'(-2728);
			32217: out = 24'(6524);
			32218: out = 24'(11188);
			32219: out = 24'(6544);
			32220: out = 24'(-3292);
			32221: out = 24'(-5640);
			32222: out = 24'(-13744);
			32223: out = 24'(-9296);
			32224: out = 24'(-836);
			32225: out = 24'(9136);
			32226: out = 24'(9624);
			32227: out = 24'(15664);
			32228: out = 24'(10804);
			32229: out = 24'(-5372);
			32230: out = 24'(-26344);
			32231: out = 24'(-18172);
			32232: out = 24'(-1420);
			32233: out = 24'(6604);
			32234: out = 24'(6256);
			32235: out = 24'(5260);
			32236: out = 24'(8888);
			32237: out = 24'(8832);
			32238: out = 24'(908);
			32239: out = 24'(-6404);
			32240: out = 24'(-9748);
			32241: out = 24'(-9928);
			32242: out = 24'(-8712);
			32243: out = 24'(976);
			32244: out = 24'(5268);
			32245: out = 24'(4832);
			32246: out = 24'(1680);
			32247: out = 24'(620);
			32248: out = 24'(304);
			32249: out = 24'(292);
			32250: out = 24'(1264);
			32251: out = 24'(5716);
			32252: out = 24'(2704);
			32253: out = 24'(104);
			32254: out = 24'(1120);
			32255: out = 24'(5476);
			32256: out = 24'(1064);
			32257: out = 24'(-2640);
			32258: out = 24'(-3828);
			32259: out = 24'(-1872);
			32260: out = 24'(-2200);
			32261: out = 24'(-444);
			32262: out = 24'(576);
			32263: out = 24'(92);
			32264: out = 24'(596);
			32265: out = 24'(896);
			32266: out = 24'(6068);
			32267: out = 24'(9448);
			32268: out = 24'(-256);
			32269: out = 24'(-1720);
			32270: out = 24'(-1480);
			32271: out = 24'(100);
			32272: out = 24'(-2748);
			32273: out = 24'(-300);
			32274: out = 24'(356);
			32275: out = 24'(3500);
			32276: out = 24'(4276);
			32277: out = 24'(-536);
			32278: out = 24'(-10980);
			32279: out = 24'(-10724);
			32280: out = 24'(1728);
			32281: out = 24'(2904);
			32282: out = 24'(5360);
			32283: out = 24'(5348);
			32284: out = 24'(4408);
			32285: out = 24'(-2416);
			32286: out = 24'(-3884);
			32287: out = 24'(-4516);
			32288: out = 24'(-4128);
			32289: out = 24'(-3884);
			32290: out = 24'(3588);
			32291: out = 24'(6404);
			32292: out = 24'(2972);
			32293: out = 24'(-2184);
			32294: out = 24'(-704);
			32295: out = 24'(656);
			32296: out = 24'(-2908);
			32297: out = 24'(-7684);
			32298: out = 24'(-648);
			32299: out = 24'(2120);
			32300: out = 24'(-544);
			32301: out = 24'(-4268);
			32302: out = 24'(-4328);
			32303: out = 24'(3520);
			32304: out = 24'(2404);
			32305: out = 24'(-7476);
			32306: out = 24'(-15408);
			32307: out = 24'(-3372);
			32308: out = 24'(2544);
			32309: out = 24'(-2296);
			32310: out = 24'(-6208);
			32311: out = 24'(4716);
			32312: out = 24'(13792);
			32313: out = 24'(12620);
			32314: out = 24'(3680);
			32315: out = 24'(-10396);
			32316: out = 24'(-8544);
			32317: out = 24'(2964);
			32318: out = 24'(10508);
			32319: out = 24'(5796);
			32320: out = 24'(-4092);
			32321: out = 24'(-8220);
			32322: out = 24'(800);
			32323: out = 24'(15364);
			32324: out = 24'(5072);
			32325: out = 24'(-9256);
			32326: out = 24'(-11476);
			32327: out = 24'(828);
			32328: out = 24'(6292);
			32329: out = 24'(3796);
			32330: out = 24'(-2152);
			32331: out = 24'(-3132);
			32332: out = 24'(4212);
			32333: out = 24'(7148);
			32334: out = 24'(5104);
			32335: out = 24'(384);
			32336: out = 24'(-2000);
			32337: out = 24'(-6844);
			32338: out = 24'(-7240);
			32339: out = 24'(-2692);
			32340: out = 24'(-112);
			32341: out = 24'(4352);
			32342: out = 24'(5888);
			32343: out = 24'(4064);
			32344: out = 24'(-168);
			32345: out = 24'(-2116);
			32346: out = 24'(-616);
			32347: out = 24'(1648);
			32348: out = 24'(-676);
			32349: out = 24'(280);
			32350: out = 24'(-580);
			32351: out = 24'(852);
			32352: out = 24'(920);
			32353: out = 24'(-3504);
			32354: out = 24'(-2536);
			32355: out = 24'(5168);
			32356: out = 24'(8908);
			32357: out = 24'(152);
			32358: out = 24'(-13052);
			32359: out = 24'(-12052);
			32360: out = 24'(3208);
			32361: out = 24'(10548);
			32362: out = 24'(9452);
			32363: out = 24'(404);
			32364: out = 24'(-580);
			32365: out = 24'(4648);
			32366: out = 24'(1232);
			32367: out = 24'(-9568);
			32368: out = 24'(-12168);
			32369: out = 24'(-44);
			32370: out = 24'(4016);
			32371: out = 24'(2908);
			32372: out = 24'(-4836);
			32373: out = 24'(-6720);
			32374: out = 24'(-676);
			32375: out = 24'(6104);
			32376: out = 24'(3256);
			32377: out = 24'(-4048);
			32378: out = 24'(-5568);
			32379: out = 24'(2644);
			32380: out = 24'(6708);
			32381: out = 24'(2784);
			32382: out = 24'(-2024);
			32383: out = 24'(-964);
			32384: out = 24'(1632);
			32385: out = 24'(216);
			32386: out = 24'(-2104);
			32387: out = 24'(-804);
			32388: out = 24'(5120);
			32389: out = 24'(3488);
			32390: out = 24'(-6372);
			32391: out = 24'(-7248);
			32392: out = 24'(-3580);
			32393: out = 24'(5964);
			32394: out = 24'(8944);
			32395: out = 24'(1836);
			32396: out = 24'(-5232);
			32397: out = 24'(-1316);
			32398: out = 24'(7316);
			32399: out = 24'(5256);
			32400: out = 24'(2104);
			32401: out = 24'(-7560);
			32402: out = 24'(-8128);
			32403: out = 24'(1264);
			32404: out = 24'(10468);
			32405: out = 24'(8160);
			32406: out = 24'(2016);
			32407: out = 24'(-392);
			32408: out = 24'(1104);
			32409: out = 24'(-5272);
			32410: out = 24'(-10244);
			32411: out = 24'(-5568);
			32412: out = 24'(4412);
			32413: out = 24'(7144);
			32414: out = 24'(3236);
			32415: out = 24'(-2200);
			32416: out = 24'(-6324);
			32417: out = 24'(-384);
			32418: out = 24'(3840);
			32419: out = 24'(3972);
			32420: out = 24'(-1344);
			32421: out = 24'(-1688);
			32422: out = 24'(-7132);
			32423: out = 24'(-6272);
			32424: out = 24'(552);
			32425: out = 24'(4696);
			32426: out = 24'(5196);
			32427: out = 24'(3716);
			32428: out = 24'(432);
			32429: out = 24'(96);
			32430: out = 24'(-7132);
			32431: out = 24'(-7832);
			32432: out = 24'(-5804);
			32433: out = 24'(-1640);
			32434: out = 24'(-1676);
			32435: out = 24'(7500);
			32436: out = 24'(8380);
			32437: out = 24'(-5636);
			32438: out = 24'(-11916);
			32439: out = 24'(-2320);
			32440: out = 24'(7652);
			32441: out = 24'(3024);
			32442: out = 24'(-6552);
			32443: out = 24'(-4128);
			32444: out = 24'(3728);
			32445: out = 24'(3668);
			32446: out = 24'(-3420);
			32447: out = 24'(-1860);
			32448: out = 24'(1724);
			32449: out = 24'(-476);
			32450: out = 24'(-5652);
			32451: out = 24'(-1680);
			32452: out = 24'(2832);
			32453: out = 24'(2592);
			32454: out = 24'(304);
			32455: out = 24'(4272);
			32456: out = 24'(4092);
			32457: out = 24'(-2112);
			32458: out = 24'(-8696);
			32459: out = 24'(-12424);
			32460: out = 24'(-8260);
			32461: out = 24'(-2848);
			32462: out = 24'(4788);
			32463: out = 24'(13748);
			32464: out = 24'(17516);
			32465: out = 24'(6936);
			32466: out = 24'(-7076);
			32467: out = 24'(-8032);
			32468: out = 24'(-8480);
			32469: out = 24'(-9360);
			32470: out = 24'(-8408);
			32471: out = 24'(-1272);
			32472: out = 24'(4788);
			32473: out = 24'(3124);
			32474: out = 24'(-84);
			32475: out = 24'(2888);
			32476: out = 24'(4944);
			32477: out = 24'(2716);
			32478: out = 24'(-2192);
			32479: out = 24'(-4080);
			32480: out = 24'(-5980);
			32481: out = 24'(-4684);
			32482: out = 24'(588);
			32483: out = 24'(10164);
			32484: out = 24'(15184);
			32485: out = 24'(5236);
			32486: out = 24'(-8204);
			32487: out = 24'(-9736);
			32488: out = 24'(92);
			32489: out = 24'(5340);
			32490: out = 24'(2008);
			32491: out = 24'(396);
			32492: out = 24'(4368);
			32493: out = 24'(15128);
			32494: out = 24'(3656);
			32495: out = 24'(-14768);
			32496: out = 24'(-21616);
			32497: out = 24'(-5856);
			32498: out = 24'(3408);
			32499: out = 24'(6304);
			32500: out = 24'(4068);
			32501: out = 24'(-1532);
			32502: out = 24'(-3148);
			32503: out = 24'(2628);
			32504: out = 24'(6360);
			32505: out = 24'(-852);
			32506: out = 24'(-10100);
			32507: out = 24'(-9176);
			32508: out = 24'(-1116);
			32509: out = 24'(1460);
			32510: out = 24'(5520);
			32511: out = 24'(9072);
			32512: out = 24'(12696);
			32513: out = 24'(8120);
			32514: out = 24'(1556);
			32515: out = 24'(-6624);
			32516: out = 24'(-8276);
			32517: out = 24'(-7980);
			32518: out = 24'(-1668);
			32519: out = 24'(-2112);
			32520: out = 24'(7764);
			32521: out = 24'(16212);
			32522: out = 24'(9348);
			32523: out = 24'(-7688);
			32524: out = 24'(-12056);
			32525: out = 24'(-1872);
			32526: out = 24'(4068);
			32527: out = 24'(-1916);
			32528: out = 24'(-5128);
			32529: out = 24'(2488);
			32530: out = 24'(9524);
			32531: out = 24'(6516);
			32532: out = 24'(-6724);
			32533: out = 24'(-12368);
			32534: out = 24'(-3832);
			32535: out = 24'(288);
			32536: out = 24'(5604);
			32537: out = 24'(508);
			32538: out = 24'(-8240);
			32539: out = 24'(-13748);
			32540: out = 24'(608);
			32541: out = 24'(7760);
			32542: out = 24'(2416);
			32543: out = 24'(-3544);
			32544: out = 24'(-8416);
			32545: out = 24'(-588);
			32546: out = 24'(8272);
			32547: out = 24'(9344);
			32548: out = 24'(1356);
			32549: out = 24'(-1072);
			32550: out = 24'(600);
			32551: out = 24'(-1508);
			32552: out = 24'(-6816);
			32553: out = 24'(-13416);
			32554: out = 24'(-9036);
			32555: out = 24'(3616);
			32556: out = 24'(11164);
			32557: out = 24'(8168);
			32558: out = 24'(700);
			32559: out = 24'(-1800);
			32560: out = 24'(1312);
			32561: out = 24'(6212);
			32562: out = 24'(4396);
			32563: out = 24'(-1116);
			32564: out = 24'(-4868);
			32565: out = 24'(-13204);
			32566: out = 24'(-11732);
			32567: out = 24'(-2736);
			32568: out = 24'(6556);
			32569: out = 24'(10180);
			32570: out = 24'(5144);
			32571: out = 24'(-892);
			32572: out = 24'(-1780);
			32573: out = 24'(-564);
			32574: out = 24'(4336);
			32575: out = 24'(2348);
			32576: out = 24'(-3696);
			32577: out = 24'(-1628);
			32578: out = 24'(2872);
			32579: out = 24'(9808);
			32580: out = 24'(9956);
			32581: out = 24'(4504);
			32582: out = 24'(-2248);
			32583: out = 24'(1368);
			32584: out = 24'(4284);
			32585: out = 24'(-2076);
			32586: out = 24'(-3784);
			32587: out = 24'(-5724);
			32588: out = 24'(-2632);
			32589: out = 24'(-900);
			32590: out = 24'(-4208);
			32591: out = 24'(-1268);
			32592: out = 24'(4004);
			32593: out = 24'(2684);
			32594: out = 24'(-6104);
			32595: out = 24'(-7548);
			32596: out = 24'(-128);
			32597: out = 24'(4888);
			32598: out = 24'(-1112);
			32599: out = 24'(-5228);
			32600: out = 24'(-4896);
			32601: out = 24'(-1032);
			32602: out = 24'(-908);
			32603: out = 24'(508);
			32604: out = 24'(244);
			32605: out = 24'(3912);
			32606: out = 24'(6096);
			32607: out = 24'(324);
			32608: out = 24'(-7648);
			32609: out = 24'(-10776);
			32610: out = 24'(-5880);
			32611: out = 24'(1440);
			32612: out = 24'(6608);
			32613: out = 24'(2960);
			32614: out = 24'(-4136);
			32615: out = 24'(-3096);
			32616: out = 24'(2928);
			32617: out = 24'(7300);
			32618: out = 24'(460);
			32619: out = 24'(-6996);
			32620: out = 24'(2636);
			32621: out = 24'(13388);
			32622: out = 24'(7704);
			32623: out = 24'(-9388);
			32624: out = 24'(-22636);
			32625: out = 24'(-4532);
			32626: out = 24'(9860);
			32627: out = 24'(3128);
			32628: out = 24'(-6464);
			32629: out = 24'(-3508);
			32630: out = 24'(5368);
			32631: out = 24'(4388);
			32632: out = 24'(-3508);
			32633: out = 24'(-1716);
			32634: out = 24'(6840);
			32635: out = 24'(8272);
			32636: out = 24'(-1616);
			32637: out = 24'(-10592);
			32638: out = 24'(-10056);
			32639: out = 24'(-968);
			32640: out = 24'(5784);
			32641: out = 24'(7336);
			32642: out = 24'(5572);
			32643: out = 24'(5524);
			32644: out = 24'(3460);
			32645: out = 24'(-3888);
			32646: out = 24'(-15660);
			32647: out = 24'(-15612);
			32648: out = 24'(-3068);
			32649: out = 24'(6752);
			32650: out = 24'(11048);
			32651: out = 24'(4904);
			32652: out = 24'(-1028);
			32653: out = 24'(768);
			32654: out = 24'(4336);
			32655: out = 24'(3224);
			32656: out = 24'(-3732);
			32657: out = 24'(-7784);
			32658: out = 24'(-8796);
			32659: out = 24'(2600);
			32660: out = 24'(7988);
			32661: out = 24'(3608);
			32662: out = 24'(-3548);
			32663: out = 24'(-4476);
			32664: out = 24'(-2204);
			32665: out = 24'(1764);
			32666: out = 24'(4924);
			32667: out = 24'(3336);
			32668: out = 24'(-4300);
			32669: out = 24'(-6520);
			32670: out = 24'(400);
			32671: out = 24'(644);
			32672: out = 24'(-2688);
			32673: out = 24'(-1416);
			32674: out = 24'(6256);
			32675: out = 24'(7136);
			32676: out = 24'(2300);
			32677: out = 24'(1184);
			32678: out = 24'(5312);
			32679: out = 24'(-108);
			32680: out = 24'(-4660);
			32681: out = 24'(-4416);
			32682: out = 24'(1084);
			32683: out = 24'(-664);
			32684: out = 24'(1700);
			32685: out = 24'(1772);
			32686: out = 24'(728);
			32687: out = 24'(-4496);
			32688: out = 24'(-500);
			32689: out = 24'(92);
			32690: out = 24'(260);
			32691: out = 24'(2408);
			32692: out = 24'(6024);
			32693: out = 24'(4796);
			32694: out = 24'(-4624);
			32695: out = 24'(-14572);
			32696: out = 24'(-10560);
			32697: out = 24'(4092);
			32698: out = 24'(12724);
			32699: out = 24'(7256);
			32700: out = 24'(-1332);
			32701: out = 24'(-588);
			32702: out = 24'(4664);
			32703: out = 24'(1912);
			32704: out = 24'(-8028);
			32705: out = 24'(-7848);
			32706: out = 24'(664);
			32707: out = 24'(4220);
			32708: out = 24'(-3732);
			32709: out = 24'(-14488);
			32710: out = 24'(-10652);
			32711: out = 24'(1824);
			32712: out = 24'(6716);
			32713: out = 24'(6440);
			32714: out = 24'(1232);
			32715: out = 24'(196);
			32716: out = 24'(-420);
			32717: out = 24'(708);
			32718: out = 24'(-8060);
			32719: out = 24'(-6304);
			32720: out = 24'(2872);
			32721: out = 24'(6492);
			32722: out = 24'(-1180);
			32723: out = 24'(-4656);
			32724: out = 24'(928);
			32725: out = 24'(4980);
			32726: out = 24'(6192);
			32727: out = 24'(2376);
			32728: out = 24'(2560);
			32729: out = 24'(5032);
			32730: out = 24'(5512);
			32731: out = 24'(-4788);
			32732: out = 24'(-14336);
			32733: out = 24'(-14464);
			32734: out = 24'(-532);
			32735: out = 24'(1992);
			32736: out = 24'(2056);
			32737: out = 24'(1504);
			32738: out = 24'(2304);
			32739: out = 24'(-1536);
			32740: out = 24'(-984);
			32741: out = 24'(-284);
			32742: out = 24'(-2076);
			32743: out = 24'(-4304);
			32744: out = 24'(-284);
			32745: out = 24'(1308);
			32746: out = 24'(-2172);
			32747: out = 24'(-300);
			32748: out = 24'(6996);
			32749: out = 24'(9744);
			32750: out = 24'(3492);
			32751: out = 24'(-3460);
			32752: out = 24'(-1892);
			32753: out = 24'(-16);
			32754: out = 24'(-4020);
			32755: out = 24'(-7664);
			32756: out = 24'(-7040);
			32757: out = 24'(-3876);
			32758: out = 24'(-1288);
			32759: out = 24'(488);
			32760: out = 24'(6216);
			32761: out = 24'(6692);
			32762: out = 24'(5436);
			32763: out = 24'(6640);
			32764: out = 24'(-2968);
			32765: out = 24'(-6344);
			32766: out = 24'(-2532);
			32767: out = 24'(6592);
			32768: out = 24'(4632);
			32769: out = 24'(5904);
			32770: out = 24'(2640);
			32771: out = 24'(-164);
			32772: out = 24'(1204);
			32773: out = 24'(772);
			32774: out = 24'(-5144);
			32775: out = 24'(-11100);
			32776: out = 24'(-7316);
			32777: out = 24'(-620);
			32778: out = 24'(5880);
			32779: out = 24'(5640);
			32780: out = 24'(940);
			32781: out = 24'(-5624);
			32782: out = 24'(-36);
			32783: out = 24'(8544);
			32784: out = 24'(8284);
			32785: out = 24'(-672);
			32786: out = 24'(-9284);
			32787: out = 24'(-6840);
			32788: out = 24'(824);
			32789: out = 24'(-300);
			32790: out = 24'(4768);
			32791: out = 24'(9932);
			32792: out = 24'(9544);
			32793: out = 24'(-880);
			32794: out = 24'(-10128);
			32795: out = 24'(-14052);
			32796: out = 24'(-9716);
			32797: out = 24'(-1472);
			32798: out = 24'(9864);
			32799: out = 24'(12996);
			32800: out = 24'(7856);
			32801: out = 24'(-2608);
			32802: out = 24'(-18896);
			32803: out = 24'(-24244);
			32804: out = 24'(-16668);
			32805: out = 24'(364);
			32806: out = 24'(10732);
			32807: out = 24'(14336);
			32808: out = 24'(3696);
			32809: out = 24'(-6020);
			32810: out = 24'(552);
			32811: out = 24'(8624);
			32812: out = 24'(6504);
			32813: out = 24'(-4548);
			32814: out = 24'(-11708);
			32815: out = 24'(-9068);
			32816: out = 24'(-4208);
			32817: out = 24'(696);
			32818: out = 24'(6624);
			32819: out = 24'(10056);
			32820: out = 24'(5012);
			32821: out = 24'(-5948);
			32822: out = 24'(-13972);
			32823: out = 24'(-8092);
			32824: out = 24'(-1112);
			32825: out = 24'(2688);
			32826: out = 24'(-620);
			32827: out = 24'(1692);
			32828: out = 24'(148);
			32829: out = 24'(7508);
			32830: out = 24'(8380);
			32831: out = 24'(444);
			32832: out = 24'(-14756);
			32833: out = 24'(-4956);
			32834: out = 24'(8400);
			32835: out = 24'(4140);
			32836: out = 24'(-2436);
			32837: out = 24'(-844);
			32838: out = 24'(1488);
			32839: out = 24'(-5496);
			32840: out = 24'(-6800);
			32841: out = 24'(-2260);
			32842: out = 24'(7012);
			32843: out = 24'(10192);
			32844: out = 24'(5652);
			32845: out = 24'(1640);
			32846: out = 24'(-2452);
			32847: out = 24'(-3260);
			32848: out = 24'(40);
			32849: out = 24'(1980);
			32850: out = 24'(-3708);
			32851: out = 24'(-6924);
			32852: out = 24'(1724);
			32853: out = 24'(9068);
			32854: out = 24'(8516);
			32855: out = 24'(4132);
			32856: out = 24'(6120);
			32857: out = 24'(4452);
			32858: out = 24'(2648);
			32859: out = 24'(-4532);
			32860: out = 24'(-7820);
			32861: out = 24'(-6832);
			32862: out = 24'(4300);
			32863: out = 24'(5552);
			32864: out = 24'(280);
			32865: out = 24'(-2292);
			32866: out = 24'(-5400);
			32867: out = 24'(-6860);
			32868: out = 24'(-2760);
			32869: out = 24'(5552);
			32870: out = 24'(9352);
			32871: out = 24'(6776);
			32872: out = 24'(4840);
			32873: out = 24'(5772);
			32874: out = 24'(36);
			32875: out = 24'(-6180);
			32876: out = 24'(-5096);
			32877: out = 24'(2416);
			32878: out = 24'(-768);
			32879: out = 24'(-1284);
			32880: out = 24'(-3000);
			32881: out = 24'(-1580);
			32882: out = 24'(-460);
			32883: out = 24'(64);
			32884: out = 24'(-460);
			32885: out = 24'(-728);
			32886: out = 24'(-2780);
			32887: out = 24'(-3428);
			32888: out = 24'(-5440);
			32889: out = 24'(-3680);
			32890: out = 24'(3128);
			32891: out = 24'(9800);
			32892: out = 24'(10964);
			32893: out = 24'(5432);
			32894: out = 24'(-1648);
			32895: out = 24'(-7676);
			32896: out = 24'(-2824);
			32897: out = 24'(748);
			32898: out = 24'(-1388);
			32899: out = 24'(-3704);
			32900: out = 24'(-3216);
			32901: out = 24'(-688);
			32902: out = 24'(0);
			32903: out = 24'(1532);
			32904: out = 24'(-5156);
			32905: out = 24'(-2764);
			32906: out = 24'(800);
			32907: out = 24'(-708);
			32908: out = 24'(-8124);
			32909: out = 24'(-4556);
			32910: out = 24'(5192);
			32911: out = 24'(8688);
			32912: out = 24'(1084);
			32913: out = 24'(-4456);
			32914: out = 24'(-5852);
			32915: out = 24'(-5240);
			32916: out = 24'(-1544);
			32917: out = 24'(472);
			32918: out = 24'(6320);
			32919: out = 24'(10148);
			32920: out = 24'(9116);
			32921: out = 24'(-6152);
			32922: out = 24'(-8244);
			32923: out = 24'(0);
			32924: out = 24'(4108);
			32925: out = 24'(-3364);
			32926: out = 24'(-9100);
			32927: out = 24'(-5988);
			32928: out = 24'(1888);
			32929: out = 24'(10644);
			32930: out = 24'(4828);
			32931: out = 24'(-5608);
			32932: out = 24'(-9868);
			32933: out = 24'(1332);
			32934: out = 24'(-452);
			32935: out = 24'(-3276);
			32936: out = 24'(-1684);
			32937: out = 24'(5492);
			32938: out = 24'(9208);
			32939: out = 24'(6212);
			32940: out = 24'(-128);
			32941: out = 24'(604);
			32942: out = 24'(-1036);
			32943: out = 24'(1360);
			32944: out = 24'(-4720);
			32945: out = 24'(-12488);
			32946: out = 24'(-6952);
			32947: out = 24'(5724);
			32948: out = 24'(9160);
			32949: out = 24'(4620);
			32950: out = 24'(4852);
			32951: out = 24'(3584);
			32952: out = 24'(-5292);
			32953: out = 24'(-12572);
			32954: out = 24'(-3348);
			32955: out = 24'(10456);
			32956: out = 24'(13120);
			32957: out = 24'(7600);
			32958: out = 24'(4376);
			32959: out = 24'(2288);
			32960: out = 24'(-9804);
			32961: out = 24'(-17544);
			32962: out = 24'(-7228);
			32963: out = 24'(-1684);
			32964: out = 24'(2432);
			32965: out = 24'(888);
			32966: out = 24'(400);
			32967: out = 24'(-228);
			32968: out = 24'(-60);
			32969: out = 24'(2800);
			32970: out = 24'(6476);
			32971: out = 24'(-504);
			32972: out = 24'(-6444);
			32973: out = 24'(-11908);
			32974: out = 24'(-7248);
			32975: out = 24'(5472);
			32976: out = 24'(7088);
			32977: out = 24'(4084);
			32978: out = 24'(2220);
			32979: out = 24'(5284);
			32980: out = 24'(424);
			32981: out = 24'(16);
			32982: out = 24'(500);
			32983: out = 24'(1584);
			32984: out = 24'(-3672);
			32985: out = 24'(-1252);
			32986: out = 24'(1668);
			32987: out = 24'(3324);
			32988: out = 24'(-248);
			32989: out = 24'(444);
			32990: out = 24'(-1276);
			32991: out = 24'(-1808);
			32992: out = 24'(-2604);
			32993: out = 24'(704);
			32994: out = 24'(-5268);
			32995: out = 24'(-8152);
			32996: out = 24'(-972);
			32997: out = 24'(10008);
			32998: out = 24'(5460);
			32999: out = 24'(-1616);
			33000: out = 24'(960);
			33001: out = 24'(5632);
			33002: out = 24'(3836);
			33003: out = 24'(0);
			33004: out = 24'(-144);
			33005: out = 24'(-2524);
			33006: out = 24'(-3800);
			33007: out = 24'(-1932);
			33008: out = 24'(2392);
			33009: out = 24'(356);
			33010: out = 24'(-6640);
			33011: out = 24'(-13112);
			33012: out = 24'(-10280);
			33013: out = 24'(-1156);
			33014: out = 24'(11956);
			33015: out = 24'(11128);
			33016: out = 24'(1624);
			33017: out = 24'(-5364);
			33018: out = 24'(580);
			33019: out = 24'(4464);
			33020: out = 24'(3032);
			33021: out = 24'(-428);
			33022: out = 24'(1068);
			33023: out = 24'(-2228);
			33024: out = 24'(-7236);
			33025: out = 24'(-8300);
			33026: out = 24'(308);
			33027: out = 24'(8676);
			33028: out = 24'(11560);
			33029: out = 24'(6468);
			33030: out = 24'(-812);
			33031: out = 24'(-16760);
			33032: out = 24'(-17184);
			33033: out = 24'(-5016);
			33034: out = 24'(5272);
			33035: out = 24'(5836);
			33036: out = 24'(4320);
			33037: out = 24'(7788);
			33038: out = 24'(9728);
			33039: out = 24'(2620);
			33040: out = 24'(-9864);
			33041: out = 24'(-10416);
			33042: out = 24'(736);
			33043: out = 24'(5656);
			33044: out = 24'(-2156);
			33045: out = 24'(-5272);
			33046: out = 24'(4804);
			33047: out = 24'(12036);
			33048: out = 24'(2336);
			33049: out = 24'(-13392);
			33050: out = 24'(-12028);
			33051: out = 24'(6192);
			33052: out = 24'(5164);
			33053: out = 24'(1408);
			33054: out = 24'(3844);
			33055: out = 24'(14668);
			33056: out = 24'(8536);
			33057: out = 24'(956);
			33058: out = 24'(-10432);
			33059: out = 24'(-11912);
			33060: out = 24'(-5216);
			33061: out = 24'(3960);
			33062: out = 24'(1376);
			33063: out = 24'(-1340);
			33064: out = 24'(5084);
			33065: out = 24'(12304);
			33066: out = 24'(7592);
			33067: out = 24'(-2376);
			33068: out = 24'(-6320);
			33069: out = 24'(-11608);
			33070: out = 24'(-11216);
			33071: out = 24'(-5948);
			33072: out = 24'(2388);
			33073: out = 24'(-272);
			33074: out = 24'(2220);
			33075: out = 24'(4280);
			33076: out = 24'(4068);
			33077: out = 24'(-268);
			33078: out = 24'(-6192);
			33079: out = 24'(-6100);
			33080: out = 24'(-632);
			33081: out = 24'(-552);
			33082: out = 24'(1988);
			33083: out = 24'(1160);
			33084: out = 24'(2856);
			33085: out = 24'(4568);
			33086: out = 24'(5380);
			33087: out = 24'(-648);
			33088: out = 24'(-6092);
			33089: out = 24'(-7476);
			33090: out = 24'(-2476);
			33091: out = 24'(-980);
			33092: out = 24'(2872);
			33093: out = 24'(5680);
			33094: out = 24'(-1820);
			33095: out = 24'(-8136);
			33096: out = 24'(-6052);
			33097: out = 24'(1924);
			33098: out = 24'(1064);
			33099: out = 24'(5040);
			33100: out = 24'(3164);
			33101: out = 24'(-152);
			33102: out = 24'(-4184);
			33103: out = 24'(-2144);
			33104: out = 24'(-2164);
			33105: out = 24'(-1184);
			33106: out = 24'(-112);
			33107: out = 24'(-4708);
			33108: out = 24'(-6076);
			33109: out = 24'(-1820);
			33110: out = 24'(4120);
			33111: out = 24'(220);
			33112: out = 24'(324);
			33113: out = 24'(2096);
			33114: out = 24'(6012);
			33115: out = 24'(4244);
			33116: out = 24'(-3408);
			33117: out = 24'(-13264);
			33118: out = 24'(-11196);
			33119: out = 24'(808);
			33120: out = 24'(12940);
			33121: out = 24'(7104);
			33122: out = 24'(-1972);
			33123: out = 24'(-764);
			33124: out = 24'(5568);
			33125: out = 24'(3492);
			33126: out = 24'(-1824);
			33127: out = 24'(-616);
			33128: out = 24'(5688);
			33129: out = 24'(6192);
			33130: out = 24'(2960);
			33131: out = 24'(1108);
			33132: out = 24'(-332);
			33133: out = 24'(52);
			33134: out = 24'(-1168);
			33135: out = 24'(-2428);
			33136: out = 24'(-2088);
			33137: out = 24'(-516);
			33138: out = 24'(184);
			33139: out = 24'(-252);
			33140: out = 24'(232);
			33141: out = 24'(-452);
			33142: out = 24'(416);
			33143: out = 24'(-1584);
			33144: out = 24'(-3600);
			33145: out = 24'(-2724);
			33146: out = 24'(5984);
			33147: out = 24'(10892);
			33148: out = 24'(10548);
			33149: out = 24'(10328);
			33150: out = 24'(7548);
			33151: out = 24'(-1584);
			33152: out = 24'(-12260);
			33153: out = 24'(-11232);
			33154: out = 24'(-9512);
			33155: out = 24'(-3480);
			33156: out = 24'(1500);
			33157: out = 24'(4684);
			33158: out = 24'(1996);
			33159: out = 24'(104);
			33160: out = 24'(-220);
			33161: out = 24'(-1436);
			33162: out = 24'(-11812);
			33163: out = 24'(-14680);
			33164: out = 24'(-7432);
			33165: out = 24'(3644);
			33166: out = 24'(4688);
			33167: out = 24'(5576);
			33168: out = 24'(2864);
			33169: out = 24'(-544);
			33170: out = 24'(72);
			33171: out = 24'(-2320);
			33172: out = 24'(1684);
			33173: out = 24'(4672);
			33174: out = 24'(-768);
			33175: out = 24'(-5984);
			33176: out = 24'(-6572);
			33177: out = 24'(116);
			33178: out = 24'(6744);
			33179: out = 24'(6924);
			33180: out = 24'(-836);
			33181: out = 24'(-9192);
			33182: out = 24'(-9732);
			33183: out = 24'(-852);
			33184: out = 24'(7692);
			33185: out = 24'(8528);
			33186: out = 24'(3456);
			33187: out = 24'(392);
			33188: out = 24'(-620);
			33189: out = 24'(-1140);
			33190: out = 24'(-2636);
			33191: out = 24'(-1776);
			33192: out = 24'(-808);
			33193: out = 24'(3688);
			33194: out = 24'(8168);
			33195: out = 24'(10072);
			33196: out = 24'(-2460);
			33197: out = 24'(-7252);
			33198: out = 24'(-7796);
			33199: out = 24'(-8124);
			33200: out = 24'(-11020);
			33201: out = 24'(-10332);
			33202: out = 24'(-5400);
			33203: out = 24'(3020);
			33204: out = 24'(10760);
			33205: out = 24'(5272);
			33206: out = 24'(-2144);
			33207: out = 24'(-2468);
			33208: out = 24'(-316);
			33209: out = 24'(6556);
			33210: out = 24'(2744);
			33211: out = 24'(2164);
			33212: out = 24'(9832);
			33213: out = 24'(11232);
			33214: out = 24'(860);
			33215: out = 24'(-7992);
			33216: out = 24'(-4248);
			33217: out = 24'(3480);
			33218: out = 24'(2276);
			33219: out = 24'(-1368);
			33220: out = 24'(368);
			33221: out = 24'(-772);
			33222: out = 24'(1364);
			33223: out = 24'(624);
			33224: out = 24'(-968);
			33225: out = 24'(-4060);
			33226: out = 24'(2780);
			33227: out = 24'(5812);
			33228: out = 24'(1644);
			33229: out = 24'(-6160);
			33230: out = 24'(-8180);
			33231: out = 24'(-748);
			33232: out = 24'(7720);
			33233: out = 24'(7832);
			33234: out = 24'(-2544);
			33235: out = 24'(-5424);
			33236: out = 24'(-1892);
			33237: out = 24'(-1860);
			33238: out = 24'(-12328);
			33239: out = 24'(-10572);
			33240: out = 24'(1320);
			33241: out = 24'(13212);
			33242: out = 24'(12740);
			33243: out = 24'(5072);
			33244: out = 24'(-4664);
			33245: out = 24'(-6172);
			33246: out = 24'(852);
			33247: out = 24'(-5888);
			33248: out = 24'(-10024);
			33249: out = 24'(-5160);
			33250: out = 24'(6060);
			33251: out = 24'(9136);
			33252: out = 24'(3928);
			33253: out = 24'(-1668);
			33254: out = 24'(1152);
			33255: out = 24'(2008);
			33256: out = 24'(8344);
			33257: out = 24'(6156);
			33258: out = 24'(-1148);
			33259: out = 24'(-7764);
			33260: out = 24'(-2340);
			33261: out = 24'(-372);
			33262: out = 24'(-4436);
			33263: out = 24'(-9020);
			33264: out = 24'(7064);
			33265: out = 24'(9076);
			33266: out = 24'(-3376);
			33267: out = 24'(-12012);
			33268: out = 24'(-1700);
			33269: out = 24'(8792);
			33270: out = 24'(2992);
			33271: out = 24'(-11236);
			33272: out = 24'(-17332);
			33273: out = 24'(408);
			33274: out = 24'(13552);
			33275: out = 24'(7348);
			33276: out = 24'(-2392);
			33277: out = 24'(1812);
			33278: out = 24'(12148);
			33279: out = 24'(8860);
			33280: out = 24'(-5788);
			33281: out = 24'(-16968);
			33282: out = 24'(-8992);
			33283: out = 24'(3152);
			33284: out = 24'(3820);
			33285: out = 24'(-3808);
			33286: out = 24'(-7812);
			33287: out = 24'(-5740);
			33288: out = 24'(-964);
			33289: out = 24'(4460);
			33290: out = 24'(8612);
			33291: out = 24'(8260);
			33292: out = 24'(2848);
			33293: out = 24'(-5380);
			33294: out = 24'(-7668);
			33295: out = 24'(-6284);
			33296: out = 24'(-2904);
			33297: out = 24'(-2436);
			33298: out = 24'(4204);
			33299: out = 24'(5040);
			33300: out = 24'(4680);
			33301: out = 24'(732);
			33302: out = 24'(5704);
			33303: out = 24'(-4288);
			33304: out = 24'(-8008);
			33305: out = 24'(1256);
			33306: out = 24'(5844);
			33307: out = 24'(2948);
			33308: out = 24'(2144);
			33309: out = 24'(3744);
			33310: out = 24'(-5292);
			33311: out = 24'(-12448);
			33312: out = 24'(-6784);
			33313: out = 24'(6260);
			33314: out = 24'(8820);
			33315: out = 24'(-2208);
			33316: out = 24'(-4644);
			33317: out = 24'(1600);
			33318: out = 24'(-1344);
			33319: out = 24'(-4020);
			33320: out = 24'(-3892);
			33321: out = 24'(4680);
			33322: out = 24'(10188);
			33323: out = 24'(6356);
			33324: out = 24'(-2832);
			33325: out = 24'(-4792);
			33326: out = 24'(1248);
			33327: out = 24'(5532);
			33328: out = 24'(-3532);
			33329: out = 24'(-16356);
			33330: out = 24'(-15960);
			33331: out = 24'(-740);
			33332: out = 24'(5688);
			33333: out = 24'(-1148);
			33334: out = 24'(-6720);
			33335: out = 24'(656);
			33336: out = 24'(12104);
			33337: out = 24'(7672);
			33338: out = 24'(-4100);
			33339: out = 24'(-5972);
			33340: out = 24'(4380);
			33341: out = 24'(4500);
			33342: out = 24'(-5984);
			33343: out = 24'(-12140);
			33344: out = 24'(-4920);
			33345: out = 24'(3512);
			33346: out = 24'(3776);
			33347: out = 24'(-284);
			33348: out = 24'(616);
			33349: out = 24'(8124);
			33350: out = 24'(12788);
			33351: out = 24'(6668);
			33352: out = 24'(-7596);
			33353: out = 24'(-8508);
			33354: out = 24'(-2692);
			33355: out = 24'(1952);
			33356: out = 24'(-240);
			33357: out = 24'(1812);
			33358: out = 24'(1640);
			33359: out = 24'(1320);
			33360: out = 24'(-512);
			33361: out = 24'(-3328);
			33362: out = 24'(-1804);
			33363: out = 24'(2764);
			33364: out = 24'(3892);
			33365: out = 24'(-3388);
			33366: out = 24'(-9776);
			33367: out = 24'(-9364);
			33368: out = 24'(-3228);
			33369: out = 24'(256);
			33370: out = 24'(4888);
			33371: out = 24'(3952);
			33372: out = 24'(1528);
			33373: out = 24'(1776);
			33374: out = 24'(-1540);
			33375: out = 24'(-1816);
			33376: out = 24'(-1888);
			33377: out = 24'(-1812);
			33378: out = 24'(-5188);
			33379: out = 24'(-512);
			33380: out = 24'(4136);
			33381: out = 24'(4432);
			33382: out = 24'(-3112);
			33383: out = 24'(-1036);
			33384: out = 24'(3396);
			33385: out = 24'(7396);
			33386: out = 24'(4544);
			33387: out = 24'(7208);
			33388: out = 24'(1192);
			33389: out = 24'(-5024);
			33390: out = 24'(-5472);
			33391: out = 24'(-652);
			33392: out = 24'(-4188);
			33393: out = 24'(-5936);
			33394: out = 24'(1676);
			33395: out = 24'(5972);
			33396: out = 24'(4128);
			33397: out = 24'(2672);
			33398: out = 24'(6948);
			33399: out = 24'(-332);
			33400: out = 24'(-932);
			33401: out = 24'(-3396);
			33402: out = 24'(-3300);
			33403: out = 24'(-2384);
			33404: out = 24'(1436);
			33405: out = 24'(1052);
			33406: out = 24'(348);
			33407: out = 24'(1788);
			33408: out = 24'(4544);
			33409: out = 24'(2644);
			33410: out = 24'(-1328);
			33411: out = 24'(-1712);
			33412: out = 24'(-796);
			33413: out = 24'(496);
			33414: out = 24'(-3100);
			33415: out = 24'(-7600);
			33416: out = 24'(-5948);
			33417: out = 24'(-1432);
			33418: out = 24'(616);
			33419: out = 24'(744);
			33420: out = 24'(4980);
			33421: out = 24'(5368);
			33422: out = 24'(1272);
			33423: out = 24'(-6100);
			33424: out = 24'(-8604);
			33425: out = 24'(-2624);
			33426: out = 24'(6536);
			33427: out = 24'(7880);
			33428: out = 24'(-776);
			33429: out = 24'(-3000);
			33430: out = 24'(-4228);
			33431: out = 24'(-2972);
			33432: out = 24'(-1228);
			33433: out = 24'(6340);
			33434: out = 24'(6728);
			33435: out = 24'(6756);
			33436: out = 24'(4916);
			33437: out = 24'(-5084);
			33438: out = 24'(-12816);
			33439: out = 24'(-13760);
			33440: out = 24'(-6608);
			33441: out = 24'(-2152);
			33442: out = 24'(4696);
			33443: out = 24'(6128);
			33444: out = 24'(7120);
			33445: out = 24'(4184);
			33446: out = 24'(3604);
			33447: out = 24'(-6624);
			33448: out = 24'(-9248);
			33449: out = 24'(1548);
			33450: out = 24'(10008);
			33451: out = 24'(2888);
			33452: out = 24'(-9428);
			33453: out = 24'(-10968);
			33454: out = 24'(3836);
			33455: out = 24'(6160);
			33456: out = 24'(2584);
			33457: out = 24'(-140);
			33458: out = 24'(-60);
			33459: out = 24'(-1336);
			33460: out = 24'(-5624);
			33461: out = 24'(-10200);
			33462: out = 24'(-5744);
			33463: out = 24'(5744);
			33464: out = 24'(15780);
			33465: out = 24'(7800);
			33466: out = 24'(-10220);
			33467: out = 24'(-15684);
			33468: out = 24'(-2284);
			33469: out = 24'(5992);
			33470: out = 24'(568);
			33471: out = 24'(628);
			33472: out = 24'(6552);
			33473: out = 24'(9724);
			33474: out = 24'(4016);
			33475: out = 24'(-5340);
			33476: out = 24'(-744);
			33477: out = 24'(1136);
			33478: out = 24'(-812);
			33479: out = 24'(196);
			33480: out = 24'(4208);
			33481: out = 24'(2412);
			33482: out = 24'(348);
			33483: out = 24'(4820);
			33484: out = 24'(-1324);
			33485: out = 24'(-7552);
			33486: out = 24'(-7068);
			33487: out = 24'(1940);
			33488: out = 24'(-4152);
			33489: out = 24'(-1504);
			33490: out = 24'(3936);
			33491: out = 24'(9400);
			33492: out = 24'(1216);
			33493: out = 24'(-1076);
			33494: out = 24'(-2192);
			33495: out = 24'(1612);
			33496: out = 24'(3892);
			33497: out = 24'(-1416);
			33498: out = 24'(-8652);
			33499: out = 24'(-6760);
			33500: out = 24'(1468);
			33501: out = 24'(6512);
			33502: out = 24'(420);
			33503: out = 24'(-5728);
			33504: out = 24'(-4840);
			33505: out = 24'(1148);
			33506: out = 24'(1716);
			33507: out = 24'(3484);
			33508: out = 24'(6140);
			33509: out = 24'(-88);
			33510: out = 24'(-1840);
			33511: out = 24'(-1400);
			33512: out = 24'(36);
			33513: out = 24'(-716);
			33514: out = 24'(-7948);
			33515: out = 24'(-5108);
			33516: out = 24'(5584);
			33517: out = 24'(8400);
			33518: out = 24'(6696);
			33519: out = 24'(-824);
			33520: out = 24'(1008);
			33521: out = 24'(9384);
			33522: out = 24'(5176);
			33523: out = 24'(-7012);
			33524: out = 24'(-17484);
			33525: out = 24'(-14980);
			33526: out = 24'(-1796);
			33527: out = 24'(4740);
			33528: out = 24'(3468);
			33529: out = 24'(1484);
			33530: out = 24'(-384);
			33531: out = 24'(536);
			33532: out = 24'(-3928);
			33533: out = 24'(-8928);
			33534: out = 24'(-10968);
			33535: out = 24'(3012);
			33536: out = 24'(4256);
			33537: out = 24'(364);
			33538: out = 24'(1008);
			33539: out = 24'(5516);
			33540: out = 24'(2976);
			33541: out = 24'(-3196);
			33542: out = 24'(-4196);
			33543: out = 24'(-424);
			33544: out = 24'(5016);
			33545: out = 24'(4600);
			33546: out = 24'(524);
			33547: out = 24'(1648);
			33548: out = 24'(840);
			33549: out = 24'(1256);
			33550: out = 24'(-1120);
			33551: out = 24'(-1248);
			33552: out = 24'(-1216);
			33553: out = 24'(6680);
			33554: out = 24'(8072);
			33555: out = 24'(-1084);
			33556: out = 24'(-3332);
			33557: out = 24'(976);
			33558: out = 24'(5972);
			33559: out = 24'(4704);
			33560: out = 24'(228);
			33561: out = 24'(-1944);
			33562: out = 24'(-3684);
			33563: out = 24'(-5468);
			33564: out = 24'(-2172);
			33565: out = 24'(-604);
			33566: out = 24'(-168);
			33567: out = 24'(712);
			33568: out = 24'(4472);
			33569: out = 24'(4512);
			33570: out = 24'(1088);
			33571: out = 24'(-5164);
			33572: out = 24'(-10676);
			33573: out = 24'(-4616);
			33574: out = 24'(-1412);
			33575: out = 24'(3056);
			33576: out = 24'(9024);
			33577: out = 24'(4608);
			33578: out = 24'(-2932);
			33579: out = 24'(-10152);
			33580: out = 24'(-8700);
			33581: out = 24'(-780);
			33582: out = 24'(4292);
			33583: out = 24'(2388);
			33584: out = 24'(132);
			33585: out = 24'(4752);
			33586: out = 24'(956);
			33587: out = 24'(-2904);
			33588: out = 24'(-5800);
			33589: out = 24'(-4652);
			33590: out = 24'(-2636);
			33591: out = 24'(504);
			33592: out = 24'(1268);
			33593: out = 24'(300);
			33594: out = 24'(56);
			33595: out = 24'(3212);
			33596: out = 24'(5340);
			33597: out = 24'(3816);
			33598: out = 24'(324);
			33599: out = 24'(-6120);
			33600: out = 24'(-10584);
			33601: out = 24'(-8044);
			33602: out = 24'(1372);
			33603: out = 24'(4700);
			33604: out = 24'(3448);
			33605: out = 24'(2176);
			33606: out = 24'(4808);
			33607: out = 24'(1156);
			33608: out = 24'(-4968);
			33609: out = 24'(-8732);
			33610: out = 24'(-3892);
			33611: out = 24'(-4208);
			33612: out = 24'(688);
			33613: out = 24'(1936);
			33614: out = 24'(2704);
			33615: out = 24'(5652);
			33616: out = 24'(7104);
			33617: out = 24'(1840);
			33618: out = 24'(-4316);
			33619: out = 24'(-5096);
			33620: out = 24'(2680);
			33621: out = 24'(3284);
			33622: out = 24'(-552);
			33623: out = 24'(1848);
			33624: out = 24'(1292);
			33625: out = 24'(136);
			33626: out = 24'(-3880);
			33627: out = 24'(-6660);
			33628: out = 24'(-4128);
			33629: out = 24'(-284);
			33630: out = 24'(2100);
			33631: out = 24'(1376);
			33632: out = 24'(-1176);
			33633: out = 24'(-1080);
			33634: out = 24'(4280);
			33635: out = 24'(8912);
			33636: out = 24'(4640);
			33637: out = 24'(-1620);
			33638: out = 24'(-2944);
			33639: out = 24'(1600);
			33640: out = 24'(4032);
			33641: out = 24'(1080);
			33642: out = 24'(1220);
			33643: out = 24'(7040);
			33644: out = 24'(8900);
			33645: out = 24'(5956);
			33646: out = 24'(-2668);
			33647: out = 24'(-4656);
			33648: out = 24'(200);
			33649: out = 24'(3924);
			33650: out = 24'(924);
			33651: out = 24'(-1200);
			33652: out = 24'(-376);
			33653: out = 24'(-424);
			33654: out = 24'(-4508);
			33655: out = 24'(-3968);
			33656: out = 24'(1276);
			33657: out = 24'(3780);
			33658: out = 24'(812);
			33659: out = 24'(-1912);
			33660: out = 24'(-1980);
			33661: out = 24'(-116);
			33662: out = 24'(544);
			33663: out = 24'(4060);
			33664: out = 24'(4112);
			33665: out = 24'(-1412);
			33666: out = 24'(-3708);
			33667: out = 24'(-4464);
			33668: out = 24'(-4096);
			33669: out = 24'(-3552);
			33670: out = 24'(-612);
			33671: out = 24'(4252);
			33672: out = 24'(3900);
			33673: out = 24'(-2716);
			33674: out = 24'(-8444);
			33675: out = 24'(-5820);
			33676: out = 24'(-932);
			33677: out = 24'(-720);
			33678: out = 24'(-1604);
			33679: out = 24'(-4148);
			33680: out = 24'(3244);
			33681: out = 24'(11664);
			33682: out = 24'(12532);
			33683: out = 24'(2536);
			33684: out = 24'(-4268);
			33685: out = 24'(-4408);
			33686: out = 24'(716);
			33687: out = 24'(3364);
			33688: out = 24'(2648);
			33689: out = 24'(-2808);
			33690: out = 24'(-4732);
			33691: out = 24'(748);
			33692: out = 24'(4176);
			33693: out = 24'(336);
			33694: out = 24'(-4588);
			33695: out = 24'(-2240);
			33696: out = 24'(-7756);
			33697: out = 24'(-9968);
			33698: out = 24'(-5016);
			33699: out = 24'(5368);
			33700: out = 24'(8396);
			33701: out = 24'(7072);
			33702: out = 24'(5476);
			33703: out = 24'(5232);
			33704: out = 24'(4504);
			33705: out = 24'(-8436);
			33706: out = 24'(-16428);
			33707: out = 24'(-8552);
			33708: out = 24'(4596);
			33709: out = 24'(9172);
			33710: out = 24'(6212);
			33711: out = 24'(3780);
			33712: out = 24'(504);
			33713: out = 24'(500);
			33714: out = 24'(-5468);
			33715: out = 24'(-9868);
			33716: out = 24'(-8492);
			33717: out = 24'(-1248);
			33718: out = 24'(272);
			33719: out = 24'(248);
			33720: out = 24'(1676);
			33721: out = 24'(1388);
			33722: out = 24'(412);
			33723: out = 24'(-1500);
			33724: out = 24'(-3744);
			33725: out = 24'(1440);
			33726: out = 24'(-312);
			33727: out = 24'(2884);
			33728: out = 24'(5804);
			33729: out = 24'(4396);
			33730: out = 24'(-5276);
			33731: out = 24'(-4456);
			33732: out = 24'(1900);
			33733: out = 24'(4096);
			33734: out = 24'(468);
			33735: out = 24'(-348);
			33736: out = 24'(-3056);
			33737: out = 24'(-8716);
			33738: out = 24'(-916);
			33739: out = 24'(6332);
			33740: out = 24'(5864);
			33741: out = 24'(-3976);
			33742: out = 24'(-2852);
			33743: out = 24'(-1968);
			33744: out = 24'(920);
			33745: out = 24'(-1408);
			33746: out = 24'(-952);
			33747: out = 24'(2728);
			33748: out = 24'(12688);
			33749: out = 24'(13412);
			33750: out = 24'(3472);
			33751: out = 24'(-7928);
			33752: out = 24'(-6152);
			33753: out = 24'(-1744);
			33754: out = 24'(-2932);
			33755: out = 24'(-7236);
			33756: out = 24'(-180);
			33757: out = 24'(4744);
			33758: out = 24'(-672);
			33759: out = 24'(-6280);
			33760: out = 24'(-2588);
			33761: out = 24'(3984);
			33762: out = 24'(2404);
			33763: out = 24'(-3260);
			33764: out = 24'(-9944);
			33765: out = 24'(-7960);
			33766: out = 24'(-744);
			33767: out = 24'(5848);
			33768: out = 24'(1288);
			33769: out = 24'(-1800);
			33770: out = 24'(112);
			33771: out = 24'(6364);
			33772: out = 24'(4492);
			33773: out = 24'(-1156);
			33774: out = 24'(-8256);
			33775: out = 24'(-7204);
			33776: out = 24'(-1600);
			33777: out = 24'(6716);
			33778: out = 24'(2440);
			33779: out = 24'(-6520);
			33780: out = 24'(-6908);
			33781: out = 24'(944);
			33782: out = 24'(1748);
			33783: out = 24'(-2548);
			33784: out = 24'(372);
			33785: out = 24'(3672);
			33786: out = 24'(2872);
			33787: out = 24'(-1384);
			33788: out = 24'(-1808);
			33789: out = 24'(-6612);
			33790: out = 24'(-7052);
			33791: out = 24'(-4768);
			33792: out = 24'(1292);
			33793: out = 24'(-188);
			33794: out = 24'(3804);
			33795: out = 24'(5200);
			33796: out = 24'(4020);
			33797: out = 24'(-1708);
			33798: out = 24'(696);
			33799: out = 24'(1656);
			33800: out = 24'(-3232);
			33801: out = 24'(-17900);
			33802: out = 24'(-12044);
			33803: out = 24'(-4564);
			33804: out = 24'(5232);
			33805: out = 24'(14644);
			33806: out = 24'(14916);
			33807: out = 24'(6972);
			33808: out = 24'(-1536);
			33809: out = 24'(-5856);
			33810: out = 24'(-11488);
			33811: out = 24'(-9628);
			33812: out = 24'(-136);
			33813: out = 24'(11104);
			33814: out = 24'(13636);
			33815: out = 24'(10960);
			33816: out = 24'(4580);
			33817: out = 24'(-1792);
			33818: out = 24'(-5024);
			33819: out = 24'(-7200);
			33820: out = 24'(-5076);
			33821: out = 24'(-3480);
			33822: out = 24'(-2952);
			33823: out = 24'(-796);
			33824: out = 24'(3724);
			33825: out = 24'(2972);
			33826: out = 24'(-1868);
			33827: out = 24'(-3808);
			33828: out = 24'(4920);
			33829: out = 24'(8724);
			33830: out = 24'(3236);
			33831: out = 24'(-1460);
			33832: out = 24'(2352);
			33833: out = 24'(4116);
			33834: out = 24'(156);
			33835: out = 24'(-1672);
			33836: out = 24'(412);
			33837: out = 24'(288);
			33838: out = 24'(-3436);
			33839: out = 24'(-5064);
			33840: out = 24'(-4152);
			33841: out = 24'(-1612);
			33842: out = 24'(2072);
			33843: out = 24'(6076);
			33844: out = 24'(6272);
			33845: out = 24'(2028);
			33846: out = 24'(-228);
			33847: out = 24'(676);
			33848: out = 24'(-4948);
			33849: out = 24'(-6024);
			33850: out = 24'(-1412);
			33851: out = 24'(5624);
			33852: out = 24'(5528);
			33853: out = 24'(1596);
			33854: out = 24'(-1020);
			33855: out = 24'(-488);
			33856: out = 24'(-2588);
			33857: out = 24'(-636);
			33858: out = 24'(-412);
			33859: out = 24'(304);
			33860: out = 24'(1736);
			33861: out = 24'(7460);
			33862: out = 24'(7076);
			33863: out = 24'(-1540);
			33864: out = 24'(-12888);
			33865: out = 24'(-6164);
			33866: out = 24'(2024);
			33867: out = 24'(6828);
			33868: out = 24'(2656);
			33869: out = 24'(532);
			33870: out = 24'(-6620);
			33871: out = 24'(-3460);
			33872: out = 24'(1808);
			33873: out = 24'(-380);
			33874: out = 24'(-4416);
			33875: out = 24'(-3304);
			33876: out = 24'(2016);
			33877: out = 24'(5792);
			33878: out = 24'(5912);
			33879: out = 24'(5056);
			33880: out = 24'(2668);
			33881: out = 24'(-856);
			33882: out = 24'(-6952);
			33883: out = 24'(-2440);
			33884: out = 24'(1092);
			33885: out = 24'(-4396);
			33886: out = 24'(-12884);
			33887: out = 24'(-8644);
			33888: out = 24'(5436);
			33889: out = 24'(14164);
			33890: out = 24'(9780);
			33891: out = 24'(-1652);
			33892: out = 24'(-7556);
			33893: out = 24'(-2244);
			33894: out = 24'(5040);
			33895: out = 24'(236);
			33896: out = 24'(-8420);
			33897: out = 24'(-7232);
			33898: out = 24'(5716);
			33899: out = 24'(9112);
			33900: out = 24'(7016);
			33901: out = 24'(1672);
			33902: out = 24'(-684);
			33903: out = 24'(-2564);
			33904: out = 24'(-4712);
			33905: out = 24'(-5756);
			33906: out = 24'(-2840);
			33907: out = 24'(-844);
			33908: out = 24'(3764);
			33909: out = 24'(2272);
			33910: out = 24'(-576);
			33911: out = 24'(1168);
			33912: out = 24'(4740);
			33913: out = 24'(3832);
			33914: out = 24'(-1556);
			33915: out = 24'(-3804);
			33916: out = 24'(-7540);
			33917: out = 24'(-4380);
			33918: out = 24'(-8);
			33919: out = 24'(4828);
			33920: out = 24'(-744);
			33921: out = 24'(1460);
			33922: out = 24'(-2724);
			33923: out = 24'(-6876);
			33924: out = 24'(-2812);
			33925: out = 24'(6992);
			33926: out = 24'(2468);
			33927: out = 24'(-9628);
			33928: out = 24'(-7984);
			33929: out = 24'(-2308);
			33930: out = 24'(1168);
			33931: out = 24'(-612);
			33932: out = 24'(292);
			33933: out = 24'(-3332);
			33934: out = 24'(-4632);
			33935: out = 24'(-3960);
			33936: out = 24'(1060);
			33937: out = 24'(1176);
			33938: out = 24'(3948);
			33939: out = 24'(6172);
			33940: out = 24'(9040);
			33941: out = 24'(5392);
			33942: out = 24'(2092);
			33943: out = 24'(-4188);
			33944: out = 24'(-8104);
			33945: out = 24'(-12508);
			33946: out = 24'(5908);
			33947: out = 24'(9964);
			33948: out = 24'(1924);
			33949: out = 24'(-6836);
			33950: out = 24'(20);
			33951: out = 24'(2024);
			33952: out = 24'(448);
			33953: out = 24'(324);
			33954: out = 24'(4000);
			33955: out = 24'(2776);
			33956: out = 24'(440);
			33957: out = 24'(-752);
			33958: out = 24'(-5156);
			33959: out = 24'(-3768);
			33960: out = 24'(2916);
			33961: out = 24'(9780);
			33962: out = 24'(9468);
			33963: out = 24'(5592);
			33964: out = 24'(2200);
			33965: out = 24'(-1212);
			33966: out = 24'(-10092);
			33967: out = 24'(-11924);
			33968: out = 24'(-12520);
			33969: out = 24'(-7352);
			33970: out = 24'(1524);
			33971: out = 24'(12484);
			33972: out = 24'(12604);
			33973: out = 24'(5604);
			33974: out = 24'(-1116);
			33975: out = 24'(-2372);
			33976: out = 24'(-4820);
			33977: out = 24'(-5160);
			33978: out = 24'(-368);
			33979: out = 24'(3284);
			33980: out = 24'(4580);
			33981: out = 24'(-6176);
			33982: out = 24'(-14224);
			33983: out = 24'(-4268);
			33984: out = 24'(6112);
			33985: out = 24'(7940);
			33986: out = 24'(1732);
			33987: out = 24'(732);
			33988: out = 24'(2868);
			33989: out = 24'(5644);
			33990: out = 24'(-760);
			33991: out = 24'(-10096);
			33992: out = 24'(-14348);
			33993: out = 24'(-4852);
			33994: out = 24'(3352);
			33995: out = 24'(3568);
			33996: out = 24'(-1592);
			33997: out = 24'(360);
			33998: out = 24'(3348);
			33999: out = 24'(4656);
			34000: out = 24'(4228);
			34001: out = 24'(-564);
			34002: out = 24'(-4576);
			34003: out = 24'(-3948);
			34004: out = 24'(76);
			34005: out = 24'(184);
			34006: out = 24'(-396);
			34007: out = 24'(2116);
			34008: out = 24'(5588);
			34009: out = 24'(608);
			34010: out = 24'(-4232);
			34011: out = 24'(-3176);
			34012: out = 24'(2216);
			34013: out = 24'(948);
			34014: out = 24'(-2360);
			34015: out = 24'(-2344);
			34016: out = 24'(2264);
			34017: out = 24'(844);
			34018: out = 24'(960);
			34019: out = 24'(-2596);
			34020: out = 24'(-2820);
			34021: out = 24'(-112);
			34022: out = 24'(228);
			34023: out = 24'(-496);
			34024: out = 24'(1872);
			34025: out = 24'(6020);
			34026: out = 24'(6056);
			34027: out = 24'(-2092);
			34028: out = 24'(-11292);
			34029: out = 24'(-13336);
			34030: out = 24'(-7408);
			34031: out = 24'(-1584);
			34032: out = 24'(2600);
			34033: out = 24'(5528);
			34034: out = 24'(6096);
			34035: out = 24'(9304);
			34036: out = 24'(10004);
			34037: out = 24'(6016);
			34038: out = 24'(-3060);
			34039: out = 24'(-13784);
			34040: out = 24'(-15796);
			34041: out = 24'(-7264);
			34042: out = 24'(2452);
			34043: out = 24'(10068);
			34044: out = 24'(6796);
			34045: out = 24'(4236);
			34046: out = 24'(3920);
			34047: out = 24'(368);
			34048: out = 24'(-7708);
			34049: out = 24'(-9752);
			34050: out = 24'(-3368);
			34051: out = 24'(-508);
			34052: out = 24'(676);
			34053: out = 24'(-888);
			34054: out = 24'(-2700);
			34055: out = 24'(-6816);
			34056: out = 24'(-924);
			34057: out = 24'(2928);
			34058: out = 24'(6360);
			34059: out = 24'(8504);
			34060: out = 24'(1400);
			34061: out = 24'(-5528);
			34062: out = 24'(-9676);
			34063: out = 24'(-7360);
			34064: out = 24'(-2696);
			34065: out = 24'(6124);
			34066: out = 24'(10484);
			34067: out = 24'(9040);
			34068: out = 24'(128);
			34069: out = 24'(3364);
			34070: out = 24'(3112);
			34071: out = 24'(-2072);
			34072: out = 24'(-6684);
			34073: out = 24'(-3556);
			34074: out = 24'(1836);
			34075: out = 24'(5512);
			34076: out = 24'(5128);
			34077: out = 24'(-3204);
			34078: out = 24'(-7120);
			34079: out = 24'(68);
			34080: out = 24'(9772);
			34081: out = 24'(1244);
			34082: out = 24'(-5788);
			34083: out = 24'(-2812);
			34084: out = 24'(6944);
			34085: out = 24'(3900);
			34086: out = 24'(-3432);
			34087: out = 24'(-9068);
			34088: out = 24'(-4940);
			34089: out = 24'(-780);
			34090: out = 24'(5424);
			34091: out = 24'(3904);
			34092: out = 24'(-260);
			34093: out = 24'(-5724);
			34094: out = 24'(-4980);
			34095: out = 24'(-6748);
			34096: out = 24'(-4524);
			34097: out = 24'(2092);
			34098: out = 24'(4624);
			34099: out = 24'(2004);
			34100: out = 24'(-436);
			34101: out = 24'(352);
			34102: out = 24'(36);
			34103: out = 24'(-1280);
			34104: out = 24'(-844);
			34105: out = 24'(1244);
			34106: out = 24'(-3764);
			34107: out = 24'(3016);
			34108: out = 24'(5476);
			34109: out = 24'(2764);
			34110: out = 24'(-3536);
			34111: out = 24'(-644);
			34112: out = 24'(504);
			34113: out = 24'(-1412);
			34114: out = 24'(-5092);
			34115: out = 24'(-364);
			34116: out = 24'(484);
			34117: out = 24'(-592);
			34118: out = 24'(-1572);
			34119: out = 24'(1180);
			34120: out = 24'(3788);
			34121: out = 24'(5084);
			34122: out = 24'(3760);
			34123: out = 24'(168);
			34124: out = 24'(-5268);
			34125: out = 24'(-7792);
			34126: out = 24'(-4900);
			34127: out = 24'(1948);
			34128: out = 24'(4316);
			34129: out = 24'(4952);
			34130: out = 24'(3528);
			34131: out = 24'(-108);
			34132: out = 24'(4116);
			34133: out = 24'(2128);
			34134: out = 24'(-2348);
			34135: out = 24'(-4924);
			34136: out = 24'(1016);
			34137: out = 24'(3612);
			34138: out = 24'(5332);
			34139: out = 24'(5064);
			34140: out = 24'(-48);
			34141: out = 24'(-2972);
			34142: out = 24'(-4812);
			34143: out = 24'(-5844);
			34144: out = 24'(-6848);
			34145: out = 24'(-1632);
			34146: out = 24'(3104);
			34147: out = 24'(4084);
			34148: out = 24'(1616);
			34149: out = 24'(5108);
			34150: out = 24'(6464);
			34151: out = 24'(2784);
			34152: out = 24'(-4860);
			34153: out = 24'(-6876);
			34154: out = 24'(-3284);
			34155: out = 24'(2616);
			34156: out = 24'(3768);
			34157: out = 24'(1920);
			34158: out = 24'(-2860);
			34159: out = 24'(-2684);
			34160: out = 24'(-468);
			34161: out = 24'(-2248);
			34162: out = 24'(-2172);
			34163: out = 24'(-976);
			34164: out = 24'(-576);
			34165: out = 24'(-3968);
			34166: out = 24'(-6448);
			34167: out = 24'(-3572);
			34168: out = 24'(2772);
			34169: out = 24'(4160);
			34170: out = 24'(6788);
			34171: out = 24'(-1496);
			34172: out = 24'(-5372);
			34173: out = 24'(-460);
			34174: out = 24'(3848);
			34175: out = 24'(2932);
			34176: out = 24'(128);
			34177: out = 24'(-440);
			34178: out = 24'(-2484);
			34179: out = 24'(-1636);
			34180: out = 24'(-3940);
			34181: out = 24'(-4980);
			34182: out = 24'(-3336);
			34183: out = 24'(4676);
			34184: out = 24'(6048);
			34185: out = 24'(3032);
			34186: out = 24'(-160);
			34187: out = 24'(1120);
			34188: out = 24'(-784);
			34189: out = 24'(-3432);
			34190: out = 24'(-5208);
			34191: out = 24'(-1940);
			34192: out = 24'(-104);
			34193: out = 24'(3388);
			34194: out = 24'(3788);
			34195: out = 24'(540);
			34196: out = 24'(-3520);
			34197: out = 24'(288);
			34198: out = 24'(4600);
			34199: out = 24'(1168);
			34200: out = 24'(-8648);
			34201: out = 24'(-5816);
			34202: out = 24'(5308);
			34203: out = 24'(7796);
			34204: out = 24'(5940);
			34205: out = 24'(-328);
			34206: out = 24'(-1996);
			34207: out = 24'(-552);
			34208: out = 24'(-100);
			34209: out = 24'(-3348);
			34210: out = 24'(-5836);
			34211: out = 24'(-3212);
			34212: out = 24'(4956);
			34213: out = 24'(5032);
			34214: out = 24'(2096);
			34215: out = 24'(1496);
			34216: out = 24'(3720);
			34217: out = 24'(5340);
			34218: out = 24'(1280);
			34219: out = 24'(-3752);
			34220: out = 24'(-4800);
			34221: out = 24'(3824);
			34222: out = 24'(2640);
			34223: out = 24'(-2496);
			34224: out = 24'(-2808);
			34225: out = 24'(2916);
			34226: out = 24'(1776);
			34227: out = 24'(-3084);
			34228: out = 24'(-4940);
			34229: out = 24'(-4108);
			34230: out = 24'(-2284);
			34231: out = 24'(-1524);
			34232: out = 24'(1072);
			34233: out = 24'(3516);
			34234: out = 24'(5688);
			34235: out = 24'(2204);
			34236: out = 24'(-1328);
			34237: out = 24'(-3956);
			34238: out = 24'(-1808);
			34239: out = 24'(-5168);
			34240: out = 24'(-4992);
			34241: out = 24'(1120);
			34242: out = 24'(11816);
			34243: out = 24'(5076);
			34244: out = 24'(-3632);
			34245: out = 24'(-4148);
			34246: out = 24'(648);
			34247: out = 24'(-884);
			34248: out = 24'(-1804);
			34249: out = 24'(180);
			34250: out = 24'(-504);
			34251: out = 24'(528);
			34252: out = 24'(2444);
			34253: out = 24'(3052);
			34254: out = 24'(-2464);
			34255: out = 24'(496);
			34256: out = 24'(1444);
			34257: out = 24'(-1916);
			34258: out = 24'(-10272);
			34259: out = 24'(-1120);
			34260: out = 24'(1884);
			34261: out = 24'(1968);
			34262: out = 24'(-772);
			34263: out = 24'(60);
			34264: out = 24'(-540);
			34265: out = 24'(172);
			34266: out = 24'(-1068);
			34267: out = 24'(-3000);
			34268: out = 24'(-1744);
			34269: out = 24'(4496);
			34270: out = 24'(6752);
			34271: out = 24'(-692);
			34272: out = 24'(-5716);
			34273: out = 24'(-3696);
			34274: out = 24'(960);
			34275: out = 24'(-884);
			34276: out = 24'(-1076);
			34277: out = 24'(-2560);
			34278: out = 24'(-772);
			34279: out = 24'(268);
			34280: out = 24'(7960);
			34281: out = 24'(2428);
			34282: out = 24'(-2900);
			34283: out = 24'(-4712);
			34284: out = 24'(1200);
			34285: out = 24'(-608);
			34286: out = 24'(2408);
			34287: out = 24'(4776);
			34288: out = 24'(-412);
			34289: out = 24'(-5560);
			34290: out = 24'(-4724);
			34291: out = 24'(-1800);
			34292: out = 24'(-5456);
			34293: out = 24'(-4524);
			34294: out = 24'(-3364);
			34295: out = 24'(-228);
			34296: out = 24'(2416);
			34297: out = 24'(10928);
			34298: out = 24'(8508);
			34299: out = 24'(-264);
			34300: out = 24'(-8648);
			34301: out = 24'(-3408);
			34302: out = 24'(-2396);
			34303: out = 24'(-524);
			34304: out = 24'(2124);
			34305: out = 24'(5556);
			34306: out = 24'(11132);
			34307: out = 24'(11264);
			34308: out = 24'(3904);
			34309: out = 24'(-5272);
			34310: out = 24'(-3340);
			34311: out = 24'(-680);
			34312: out = 24'(-2752);
			34313: out = 24'(-6196);
			34314: out = 24'(2500);
			34315: out = 24'(7244);
			34316: out = 24'(4960);
			34317: out = 24'(-1236);
			34318: out = 24'(-308);
			34319: out = 24'(-636);
			34320: out = 24'(-1124);
			34321: out = 24'(-2532);
			34322: out = 24'(-2176);
			34323: out = 24'(-1272);
			34324: out = 24'(-532);
			34325: out = 24'(-816);
			34326: out = 24'(-16);
			34327: out = 24'(2760);
			34328: out = 24'(4976);
			34329: out = 24'(3856);
			34330: out = 24'(272);
			34331: out = 24'(-6116);
			34332: out = 24'(-5764);
			34333: out = 24'(-1808);
			34334: out = 24'(400);
			34335: out = 24'(-1844);
			34336: out = 24'(-440);
			34337: out = 24'(2720);
			34338: out = 24'(3204);
			34339: out = 24'(1368);
			34340: out = 24'(-4060);
			34341: out = 24'(-3068);
			34342: out = 24'(3352);
			34343: out = 24'(8420);
			34344: out = 24'(5136);
			34345: out = 24'(808);
			34346: out = 24'(-1252);
			34347: out = 24'(-2752);
			34348: out = 24'(-5088);
			34349: out = 24'(-4188);
			34350: out = 24'(-1060);
			34351: out = 24'(-848);
			34352: out = 24'(-40);
			34353: out = 24'(-2088);
			34354: out = 24'(-1336);
			34355: out = 24'(-836);
			34356: out = 24'(-1700);
			34357: out = 24'(-7424);
			34358: out = 24'(-4780);
			34359: out = 24'(3488);
			34360: out = 24'(7324);
			34361: out = 24'(1780);
			34362: out = 24'(-2924);
			34363: out = 24'(-2932);
			34364: out = 24'(-124);
			34365: out = 24'(-612);
			34366: out = 24'(112);
			34367: out = 24'(-1980);
			34368: out = 24'(-4684);
			34369: out = 24'(-1184);
			34370: out = 24'(8584);
			34371: out = 24'(11320);
			34372: out = 24'(2364);
			34373: out = 24'(-5792);
			34374: out = 24'(-5796);
			34375: out = 24'(-1428);
			34376: out = 24'(-756);
			34377: out = 24'(88);
			34378: out = 24'(-1024);
			34379: out = 24'(2840);
			34380: out = 24'(3968);
			34381: out = 24'(-2868);
			34382: out = 24'(-4716);
			34383: out = 24'(-4940);
			34384: out = 24'(-2344);
			34385: out = 24'(84);
			34386: out = 24'(4784);
			34387: out = 24'(5328);
			34388: out = 24'(4772);
			34389: out = 24'(2948);
			34390: out = 24'(-116);
			34391: out = 24'(-2204);
			34392: out = 24'(-1516);
			34393: out = 24'(-744);
			34394: out = 24'(-2224);
			34395: out = 24'(-4872);
			34396: out = 24'(-3212);
			34397: out = 24'(1132);
			34398: out = 24'(3692);
			34399: out = 24'(3944);
			34400: out = 24'(2388);
			34401: out = 24'(-2056);
			34402: out = 24'(-8792);
			34403: out = 24'(-4164);
			34404: out = 24'(-1468);
			34405: out = 24'(1364);
			34406: out = 24'(4372);
			34407: out = 24'(3632);
			34408: out = 24'(4256);
			34409: out = 24'(1364);
			34410: out = 24'(-3156);
			34411: out = 24'(-5216);
			34412: out = 24'(-548);
			34413: out = 24'(1092);
			34414: out = 24'(-956);
			34415: out = 24'(72);
			34416: out = 24'(-704);
			34417: out = 24'(-776);
			34418: out = 24'(-3844);
			34419: out = 24'(-6296);
			34420: out = 24'(-3068);
			34421: out = 24'(2304);
			34422: out = 24'(3580);
			34423: out = 24'(936);
			34424: out = 24'(1180);
			34425: out = 24'(-2468);
			34426: out = 24'(-9064);
			34427: out = 24'(-11972);
			34428: out = 24'(-2136);
			34429: out = 24'(3308);
			34430: out = 24'(2840);
			34431: out = 24'(-836);
			34432: out = 24'(692);
			34433: out = 24'(7300);
			34434: out = 24'(8156);
			34435: out = 24'(380);
			34436: out = 24'(-4112);
			34437: out = 24'(-5036);
			34438: out = 24'(2372);
			34439: out = 24'(976);
			34440: out = 24'(-6612);
			34441: out = 24'(-4128);
			34442: out = 24'(7036);
			34443: out = 24'(11740);
			34444: out = 24'(6012);
			34445: out = 24'(184);
			34446: out = 24'(-4804);
			34447: out = 24'(-11836);
			34448: out = 24'(-15432);
			34449: out = 24'(-2500);
			34450: out = 24'(2708);
			34451: out = 24'(5276);
			34452: out = 24'(4232);
			34453: out = 24'(6064);
			34454: out = 24'(7352);
			34455: out = 24'(7152);
			34456: out = 24'(1832);
			34457: out = 24'(-5780);
			34458: out = 24'(-6348);
			34459: out = 24'(-8088);
			34460: out = 24'(-5652);
			34461: out = 24'(1652);
			34462: out = 24'(8656);
			34463: out = 24'(6316);
			34464: out = 24'(1452);
			34465: out = 24'(-84);
			34466: out = 24'(-492);
			34467: out = 24'(304);
			34468: out = 24'(-2824);
			34469: out = 24'(-4172);
			34470: out = 24'(1744);
			34471: out = 24'(7568);
			34472: out = 24'(10148);
			34473: out = 24'(5988);
			34474: out = 24'(-1280);
			34475: out = 24'(-7816);
			34476: out = 24'(-7120);
			34477: out = 24'(-3072);
			34478: out = 24'(-44);
			34479: out = 24'(-332);
			34480: out = 24'(648);
			34481: out = 24'(2208);
			34482: out = 24'(4236);
			34483: out = 24'(3284);
			34484: out = 24'(-4560);
			34485: out = 24'(-13480);
			34486: out = 24'(-11796);
			34487: out = 24'(-4);
			34488: out = 24'(8536);
			34489: out = 24'(4384);
			34490: out = 24'(-1304);
			34491: out = 24'(1352);
			34492: out = 24'(1208);
			34493: out = 24'(-1604);
			34494: out = 24'(-2764);
			34495: out = 24'(1288);
			34496: out = 24'(-2048);
			34497: out = 24'(-2004);
			34498: out = 24'(-672);
			34499: out = 24'(1468);
			34500: out = 24'(-196);
			34501: out = 24'(820);
			34502: out = 24'(2696);
			34503: out = 24'(3704);
			34504: out = 24'(1028);
			34505: out = 24'(-1408);
			34506: out = 24'(-2276);
			34507: out = 24'(-2352);
			34508: out = 24'(-3616);
			34509: out = 24'(-4852);
			34510: out = 24'(-3144);
			34511: out = 24'(-2332);
			34512: out = 24'(-4668);
			34513: out = 24'(808);
			34514: out = 24'(5724);
			34515: out = 24'(9064);
			34516: out = 24'(6680);
			34517: out = 24'(1816);
			34518: out = 24'(664);
			34519: out = 24'(56);
			34520: out = 24'(-6860);
			34521: out = 24'(-15704);
			34522: out = 24'(-15368);
			34523: out = 24'(-2640);
			34524: out = 24'(7876);
			34525: out = 24'(8156);
			34526: out = 24'(5848);
			34527: out = 24'(7236);
			34528: out = 24'(6036);
			34529: out = 24'(-1668);
			34530: out = 24'(-13224);
			34531: out = 24'(-12784);
			34532: out = 24'(-6140);
			34533: out = 24'(-372);
			34534: out = 24'(3976);
			34535: out = 24'(10120);
			34536: out = 24'(9916);
			34537: out = 24'(3888);
			34538: out = 24'(1672);
			34539: out = 24'(-228);
			34540: out = 24'(-956);
			34541: out = 24'(-2896);
			34542: out = 24'(-5096);
			34543: out = 24'(-4948);
			34544: out = 24'(-2776);
			34545: out = 24'(3392);
			34546: out = 24'(9116);
			34547: out = 24'(10008);
			34548: out = 24'(844);
			34549: out = 24'(-3348);
			34550: out = 24'(1812);
			34551: out = 24'(-620);
			34552: out = 24'(-4368);
			34553: out = 24'(-6732);
			34554: out = 24'(-1452);
			34555: out = 24'(3348);
			34556: out = 24'(7584);
			34557: out = 24'(6152);
			34558: out = 24'(1568);
			34559: out = 24'(-7096);
			34560: out = 24'(-6812);
			34561: out = 24'(-4888);
			34562: out = 24'(1596);
			34563: out = 24'(9364);
			34564: out = 24'(9288);
			34565: out = 24'(5796);
			34566: out = 24'(2012);
			34567: out = 24'(-1448);
			34568: out = 24'(-6312);
			34569: out = 24'(-9756);
			34570: out = 24'(-7412);
			34571: out = 24'(-872);
			34572: out = 24'(-564);
			34573: out = 24'(3052);
			34574: out = 24'(4368);
			34575: out = 24'(2772);
			34576: out = 24'(-2164);
			34577: out = 24'(-680);
			34578: out = 24'(-212);
			34579: out = 24'(-528);
			34580: out = 24'(-132);
			34581: out = 24'(752);
			34582: out = 24'(576);
			34583: out = 24'(-1348);
			34584: out = 24'(-1784);
			34585: out = 24'(-820);
			34586: out = 24'(300);
			34587: out = 24'(-2916);
			34588: out = 24'(-7032);
			34589: out = 24'(-8416);
			34590: out = 24'(1788);
			34591: out = 24'(4788);
			34592: out = 24'(-3460);
			34593: out = 24'(-12056);
			34594: out = 24'(-7524);
			34595: out = 24'(-680);
			34596: out = 24'(-768);
			34597: out = 24'(-2168);
			34598: out = 24'(176);
			34599: out = 24'(9224);
			34600: out = 24'(11928);
			34601: out = 24'(4044);
			34602: out = 24'(-3332);
			34603: out = 24'(-9444);
			34604: out = 24'(-11720);
			34605: out = 24'(-9340);
			34606: out = 24'(-292);
			34607: out = 24'(7592);
			34608: out = 24'(9056);
			34609: out = 24'(4188);
			34610: out = 24'(400);
			34611: out = 24'(692);
			34612: out = 24'(3408);
			34613: out = 24'(3412);
			34614: out = 24'(-116);
			34615: out = 24'(1044);
			34616: out = 24'(-1904);
			34617: out = 24'(-5216);
			34618: out = 24'(-600);
			34619: out = 24'(-1136);
			34620: out = 24'(3832);
			34621: out = 24'(920);
			34622: out = 24'(-4256);
			34623: out = 24'(3264);
			34624: out = 24'(8000);
			34625: out = 24'(3340);
			34626: out = 24'(-3816);
			34627: out = 24'(972);
			34628: out = 24'(6552);
			34629: out = 24'(5376);
			34630: out = 24'(-120);
			34631: out = 24'(-172);
			34632: out = 24'(-380);
			34633: out = 24'(-2956);
			34634: out = 24'(-4584);
			34635: out = 24'(312);
			34636: out = 24'(-464);
			34637: out = 24'(-2084);
			34638: out = 24'(-3656);
			34639: out = 24'(-1432);
			34640: out = 24'(-856);
			34641: out = 24'(2612);
			34642: out = 24'(5952);
			34643: out = 24'(6968);
			34644: out = 24'(-172);
			34645: out = 24'(-1968);
			34646: out = 24'(-888);
			34647: out = 24'(1224);
			34648: out = 24'(-768);
			34649: out = 24'(-3992);
			34650: out = 24'(-4588);
			34651: out = 24'(608);
			34652: out = 24'(4776);
			34653: out = 24'(2340);
			34654: out = 24'(-3952);
			34655: out = 24'(-7620);
			34656: out = 24'(-8276);
			34657: out = 24'(-7892);
			34658: out = 24'(-5604);
			34659: out = 24'(1888);
			34660: out = 24'(9044);
			34661: out = 24'(9428);
			34662: out = 24'(2524);
			34663: out = 24'(-876);
			34664: out = 24'(-604);
			34665: out = 24'(-5320);
			34666: out = 24'(-9844);
			34667: out = 24'(-9092);
			34668: out = 24'(-1304);
			34669: out = 24'(4068);
			34670: out = 24'(5172);
			34671: out = 24'(1400);
			34672: out = 24'(1504);
			34673: out = 24'(5904);
			34674: out = 24'(4200);
			34675: out = 24'(-212);
			34676: out = 24'(-6988);
			34677: out = 24'(-11960);
			34678: out = 24'(-16248);
			34679: out = 24'(-7432);
			34680: out = 24'(2796);
			34681: out = 24'(8292);
			34682: out = 24'(9660);
			34683: out = 24'(9980);
			34684: out = 24'(5420);
			34685: out = 24'(-3848);
			34686: out = 24'(-12872);
			34687: out = 24'(-17784);
			34688: out = 24'(-12976);
			34689: out = 24'(-2716);
			34690: out = 24'(5560);
			34691: out = 24'(8548);
			34692: out = 24'(10976);
			34693: out = 24'(12120);
			34694: out = 24'(7392);
			34695: out = 24'(-3232);
			34696: out = 24'(-11392);
			34697: out = 24'(-10600);
			34698: out = 24'(-4380);
			34699: out = 24'(448);
			34700: out = 24'(3856);
			34701: out = 24'(4236);
			34702: out = 24'(-172);
			34703: out = 24'(-3420);
			34704: out = 24'(-1696);
			34705: out = 24'(8276);
			34706: out = 24'(9492);
			34707: out = 24'(-368);
			34708: out = 24'(-5880);
			34709: out = 24'(1000);
			34710: out = 24'(6676);
			34711: out = 24'(3592);
			34712: out = 24'(280);
			34713: out = 24'(6712);
			34714: out = 24'(5852);
			34715: out = 24'(-6256);
			34716: out = 24'(-9948);
			34717: out = 24'(-4076);
			34718: out = 24'(5684);
			34719: out = 24'(6884);
			34720: out = 24'(1232);
			34721: out = 24'(-1480);
			34722: out = 24'(-980);
			34723: out = 24'(656);
			34724: out = 24'(1304);
			34725: out = 24'(4168);
			34726: out = 24'(2120);
			34727: out = 24'(1752);
			34728: out = 24'(3828);
			34729: out = 24'(1464);
			34730: out = 24'(-4536);
			34731: out = 24'(-5008);
			34732: out = 24'(784);
			34733: out = 24'(-556);
			34734: out = 24'(-1100);
			34735: out = 24'(-1636);
			34736: out = 24'(1116);
			34737: out = 24'(3596);
			34738: out = 24'(-4728);
			34739: out = 24'(-11452);
			34740: out = 24'(-7196);
			34741: out = 24'(4804);
			34742: out = 24'(8108);
			34743: out = 24'(3956);
			34744: out = 24'(-2336);
			34745: out = 24'(-4744);
			34746: out = 24'(-8060);
			34747: out = 24'(-4008);
			34748: out = 24'(-152);
			34749: out = 24'(-104);
			34750: out = 24'(-2724);
			34751: out = 24'(-1140);
			34752: out = 24'(816);
			34753: out = 24'(-20);
			34754: out = 24'(728);
			34755: out = 24'(-188);
			34756: out = 24'(3240);
			34757: out = 24'(5924);
			34758: out = 24'(4072);
			34759: out = 24'(988);
			34760: out = 24'(-3168);
			34761: out = 24'(-9204);
			34762: out = 24'(-13972);
			34763: out = 24'(-7496);
			34764: out = 24'(3444);
			34765: out = 24'(11276);
			34766: out = 24'(10432);
			34767: out = 24'(-364);
			34768: out = 24'(-4316);
			34769: out = 24'(-3564);
			34770: out = 24'(-820);
			34771: out = 24'(92);
			34772: out = 24'(1868);
			34773: out = 24'(136);
			34774: out = 24'(-532);
			34775: out = 24'(4812);
			34776: out = 24'(8656);
			34777: out = 24'(7948);
			34778: out = 24'(3780);
			34779: out = 24'(1408);
			34780: out = 24'(876);
			34781: out = 24'(-3052);
			34782: out = 24'(-9580);
			34783: out = 24'(-12408);
			34784: out = 24'(-8736);
			34785: out = 24'(508);
			34786: out = 24'(7500);
			34787: out = 24'(9488);
			34788: out = 24'(8244);
			34789: out = 24'(3356);
			34790: out = 24'(-1856);
			34791: out = 24'(-5688);
			34792: out = 24'(-6228);
			34793: out = 24'(-1640);
			34794: out = 24'(2840);
			34795: out = 24'(3472);
			34796: out = 24'(-172);
			34797: out = 24'(948);
			34798: out = 24'(1008);
			34799: out = 24'(708);
			34800: out = 24'(-116);
			34801: out = 24'(-164);
			34802: out = 24'(736);
			34803: out = 24'(1064);
			34804: out = 24'(-436);
			34805: out = 24'(1312);
			34806: out = 24'(-5740);
			34807: out = 24'(-7284);
			34808: out = 24'(-1672);
			34809: out = 24'(-644);
			34810: out = 24'(4024);
			34811: out = 24'(2180);
			34812: out = 24'(-592);
			34813: out = 24'(-1908);
			34814: out = 24'(-412);
			34815: out = 24'(-2128);
			34816: out = 24'(-2668);
			34817: out = 24'(664);
			34818: out = 24'(3760);
			34819: out = 24'(4436);
			34820: out = 24'(4448);
			34821: out = 24'(5108);
			34822: out = 24'(1284);
			34823: out = 24'(-980);
			34824: out = 24'(-3636);
			34825: out = 24'(-5140);
			34826: out = 24'(-3432);
			34827: out = 24'(-3572);
			34828: out = 24'(-1652);
			34829: out = 24'(300);
			34830: out = 24'(-4);
			34831: out = 24'(968);
			34832: out = 24'(812);
			34833: out = 24'(-1152);
			34834: out = 24'(-2880);
			34835: out = 24'(3160);
			34836: out = 24'(7276);
			34837: out = 24'(6068);
			34838: out = 24'(8);
			34839: out = 24'(-5952);
			34840: out = 24'(-2244);
			34841: out = 24'(3516);
			34842: out = 24'(2820);
			34843: out = 24'(-1340);
			34844: out = 24'(-5012);
			34845: out = 24'(-3856);
			34846: out = 24'(-4984);
			34847: out = 24'(-10868);
			34848: out = 24'(-9280);
			34849: out = 24'(1120);
			34850: out = 24'(11176);
			34851: out = 24'(10600);
			34852: out = 24'(756);
			34853: out = 24'(-5004);
			34854: out = 24'(-2752);
			34855: out = 24'(-376);
			34856: out = 24'(-3792);
			34857: out = 24'(-8692);
			34858: out = 24'(-6052);
			34859: out = 24'(2552);
			34860: out = 24'(7896);
			34861: out = 24'(7160);
			34862: out = 24'(2988);
			34863: out = 24'(-1484);
			34864: out = 24'(-7960);
			34865: out = 24'(-7900);
			34866: out = 24'(-5632);
			34867: out = 24'(-948);
			34868: out = 24'(2168);
			34869: out = 24'(11148);
			34870: out = 24'(8312);
			34871: out = 24'(844);
			34872: out = 24'(-5256);
			34873: out = 24'(-7576);
			34874: out = 24'(-7144);
			34875: out = 24'(-3408);
			34876: out = 24'(1140);
			34877: out = 24'(1804);
			34878: out = 24'(956);
			34879: out = 24'(804);
			34880: out = 24'(2320);
			34881: out = 24'(4204);
			34882: out = 24'(4192);
			34883: out = 24'(4120);
			34884: out = 24'(3320);
			34885: out = 24'(1108);
			34886: out = 24'(-3572);
			34887: out = 24'(-3304);
			34888: out = 24'(-244);
			34889: out = 24'(1864);
			34890: out = 24'(7012);
			34891: out = 24'(7792);
			34892: out = 24'(4856);
			34893: out = 24'(-1780);
			34894: out = 24'(-5316);
			34895: out = 24'(-7012);
			34896: out = 24'(-2076);
			34897: out = 24'(3552);
			34898: out = 24'(4976);
			34899: out = 24'(4008);
			34900: out = 24'(3808);
			34901: out = 24'(2212);
			34902: out = 24'(-3428);
			34903: out = 24'(-5748);
			34904: out = 24'(-3940);
			34905: out = 24'(-1020);
			34906: out = 24'(-1868);
			34907: out = 24'(212);
			34908: out = 24'(-160);
			34909: out = 24'(-1364);
			34910: out = 24'(-4868);
			34911: out = 24'(-2332);
			34912: out = 24'(-1508);
			34913: out = 24'(4056);
			34914: out = 24'(6980);
			34915: out = 24'(4172);
			34916: out = 24'(-8292);
			34917: out = 24'(-11904);
			34918: out = 24'(-5868);
			34919: out = 24'(1600);
			34920: out = 24'(1536);
			34921: out = 24'(3768);
			34922: out = 24'(4484);
			34923: out = 24'(-772);
			34924: out = 24'(-7364);
			34925: out = 24'(-7020);
			34926: out = 24'(-528);
			34927: out = 24'(4104);
			34928: out = 24'(624);
			34929: out = 24'(-792);
			34930: out = 24'(-2108);
			34931: out = 24'(-1868);
			34932: out = 24'(4024);
			34933: out = 24'(4500);
			34934: out = 24'(2144);
			34935: out = 24'(752);
			34936: out = 24'(5272);
			34937: out = 24'(2144);
			34938: out = 24'(-3300);
			34939: out = 24'(-8616);
			34940: out = 24'(-8196);
			34941: out = 24'(-10212);
			34942: out = 24'(-4112);
			34943: out = 24'(5204);
			34944: out = 24'(12412);
			34945: out = 24'(8028);
			34946: out = 24'(5372);
			34947: out = 24'(2576);
			34948: out = 24'(916);
			34949: out = 24'(-332);
			34950: out = 24'(916);
			34951: out = 24'(1300);
			34952: out = 24'(576);
			34953: out = 24'(-1776);
			34954: out = 24'(3608);
			34955: out = 24'(5416);
			34956: out = 24'(3892);
			34957: out = 24'(748);
			34958: out = 24'(36);
			34959: out = 24'(-1520);
			34960: out = 24'(-1540);
			34961: out = 24'(-16);
			34962: out = 24'(4532);
			34963: out = 24'(1580);
			34964: out = 24'(-648);
			34965: out = 24'(848);
			34966: out = 24'(-464);
			34967: out = 24'(444);
			34968: out = 24'(756);
			34969: out = 24'(-1824);
			34970: out = 24'(-5604);
			34971: out = 24'(-6172);
			34972: out = 24'(1688);
			34973: out = 24'(6552);
			34974: out = 24'(-896);
			34975: out = 24'(-8924);
			34976: out = 24'(-4792);
			34977: out = 24'(6208);
			34978: out = 24'(7252);
			34979: out = 24'(8304);
			34980: out = 24'(1680);
			34981: out = 24'(-1128);
			34982: out = 24'(-2940);
			34983: out = 24'(-5624);
			34984: out = 24'(-7312);
			34985: out = 24'(-1912);
			34986: out = 24'(4212);
			34987: out = 24'(3532);
			34988: out = 24'(-1760);
			34989: out = 24'(-2500);
			34990: out = 24'(-136);
			34991: out = 24'(-3872);
			34992: out = 24'(-8708);
			34993: out = 24'(-8836);
			34994: out = 24'(268);
			34995: out = 24'(8528);
			34996: out = 24'(12104);
			34997: out = 24'(4644);
			34998: out = 24'(-3580);
			34999: out = 24'(-8216);
			35000: out = 24'(-10008);
			35001: out = 24'(-8264);
			35002: out = 24'(-972);
			35003: out = 24'(5620);
			35004: out = 24'(4052);
			35005: out = 24'(788);
			35006: out = 24'(1456);
			35007: out = 24'(3572);
			35008: out = 24'(-304);
			35009: out = 24'(-152);
			35010: out = 24'(-12);
			35011: out = 24'(-956);
			35012: out = 24'(-3028);
			35013: out = 24'(-2380);
			35014: out = 24'(1932);
			35015: out = 24'(2964);
			35016: out = 24'(-64);
			35017: out = 24'(3104);
			35018: out = 24'(6656);
			35019: out = 24'(3668);
			35020: out = 24'(-4096);
			35021: out = 24'(-132);
			35022: out = 24'(-236);
			35023: out = 24'(-2096);
			35024: out = 24'(-4568);
			35025: out = 24'(204);
			35026: out = 24'(5312);
			35027: out = 24'(6484);
			35028: out = 24'(1488);
			35029: out = 24'(236);
			35030: out = 24'(-2716);
			35031: out = 24'(1576);
			35032: out = 24'(2236);
			35033: out = 24'(-2520);
			35034: out = 24'(-3484);
			35035: out = 24'(-1332);
			35036: out = 24'(-1116);
			35037: out = 24'(-3328);
			35038: out = 24'(612);
			35039: out = 24'(196);
			35040: out = 24'(-624);
			35041: out = 24'(720);
			35042: out = 24'(4268);
			35043: out = 24'(5336);
			35044: out = 24'(-20);
			35045: out = 24'(-5672);
			35046: out = 24'(-2988);
			35047: out = 24'(-2580);
			35048: out = 24'(-232);
			35049: out = 24'(1976);
			35050: out = 24'(3156);
			35051: out = 24'(-940);
			35052: out = 24'(-6176);
			35053: out = 24'(-5696);
			35054: out = 24'(740);
			35055: out = 24'(-548);
			35056: out = 24'(104);
			35057: out = 24'(-348);
			35058: out = 24'(-276);
			35059: out = 24'(-3316);
			35060: out = 24'(-996);
			35061: out = 24'(-104);
			35062: out = 24'(152);
			35063: out = 24'(1172);
			35064: out = 24'(-1132);
			35065: out = 24'(-780);
			35066: out = 24'(1432);
			35067: out = 24'(-640);
			35068: out = 24'(3904);
			35069: out = 24'(916);
			35070: out = 24'(832);
			35071: out = 24'(4016);
			35072: out = 24'(8240);
			35073: out = 24'(-300);
			35074: out = 24'(-7476);
			35075: out = 24'(-6500);
			35076: out = 24'(768);
			35077: out = 24'(1052);
			35078: out = 24'(2660);
			35079: out = 24'(4888);
			35080: out = 24'(3380);
			35081: out = 24'(-992);
			35082: out = 24'(-2352);
			35083: out = 24'(-2948);
			35084: out = 24'(-6300);
			35085: out = 24'(-6352);
			35086: out = 24'(-2352);
			35087: out = 24'(396);
			35088: out = 24'(516);
			35089: out = 24'(6524);
			35090: out = 24'(10840);
			35091: out = 24'(8036);
			35092: out = 24'(-1076);
			35093: out = 24'(-5764);
			35094: out = 24'(-7644);
			35095: out = 24'(-8500);
			35096: out = 24'(-7664);
			35097: out = 24'(1152);
			35098: out = 24'(6124);
			35099: out = 24'(6296);
			35100: out = 24'(2028);
			35101: out = 24'(-216);
			35102: out = 24'(-4304);
			35103: out = 24'(-3492);
			35104: out = 24'(-552);
			35105: out = 24'(1168);
			35106: out = 24'(3564);
			35107: out = 24'(3448);
			35108: out = 24'(3892);
			35109: out = 24'(2164);
			35110: out = 24'(-3928);
			35111: out = 24'(-9972);
			35112: out = 24'(-6628);
			35113: out = 24'(1180);
			35114: out = 24'(744);
			35115: out = 24'(1380);
			35116: out = 24'(2252);
			35117: out = 24'(3528);
			35118: out = 24'(728);
			35119: out = 24'(112);
			35120: out = 24'(44);
			35121: out = 24'(876);
			35122: out = 24'(-712);
			35123: out = 24'(-2696);
			35124: out = 24'(-3744);
			35125: out = 24'(-1916);
			35126: out = 24'(0);
			35127: out = 24'(-68);
			35128: out = 24'(2356);
			35129: out = 24'(4380);
			35130: out = 24'(2640);
			35131: out = 24'(240);
			35132: out = 24'(-5184);
			35133: out = 24'(-3212);
			35134: out = 24'(2692);
			35135: out = 24'(3104);
			35136: out = 24'(780);
			35137: out = 24'(-2788);
			35138: out = 24'(-2368);
			35139: out = 24'(-172);
			35140: out = 24'(1132);
			35141: out = 24'(204);
			35142: out = 24'(-252);
			35143: out = 24'(-356);
			35144: out = 24'(4);
			35145: out = 24'(-504);
			35146: out = 24'(548);
			35147: out = 24'(-368);
			35148: out = 24'(-5556);
			35149: out = 24'(-9996);
			35150: out = 24'(-5584);
			35151: out = 24'(4516);
			35152: out = 24'(10228);
			35153: out = 24'(9444);
			35154: out = 24'(4428);
			35155: out = 24'(-1064);
			35156: out = 24'(-4924);
			35157: out = 24'(-10128);
			35158: out = 24'(-8252);
			35159: out = 24'(-4164);
			35160: out = 24'(-1088);
			35161: out = 24'(-328);
			35162: out = 24'(9988);
			35163: out = 24'(15484);
			35164: out = 24'(8212);
			35165: out = 24'(-3308);
			35166: out = 24'(-8280);
			35167: out = 24'(-4732);
			35168: out = 24'(-2044);
			35169: out = 24'(-2860);
			35170: out = 24'(-3648);
			35171: out = 24'(1304);
			35172: out = 24'(5536);
			35173: out = 24'(3316);
			35174: out = 24'(484);
			35175: out = 24'(1664);
			35176: out = 24'(3728);
			35177: out = 24'(-196);
			35178: out = 24'(-4780);
			35179: out = 24'(-8088);
			35180: out = 24'(-5036);
			35181: out = 24'(-1200);
			35182: out = 24'(1608);
			35183: out = 24'(-104);
			35184: out = 24'(3348);
			35185: out = 24'(7100);
			35186: out = 24'(1004);
			35187: out = 24'(-1160);
			35188: out = 24'(-1256);
			35189: out = 24'(152);
			35190: out = 24'(-320);
			35191: out = 24'(-2636);
			35192: out = 24'(-1780);
			35193: out = 24'(532);
			35194: out = 24'(-504);
			35195: out = 24'(152);
			35196: out = 24'(-740);
			35197: out = 24'(2668);
			35198: out = 24'(7408);
			35199: out = 24'(3660);
			35200: out = 24'(1868);
			35201: out = 24'(-404);
			35202: out = 24'(-1956);
			35203: out = 24'(-220);
			35204: out = 24'(-444);
			35205: out = 24'(304);
			35206: out = 24'(1088);
			35207: out = 24'(868);
			35208: out = 24'(-1320);
			35209: out = 24'(-2400);
			35210: out = 24'(-1128);
			35211: out = 24'(616);
			35212: out = 24'(84);
			35213: out = 24'(-568);
			35214: out = 24'(1036);
			35215: out = 24'(3444);
			35216: out = 24'(1232);
			35217: out = 24'(-1168);
			35218: out = 24'(-1844);
			35219: out = 24'(-560);
			35220: out = 24'(-2200);
			35221: out = 24'(-572);
			35222: out = 24'(-228);
			35223: out = 24'(-336);
			35224: out = 24'(-348);
			35225: out = 24'(-212);
			35226: out = 24'(-388);
			35227: out = 24'(648);
			35228: out = 24'(3300);
			35229: out = 24'(-3352);
			35230: out = 24'(-6304);
			35231: out = 24'(-4064);
			35232: out = 24'(1560);
			35233: out = 24'(4372);
			35234: out = 24'(5120);
			35235: out = 24'(3344);
			35236: out = 24'(-720);
			35237: out = 24'(-7260);
			35238: out = 24'(-8120);
			35239: out = 24'(-5684);
			35240: out = 24'(-2048);
			35241: out = 24'(1168);
			35242: out = 24'(1260);
			35243: out = 24'(-364);
			35244: out = 24'(-1724);
			35245: out = 24'(592);
			35246: out = 24'(3508);
			35247: out = 24'(7808);
			35248: out = 24'(6260);
			35249: out = 24'(-264);
			35250: out = 24'(-11108);
			35251: out = 24'(-7524);
			35252: out = 24'(-328);
			35253: out = 24'(444);
			35254: out = 24'(-3816);
			35255: out = 24'(-2172);
			35256: out = 24'(3604);
			35257: out = 24'(7824);
			35258: out = 24'(6896);
			35259: out = 24'(-1048);
			35260: out = 24'(-10580);
			35261: out = 24'(-10704);
			35262: out = 24'(4412);
			35263: out = 24'(4920);
			35264: out = 24'(3016);
			35265: out = 24'(312);
			35266: out = 24'(1508);
			35267: out = 24'(552);
			35268: out = 24'(404);
			35269: out = 24'(-268);
			35270: out = 24'(1520);
			35271: out = 24'(616);
			35272: out = 24'(768);
			35273: out = 24'(-2612);
			35274: out = 24'(-4352);
			35275: out = 24'(-3772);
			35276: out = 24'(-60);
			35277: out = 24'(-2952);
			35278: out = 24'(-5476);
			35279: out = 24'(-1492);
			35280: out = 24'(6272);
			35281: out = 24'(3444);
			35282: out = 24'(-4088);
			35283: out = 24'(-5008);
			35284: out = 24'(3336);
			35285: out = 24'(5996);
			35286: out = 24'(3008);
			35287: out = 24'(-460);
			35288: out = 24'(16);
			35289: out = 24'(-676);
			35290: out = 24'(2688);
			35291: out = 24'(7284);
			35292: out = 24'(3456);
			35293: out = 24'(468);
			35294: out = 24'(-564);
			35295: out = 24'(-1736);
			35296: out = 24'(-7648);
			35297: out = 24'(-3880);
			35298: out = 24'(5088);
			35299: out = 24'(9988);
			35300: out = 24'(1864);
			35301: out = 24'(-8028);
			35302: out = 24'(-12516);
			35303: out = 24'(-6352);
			35304: out = 24'(1524);
			35305: out = 24'(1472);
			35306: out = 24'(848);
			35307: out = 24'(2044);
			35308: out = 24'(4392);
			35309: out = 24'(8156);
			35310: out = 24'(3280);
			35311: out = 24'(-3220);
			35312: out = 24'(-6020);
			35313: out = 24'(-1812);
			35314: out = 24'(-3108);
			35315: out = 24'(-3384);
			35316: out = 24'(-2656);
			35317: out = 24'(300);
			35318: out = 24'(-620);
			35319: out = 24'(4452);
			35320: out = 24'(6108);
			35321: out = 24'(-1784);
			35322: out = 24'(-4716);
			35323: out = 24'(-10676);
			35324: out = 24'(-10768);
			35325: out = 24'(-5552);
			35326: out = 24'(3700);
			35327: out = 24'(6792);
			35328: out = 24'(8040);
			35329: out = 24'(6188);
			35330: out = 24'(1100);
			35331: out = 24'(-5856);
			35332: out = 24'(-7556);
			35333: out = 24'(-4628);
			35334: out = 24'(-1588);
			35335: out = 24'(-2624);
			35336: out = 24'(-1320);
			35337: out = 24'(1668);
			35338: out = 24'(3680);
			35339: out = 24'(-3332);
			35340: out = 24'(-3952);
			35341: out = 24'(-1336);
			35342: out = 24'(364);
			35343: out = 24'(276);
			35344: out = 24'(112);
			35345: out = 24'(-632);
			35346: out = 24'(-1240);
			35347: out = 24'(332);
			35348: out = 24'(1132);
			35349: out = 24'(940);
			35350: out = 24'(264);
			35351: out = 24'(1724);
			35352: out = 24'(376);
			35353: out = 24'(848);
			35354: out = 24'(1460);
			35355: out = 24'(-32);
			35356: out = 24'(236);
			35357: out = 24'(-1316);
			35358: out = 24'(360);
			35359: out = 24'(4328);
			35360: out = 24'(1448);
			35361: out = 24'(1312);
			35362: out = 24'(956);
			35363: out = 24'(1044);
			35364: out = 24'(92);
			35365: out = 24'(860);
			35366: out = 24'(56);
			35367: out = 24'(-2872);
			35368: out = 24'(-5492);
			35369: out = 24'(-3892);
			35370: out = 24'(-100);
			35371: out = 24'(1764);
			35372: out = 24'(1488);
			35373: out = 24'(-1340);
			35374: out = 24'(1724);
			35375: out = 24'(4684);
			35376: out = 24'(3096);
			35377: out = 24'(-2272);
			35378: out = 24'(-1652);
			35379: out = 24'(2516);
			35380: out = 24'(4568);
			35381: out = 24'(208);
			35382: out = 24'(2304);
			35383: out = 24'(5888);
			35384: out = 24'(6248);
			35385: out = 24'(760);
			35386: out = 24'(-4468);
			35387: out = 24'(-7200);
			35388: out = 24'(-3080);
			35389: out = 24'(4980);
			35390: out = 24'(4132);
			35391: out = 24'(1728);
			35392: out = 24'(1448);
			35393: out = 24'(3712);
			35394: out = 24'(4660);
			35395: out = 24'(-1892);
			35396: out = 24'(-9316);
			35397: out = 24'(-9132);
			35398: out = 24'(-1168);
			35399: out = 24'(4188);
			35400: out = 24'(2920);
			35401: out = 24'(-300);
			35402: out = 24'(3932);
			35403: out = 24'(3068);
			35404: out = 24'(4544);
			35405: out = 24'(2832);
			35406: out = 24'(-3768);
			35407: out = 24'(-7452);
			35408: out = 24'(-4864);
			35409: out = 24'(-1456);
			35410: out = 24'(-3548);
			35411: out = 24'(1164);
			35412: out = 24'(244);
			35413: out = 24'(212);
			35414: out = 24'(1544);
			35415: out = 24'(4640);
			35416: out = 24'(1604);
			35417: out = 24'(-4416);
			35418: out = 24'(-9688);
			35419: out = 24'(-6948);
			35420: out = 24'(-2516);
			35421: out = 24'(5140);
			35422: out = 24'(7912);
			35423: out = 24'(3600);
			35424: out = 24'(-2092);
			35425: out = 24'(-1988);
			35426: out = 24'(396);
			35427: out = 24'(-740);
			35428: out = 24'(-7656);
			35429: out = 24'(-7952);
			35430: out = 24'(-3220);
			35431: out = 24'(400);
			35432: out = 24'(1288);
			35433: out = 24'(356);
			35434: out = 24'(-756);
			35435: out = 24'(-1316);
			35436: out = 24'(152);
			35437: out = 24'(2972);
			35438: out = 24'(4444);
			35439: out = 24'(3012);
			35440: out = 24'(-32);
			35441: out = 24'(704);
			35442: out = 24'(1208);
			35443: out = 24'(896);
			35444: out = 24'(-572);
			35445: out = 24'(-4796);
			35446: out = 24'(-7804);
			35447: out = 24'(-3840);
			35448: out = 24'(4708);
			35449: out = 24'(3824);
			35450: out = 24'(1644);
			35451: out = 24'(-568);
			35452: out = 24'(736);
			35453: out = 24'(3404);
			35454: out = 24'(464);
			35455: out = 24'(-3348);
			35456: out = 24'(-1444);
			35457: out = 24'(3412);
			35458: out = 24'(5384);
			35459: out = 24'(2680);
			35460: out = 24'(1628);
			35461: out = 24'(3244);
			35462: out = 24'(840);
			35463: out = 24'(-4244);
			35464: out = 24'(-4964);
			35465: out = 24'(-288);
			35466: out = 24'(72);
			35467: out = 24'(-3256);
			35468: out = 24'(-3028);
			35469: out = 24'(2376);
			35470: out = 24'(6872);
			35471: out = 24'(2304);
			35472: out = 24'(-1264);
			35473: out = 24'(228);
			35474: out = 24'(-616);
			35475: out = 24'(-116);
			35476: out = 24'(-376);
			35477: out = 24'(-200);
			35478: out = 24'(-232);
			35479: out = 24'(-432);
			35480: out = 24'(560);
			35481: out = 24'(-8);
			35482: out = 24'(-1932);
			35483: out = 24'(-3580);
			35484: out = 24'(3304);
			35485: out = 24'(7576);
			35486: out = 24'(3388);
			35487: out = 24'(68);
			35488: out = 24'(-2180);
			35489: out = 24'(-1784);
			35490: out = 24'(-2744);
			35491: out = 24'(-4568);
			35492: out = 24'(-6076);
			35493: out = 24'(-4424);
			35494: out = 24'(-16);
			35495: out = 24'(3548);
			35496: out = 24'(4132);
			35497: out = 24'(1292);
			35498: out = 24'(452);
			35499: out = 24'(3548);
			35500: out = 24'(420);
			35501: out = 24'(-4888);
			35502: out = 24'(-8044);
			35503: out = 24'(-5428);
			35504: out = 24'(-6336);
			35505: out = 24'(600);
			35506: out = 24'(6684);
			35507: out = 24'(7944);
			35508: out = 24'(3960);
			35509: out = 24'(-488);
			35510: out = 24'(-3088);
			35511: out = 24'(-2752);
			35512: out = 24'(-100);
			35513: out = 24'(-1472);
			35514: out = 24'(-1976);
			35515: out = 24'(-1296);
			35516: out = 24'(1752);
			35517: out = 24'(2856);
			35518: out = 24'(6436);
			35519: out = 24'(4960);
			35520: out = 24'(-940);
			35521: out = 24'(-2016);
			35522: out = 24'(84);
			35523: out = 24'(-1196);
			35524: out = 24'(-7328);
			35525: out = 24'(-7164);
			35526: out = 24'(-2976);
			35527: out = 24'(4196);
			35528: out = 24'(6540);
			35529: out = 24'(956);
			35530: out = 24'(-1136);
			35531: out = 24'(-3060);
			35532: out = 24'(-2208);
			35533: out = 24'(1420);
			35534: out = 24'(4324);
			35535: out = 24'(4392);
			35536: out = 24'(3008);
			35537: out = 24'(1916);
			35538: out = 24'(-1568);
			35539: out = 24'(-1588);
			35540: out = 24'(1916);
			35541: out = 24'(3988);
			35542: out = 24'(-1492);
			35543: out = 24'(-6760);
			35544: out = 24'(-4600);
			35545: out = 24'(2560);
			35546: out = 24'(2984);
			35547: out = 24'(900);
			35548: out = 24'(-1608);
			35549: out = 24'(1028);
			35550: out = 24'(3632);
			35551: out = 24'(1068);
			35552: out = 24'(-4956);
			35553: out = 24'(-5632);
			35554: out = 24'(384);
			35555: out = 24'(3672);
			35556: out = 24'(1760);
			35557: out = 24'(-1984);
			35558: out = 24'(-3044);
			35559: out = 24'(-3276);
			35560: out = 24'(-2184);
			35561: out = 24'(-1132);
			35562: out = 24'(12);
			35563: out = 24'(-400);
			35564: out = 24'(8);
			35565: out = 24'(-1476);
			35566: out = 24'(-4180);
			35567: out = 24'(-8028);
			35568: out = 24'(-1860);
			35569: out = 24'(2328);
			35570: out = 24'(3668);
			35571: out = 24'(3332);
			35572: out = 24'(1392);
			35573: out = 24'(812);
			35574: out = 24'(128);
			35575: out = 24'(-2256);
			35576: out = 24'(-4976);
			35577: out = 24'(-4208);
			35578: out = 24'(232);
			35579: out = 24'(4224);
			35580: out = 24'(6704);
			35581: out = 24'(2512);
			35582: out = 24'(1584);
			35583: out = 24'(3276);
			35584: out = 24'(-740);
			35585: out = 24'(8);
			35586: out = 24'(-2188);
			35587: out = 24'(-2368);
			35588: out = 24'(-52);
			35589: out = 24'(-100);
			35590: out = 24'(224);
			35591: out = 24'(2232);
			35592: out = 24'(4016);
			35593: out = 24'(-60);
			35594: out = 24'(-3412);
			35595: out = 24'(-3312);
			35596: out = 24'(24);
			35597: out = 24'(-516);
			35598: out = 24'(-864);
			35599: out = 24'(-2796);
			35600: out = 24'(-1536);
			35601: out = 24'(4392);
			35602: out = 24'(7112);
			35603: out = 24'(5600);
			35604: out = 24'(1608);
			35605: out = 24'(-388);
			35606: out = 24'(-1952);
			35607: out = 24'(-1268);
			35608: out = 24'(-660);
			35609: out = 24'(-116);
			35610: out = 24'(2576);
			35611: out = 24'(3416);
			35612: out = 24'(660);
			35613: out = 24'(-3956);
			35614: out = 24'(-4288);
			35615: out = 24'(-3884);
			35616: out = 24'(-1808);
			35617: out = 24'(816);
			35618: out = 24'(6420);
			35619: out = 24'(2124);
			35620: out = 24'(-208);
			35621: out = 24'(-1024);
			35622: out = 24'(-1876);
			35623: out = 24'(380);
			35624: out = 24'(1068);
			35625: out = 24'(-24);
			35626: out = 24'(-2012);
			35627: out = 24'(-3192);
			35628: out = 24'(-760);
			35629: out = 24'(728);
			35630: out = 24'(-472);
			35631: out = 24'(756);
			35632: out = 24'(1988);
			35633: out = 24'(4912);
			35634: out = 24'(5300);
			35635: out = 24'(-500);
			35636: out = 24'(-3708);
			35637: out = 24'(-3988);
			35638: out = 24'(-200);
			35639: out = 24'(3800);
			35640: out = 24'(1480);
			35641: out = 24'(-2300);
			35642: out = 24'(-1772);
			35643: out = 24'(3100);
			35644: out = 24'(-108);
			35645: out = 24'(-1792);
			35646: out = 24'(-520);
			35647: out = 24'(2848);
			35648: out = 24'(-3052);
			35649: out = 24'(-4320);
			35650: out = 24'(-3216);
			35651: out = 24'(628);
			35652: out = 24'(2536);
			35653: out = 24'(1088);
			35654: out = 24'(-2980);
			35655: out = 24'(-3444);
			35656: out = 24'(156);
			35657: out = 24'(564);
			35658: out = 24'(-4308);
			35659: out = 24'(-5800);
			35660: out = 24'(0);
			35661: out = 24'(100);
			35662: out = 24'(-4892);
			35663: out = 24'(-7432);
			35664: out = 24'(56);
			35665: out = 24'(3352);
			35666: out = 24'(4880);
			35667: out = 24'(784);
			35668: out = 24'(-1204);
			35669: out = 24'(-620);
			35670: out = 24'(3652);
			35671: out = 24'(2612);
			35672: out = 24'(-1964);
			35673: out = 24'(-9404);
			35674: out = 24'(488);
			35675: out = 24'(4940);
			35676: out = 24'(3172);
			35677: out = 24'(-464);
			35678: out = 24'(84);
			35679: out = 24'(-4112);
			35680: out = 24'(-6232);
			35681: out = 24'(-584);
			35682: out = 24'(2548);
			35683: out = 24'(2472);
			35684: out = 24'(16);
			35685: out = 24'(256);
			35686: out = 24'(328);
			35687: out = 24'(1108);
			35688: out = 24'(-584);
			35689: out = 24'(-1728);
			35690: out = 24'(-1744);
			35691: out = 24'(2164);
			35692: out = 24'(3780);
			35693: out = 24'(1616);
			35694: out = 24'(-4288);
			35695: out = 24'(-3440);
			35696: out = 24'(760);
			35697: out = 24'(6260);
			35698: out = 24'(6424);
			35699: out = 24'(1332);
			35700: out = 24'(-5500);
			35701: out = 24'(-5096);
			35702: out = 24'(392);
			35703: out = 24'(4196);
			35704: out = 24'(832);
			35705: out = 24'(1712);
			35706: out = 24'(6628);
			35707: out = 24'(2576);
			35708: out = 24'(-1364);
			35709: out = 24'(-5336);
			35710: out = 24'(-5628);
			35711: out = 24'(-4392);
			35712: out = 24'(-1400);
			35713: out = 24'(3936);
			35714: out = 24'(7964);
			35715: out = 24'(5412);
			35716: out = 24'(3736);
			35717: out = 24'(-1152);
			35718: out = 24'(-4848);
			35719: out = 24'(-5608);
			35720: out = 24'(-1032);
			35721: out = 24'(-272);
			35722: out = 24'(-1196);
			35723: out = 24'(-1808);
			35724: out = 24'(-596);
			35725: out = 24'(508);
			35726: out = 24'(240);
			35727: out = 24'(-368);
			35728: out = 24'(740);
			35729: out = 24'(2532);
			35730: out = 24'(1488);
			35731: out = 24'(-1984);
			35732: out = 24'(-4516);
			35733: out = 24'(-5932);
			35734: out = 24'(-3048);
			35735: out = 24'(3096);
			35736: out = 24'(9036);
			35737: out = 24'(268);
			35738: out = 24'(-2592);
			35739: out = 24'(-3496);
			35740: out = 24'(-3844);
			35741: out = 24'(-9564);
			35742: out = 24'(-6116);
			35743: out = 24'(-1440);
			35744: out = 24'(1856);
			35745: out = 24'(3200);
			35746: out = 24'(3692);
			35747: out = 24'(1480);
			35748: out = 24'(-300);
			35749: out = 24'(512);
			35750: out = 24'(-4456);
			35751: out = 24'(-7024);
			35752: out = 24'(-4464);
			35753: out = 24'(1740);
			35754: out = 24'(3308);
			35755: out = 24'(-872);
			35756: out = 24'(-5660);
			35757: out = 24'(-4164);
			35758: out = 24'(-664);
			35759: out = 24'(3208);
			35760: out = 24'(2136);
			35761: out = 24'(-160);
			35762: out = 24'(-84);
			35763: out = 24'(208);
			35764: out = 24'(-788);
			35765: out = 24'(-1448);
			35766: out = 24'(-1524);
			35767: out = 24'(3984);
			35768: out = 24'(3012);
			35769: out = 24'(416);
			35770: out = 24'(-124);
			35771: out = 24'(32);
			35772: out = 24'(-2636);
			35773: out = 24'(-3792);
			35774: out = 24'(-856);
			35775: out = 24'(-300);
			35776: out = 24'(2492);
			35777: out = 24'(3932);
			35778: out = 24'(2432);
			35779: out = 24'(-1220);
			35780: out = 24'(-4164);
			35781: out = 24'(-480);
			35782: out = 24'(3612);
			35783: out = 24'(-684);
			35784: out = 24'(-1944);
			35785: out = 24'(-3376);
			35786: out = 24'(-1752);
			35787: out = 24'(308);
			35788: out = 24'(4068);
			35789: out = 24'(4296);
			35790: out = 24'(2068);
			35791: out = 24'(-308);
			35792: out = 24'(-156);
			35793: out = 24'(-1812);
			35794: out = 24'(-4392);
			35795: out = 24'(-4272);
			35796: out = 24'(3244);
			35797: out = 24'(4616);
			35798: out = 24'(2420);
			35799: out = 24'(-704);
			35800: out = 24'(112);
			35801: out = 24'(-360);
			35802: out = 24'(-60);
			35803: out = 24'(-40);
			35804: out = 24'(1232);
			35805: out = 24'(2764);
			35806: out = 24'(3880);
			35807: out = 24'(1128);
			35808: out = 24'(-2924);
			35809: out = 24'(660);
			35810: out = 24'(4664);
			35811: out = 24'(6448);
			35812: out = 24'(2288);
			35813: out = 24'(-5012);
			35814: out = 24'(-8360);
			35815: out = 24'(-6020);
			35816: out = 24'(-1968);
			35817: out = 24'(-72);
			35818: out = 24'(2560);
			35819: out = 24'(3912);
			35820: out = 24'(1100);
			35821: out = 24'(-5668);
			35822: out = 24'(-3476);
			35823: out = 24'(-1060);
			35824: out = 24'(404);
			35825: out = 24'(1404);
			35826: out = 24'(2972);
			35827: out = 24'(3784);
			35828: out = 24'(1028);
			35829: out = 24'(-3984);
			35830: out = 24'(-7840);
			35831: out = 24'(-6548);
			35832: out = 24'(-2588);
			35833: out = 24'(2244);
			35834: out = 24'(3012);
			35835: out = 24'(1712);
			35836: out = 24'(-4696);
			35837: out = 24'(-7140);
			35838: out = 24'(-2320);
			35839: out = 24'(4116);
			35840: out = 24'(2240);
			35841: out = 24'(928);
			35842: out = 24'(5004);
			35843: out = 24'(4824);
			35844: out = 24'(-3172);
			35845: out = 24'(-8832);
			35846: out = 24'(-3252);
			35847: out = 24'(2500);
			35848: out = 24'(3012);
			35849: out = 24'(-664);
			35850: out = 24'(-656);
			35851: out = 24'(-420);
			35852: out = 24'(720);
			35853: out = 24'(-1620);
			35854: out = 24'(-1444);
			35855: out = 24'(2360);
			35856: out = 24'(4788);
			35857: out = 24'(2056);
			35858: out = 24'(-80);
			35859: out = 24'(1136);
			35860: out = 24'(3380);
			35861: out = 24'(560);
			35862: out = 24'(-2580);
			35863: out = 24'(-2420);
			35864: out = 24'(1044);
			35865: out = 24'(-2132);
			35866: out = 24'(-4280);
			35867: out = 24'(-1836);
			35868: out = 24'(-108);
			35869: out = 24'(1028);
			35870: out = 24'(2716);
			35871: out = 24'(4908);
			35872: out = 24'(2968);
			35873: out = 24'(932);
			35874: out = 24'(-2572);
			35875: out = 24'(-4628);
			35876: out = 24'(-5288);
			35877: out = 24'(-1956);
			35878: out = 24'(-376);
			35879: out = 24'(244);
			35880: out = 24'(416);
			35881: out = 24'(4428);
			35882: out = 24'(1868);
			35883: out = 24'(-1904);
			35884: out = 24'(-3824);
			35885: out = 24'(-1432);
			35886: out = 24'(-1408);
			35887: out = 24'(-752);
			35888: out = 24'(1292);
			35889: out = 24'(6812);
			35890: out = 24'(1424);
			35891: out = 24'(-668);
			35892: out = 24'(860);
			35893: out = 24'(3344);
			35894: out = 24'(252);
			35895: out = 24'(268);
			35896: out = 24'(612);
			35897: out = 24'(-312);
			35898: out = 24'(4016);
			35899: out = 24'(4148);
			35900: out = 24'(452);
			35901: out = 24'(-4652);
			35902: out = 24'(-1692);
			35903: out = 24'(-604);
			35904: out = 24'(-96);
			35905: out = 24'(232);
			35906: out = 24'(3248);
			35907: out = 24'(688);
			35908: out = 24'(-2448);
			35909: out = 24'(-4224);
			35910: out = 24'(-1520);
			35911: out = 24'(-6304);
			35912: out = 24'(-3120);
			35913: out = 24'(3868);
			35914: out = 24'(6980);
			35915: out = 24'(1180);
			35916: out = 24'(-2660);
			35917: out = 24'(-1732);
			35918: out = 24'(-232);
			35919: out = 24'(312);
			35920: out = 24'(-4104);
			35921: out = 24'(-3620);
			35922: out = 24'(868);
			35923: out = 24'(864);
			35924: out = 24'(-2212);
			35925: out = 24'(-6024);
			35926: out = 24'(-4984);
			35927: out = 24'(1388);
			35928: out = 24'(348);
			35929: out = 24'(364);
			35930: out = 24'(-208);
			35931: out = 24'(-1048);
			35932: out = 24'(592);
			35933: out = 24'(3732);
			35934: out = 24'(4508);
			35935: out = 24'(3588);
			35936: out = 24'(4292);
			35937: out = 24'(2808);
			35938: out = 24'(-2984);
			35939: out = 24'(-8452);
			35940: out = 24'(-6812);
			35941: out = 24'(-676);
			35942: out = 24'(1056);
			35943: out = 24'(1136);
			35944: out = 24'(6880);
			35945: out = 24'(4456);
			35946: out = 24'(-1972);
			35947: out = 24'(-7876);
			35948: out = 24'(-5976);
			35949: out = 24'(-3496);
			35950: out = 24'(-692);
			35951: out = 24'(1592);
			35952: out = 24'(5308);
			35953: out = 24'(6488);
			35954: out = 24'(4948);
			35955: out = 24'(1588);
			35956: out = 24'(-384);
			35957: out = 24'(-1688);
			35958: out = 24'(-4300);
			35959: out = 24'(-5460);
			35960: out = 24'(-2588);
			35961: out = 24'(972);
			35962: out = 24'(1688);
			35963: out = 24'(-292);
			35964: out = 24'(-1192);
			35965: out = 24'(260);
			35966: out = 24'(4036);
			35967: out = 24'(2512);
			35968: out = 24'(-2252);
			35969: out = 24'(-5224);
			35970: out = 24'(-4340);
			35971: out = 24'(-1048);
			35972: out = 24'(508);
			35973: out = 24'(12);
			35974: out = 24'(40);
			35975: out = 24'(2412);
			35976: out = 24'(4324);
			35977: out = 24'(1368);
			35978: out = 24'(-7500);
			35979: out = 24'(-3788);
			35980: out = 24'(4256);
			35981: out = 24'(6756);
			35982: out = 24'(-372);
			35983: out = 24'(908);
			35984: out = 24'(492);
			35985: out = 24'(-860);
			35986: out = 24'(-2824);
			35987: out = 24'(-1736);
			35988: out = 24'(-572);
			35989: out = 24'(-168);
			35990: out = 24'(824);
			35991: out = 24'(6256);
			35992: out = 24'(5088);
			35993: out = 24'(-692);
			35994: out = 24'(-6072);
			35995: out = 24'(-5280);
			35996: out = 24'(-596);
			35997: out = 24'(1196);
			35998: out = 24'(-352);
			35999: out = 24'(324);
			36000: out = 24'(-248);
			36001: out = 24'(324);
			36002: out = 24'(-528);
			36003: out = 24'(-1240);
			36004: out = 24'(-204);
			36005: out = 24'(-1056);
			36006: out = 24'(-5028);
			36007: out = 24'(-7124);
			36008: out = 24'(-456);
			36009: out = 24'(3948);
			36010: out = 24'(3724);
			36011: out = 24'(932);
			36012: out = 24'(1480);
			36013: out = 24'(1064);
			36014: out = 24'(716);
			36015: out = 24'(-740);
			36016: out = 24'(-4060);
			36017: out = 24'(-4936);
			36018: out = 24'(-3572);
			36019: out = 24'(812);
			36020: out = 24'(3256);
			36021: out = 24'(1356);
			36022: out = 24'(-3788);
			36023: out = 24'(-2524);
			36024: out = 24'(4612);
			36025: out = 24'(6692);
			36026: out = 24'(3148);
			36027: out = 24'(68);
			36028: out = 24'(36);
			36029: out = 24'(120);
			36030: out = 24'(-5072);
			36031: out = 24'(-4128);
			36032: out = 24'(3348);
			36033: out = 24'(6148);
			36034: out = 24'(2780);
			36035: out = 24'(-1820);
			36036: out = 24'(-1816);
			36037: out = 24'(1336);
			36038: out = 24'(136);
			36039: out = 24'(-36);
			36040: out = 24'(-64);
			36041: out = 24'(372);
			36042: out = 24'(2976);
			36043: out = 24'(2556);
			36044: out = 24'(-1776);
			36045: out = 24'(-4752);
			36046: out = 24'(704);
			36047: out = 24'(5668);
			36048: out = 24'(4592);
			36049: out = 24'(148);
			36050: out = 24'(-28);
			36051: out = 24'(-2176);
			36052: out = 24'(-5932);
			36053: out = 24'(-7256);
			36054: out = 24'(-784);
			36055: out = 24'(2588);
			36056: out = 24'(2676);
			36057: out = 24'(-500);
			36058: out = 24'(-1124);
			36059: out = 24'(-504);
			36060: out = 24'(348);
			36061: out = 24'(-928);
			36062: out = 24'(-720);
			36063: out = 24'(3972);
			36064: out = 24'(4372);
			36065: out = 24'(360);
			36066: out = 24'(-3572);
			36067: out = 24'(-5568);
			36068: out = 24'(-3140);
			36069: out = 24'(-2936);
			36070: out = 24'(-1100);
			36071: out = 24'(3696);
			36072: out = 24'(6588);
			36073: out = 24'(3132);
			36074: out = 24'(-1392);
			36075: out = 24'(-2996);
			36076: out = 24'(-6088);
			36077: out = 24'(-5040);
			36078: out = 24'(1468);
			36079: out = 24'(6560);
			36080: out = 24'(4332);
			36081: out = 24'(-5816);
			36082: out = 24'(-7268);
			36083: out = 24'(124);
			36084: out = 24'(-308);
			36085: out = 24'(-588);
			36086: out = 24'(-888);
			36087: out = 24'(628);
			36088: out = 24'(184);
			36089: out = 24'(1052);
			36090: out = 24'(2964);
			36091: out = 24'(1700);
			36092: out = 24'(-5612);
			36093: out = 24'(-6356);
			36094: out = 24'(-2548);
			36095: out = 24'(1516);
			36096: out = 24'(816);
			36097: out = 24'(672);
			36098: out = 24'(88);
			36099: out = 24'(752);
			36100: out = 24'(1224);
			36101: out = 24'(124);
			36102: out = 24'(2936);
			36103: out = 24'(2020);
			36104: out = 24'(-2928);
			36105: out = 24'(-6088);
			36106: out = 24'(-3752);
			36107: out = 24'(1024);
			36108: out = 24'(5360);
			36109: out = 24'(7712);
			36110: out = 24'(5488);
			36111: out = 24'(216);
			36112: out = 24'(-3780);
			36113: out = 24'(-3600);
			36114: out = 24'(-1760);
			36115: out = 24'(-2032);
			36116: out = 24'(-1960);
			36117: out = 24'(1368);
			36118: out = 24'(6256);
			36119: out = 24'(1792);
			36120: out = 24'(-4884);
			36121: out = 24'(-5204);
			36122: out = 24'(-152);
			36123: out = 24'(708);
			36124: out = 24'(-1064);
			36125: out = 24'(396);
			36126: out = 24'(4572);
			36127: out = 24'(5348);
			36128: out = 24'(-348);
			36129: out = 24'(-4248);
			36130: out = 24'(-2224);
			36131: out = 24'(1132);
			36132: out = 24'(-1212);
			36133: out = 24'(-1032);
			36134: out = 24'(4456);
			36135: out = 24'(4332);
			36136: out = 24'(1688);
			36137: out = 24'(-760);
			36138: out = 24'(664);
			36139: out = 24'(1888);
			36140: out = 24'(-1916);
			36141: out = 24'(-6320);
			36142: out = 24'(-5144);
			36143: out = 24'(240);
			36144: out = 24'(3056);
			36145: out = 24'(4260);
			36146: out = 24'(4384);
			36147: out = 24'(3156);
			36148: out = 24'(1332);
			36149: out = 24'(-2952);
			36150: out = 24'(-7092);
			36151: out = 24'(-7040);
			36152: out = 24'(-148);
			36153: out = 24'(5492);
			36154: out = 24'(6192);
			36155: out = 24'(3884);
			36156: out = 24'(956);
			36157: out = 24'(476);
			36158: out = 24'(-3832);
			36159: out = 24'(-8348);
			36160: out = 24'(-3460);
			36161: out = 24'(2632);
			36162: out = 24'(5288);
			36163: out = 24'(624);
			36164: out = 24'(-5088);
			36165: out = 24'(-2636);
			36166: out = 24'(2100);
			36167: out = 24'(2688);
			36168: out = 24'(-460);
			36169: out = 24'(-2644);
			36170: out = 24'(-1100);
			36171: out = 24'(724);
			36172: out = 24'(80);
			36173: out = 24'(-6492);
			36174: out = 24'(1156);
			36175: out = 24'(7012);
			36176: out = 24'(4212);
			36177: out = 24'(-5200);
			36178: out = 24'(-7008);
			36179: out = 24'(-4556);
			36180: out = 24'(-3128);
			36181: out = 24'(-6644);
			36182: out = 24'(-856);
			36183: out = 24'(4636);
			36184: out = 24'(9288);
			36185: out = 24'(5760);
			36186: out = 24'(-3776);
			36187: out = 24'(-17112);
			36188: out = 24'(-14304);
			36189: out = 24'(1984);
			36190: out = 24'(7336);
			36191: out = 24'(6600);
			36192: out = 24'(3096);
			36193: out = 24'(1308);
			36194: out = 24'(1312);
			36195: out = 24'(-1996);
			36196: out = 24'(-1172);
			36197: out = 24'(-224);
			36198: out = 24'(-3708);
			36199: out = 24'(-1952);
			36200: out = 24'(2300);
			36201: out = 24'(1720);
			36202: out = 24'(-5188);
			36203: out = 24'(-356);
			36204: out = 24'(5084);
			36205: out = 24'(4936);
			36206: out = 24'(-2224);
			36207: out = 24'(212);
			36208: out = 24'(16);
			36209: out = 24'(-300);
			36210: out = 24'(-580);
			36211: out = 24'(4816);
			36212: out = 24'(6496);
			36213: out = 24'(3368);
			36214: out = 24'(-3532);
			36215: out = 24'(-4792);
			36216: out = 24'(-8260);
			36217: out = 24'(-4308);
			36218: out = 24'(672);
			36219: out = 24'(3908);
			36220: out = 24'(5832);
			36221: out = 24'(6472);
			36222: out = 24'(4932);
			36223: out = 24'(2272);
			36224: out = 24'(-3344);
			36225: out = 24'(-3244);
			36226: out = 24'(-1420);
			36227: out = 24'(284);
			36228: out = 24'(-268);
			36229: out = 24'(3320);
			36230: out = 24'(2456);
			36231: out = 24'(-1280);
			36232: out = 24'(-3536);
			36233: out = 24'(-1060);
			36234: out = 24'(-568);
			36235: out = 24'(-1468);
			36236: out = 24'(-108);
			36237: out = 24'(-1356);
			36238: out = 24'(-652);
			36239: out = 24'(2212);
			36240: out = 24'(7364);
			36241: out = 24'(3740);
			36242: out = 24'(1660);
			36243: out = 24'(-3332);
			36244: out = 24'(-5592);
			36245: out = 24'(-1852);
			36246: out = 24'(3164);
			36247: out = 24'(2348);
			36248: out = 24'(-836);
			36249: out = 24'(-1444);
			36250: out = 24'(-108);
			36251: out = 24'(-2540);
			36252: out = 24'(-4868);
			36253: out = 24'(-1728);
			36254: out = 24'(4832);
			36255: out = 24'(3960);
			36256: out = 24'(-1184);
			36257: out = 24'(-1812);
			36258: out = 24'(-856);
			36259: out = 24'(2684);
			36260: out = 24'(620);
			36261: out = 24'(-4380);
			36262: out = 24'(-4552);
			36263: out = 24'(-1524);
			36264: out = 24'(1136);
			36265: out = 24'(428);
			36266: out = 24'(-872);
			36267: out = 24'(2488);
			36268: out = 24'(6004);
			36269: out = 24'(3496);
			36270: out = 24'(-3844);
			36271: out = 24'(-5076);
			36272: out = 24'(-2544);
			36273: out = 24'(-1864);
			36274: out = 24'(-3076);
			36275: out = 24'(2308);
			36276: out = 24'(5792);
			36277: out = 24'(3144);
			36278: out = 24'(-3532);
			36279: out = 24'(-5700);
			36280: out = 24'(-2160);
			36281: out = 24'(712);
			36282: out = 24'(-248);
			36283: out = 24'(404);
			36284: out = 24'(-220);
			36285: out = 24'(48);
			36286: out = 24'(40);
			36287: out = 24'(20);
			36288: out = 24'(-1856);
			36289: out = 24'(-1524);
			36290: out = 24'(2360);
			36291: out = 24'(5484);
			36292: out = 24'(1296);
			36293: out = 24'(-5808);
			36294: out = 24'(-6652);
			36295: out = 24'(76);
			36296: out = 24'(3696);
			36297: out = 24'(3816);
			36298: out = 24'(2964);
			36299: out = 24'(2904);
			36300: out = 24'(1020);
			36301: out = 24'(-3544);
			36302: out = 24'(-2824);
			36303: out = 24'(3280);
			36304: out = 24'(6164);
			36305: out = 24'(2532);
			36306: out = 24'(-3224);
			36307: out = 24'(-3812);
			36308: out = 24'(320);
			36309: out = 24'(3428);
			36310: out = 24'(3712);
			36311: out = 24'(1712);
			36312: out = 24'(-348);
			36313: out = 24'(616);
			36314: out = 24'(-2940);
			36315: out = 24'(-6304);
			36316: out = 24'(-4528);
			36317: out = 24'(2408);
			36318: out = 24'(5812);
			36319: out = 24'(4316);
			36320: out = 24'(3500);
			36321: out = 24'(6212);
			36322: out = 24'(1492);
			36323: out = 24'(-7024);
			36324: out = 24'(-10188);
			36325: out = 24'(-1828);
			36326: out = 24'(136);
			36327: out = 24'(1376);
			36328: out = 24'(392);
			36329: out = 24'(-80);
			36330: out = 24'(-188);
			36331: out = 24'(412);
			36332: out = 24'(1548);
			36333: out = 24'(2764);
			36334: out = 24'(-396);
			36335: out = 24'(-1264);
			36336: out = 24'(-1156);
			36337: out = 24'(224);
			36338: out = 24'(592);
			36339: out = 24'(876);
			36340: out = 24'(-692);
			36341: out = 24'(-1948);
			36342: out = 24'(-2704);
			36343: out = 24'(208);
			36344: out = 24'(-1024);
			36345: out = 24'(-2944);
			36346: out = 24'(-868);
			36347: out = 24'(-664);
			36348: out = 24'(2368);
			36349: out = 24'(1904);
			36350: out = 24'(-312);
			36351: out = 24'(-276);
			36352: out = 24'(2168);
			36353: out = 24'(1896);
			36354: out = 24'(-652);
			36355: out = 24'(764);
			36356: out = 24'(-1172);
			36357: out = 24'(-2296);
			36358: out = 24'(-2308);
			36359: out = 24'(100);
			36360: out = 24'(2224);
			36361: out = 24'(3296);
			36362: out = 24'(1772);
			36363: out = 24'(-388);
			36364: out = 24'(-344);
			36365: out = 24'(-960);
			36366: out = 24'(-2056);
			36367: out = 24'(-1216);
			36368: out = 24'(-636);
			36369: out = 24'(2860);
			36370: out = 24'(3000);
			36371: out = 24'(-884);
			36372: out = 24'(-6012);
			36373: out = 24'(-3912);
			36374: out = 24'(-752);
			36375: out = 24'(852);
			36376: out = 24'(928);
			36377: out = 24'(3348);
			36378: out = 24'(2604);
			36379: out = 24'(-944);
			36380: out = 24'(-2396);
			36381: out = 24'(-232);
			36382: out = 24'(2940);
			36383: out = 24'(3524);
			36384: out = 24'(2276);
			36385: out = 24'(-2580);
			36386: out = 24'(-2288);
			36387: out = 24'(-1596);
			36388: out = 24'(-2064);
			36389: out = 24'(-5076);
			36390: out = 24'(-704);
			36391: out = 24'(1400);
			36392: out = 24'(468);
			36393: out = 24'(-104);
			36394: out = 24'(-208);
			36395: out = 24'(-1420);
			36396: out = 24'(-2828);
			36397: out = 24'(-1028);
			36398: out = 24'(2120);
			36399: out = 24'(3532);
			36400: out = 24'(992);
			36401: out = 24'(-2876);
			36402: out = 24'(-1664);
			36403: out = 24'(-164);
			36404: out = 24'(972);
			36405: out = 24'(580);
			36406: out = 24'(-112);
			36407: out = 24'(336);
			36408: out = 24'(724);
			36409: out = 24'(-1260);
			36410: out = 24'(-3440);
			36411: out = 24'(-2756);
			36412: out = 24'(2692);
			36413: out = 24'(5604);
			36414: out = 24'(2556);
			36415: out = 24'(104);
			36416: out = 24'(-1028);
			36417: out = 24'(-3264);
			36418: out = 24'(-6124);
			36419: out = 24'(-4496);
			36420: out = 24'(3116);
			36421: out = 24'(7784);
			36422: out = 24'(5444);
			36423: out = 24'(80);
			36424: out = 24'(-116);
			36425: out = 24'(192);
			36426: out = 24'(-152);
			36427: out = 24'(2596);
			36428: out = 24'(436);
			36429: out = 24'(-3116);
			36430: out = 24'(-5092);
			36431: out = 24'(-2484);
			36432: out = 24'(5048);
			36433: out = 24'(5340);
			36434: out = 24'(116);
			36435: out = 24'(-4032);
			36436: out = 24'(-2140);
			36437: out = 24'(-4292);
			36438: out = 24'(-6840);
			36439: out = 24'(-3632);
			36440: out = 24'(1912);
			36441: out = 24'(4544);
			36442: out = 24'(860);
			36443: out = 24'(-2284);
			36444: out = 24'(2780);
			36445: out = 24'(5232);
			36446: out = 24'(3260);
			36447: out = 24'(-1840);
			36448: out = 24'(-2264);
			36449: out = 24'(-1536);
			36450: out = 24'(2004);
			36451: out = 24'(1492);
			36452: out = 24'(-1952);
			36453: out = 24'(-6212);
			36454: out = 24'(-2784);
			36455: out = 24'(540);
			36456: out = 24'(488);
			36457: out = 24'(-352);
			36458: out = 24'(2616);
			36459: out = 24'(2628);
			36460: out = 24'(-796);
			36461: out = 24'(864);
			36462: out = 24'(2112);
			36463: out = 24'(1728);
			36464: out = 24'(-1724);
			36465: out = 24'(-3560);
			36466: out = 24'(-1484);
			36467: out = 24'(1748);
			36468: out = 24'(2292);
			36469: out = 24'(232);
			36470: out = 24'(-1496);
			36471: out = 24'(-1328);
			36472: out = 24'(0);
			36473: out = 24'(496);
			36474: out = 24'(-128);
			36475: out = 24'(-868);
			36476: out = 24'(2232);
			36477: out = 24'(6296);
			36478: out = 24'(-696);
			36479: out = 24'(-2128);
			36480: out = 24'(-3992);
			36481: out = 24'(-3460);
			36482: out = 24'(-2028);
			36483: out = 24'(2152);
			36484: out = 24'(1888);
			36485: out = 24'(360);
			36486: out = 24'(368);
			36487: out = 24'(-168);
			36488: out = 24'(-1448);
			36489: out = 24'(-584);
			36490: out = 24'(2980);
			36491: out = 24'(2696);
			36492: out = 24'(-220);
			36493: out = 24'(-1828);
			36494: out = 24'(1444);
			36495: out = 24'(4836);
			36496: out = 24'(4828);
			36497: out = 24'(-280);
			36498: out = 24'(-4576);
			36499: out = 24'(-1940);
			36500: out = 24'(-4532);
			36501: out = 24'(-6900);
			36502: out = 24'(-6768);
			36503: out = 24'(-1140);
			36504: out = 24'(-864);
			36505: out = 24'(2400);
			36506: out = 24'(3016);
			36507: out = 24'(-796);
			36508: out = 24'(-1340);
			36509: out = 24'(-1852);
			36510: out = 24'(-1864);
			36511: out = 24'(-2936);
			36512: out = 24'(-2552);
			36513: out = 24'(-2036);
			36514: out = 24'(-308);
			36515: out = 24'(1548);
			36516: out = 24'(3984);
			36517: out = 24'(916);
			36518: out = 24'(-656);
			36519: out = 24'(676);
			36520: out = 24'(2620);
			36521: out = 24'(-360);
			36522: out = 24'(-5188);
			36523: out = 24'(-6768);
			36524: out = 24'(-1796);
			36525: out = 24'(-684);
			36526: out = 24'(2768);
			36527: out = 24'(4084);
			36528: out = 24'(2408);
			36529: out = 24'(-2112);
			36530: out = 24'(-2880);
			36531: out = 24'(-2048);
			36532: out = 24'(-1104);
			36533: out = 24'(-36);
			36534: out = 24'(2260);
			36535: out = 24'(3360);
			36536: out = 24'(2424);
			36537: out = 24'(1076);
			36538: out = 24'(3040);
			36539: out = 24'(5276);
			36540: out = 24'(4272);
			36541: out = 24'(-920);
			36542: out = 24'(-2348);
			36543: out = 24'(-3292);
			36544: out = 24'(-1900);
			36545: out = 24'(36);
			36546: out = 24'(3528);
			36547: out = 24'(1244);
			36548: out = 24'(-2080);
			36549: out = 24'(-4196);
			36550: out = 24'(-4904);
			36551: out = 24'(-1908);
			36552: out = 24'(2944);
			36553: out = 24'(5580);
			36554: out = 24'(2688);
			36555: out = 24'(-732);
			36556: out = 24'(-1144);
			36557: out = 24'(1504);
			36558: out = 24'(2344);
			36559: out = 24'(404);
			36560: out = 24'(-1600);
			36561: out = 24'(-1192);
			36562: out = 24'(-316);
			36563: out = 24'(2624);
			36564: out = 24'(16);
			36565: out = 24'(-2276);
			36566: out = 24'(-1836);
			36567: out = 24'(-5156);
			36568: out = 24'(-1088);
			36569: out = 24'(2228);
			36570: out = 24'(2084);
			36571: out = 24'(-1468);
			36572: out = 24'(-1964);
			36573: out = 24'(-728);
			36574: out = 24'(-492);
			36575: out = 24'(-1556);
			36576: out = 24'(-1848);
			36577: out = 24'(968);
			36578: out = 24'(2912);
			36579: out = 24'(356);
			36580: out = 24'(824);
			36581: out = 24'(-80);
			36582: out = 24'(-952);
			36583: out = 24'(-3228);
			36584: out = 24'(-3464);
			36585: out = 24'(-4208);
			36586: out = 24'(-2052);
			36587: out = 24'(396);
			36588: out = 24'(3100);
			36589: out = 24'(2804);
			36590: out = 24'(3228);
			36591: out = 24'(1944);
			36592: out = 24'(-120);
			36593: out = 24'(-5520);
			36594: out = 24'(-4048);
			36595: out = 24'(-520);
			36596: out = 24'(800);
			36597: out = 24'(660);
			36598: out = 24'(2596);
			36599: out = 24'(632);
			36600: out = 24'(-5316);
			36601: out = 24'(-3932);
			36602: out = 24'(1372);
			36603: out = 24'(4452);
			36604: out = 24'(2500);
			36605: out = 24'(3020);
			36606: out = 24'(784);
			36607: out = 24'(-3708);
			36608: out = 24'(-7380);
			36609: out = 24'(-2280);
			36610: out = 24'(-56);
			36611: out = 24'(56);
			36612: out = 24'(-1980);
			36613: out = 24'(-1084);
			36614: out = 24'(-1652);
			36615: out = 24'(-408);
			36616: out = 24'(292);
			36617: out = 24'(1076);
			36618: out = 24'(-256);
			36619: out = 24'(-952);
			36620: out = 24'(-1592);
			36621: out = 24'(-1024);
			36622: out = 24'(604);
			36623: out = 24'(440);
			36624: out = 24'(80);
			36625: out = 24'(1508);
			36626: out = 24'(2780);
			36627: out = 24'(5672);
			36628: out = 24'(3192);
			36629: out = 24'(-2640);
			36630: out = 24'(-8400);
			36631: out = 24'(-820);
			36632: out = 24'(1504);
			36633: out = 24'(-312);
			36634: out = 24'(-1220);
			36635: out = 24'(-276);
			36636: out = 24'(-620);
			36637: out = 24'(-2148);
			36638: out = 24'(-2096);
			36639: out = 24'(-244);
			36640: out = 24'(1728);
			36641: out = 24'(1376);
			36642: out = 24'(-520);
			36643: out = 24'(-1196);
			36644: out = 24'(-1556);
			36645: out = 24'(-616);
			36646: out = 24'(292);
			36647: out = 24'(1212);
			36648: out = 24'(3648);
			36649: out = 24'(2308);
			36650: out = 24'(-2184);
			36651: out = 24'(-3908);
			36652: out = 24'(1556);
			36653: out = 24'(8148);
			36654: out = 24'(6124);
			36655: out = 24'(-3216);
			36656: out = 24'(-7836);
			36657: out = 24'(-4332);
			36658: out = 24'(736);
			36659: out = 24'(424);
			36660: out = 24'(564);
			36661: out = 24'(68);
			36662: out = 24'(3920);
			36663: out = 24'(5428);
			36664: out = 24'(2692);
			36665: out = 24'(-4680);
			36666: out = 24'(-6280);
			36667: out = 24'(-3712);
			36668: out = 24'(-1264);
			36669: out = 24'(-208);
			36670: out = 24'(1836);
			36671: out = 24'(3432);
			36672: out = 24'(2672);
			36673: out = 24'(936);
			36674: out = 24'(656);
			36675: out = 24'(664);
			36676: out = 24'(-412);
			36677: out = 24'(1048);
			36678: out = 24'(-3440);
			36679: out = 24'(-6668);
			36680: out = 24'(-5988);
			36681: out = 24'(1472);
			36682: out = 24'(-76);
			36683: out = 24'(1784);
			36684: out = 24'(3256);
			36685: out = 24'(2892);
			36686: out = 24'(-1036);
			36687: out = 24'(-760);
			36688: out = 24'(-32);
			36689: out = 24'(-96);
			36690: out = 24'(-304);
			36691: out = 24'(240);
			36692: out = 24'(-2452);
			36693: out = 24'(-6508);
			36694: out = 24'(-5924);
			36695: out = 24'(-1492);
			36696: out = 24'(1080);
			36697: out = 24'(1616);
			36698: out = 24'(4300);
			36699: out = 24'(3444);
			36700: out = 24'(948);
			36701: out = 24'(-2552);
			36702: out = 24'(-4656);
			36703: out = 24'(-3748);
			36704: out = 24'(-1504);
			36705: out = 24'(2500);
			36706: out = 24'(5848);
			36707: out = 24'(908);
			36708: out = 24'(-2840);
			36709: out = 24'(-1824);
			36710: out = 24'(1360);
			36711: out = 24'(280);
			36712: out = 24'(-4308);
			36713: out = 24'(-4500);
			36714: out = 24'(-60);
			36715: out = 24'(-76);
			36716: out = 24'(1300);
			36717: out = 24'(1696);
			36718: out = 24'(2312);
			36719: out = 24'(960);
			36720: out = 24'(456);
			36721: out = 24'(-124);
			36722: out = 24'(224);
			36723: out = 24'(96);
			36724: out = 24'(1024);
			36725: out = 24'(2420);
			36726: out = 24'(2788);
			36727: out = 24'(436);
			36728: out = 24'(164);
			36729: out = 24'(-3712);
			36730: out = 24'(-5008);
			36731: out = 24'(-4192);
			36732: out = 24'(-1020);
			36733: out = 24'(-364);
			36734: out = 24'(3624);
			36735: out = 24'(7588);
			36736: out = 24'(5504);
			36737: out = 24'(3856);
			36738: out = 24'(964);
			36739: out = 24'(-904);
			36740: out = 24'(-3072);
			36741: out = 24'(-6656);
			36742: out = 24'(-5784);
			36743: out = 24'(-628);
			36744: out = 24'(3592);
			36745: out = 24'(6952);
			36746: out = 24'(4220);
			36747: out = 24'(2000);
			36748: out = 24'(-440);
			36749: out = 24'(-4616);
			36750: out = 24'(-10788);
			36751: out = 24'(-10852);
			36752: out = 24'(-4284);
			36753: out = 24'(3456);
			36754: out = 24'(7948);
			36755: out = 24'(8120);
			36756: out = 24'(3340);
			36757: out = 24'(-2548);
			36758: out = 24'(-7080);
			36759: out = 24'(-3672);
			36760: out = 24'(-964);
			36761: out = 24'(-2116);
			36762: out = 24'(928);
			36763: out = 24'(3656);
			36764: out = 24'(2120);
			36765: out = 24'(-3040);
			36766: out = 24'(-2024);
			36767: out = 24'(-2344);
			36768: out = 24'(-2824);
			36769: out = 24'(-2232);
			36770: out = 24'(3548);
			36771: out = 24'(5800);
			36772: out = 24'(4012);
			36773: out = 24'(-120);
			36774: out = 24'(536);
			36775: out = 24'(-1480);
			36776: out = 24'(-312);
			36777: out = 24'(192);
			36778: out = 24'(764);
			36779: out = 24'(-4448);
			36780: out = 24'(-1840);
			36781: out = 24'(1644);
			36782: out = 24'(3412);
			36783: out = 24'(2980);
			36784: out = 24'(4040);
			36785: out = 24'(2032);
			36786: out = 24'(-3552);
			36787: out = 24'(-10620);
			36788: out = 24'(-6856);
			36789: out = 24'(232);
			36790: out = 24'(5420);
			36791: out = 24'(5636);
			36792: out = 24'(3260);
			36793: out = 24'(-2132);
			36794: out = 24'(-5032);
			36795: out = 24'(-3316);
			36796: out = 24'(-3628);
			36797: out = 24'(-2156);
			36798: out = 24'(868);
			36799: out = 24'(4972);
			36800: out = 24'(6740);
			36801: out = 24'(4720);
			36802: out = 24'(1340);
			36803: out = 24'(-740);
			36804: out = 24'(-4804);
			36805: out = 24'(-2280);
			36806: out = 24'(-140);
			36807: out = 24'(1100);
			36808: out = 24'(1000);
			36809: out = 24'(364);
			36810: out = 24'(-884);
			36811: out = 24'(-1060);
			36812: out = 24'(232);
			36813: out = 24'(2792);
			36814: out = 24'(876);
			36815: out = 24'(-3540);
			36816: out = 24'(-5552);
			36817: out = 24'(-1832);
			36818: out = 24'(2704);
			36819: out = 24'(4660);
			36820: out = 24'(3244);
			36821: out = 24'(-1168);
			36822: out = 24'(-2432);
			36823: out = 24'(-2504);
			36824: out = 24'(-2508);
			36825: out = 24'(-2316);
			36826: out = 24'(-420);
			36827: out = 24'(832);
			36828: out = 24'(1544);
			36829: out = 24'(3424);
			36830: out = 24'(3016);
			36831: out = 24'(3232);
			36832: out = 24'(2248);
			36833: out = 24'(832);
			36834: out = 24'(-252);
			36835: out = 24'(-56);
			36836: out = 24'(-2204);
			36837: out = 24'(-5084);
			36838: out = 24'(-3688);
			36839: out = 24'(1768);
			36840: out = 24'(5756);
			36841: out = 24'(4724);
			36842: out = 24'(-204);
			36843: out = 24'(456);
			36844: out = 24'(-888);
			36845: out = 24'(-3244);
			36846: out = 24'(-2144);
			36847: out = 24'(-20);
			36848: out = 24'(4220);
			36849: out = 24'(5420);
			36850: out = 24'(1916);
			36851: out = 24'(-2988);
			36852: out = 24'(-5320);
			36853: out = 24'(-3196);
			36854: out = 24'(612);
			36855: out = 24'(3688);
			36856: out = 24'(3252);
			36857: out = 24'(1972);
			36858: out = 24'(140);
			36859: out = 24'(-1484);
			36860: out = 24'(-4512);
			36861: out = 24'(-4228);
			36862: out = 24'(-1688);
			36863: out = 24'(852);
			36864: out = 24'(2464);
			36865: out = 24'(3756);
			36866: out = 24'(2940);
			36867: out = 24'(132);
			36868: out = 24'(-7780);
			36869: out = 24'(-5668);
			36870: out = 24'(392);
			36871: out = 24'(4132);
			36872: out = 24'(3816);
			36873: out = 24'(3380);
			36874: out = 24'(900);
			36875: out = 24'(-2180);
			36876: out = 24'(-2788);
			36877: out = 24'(-1856);
			36878: out = 24'(-2140);
			36879: out = 24'(-2132);
			36880: out = 24'(672);
			36881: out = 24'(-1064);
			36882: out = 24'(-1856);
			36883: out = 24'(-28);
			36884: out = 24'(2768);
			36885: out = 24'(664);
			36886: out = 24'(-5444);
			36887: out = 24'(-8164);
			36888: out = 24'(-3448);
			36889: out = 24'(84);
			36890: out = 24'(4892);
			36891: out = 24'(7452);
			36892: out = 24'(7352);
			36893: out = 24'(792);
			36894: out = 24'(-1704);
			36895: out = 24'(-1812);
			36896: out = 24'(276);
			36897: out = 24'(-744);
			36898: out = 24'(-2168);
			36899: out = 24'(-5824);
			36900: out = 24'(-4684);
			36901: out = 24'(1112);
			36902: out = 24'(5700);
			36903: out = 24'(2672);
			36904: out = 24'(-976);
			36905: out = 24'(324);
			36906: out = 24'(-520);
			36907: out = 24'(-488);
			36908: out = 24'(-2556);
			36909: out = 24'(-2816);
			36910: out = 24'(-1632);
			36911: out = 24'(2568);
			36912: out = 24'(3400);
			36913: out = 24'(2040);
			36914: out = 24'(-320);
			36915: out = 24'(824);
			36916: out = 24'(-1388);
			36917: out = 24'(-3392);
			36918: out = 24'(-836);
			36919: out = 24'(4184);
			36920: out = 24'(4296);
			36921: out = 24'(476);
			36922: out = 24'(-2696);
			36923: out = 24'(-5344);
			36924: out = 24'(-2368);
			36925: out = 24'(2404);
			36926: out = 24'(5092);
			36927: out = 24'(3500);
			36928: out = 24'(-780);
			36929: out = 24'(-3896);
			36930: out = 24'(-4228);
			36931: out = 24'(-3320);
			36932: out = 24'(-872);
			36933: out = 24'(1592);
			36934: out = 24'(2240);
			36935: out = 24'(-320);
			36936: out = 24'(-32);
			36937: out = 24'(280);
			36938: out = 24'(1464);
			36939: out = 24'(2588);
			36940: out = 24'(3396);
			36941: out = 24'(1196);
			36942: out = 24'(-1468);
			36943: out = 24'(-2600);
			36944: out = 24'(-4552);
			36945: out = 24'(-3036);
			36946: out = 24'(-1140);
			36947: out = 24'(1328);
			36948: out = 24'(2176);
			36949: out = 24'(1052);
			36950: out = 24'(-3728);
			36951: out = 24'(-6272);
			36952: out = 24'(-2992);
			36953: out = 24'(1864);
			36954: out = 24'(1640);
			36955: out = 24'(-628);
			36956: out = 24'(508);
			36957: out = 24'(5200);
			36958: out = 24'(4548);
			36959: out = 24'(0);
			36960: out = 24'(-3340);
			36961: out = 24'(-696);
			36962: out = 24'(-1468);
			36963: out = 24'(-3560);
			36964: out = 24'(-3564);
			36965: out = 24'(568);
			36966: out = 24'(1016);
			36967: out = 24'(416);
			36968: out = 24'(336);
			36969: out = 24'(2764);
			36970: out = 24'(276);
			36971: out = 24'(-124);
			36972: out = 24'(-660);
			36973: out = 24'(-2412);
			36974: out = 24'(-5088);
			36975: out = 24'(-868);
			36976: out = 24'(4992);
			36977: out = 24'(5068);
			36978: out = 24'(908);
			36979: out = 24'(-4900);
			36980: out = 24'(-5948);
			36981: out = 24'(-3592);
			36982: out = 24'(-1136);
			36983: out = 24'(-320);
			36984: out = 24'(2776);
			36985: out = 24'(6912);
			36986: out = 24'(5472);
			36987: out = 24'(808);
			36988: out = 24'(-4124);
			36989: out = 24'(-1848);
			36990: out = 24'(5120);
			36991: out = 24'(3360);
			36992: out = 24'(-1304);
			36993: out = 24'(-2920);
			36994: out = 24'(96);
			36995: out = 24'(-1316);
			36996: out = 24'(-1504);
			36997: out = 24'(304);
			36998: out = 24'(3788);
			36999: out = 24'(2348);
			37000: out = 24'(-1296);
			37001: out = 24'(-4800);
			37002: out = 24'(-3244);
			37003: out = 24'(-484);
			37004: out = 24'(2548);
			37005: out = 24'(1032);
			37006: out = 24'(464);
			37007: out = 24'(3448);
			37008: out = 24'(2852);
			37009: out = 24'(172);
			37010: out = 24'(-1524);
			37011: out = 24'(-212);
			37012: out = 24'(-3164);
			37013: out = 24'(-2520);
			37014: out = 24'(372);
			37015: out = 24'(2256);
			37016: out = 24'(-1020);
			37017: out = 24'(-3220);
			37018: out = 24'(-1052);
			37019: out = 24'(2904);
			37020: out = 24'(-460);
			37021: out = 24'(2064);
			37022: out = 24'(1624);
			37023: out = 24'(-2236);
			37024: out = 24'(-8364);
			37025: out = 24'(-3032);
			37026: out = 24'(2208);
			37027: out = 24'(2100);
			37028: out = 24'(-3356);
			37029: out = 24'(128);
			37030: out = 24'(3600);
			37031: out = 24'(4952);
			37032: out = 24'(1956);
			37033: out = 24'(2940);
			37034: out = 24'(-444);
			37035: out = 24'(-2228);
			37036: out = 24'(-3868);
			37037: out = 24'(-2892);
			37038: out = 24'(-3968);
			37039: out = 24'(116);
			37040: out = 24'(3740);
			37041: out = 24'(2576);
			37042: out = 24'(-3964);
			37043: out = 24'(-3856);
			37044: out = 24'(-520);
			37045: out = 24'(-1576);
			37046: out = 24'(-2784);
			37047: out = 24'(-1116);
			37048: out = 24'(2180);
			37049: out = 24'(2540);
			37050: out = 24'(3648);
			37051: out = 24'(2876);
			37052: out = 24'(1632);
			37053: out = 24'(-280);
			37054: out = 24'(2564);
			37055: out = 24'(-1680);
			37056: out = 24'(-4464);
			37057: out = 24'(-3508);
			37058: out = 24'(-300);
			37059: out = 24'(172);
			37060: out = 24'(-336);
			37061: out = 24'(680);
			37062: out = 24'(2388);
			37063: out = 24'(744);
			37064: out = 24'(-4076);
			37065: out = 24'(-6132);
			37066: out = 24'(-2376);
			37067: out = 24'(2056);
			37068: out = 24'(3172);
			37069: out = 24'(2516);
			37070: out = 24'(2560);
			37071: out = 24'(-188);
			37072: out = 24'(-856);
			37073: out = 24'(-1548);
			37074: out = 24'(-1116);
			37075: out = 24'(-1468);
			37076: out = 24'(2568);
			37077: out = 24'(3464);
			37078: out = 24'(1544);
			37079: out = 24'(-1492);
			37080: out = 24'(-1448);
			37081: out = 24'(-836);
			37082: out = 24'(728);
			37083: out = 24'(2560);
			37084: out = 24'(2608);
			37085: out = 24'(756);
			37086: out = 24'(-320);
			37087: out = 24'(408);
			37088: out = 24'(-4420);
			37089: out = 24'(-1696);
			37090: out = 24'(1324);
			37091: out = 24'(2164);
			37092: out = 24'(-216);
			37093: out = 24'(1700);
			37094: out = 24'(3220);
			37095: out = 24'(1968);
			37096: out = 24'(-3620);
			37097: out = 24'(-1044);
			37098: out = 24'(1732);
			37099: out = 24'(3108);
			37100: out = 24'(-324);
			37101: out = 24'(-2400);
			37102: out = 24'(-5896);
			37103: out = 24'(-1976);
			37104: out = 24'(5612);
			37105: out = 24'(5864);
			37106: out = 24'(-3132);
			37107: out = 24'(-9476);
			37108: out = 24'(-5444);
			37109: out = 24'(1832);
			37110: out = 24'(3848);
			37111: out = 24'(2688);
			37112: out = 24'(2220);
			37113: out = 24'(-808);
			37114: out = 24'(176);
			37115: out = 24'(-2924);
			37116: out = 24'(-4228);
			37117: out = 24'(-2192);
			37118: out = 24'(2116);
			37119: out = 24'(1060);
			37120: out = 24'(-620);
			37121: out = 24'(300);
			37122: out = 24'(5436);
			37123: out = 24'(1396);
			37124: out = 24'(-3756);
			37125: out = 24'(-3516);
			37126: out = 24'(2088);
			37127: out = 24'(2720);
			37128: out = 24'(1436);
			37129: out = 24'(-228);
			37130: out = 24'(-1484);
			37131: out = 24'(-1720);
			37132: out = 24'(-848);
			37133: out = 24'(-348);
			37134: out = 24'(-128);
			37135: out = 24'(212);
			37136: out = 24'(1004);
			37137: out = 24'(-1984);
			37138: out = 24'(-6564);
			37139: out = 24'(-2040);
			37140: out = 24'(1616);
			37141: out = 24'(2028);
			37142: out = 24'(812);
			37143: out = 24'(2376);
			37144: out = 24'(2804);
			37145: out = 24'(48);
			37146: out = 24'(-2472);
			37147: out = 24'(-616);
			37148: out = 24'(-984);
			37149: out = 24'(-3304);
			37150: out = 24'(-3560);
			37151: out = 24'(-148);
			37152: out = 24'(944);
			37153: out = 24'(-2684);
			37154: out = 24'(-2048);
			37155: out = 24'(6124);
			37156: out = 24'(6952);
			37157: out = 24'(3508);
			37158: out = 24'(-1704);
			37159: out = 24'(-3744);
			37160: out = 24'(-5588);
			37161: out = 24'(-4308);
			37162: out = 24'(248);
			37163: out = 24'(6176);
			37164: out = 24'(5212);
			37165: out = 24'(64);
			37166: out = 24'(-5356);
			37167: out = 24'(-3276);
			37168: out = 24'(3256);
			37169: out = 24'(3740);
			37170: out = 24'(392);
			37171: out = 24'(-1828);
			37172: out = 24'(-1472);
			37173: out = 24'(-184);
			37174: out = 24'(-1276);
			37175: out = 24'(-40);
			37176: out = 24'(3980);
			37177: out = 24'(5432);
			37178: out = 24'(4164);
			37179: out = 24'(1392);
			37180: out = 24'(-1456);
			37181: out = 24'(-4512);
			37182: out = 24'(-5892);
			37183: out = 24'(-3284);
			37184: out = 24'(744);
			37185: out = 24'(2204);
			37186: out = 24'(1008);
			37187: out = 24'(-48);
			37188: out = 24'(-876);
			37189: out = 24'(-2688);
			37190: out = 24'(-3364);
			37191: out = 24'(-1248);
			37192: out = 24'(2132);
			37193: out = 24'(2948);
			37194: out = 24'(1052);
			37195: out = 24'(-2240);
			37196: out = 24'(-4192);
			37197: out = 24'(-4084);
			37198: out = 24'(-1412);
			37199: out = 24'(-396);
			37200: out = 24'(80);
			37201: out = 24'(-724);
			37202: out = 24'(-3124);
			37203: out = 24'(-904);
			37204: out = 24'(1692);
			37205: out = 24'(2760);
			37206: out = 24'(2528);
			37207: out = 24'(92);
			37208: out = 24'(-128);
			37209: out = 24'(-1104);
			37210: out = 24'(-3644);
			37211: out = 24'(-4232);
			37212: out = 24'(-1376);
			37213: out = 24'(2384);
			37214: out = 24'(3132);
			37215: out = 24'(824);
			37216: out = 24'(-36);
			37217: out = 24'(-540);
			37218: out = 24'(-2216);
			37219: out = 24'(-5168);
			37220: out = 24'(-4084);
			37221: out = 24'(-52);
			37222: out = 24'(3040);
			37223: out = 24'(388);
			37224: out = 24'(412);
			37225: out = 24'(-2352);
			37226: out = 24'(-2160);
			37227: out = 24'(1292);
			37228: out = 24'(2552);
			37229: out = 24'(3340);
			37230: out = 24'(2888);
			37231: out = 24'(0);
			37232: out = 24'(-672);
			37233: out = 24'(-5504);
			37234: out = 24'(-4664);
			37235: out = 24'(-224);
			37236: out = 24'(2760);
			37237: out = 24'(396);
			37238: out = 24'(1180);
			37239: out = 24'(2464);
			37240: out = 24'(772);
			37241: out = 24'(-2080);
			37242: out = 24'(396);
			37243: out = 24'(2424);
			37244: out = 24'(-592);
			37245: out = 24'(-3000);
			37246: out = 24'(120);
			37247: out = 24'(3412);
			37248: out = 24'(1752);
			37249: out = 24'(-2840);
			37250: out = 24'(-1012);
			37251: out = 24'(964);
			37252: out = 24'(-616);
			37253: out = 24'(104);
			37254: out = 24'(-256);
			37255: out = 24'(-104);
			37256: out = 24'(284);
			37257: out = 24'(2596);
			37258: out = 24'(1256);
			37259: out = 24'(-2004);
			37260: out = 24'(-4864);
			37261: out = 24'(-2644);
			37262: out = 24'(-52);
			37263: out = 24'(3872);
			37264: out = 24'(4924);
			37265: out = 24'(2504);
			37266: out = 24'(-3640);
			37267: out = 24'(-4468);
			37268: out = 24'(-532);
			37269: out = 24'(4144);
			37270: out = 24'(4804);
			37271: out = 24'(1500);
			37272: out = 24'(-2712);
			37273: out = 24'(-4136);
			37274: out = 24'(-1456);
			37275: out = 24'(-308);
			37276: out = 24'(-196);
			37277: out = 24'(440);
			37278: out = 24'(2572);
			37279: out = 24'(132);
			37280: out = 24'(-1972);
			37281: out = 24'(-4380);
			37282: out = 24'(-5028);
			37283: out = 24'(-1932);
			37284: out = 24'(1852);
			37285: out = 24'(1928);
			37286: out = 24'(-572);
			37287: out = 24'(-2004);
			37288: out = 24'(-1696);
			37289: out = 24'(-196);
			37290: out = 24'(1480);
			37291: out = 24'(2532);
			37292: out = 24'(2912);
			37293: out = 24'(1180);
			37294: out = 24'(-712);
			37295: out = 24'(-2516);
			37296: out = 24'(-1248);
			37297: out = 24'(-3132);
			37298: out = 24'(-3264);
			37299: out = 24'(1388);
			37300: out = 24'(3100);
			37301: out = 24'(1800);
			37302: out = 24'(-2132);
			37303: out = 24'(-3932);
			37304: out = 24'(-1452);
			37305: out = 24'(1676);
			37306: out = 24'(3468);
			37307: out = 24'(2988);
			37308: out = 24'(-92);
			37309: out = 24'(-3228);
			37310: out = 24'(-4888);
			37311: out = 24'(-3060);
			37312: out = 24'(116);
			37313: out = 24'(2436);
			37314: out = 24'(2868);
			37315: out = 24'(2108);
			37316: out = 24'(-468);
			37317: out = 24'(128);
			37318: out = 24'(-3024);
			37319: out = 24'(-3688);
			37320: out = 24'(-140);
			37321: out = 24'(5708);
			37322: out = 24'(4072);
			37323: out = 24'(1368);
			37324: out = 24'(464);
			37325: out = 24'(-156);
			37326: out = 24'(-1060);
			37327: out = 24'(-956);
			37328: out = 24'(544);
			37329: out = 24'(2564);
			37330: out = 24'(1028);
			37331: out = 24'(160);
			37332: out = 24'(-688);
			37333: out = 24'(-1272);
			37334: out = 24'(-1756);
			37335: out = 24'(1264);
			37336: out = 24'(1632);
			37337: out = 24'(-1888);
			37338: out = 24'(-2220);
			37339: out = 24'(-1776);
			37340: out = 24'(-1328);
			37341: out = 24'(-360);
			37342: out = 24'(4936);
			37343: out = 24'(6136);
			37344: out = 24'(2212);
			37345: out = 24'(-3384);
			37346: out = 24'(-936);
			37347: out = 24'(-2824);
			37348: out = 24'(-624);
			37349: out = 24'(1240);
			37350: out = 24'(2540);
			37351: out = 24'(616);
			37352: out = 24'(368);
			37353: out = 24'(164);
			37354: out = 24'(-512);
			37355: out = 24'(-3296);
			37356: out = 24'(-2308);
			37357: out = 24'(-724);
			37358: out = 24'(-112);
			37359: out = 24'(-332);
			37360: out = 24'(488);
			37361: out = 24'(-340);
			37362: out = 24'(-1332);
			37363: out = 24'(-120);
			37364: out = 24'(452);
			37365: out = 24'(-320);
			37366: out = 24'(-1892);
			37367: out = 24'(-2312);
			37368: out = 24'(-4108);
			37369: out = 24'(-2856);
			37370: out = 24'(464);
			37371: out = 24'(2564);
			37372: out = 24'(1272);
			37373: out = 24'(-1396);
			37374: out = 24'(-1292);
			37375: out = 24'(776);
			37376: out = 24'(-3144);
			37377: out = 24'(-6132);
			37378: out = 24'(-6644);
			37379: out = 24'(-2512);
			37380: out = 24'(-192);
			37381: out = 24'(3724);
			37382: out = 24'(1944);
			37383: out = 24'(596);
			37384: out = 24'(2872);
			37385: out = 24'(868);
			37386: out = 24'(-2572);
			37387: out = 24'(-3260);
			37388: out = 24'(1040);
			37389: out = 24'(5528);
			37390: out = 24'(4700);
			37391: out = 24'(496);
			37392: out = 24'(-2048);
			37393: out = 24'(-164);
			37394: out = 24'(120);
			37395: out = 24'(132);
			37396: out = 24'(868);
			37397: out = 24'(-176);
			37398: out = 24'(160);
			37399: out = 24'(-692);
			37400: out = 24'(-1708);
			37401: out = 24'(-4292);
			37402: out = 24'(64);
			37403: out = 24'(752);
			37404: out = 24'(-568);
			37405: out = 24'(-1956);
			37406: out = 24'(3196);
			37407: out = 24'(3280);
			37408: out = 24'(2648);
			37409: out = 24'(2608);
			37410: out = 24'(2840);
			37411: out = 24'(-244);
			37412: out = 24'(-1316);
			37413: out = 24'(-92);
			37414: out = 24'(-96);
			37415: out = 24'(-3200);
			37416: out = 24'(-3000);
			37417: out = 24'(1388);
			37418: out = 24'(5088);
			37419: out = 24'(3256);
			37420: out = 24'(2344);
			37421: out = 24'(2060);
			37422: out = 24'(-1000);
			37423: out = 24'(-5368);
			37424: out = 24'(-6912);
			37425: out = 24'(-2128);
			37426: out = 24'(3836);
			37427: out = 24'(3592);
			37428: out = 24'(1004);
			37429: out = 24'(-512);
			37430: out = 24'(-160);
			37431: out = 24'(-1432);
			37432: out = 24'(-1332);
			37433: out = 24'(-1788);
			37434: out = 24'(-2040);
			37435: out = 24'(40);
			37436: out = 24'(-200);
			37437: out = 24'(156);
			37438: out = 24'(-564);
			37439: out = 24'(-992);
			37440: out = 24'(-492);
			37441: out = 24'(1932);
			37442: out = 24'(1676);
			37443: out = 24'(-1640);
			37444: out = 24'(-3124);
			37445: out = 24'(-804);
			37446: out = 24'(1312);
			37447: out = 24'(444);
			37448: out = 24'(-2064);
			37449: out = 24'(-676);
			37450: out = 24'(-96);
			37451: out = 24'(-1860);
			37452: out = 24'(-3968);
			37453: out = 24'(-372);
			37454: out = 24'(2548);
			37455: out = 24'(2160);
			37456: out = 24'(-60);
			37457: out = 24'(-1016);
			37458: out = 24'(-604);
			37459: out = 24'(512);
			37460: out = 24'(644);
			37461: out = 24'(-616);
			37462: out = 24'(-3444);
			37463: out = 24'(-3020);
			37464: out = 24'(400);
			37465: out = 24'(872);
			37466: out = 24'(556);
			37467: out = 24'(-56);
			37468: out = 24'(-200);
			37469: out = 24'(-2964);
			37470: out = 24'(-752);
			37471: out = 24'(2116);
			37472: out = 24'(3336);
			37473: out = 24'(-132);
			37474: out = 24'(840);
			37475: out = 24'(336);
			37476: out = 24'(212);
			37477: out = 24'(972);
			37478: out = 24'(156);
			37479: out = 24'(-112);
			37480: out = 24'(320);
			37481: out = 24'(936);
			37482: out = 24'(-12);
			37483: out = 24'(460);
			37484: out = 24'(620);
			37485: out = 24'(-584);
			37486: out = 24'(-2984);
			37487: out = 24'(-1212);
			37488: out = 24'(2136);
			37489: out = 24'(2756);
			37490: out = 24'(-2268);
			37491: out = 24'(-104);
			37492: out = 24'(2464);
			37493: out = 24'(2904);
			37494: out = 24'(-436);
			37495: out = 24'(40);
			37496: out = 24'(-1400);
			37497: out = 24'(-2940);
			37498: out = 24'(-2948);
			37499: out = 24'(-472);
			37500: out = 24'(2408);
			37501: out = 24'(3572);
			37502: out = 24'(1972);
			37503: out = 24'(116);
			37504: out = 24'(-528);
			37505: out = 24'(364);
			37506: out = 24'(-168);
			37507: out = 24'(-2164);
			37508: out = 24'(-1012);
			37509: out = 24'(1556);
			37510: out = 24'(2096);
			37511: out = 24'(448);
			37512: out = 24'(-3148);
			37513: out = 24'(-1308);
			37514: out = 24'(808);
			37515: out = 24'(-400);
			37516: out = 24'(-172);
			37517: out = 24'(1616);
			37518: out = 24'(1976);
			37519: out = 24'(-512);
			37520: out = 24'(2696);
			37521: out = 24'(480);
			37522: out = 24'(-980);
			37523: out = 24'(-976);
			37524: out = 24'(2480);
			37525: out = 24'(1020);
			37526: out = 24'(76);
			37527: out = 24'(-412);
			37528: out = 24'(-360);
			37529: out = 24'(-1408);
			37530: out = 24'(-952);
			37531: out = 24'(152);
			37532: out = 24'(396);
			37533: out = 24'(-1148);
			37534: out = 24'(-3588);
			37535: out = 24'(-4140);
			37536: out = 24'(-1796);
			37537: out = 24'(-536);
			37538: out = 24'(148);
			37539: out = 24'(-792);
			37540: out = 24'(-1068);
			37541: out = 24'(-268);
			37542: out = 24'(2176);
			37543: out = 24'(1464);
			37544: out = 24'(-716);
			37545: out = 24'(-1280);
			37546: out = 24'(288);
			37547: out = 24'(-1316);
			37548: out = 24'(-3736);
			37549: out = 24'(-1592);
			37550: out = 24'(-712);
			37551: out = 24'(1028);
			37552: out = 24'(-316);
			37553: out = 24'(-780);
			37554: out = 24'(-548);
			37555: out = 24'(4088);
			37556: out = 24'(3788);
			37557: out = 24'(-380);
			37558: out = 24'(-3216);
			37559: out = 24'(-1724);
			37560: out = 24'(-1864);
			37561: out = 24'(-2572);
			37562: out = 24'(128);
			37563: out = 24'(2088);
			37564: out = 24'(1572);
			37565: out = 24'(1112);
			37566: out = 24'(3052);
			37567: out = 24'(2552);
			37568: out = 24'(-1552);
			37569: out = 24'(-3500);
			37570: out = 24'(604);
			37571: out = 24'(156);
			37572: out = 24'(860);
			37573: out = 24'(8);
			37574: out = 24'(-216);
			37575: out = 24'(-2212);
			37576: out = 24'(-236);
			37577: out = 24'(1388);
			37578: out = 24'(2420);
			37579: out = 24'(1940);
			37580: out = 24'(420);
			37581: out = 24'(-1188);
			37582: out = 24'(-972);
			37583: out = 24'(-212);
			37584: out = 24'(2668);
			37585: out = 24'(1156);
			37586: out = 24'(-972);
			37587: out = 24'(-1184);
			37588: out = 24'(376);
			37589: out = 24'(-1008);
			37590: out = 24'(-3564);
			37591: out = 24'(-4528);
			37592: out = 24'(-1340);
			37593: out = 24'(1292);
			37594: out = 24'(3084);
			37595: out = 24'(1912);
			37596: out = 24'(-2008);
			37597: out = 24'(-5292);
			37598: out = 24'(-4100);
			37599: out = 24'(-896);
			37600: out = 24'(708);
			37601: out = 24'(2040);
			37602: out = 24'(3852);
			37603: out = 24'(3652);
			37604: out = 24'(88);
			37605: out = 24'(576);
			37606: out = 24'(16);
			37607: out = 24'(-1028);
			37608: out = 24'(-3316);
			37609: out = 24'(-2672);
			37610: out = 24'(-708);
			37611: out = 24'(3128);
			37612: out = 24'(5324);
			37613: out = 24'(5040);
			37614: out = 24'(960);
			37615: out = 24'(-1288);
			37616: out = 24'(-884);
			37617: out = 24'(456);
			37618: out = 24'(-1776);
			37619: out = 24'(-1468);
			37620: out = 24'(924);
			37621: out = 24'(2588);
			37622: out = 24'(124);
			37623: out = 24'(-1676);
			37624: out = 24'(-2360);
			37625: out = 24'(-1980);
			37626: out = 24'(-348);
			37627: out = 24'(280);
			37628: out = 24'(188);
			37629: out = 24'(-332);
			37630: out = 24'(-188);
			37631: out = 24'(380);
			37632: out = 24'(384);
			37633: out = 24'(-516);
			37634: out = 24'(-32);
			37635: out = 24'(208);
			37636: out = 24'(1668);
			37637: out = 24'(1736);
			37638: out = 24'(448);
			37639: out = 24'(-1260);
			37640: out = 24'(-208);
			37641: out = 24'(644);
			37642: out = 24'(196);
			37643: out = 24'(-3792);
			37644: out = 24'(-2300);
			37645: out = 24'(-1284);
			37646: out = 24'(-2128);
			37647: out = 24'(-312);
			37648: out = 24'(3640);
			37649: out = 24'(5476);
			37650: out = 24'(2868);
			37651: out = 24'(-1264);
			37652: out = 24'(-4440);
			37653: out = 24'(-5140);
			37654: out = 24'(-4036);
			37655: out = 24'(-720);
			37656: out = 24'(4084);
			37657: out = 24'(5788);
			37658: out = 24'(3184);
			37659: out = 24'(-1028);
			37660: out = 24'(-3776);
			37661: out = 24'(-3000);
			37662: out = 24'(-1664);
			37663: out = 24'(-1108);
			37664: out = 24'(-276);
			37665: out = 24'(2060);
			37666: out = 24'(3000);
			37667: out = 24'(1232);
			37668: out = 24'(-1152);
			37669: out = 24'(-820);
			37670: out = 24'(1156);
			37671: out = 24'(1524);
			37672: out = 24'(-1556);
			37673: out = 24'(1636);
			37674: out = 24'(548);
			37675: out = 24'(-3224);
			37676: out = 24'(-5416);
			37677: out = 24'(-308);
			37678: out = 24'(3480);
			37679: out = 24'(3348);
			37680: out = 24'(-192);
			37681: out = 24'(-1744);
			37682: out = 24'(-3816);
			37683: out = 24'(-2524);
			37684: out = 24'(488);
			37685: out = 24'(2012);
			37686: out = 24'(-200);
			37687: out = 24'(-2604);
			37688: out = 24'(-2620);
			37689: out = 24'(-1192);
			37690: out = 24'(1796);
			37691: out = 24'(1576);
			37692: out = 24'(-788);
			37693: out = 24'(-2828);
			37694: out = 24'(164);
			37695: out = 24'(3044);
			37696: out = 24'(4888);
			37697: out = 24'(3528);
			37698: out = 24'(924);
			37699: out = 24'(-3180);
			37700: out = 24'(-2868);
			37701: out = 24'(68);
			37702: out = 24'(-488);
			37703: out = 24'(-980);
			37704: out = 24'(-1524);
			37705: out = 24'(-1052);
			37706: out = 24'(-152);
			37707: out = 24'(1500);
			37708: out = 24'(2964);
			37709: out = 24'(1316);
			37710: out = 24'(-3192);
			37711: out = 24'(-1072);
			37712: out = 24'(3076);
			37713: out = 24'(4664);
			37714: out = 24'(1232);
			37715: out = 24'(652);
			37716: out = 24'(-1792);
			37717: out = 24'(-2472);
			37718: out = 24'(-2104);
			37719: out = 24'(-420);
			37720: out = 24'(-396);
			37721: out = 24'(-336);
			37722: out = 24'(-520);
			37723: out = 24'(-1356);
			37724: out = 24'(-656);
			37725: out = 24'(864);
			37726: out = 24'(2352);
			37727: out = 24'(1716);
			37728: out = 24'(2268);
			37729: out = 24'(-172);
			37730: out = 24'(-1880);
			37731: out = 24'(-1184);
			37732: out = 24'(1716);
			37733: out = 24'(508);
			37734: out = 24'(-820);
			37735: out = 24'(-60);
			37736: out = 24'(1728);
			37737: out = 24'(392);
			37738: out = 24'(-1580);
			37739: out = 24'(-2064);
			37740: out = 24'(200);
			37741: out = 24'(1496);
			37742: out = 24'(2228);
			37743: out = 24'(1132);
			37744: out = 24'(-424);
			37745: out = 24'(-1640);
			37746: out = 24'(-360);
			37747: out = 24'(-132);
			37748: out = 24'(-1504);
			37749: out = 24'(-768);
			37750: out = 24'(1348);
			37751: out = 24'(592);
			37752: out = 24'(-3144);
			37753: out = 24'(-5756);
			37754: out = 24'(-2384);
			37755: out = 24'(1264);
			37756: out = 24'(2048);
			37757: out = 24'(2004);
			37758: out = 24'(2696);
			37759: out = 24'(952);
			37760: out = 24'(-2628);
			37761: out = 24'(-3752);
			37762: out = 24'(-692);
			37763: out = 24'(2248);
			37764: out = 24'(1960);
			37765: out = 24'(-720);
			37766: out = 24'(-2092);
			37767: out = 24'(-1988);
			37768: out = 24'(-840);
			37769: out = 24'(-340);
			37770: out = 24'(2092);
			37771: out = 24'(260);
			37772: out = 24'(-508);
			37773: out = 24'(-624);
			37774: out = 24'(-1288);
			37775: out = 24'(-4400);
			37776: out = 24'(-2820);
			37777: out = 24'(1204);
			37778: out = 24'(232);
			37779: out = 24'(768);
			37780: out = 24'(-60);
			37781: out = 24'(-96);
			37782: out = 24'(260);
			37783: out = 24'(-2744);
			37784: out = 24'(-1624);
			37785: out = 24'(456);
			37786: out = 24'(328);
			37787: out = 24'(-28);
			37788: out = 24'(-400);
			37789: out = 24'(-136);
			37790: out = 24'(-264);
			37791: out = 24'(500);
			37792: out = 24'(452);
			37793: out = 24'(324);
			37794: out = 24'(-768);
			37795: out = 24'(-1920);
			37796: out = 24'(-928);
			37797: out = 24'(1768);
			37798: out = 24'(2388);
			37799: out = 24'(-848);
			37800: out = 24'(-3352);
			37801: out = 24'(-2860);
			37802: out = 24'(376);
			37803: out = 24'(2308);
			37804: out = 24'(4456);
			37805: out = 24'(1840);
			37806: out = 24'(-140);
			37807: out = 24'(-24);
			37808: out = 24'(1952);
			37809: out = 24'(1016);
			37810: out = 24'(-764);
			37811: out = 24'(-3036);
			37812: out = 24'(-4716);
			37813: out = 24'(-2540);
			37814: out = 24'(2108);
			37815: out = 24'(4220);
			37816: out = 24'(1636);
			37817: out = 24'(-2976);
			37818: out = 24'(-3632);
			37819: out = 24'(-476);
			37820: out = 24'(2292);
			37821: out = 24'(4200);
			37822: out = 24'(3036);
			37823: out = 24'(1024);
			37824: out = 24'(208);
			37825: out = 24'(-548);
			37826: out = 24'(276);
			37827: out = 24'(-772);
			37828: out = 24'(-2436);
			37829: out = 24'(-1444);
			37830: out = 24'(-504);
			37831: out = 24'(-928);
			37832: out = 24'(-780);
			37833: out = 24'(2180);
			37834: out = 24'(2072);
			37835: out = 24'(176);
			37836: out = 24'(-2160);
			37837: out = 24'(-2020);
			37838: out = 24'(-728);
			37839: out = 24'(-124);
			37840: out = 24'(-404);
			37841: out = 24'(712);
			37842: out = 24'(1688);
			37843: out = 24'(1228);
			37844: out = 24'(-2240);
			37845: out = 24'(-4776);
			37846: out = 24'(-1464);
			37847: out = 24'(-460);
			37848: out = 24'(-1028);
			37849: out = 24'(-2600);
			37850: out = 24'(-2796);
			37851: out = 24'(-900);
			37852: out = 24'(1756);
			37853: out = 24'(3004);
			37854: out = 24'(1804);
			37855: out = 24'(200);
			37856: out = 24'(-1752);
			37857: out = 24'(-1528);
			37858: out = 24'(600);
			37859: out = 24'(216);
			37860: out = 24'(-708);
			37861: out = 24'(-1592);
			37862: out = 24'(-828);
			37863: out = 24'(204);
			37864: out = 24'(1996);
			37865: out = 24'(1116);
			37866: out = 24'(-524);
			37867: out = 24'(-68);
			37868: out = 24'(1504);
			37869: out = 24'(2556);
			37870: out = 24'(460);
			37871: out = 24'(-4140);
			37872: out = 24'(-3232);
			37873: out = 24'(-1380);
			37874: out = 24'(344);
			37875: out = 24'(384);
			37876: out = 24'(12);
			37877: out = 24'(-20);
			37878: out = 24'(580);
			37879: out = 24'(152);
			37880: out = 24'(648);
			37881: out = 24'(-476);
			37882: out = 24'(1292);
			37883: out = 24'(2552);
			37884: out = 24'(364);
			37885: out = 24'(-2764);
			37886: out = 24'(-1356);
			37887: out = 24'(360);
			37888: out = 24'(-2416);
			37889: out = 24'(-2308);
			37890: out = 24'(616);
			37891: out = 24'(3620);
			37892: out = 24'(2216);
			37893: out = 24'(236);
			37894: out = 24'(-1792);
			37895: out = 24'(-2564);
			37896: out = 24'(-2848);
			37897: out = 24'(460);
			37898: out = 24'(2216);
			37899: out = 24'(2892);
			37900: out = 24'(1268);
			37901: out = 24'(-1096);
			37902: out = 24'(-3044);
			37903: out = 24'(-1828);
			37904: out = 24'(476);
			37905: out = 24'(2012);
			37906: out = 24'(-560);
			37907: out = 24'(-3040);
			37908: out = 24'(-3712);
			37909: out = 24'(-1720);
			37910: out = 24'(-596);
			37911: out = 24'(272);
			37912: out = 24'(-1332);
			37913: out = 24'(-2504);
			37914: out = 24'(-612);
			37915: out = 24'(3948);
			37916: out = 24'(3500);
			37917: out = 24'(-1412);
			37918: out = 24'(-2580);
			37919: out = 24'(-672);
			37920: out = 24'(1972);
			37921: out = 24'(1660);
			37922: out = 24'(-120);
			37923: out = 24'(-476);
			37924: out = 24'(-788);
			37925: out = 24'(-1020);
			37926: out = 24'(1040);
			37927: out = 24'(1700);
			37928: out = 24'(2608);
			37929: out = 24'(840);
			37930: out = 24'(-1624);
			37931: out = 24'(-4796);
			37932: out = 24'(-440);
			37933: out = 24'(4116);
			37934: out = 24'(4304);
			37935: out = 24'(-112);
			37936: out = 24'(-1772);
			37937: out = 24'(-3036);
			37938: out = 24'(-4448);
			37939: out = 24'(-5620);
			37940: out = 24'(-1432);
			37941: out = 24'(1652);
			37942: out = 24'(1788);
			37943: out = 24'(-120);
			37944: out = 24'(1932);
			37945: out = 24'(1116);
			37946: out = 24'(-1364);
			37947: out = 24'(-2752);
			37948: out = 24'(-520);
			37949: out = 24'(1424);
			37950: out = 24'(2724);
			37951: out = 24'(2604);
			37952: out = 24'(652);
			37953: out = 24'(-892);
			37954: out = 24'(-1536);
			37955: out = 24'(-1268);
			37956: out = 24'(-1388);
			37957: out = 24'(116);
			37958: out = 24'(428);
			37959: out = 24'(-1040);
			37960: out = 24'(-2960);
			37961: out = 24'(-1804);
			37962: out = 24'(992);
			37963: out = 24'(2080);
			37964: out = 24'(464);
			37965: out = 24'(2872);
			37966: out = 24'(1064);
			37967: out = 24'(-1620);
			37968: out = 24'(-2876);
			37969: out = 24'(-1500);
			37970: out = 24'(224);
			37971: out = 24'(32);
			37972: out = 24'(-1864);
			37973: out = 24'(-3724);
			37974: out = 24'(-2596);
			37975: out = 24'(-1020);
			37976: out = 24'(964);
			37977: out = 24'(4652);
			37978: out = 24'(2668);
			37979: out = 24'(740);
			37980: out = 24'(-284);
			37981: out = 24'(724);
			37982: out = 24'(-340);
			37983: out = 24'(-1148);
			37984: out = 24'(-3168);
			37985: out = 24'(-3372);
			37986: out = 24'(-600);
			37987: out = 24'(1912);
			37988: out = 24'(1292);
			37989: out = 24'(-424);
			37990: out = 24'(656);
			37991: out = 24'(2504);
			37992: out = 24'(1668);
			37993: out = 24'(-576);
			37994: out = 24'(800);
			37995: out = 24'(-272);
			37996: out = 24'(-784);
			37997: out = 24'(-1072);
			37998: out = 24'(988);
			37999: out = 24'(1688);
			38000: out = 24'(1316);
			38001: out = 24'(-3436);
			38002: out = 24'(-8660);
			38003: out = 24'(-4172);
			38004: out = 24'(-716);
			38005: out = 24'(1628);
			38006: out = 24'(2172);
			38007: out = 24'(-48);
			38008: out = 24'(1748);
			38009: out = 24'(2448);
			38010: out = 24'(2216);
			38011: out = 24'(2136);
			38012: out = 24'(1012);
			38013: out = 24'(-952);
			38014: out = 24'(-2424);
			38015: out = 24'(-2004);
			38016: out = 24'(-416);
			38017: out = 24'(-136);
			38018: out = 24'(-192);
			38019: out = 24'(-224);
			38020: out = 24'(8);
			38021: out = 24'(-2756);
			38022: out = 24'(-3552);
			38023: out = 24'(-1388);
			38024: out = 24'(-240);
			38025: out = 24'(40);
			38026: out = 24'(880);
			38027: out = 24'(2780);
			38028: out = 24'(1908);
			38029: out = 24'(-584);
			38030: out = 24'(-5328);
			38031: out = 24'(-7260);
			38032: out = 24'(-3832);
			38033: out = 24'(3216);
			38034: out = 24'(6136);
			38035: out = 24'(3412);
			38036: out = 24'(-312);
			38037: out = 24'(-3588);
			38038: out = 24'(-2000);
			38039: out = 24'(-912);
			38040: out = 24'(-848);
			38041: out = 24'(-68);
			38042: out = 24'(3488);
			38043: out = 24'(4184);
			38044: out = 24'(1144);
			38045: out = 24'(-1780);
			38046: out = 24'(-1512);
			38047: out = 24'(-864);
			38048: out = 24'(-1060);
			38049: out = 24'(284);
			38050: out = 24'(-196);
			38051: out = 24'(280);
			38052: out = 24'(-404);
			38053: out = 24'(-788);
			38054: out = 24'(-384);
			38055: out = 24'(3580);
			38056: out = 24'(4928);
			38057: out = 24'(1252);
			38058: out = 24'(-1412);
			38059: out = 24'(-3840);
			38060: out = 24'(-2168);
			38061: out = 24'(304);
			38062: out = 24'(688);
			38063: out = 24'(-1860);
			38064: out = 24'(-3128);
			38065: out = 24'(-2396);
			38066: out = 24'(-1968);
			38067: out = 24'(-3092);
			38068: out = 24'(-2088);
			38069: out = 24'(2820);
			38070: out = 24'(7260);
			38071: out = 24'(5316);
			38072: out = 24'(872);
			38073: out = 24'(-2096);
			38074: out = 24'(-2660);
			38075: out = 24'(-108);
			38076: out = 24'(1392);
			38077: out = 24'(3992);
			38078: out = 24'(4292);
			38079: out = 24'(172);
			38080: out = 24'(-4732);
			38081: out = 24'(-4064);
			38082: out = 24'(-232);
			38083: out = 24'(600);
			38084: out = 24'(-708);
			38085: out = 24'(-304);
			38086: out = 24'(972);
			38087: out = 24'(412);
			38088: out = 24'(-972);
			38089: out = 24'(884);
			38090: out = 24'(2660);
			38091: out = 24'(1916);
			38092: out = 24'(712);
			38093: out = 24'(336);
			38094: out = 24'(-48);
			38095: out = 24'(-2024);
			38096: out = 24'(-6432);
			38097: out = 24'(-2800);
			38098: out = 24'(8);
			38099: out = 24'(-292);
			38100: out = 24'(-904);
			38101: out = 24'(224);
			38102: out = 24'(4);
			38103: out = 24'(-1112);
			38104: out = 24'(552);
			38105: out = 24'(4240);
			38106: out = 24'(5992);
			38107: out = 24'(3312);
			38108: out = 24'(-616);
			38109: out = 24'(-3540);
			38110: out = 24'(-4552);
			38111: out = 24'(-4320);
			38112: out = 24'(-1760);
			38113: out = 24'(2600);
			38114: out = 24'(3276);
			38115: out = 24'(-512);
			38116: out = 24'(-3888);
			38117: out = 24'(-1780);
			38118: out = 24'(2016);
			38119: out = 24'(3248);
			38120: out = 24'(1460);
			38121: out = 24'(-16);
			38122: out = 24'(476);
			38123: out = 24'(-76);
			38124: out = 24'(-2032);
			38125: out = 24'(-2528);
			38126: out = 24'(-4);
			38127: out = 24'(2444);
			38128: out = 24'(2952);
			38129: out = 24'(1668);
			38130: out = 24'(-2572);
			38131: out = 24'(-3740);
			38132: out = 24'(-3248);
			38133: out = 24'(-1104);
			38134: out = 24'(2248);
			38135: out = 24'(4700);
			38136: out = 24'(4484);
			38137: out = 24'(1676);
			38138: out = 24'(-1180);
			38139: out = 24'(-2248);
			38140: out = 24'(-1056);
			38141: out = 24'(-116);
			38142: out = 24'(-196);
			38143: out = 24'(-268);
			38144: out = 24'(-144);
			38145: out = 24'(-624);
			38146: out = 24'(-1248);
			38147: out = 24'(-2168);
			38148: out = 24'(-628);
			38149: out = 24'(-464);
			38150: out = 24'(-1040);
			38151: out = 24'(-136);
			38152: out = 24'(3948);
			38153: out = 24'(4392);
			38154: out = 24'(952);
			38155: out = 24'(-1044);
			38156: out = 24'(-704);
			38157: out = 24'(-768);
			38158: out = 24'(-3732);
			38159: out = 24'(-6352);
			38160: out = 24'(-4536);
			38161: out = 24'(212);
			38162: out = 24'(2896);
			38163: out = 24'(2248);
			38164: out = 24'(3088);
			38165: out = 24'(2560);
			38166: out = 24'(1292);
			38167: out = 24'(-528);
			38168: out = 24'(-1116);
			38169: out = 24'(-1436);
			38170: out = 24'(-688);
			38171: out = 24'(312);
			38172: out = 24'(2192);
			38173: out = 24'(288);
			38174: out = 24'(-432);
			38175: out = 24'(-304);
			38176: out = 24'(-228);
			38177: out = 24'(388);
			38178: out = 24'(-1384);
			38179: out = 24'(-3768);
			38180: out = 24'(-3320);
			38181: out = 24'(-764);
			38182: out = 24'(1896);
			38183: out = 24'(1688);
			38184: out = 24'(664);
			38185: out = 24'(460);
			38186: out = 24'(984);
			38187: out = 24'(-1536);
			38188: out = 24'(-3400);
			38189: out = 24'(568);
			38190: out = 24'(3724);
			38191: out = 24'(2656);
			38192: out = 24'(-1776);
			38193: out = 24'(-3528);
			38194: out = 24'(-3448);
			38195: out = 24'(-2580);
			38196: out = 24'(-2960);
			38197: out = 24'(-1376);
			38198: out = 24'(-648);
			38199: out = 24'(3324);
			38200: out = 24'(4160);
			38201: out = 24'(1812);
			38202: out = 24'(-56);
			38203: out = 24'(-236);
			38204: out = 24'(-780);
			38205: out = 24'(-944);
			38206: out = 24'(464);
			38207: out = 24'(236);
			38208: out = 24'(-1164);
			38209: out = 24'(-2068);
			38210: out = 24'(-2024);
			38211: out = 24'(-356);
			38212: out = 24'(-284);
			38213: out = 24'(1412);
			38214: out = 24'(4228);
			38215: out = 24'(816);
			38216: out = 24'(-4064);
			38217: out = 24'(-4096);
			38218: out = 24'(1864);
			38219: out = 24'(4036);
			38220: out = 24'(1800);
			38221: out = 24'(-1856);
			38222: out = 24'(-2936);
			38223: out = 24'(-3960);
			38224: out = 24'(-3724);
			38225: out = 24'(-2212);
			38226: out = 24'(1316);
			38227: out = 24'(2936);
			38228: out = 24'(4712);
			38229: out = 24'(2188);
			38230: out = 24'(-1476);
			38231: out = 24'(-4124);
			38232: out = 24'(-3384);
			38233: out = 24'(-2288);
			38234: out = 24'(-688);
			38235: out = 24'(1196);
			38236: out = 24'(4268);
			38237: out = 24'(1888);
			38238: out = 24'(-2200);
			38239: out = 24'(-3480);
			38240: out = 24'(-116);
			38241: out = 24'(1696);
			38242: out = 24'(1380);
			38243: out = 24'(-864);
			38244: out = 24'(-2956);
			38245: out = 24'(-736);
			38246: out = 24'(1416);
			38247: out = 24'(1824);
			38248: out = 24'(604);
			38249: out = 24'(0);
			38250: out = 24'(1008);
			38251: out = 24'(2324);
			38252: out = 24'(1492);
			38253: out = 24'(-548);
			38254: out = 24'(-2328);
			38255: out = 24'(-1940);
			38256: out = 24'(-584);
			38257: out = 24'(1980);
			38258: out = 24'(504);
			38259: out = 24'(-608);
			38260: out = 24'(-840);
			38261: out = 24'(860);
			38262: out = 24'(1296);
			38263: out = 24'(4388);
			38264: out = 24'(5428);
			38265: out = 24'(1952);
			38266: out = 24'(-3252);
			38267: out = 24'(-3792);
			38268: out = 24'(-1876);
			38269: out = 24'(-1092);
			38270: out = 24'(-264);
			38271: out = 24'(1204);
			38272: out = 24'(1112);
			38273: out = 24'(-1656);
			38274: out = 24'(-2264);
			38275: out = 24'(-1128);
			38276: out = 24'(1064);
			38277: out = 24'(1884);
			38278: out = 24'(1880);
			38279: out = 24'(256);
			38280: out = 24'(-1704);
			38281: out = 24'(-4012);
			38282: out = 24'(-4516);
			38283: out = 24'(-1196);
			38284: out = 24'(2636);
			38285: out = 24'(3668);
			38286: out = 24'(2132);
			38287: out = 24'(-1968);
			38288: out = 24'(-3220);
			38289: out = 24'(-3268);
			38290: out = 24'(-3108);
			38291: out = 24'(-3204);
			38292: out = 24'(432);
			38293: out = 24'(2920);
			38294: out = 24'(1972);
			38295: out = 24'(-628);
			38296: out = 24'(-1204);
			38297: out = 24'(-244);
			38298: out = 24'(-16);
			38299: out = 24'(0);
			38300: out = 24'(-120);
			38301: out = 24'(144);
			38302: out = 24'(-176);
			38303: out = 24'(220);
			38304: out = 24'(-376);
			38305: out = 24'(1500);
			38306: out = 24'(964);
			38307: out = 24'(-1960);
			38308: out = 24'(-1652);
			38309: out = 24'(-560);
			38310: out = 24'(120);
			38311: out = 24'(24);
			38312: out = 24'(484);
			38313: out = 24'(3500);
			38314: out = 24'(3852);
			38315: out = 24'(32);
			38316: out = 24'(-5344);
			38317: out = 24'(-2228);
			38318: out = 24'(508);
			38319: out = 24'(-88);
			38320: out = 24'(-484);
			38321: out = 24'(1296);
			38322: out = 24'(3952);
			38323: out = 24'(3092);
			38324: out = 24'(-540);
			38325: out = 24'(-1584);
			38326: out = 24'(472);
			38327: out = 24'(2380);
			38328: out = 24'(1272);
			38329: out = 24'(176);
			38330: out = 24'(-184);
			38331: out = 24'(2444);
			38332: out = 24'(3756);
			38333: out = 24'(140);
			38334: out = 24'(-996);
			38335: out = 24'(-784);
			38336: out = 24'(-648);
			38337: out = 24'(-2900);
			38338: out = 24'(-3140);
			38339: out = 24'(-2320);
			38340: out = 24'(144);
			38341: out = 24'(1932);
			38342: out = 24'(3676);
			38343: out = 24'(1704);
			38344: out = 24'(-680);
			38345: out = 24'(-1568);
			38346: out = 24'(1572);
			38347: out = 24'(396);
			38348: out = 24'(-876);
			38349: out = 24'(-1036);
			38350: out = 24'(-424);
			38351: out = 24'(-448);
			38352: out = 24'(772);
			38353: out = 24'(1548);
			38354: out = 24'(-536);
			38355: out = 24'(-2156);
			38356: out = 24'(-2516);
			38357: out = 24'(-1356);
			38358: out = 24'(-1184);
			38359: out = 24'(308);
			38360: out = 24'(-24);
			38361: out = 24'(-176);
			38362: out = 24'(-120);
			38363: out = 24'(1836);
			38364: out = 24'(1720);
			38365: out = 24'(1488);
			38366: out = 24'(-592);
			38367: out = 24'(-3640);
			38368: out = 24'(-6544);
			38369: out = 24'(-2388);
			38370: out = 24'(3784);
			38371: out = 24'(3868);
			38372: out = 24'(348);
			38373: out = 24'(-1720);
			38374: out = 24'(-416);
			38375: out = 24'(-452);
			38376: out = 24'(52);
			38377: out = 24'(-820);
			38378: out = 24'(-1004);
			38379: out = 24'(-1020);
			38380: out = 24'(568);
			38381: out = 24'(40);
			38382: out = 24'(0);
			38383: out = 24'(708);
			38384: out = 24'(1792);
			38385: out = 24'(-76);
			38386: out = 24'(-2028);
			38387: out = 24'(-1880);
			38388: out = 24'(1860);
			38389: out = 24'(900);
			38390: out = 24'(-4);
			38391: out = 24'(200);
			38392: out = 24'(1904);
			38393: out = 24'(4);
			38394: out = 24'(-300);
			38395: out = 24'(-472);
			38396: out = 24'(-1060);
			38397: out = 24'(-492);
			38398: out = 24'(320);
			38399: out = 24'(228);
			38400: out = 24'(-396);
			38401: out = 24'(-980);
			38402: out = 24'(-532);
			38403: out = 24'(112);
			38404: out = 24'(288);
			38405: out = 24'(-416);
			38406: out = 24'(-132);
			38407: out = 24'(-784);
			38408: out = 24'(-888);
			38409: out = 24'(-324);
			38410: out = 24'(2080);
			38411: out = 24'(2000);
			38412: out = 24'(2348);
			38413: out = 24'(3864);
			38414: out = 24'(364);
			38415: out = 24'(-4644);
			38416: out = 24'(-5672);
			38417: out = 24'(-168);
			38418: out = 24'(1724);
			38419: out = 24'(2468);
			38420: out = 24'(228);
			38421: out = 24'(-1364);
			38422: out = 24'(-2104);
			38423: out = 24'(-1300);
			38424: out = 24'(-1320);
			38425: out = 24'(-828);
			38426: out = 24'(-256);
			38427: out = 24'(1972);
			38428: out = 24'(1592);
			38429: out = 24'(-1336);
			38430: out = 24'(-4964);
			38431: out = 24'(-1012);
			38432: out = 24'(0);
			38433: out = 24'(-280);
			38434: out = 24'(-32);
			38435: out = 24'(1652);
			38436: out = 24'(980);
			38437: out = 24'(-664);
			38438: out = 24'(-2040);
			38439: out = 24'(-1712);
			38440: out = 24'(-584);
			38441: out = 24'(2492);
			38442: out = 24'(3892);
			38443: out = 24'(228);
			38444: out = 24'(-1472);
			38445: out = 24'(-2036);
			38446: out = 24'(-2048);
			38447: out = 24'(-2460);
			38448: out = 24'(-676);
			38449: out = 24'(2384);
			38450: out = 24'(3112);
			38451: out = 24'(-440);
			38452: out = 24'(-2796);
			38453: out = 24'(-1840);
			38454: out = 24'(1252);
			38455: out = 24'(1144);
			38456: out = 24'(-544);
			38457: out = 24'(-3288);
			38458: out = 24'(-988);
			38459: out = 24'(2264);
			38460: out = 24'(1748);
			38461: out = 24'(-444);
			38462: out = 24'(-620);
			38463: out = 24'(1084);
			38464: out = 24'(1616);
			38465: out = 24'(-632);
			38466: out = 24'(-2128);
			38467: out = 24'(-2920);
			38468: out = 24'(-3056);
			38469: out = 24'(-532);
			38470: out = 24'(1820);
			38471: out = 24'(1868);
			38472: out = 24'(-572);
			38473: out = 24'(0);
			38474: out = 24'(-1368);
			38475: out = 24'(-2268);
			38476: out = 24'(-2072);
			38477: out = 24'(-100);
			38478: out = 24'(1524);
			38479: out = 24'(1136);
			38480: out = 24'(-512);
			38481: out = 24'(100);
			38482: out = 24'(172);
			38483: out = 24'(492);
			38484: out = 24'(-1128);
			38485: out = 24'(-2352);
			38486: out = 24'(-3536);
			38487: out = 24'(172);
			38488: out = 24'(2452);
			38489: out = 24'(1700);
			38490: out = 24'(492);
			38491: out = 24'(608);
			38492: out = 24'(-844);
			38493: out = 24'(-4008);
			38494: out = 24'(-5304);
			38495: out = 24'(-2272);
			38496: out = 24'(1140);
			38497: out = 24'(2060);
			38498: out = 24'(2164);
			38499: out = 24'(2440);
			38500: out = 24'(2856);
			38501: out = 24'(1616);
			38502: out = 24'(-1392);
			38503: out = 24'(-3588);
			38504: out = 24'(-2036);
			38505: out = 24'(2132);
			38506: out = 24'(4088);
			38507: out = 24'(1100);
			38508: out = 24'(-2400);
			38509: out = 24'(-2204);
			38510: out = 24'(416);
			38511: out = 24'(492);
			38512: out = 24'(164);
			38513: out = 24'(-136);
			38514: out = 24'(-244);
			38515: out = 24'(-1700);
			38516: out = 24'(-408);
			38517: out = 24'(1196);
			38518: out = 24'(1784);
			38519: out = 24'(296);
			38520: out = 24'(92);
			38521: out = 24'(-624);
			38522: out = 24'(-1952);
			38523: out = 24'(-3936);
			38524: out = 24'(-1028);
			38525: out = 24'(968);
			38526: out = 24'(3064);
			38527: out = 24'(3544);
			38528: out = 24'(2072);
			38529: out = 24'(308);
			38530: out = 24'(-876);
			38531: out = 24'(-2404);
			38532: out = 24'(-3848);
			38533: out = 24'(-2516);
			38534: out = 24'(608);
			38535: out = 24'(1684);
			38536: out = 24'(-172);
			38537: out = 24'(-1504);
			38538: out = 24'(-444);
			38539: out = 24'(352);
			38540: out = 24'(-1068);
			38541: out = 24'(40);
			38542: out = 24'(324);
			38543: out = 24'(96);
			38544: out = 24'(-1092);
			38545: out = 24'(-744);
			38546: out = 24'(-376);
			38547: out = 24'(304);
			38548: out = 24'(892);
			38549: out = 24'(2628);
			38550: out = 24'(600);
			38551: out = 24'(-1600);
			38552: out = 24'(-3684);
			38553: out = 24'(-3568);
			38554: out = 24'(-804);
			38555: out = 24'(1620);
			38556: out = 24'(1636);
			38557: out = 24'(-196);
			38558: out = 24'(-2072);
			38559: out = 24'(-1544);
			38560: out = 24'(-20);
			38561: out = 24'(900);
			38562: out = 24'(1988);
			38563: out = 24'(2560);
			38564: out = 24'(1996);
			38565: out = 24'(264);
			38566: out = 24'(692);
			38567: out = 24'(-1960);
			38568: out = 24'(-1524);
			38569: out = 24'(1096);
			38570: out = 24'(4408);
			38571: out = 24'(2948);
			38572: out = 24'(1044);
			38573: out = 24'(-908);
			38574: out = 24'(-1812);
			38575: out = 24'(-4748);
			38576: out = 24'(-1756);
			38577: out = 24'(1864);
			38578: out = 24'(2352);
			38579: out = 24'(2664);
			38580: out = 24'(664);
			38581: out = 24'(-1052);
			38582: out = 24'(-1676);
			38583: out = 24'(-256);
			38584: out = 24'(1796);
			38585: out = 24'(1920);
			38586: out = 24'(-704);
			38587: out = 24'(-2288);
			38588: out = 24'(-1728);
			38589: out = 24'(1008);
			38590: out = 24'(2612);
			38591: out = 24'(2300);
			38592: out = 24'(36);
			38593: out = 24'(-452);
			38594: out = 24'(-160);
			38595: out = 24'(236);
			38596: out = 24'(-3244);
			38597: out = 24'(-1512);
			38598: out = 24'(852);
			38599: out = 24'(1656);
			38600: out = 24'(340);
			38601: out = 24'(572);
			38602: out = 24'(-848);
			38603: out = 24'(-3192);
			38604: out = 24'(-4056);
			38605: out = 24'(-2308);
			38606: out = 24'(-888);
			38607: out = 24'(516);
			38608: out = 24'(1588);
			38609: out = 24'(-1360);
			38610: out = 24'(-5808);
			38611: out = 24'(-5508);
			38612: out = 24'(808);
			38613: out = 24'(4032);
			38614: out = 24'(2100);
			38615: out = 24'(-1304);
			38616: out = 24'(-1160);
			38617: out = 24'(100);
			38618: out = 24'(428);
			38619: out = 24'(-380);
			38620: out = 24'(352);
			38621: out = 24'(184);
			38622: out = 24'(768);
			38623: out = 24'(-792);
			38624: out = 24'(-1592);
			38625: out = 24'(-860);
			38626: out = 24'(1600);
			38627: out = 24'(1376);
			38628: out = 24'(384);
			38629: out = 24'(604);
			38630: out = 24'(-848);
			38631: out = 24'(-1124);
			38632: out = 24'(-672);
			38633: out = 24'(32);
			38634: out = 24'(564);
			38635: out = 24'(108);
			38636: out = 24'(-208);
			38637: out = 24'(-76);
			38638: out = 24'(-60);
			38639: out = 24'(316);
			38640: out = 24'(1256);
			38641: out = 24'(1756);
			38642: out = 24'(476);
			38643: out = 24'(472);
			38644: out = 24'(1248);
			38645: out = 24'(1504);
			38646: out = 24'(-500);
			38647: out = 24'(-828);
			38648: out = 24'(-800);
			38649: out = 24'(884);
			38650: out = 24'(2192);
			38651: out = 24'(104);
			38652: out = 24'(-2512);
			38653: out = 24'(-2800);
			38654: out = 24'(-284);
			38655: out = 24'(2264);
			38656: out = 24'(2720);
			38657: out = 24'(1180);
			38658: out = 24'(-908);
			38659: out = 24'(-1768);
			38660: out = 24'(-2720);
			38661: out = 24'(-428);
			38662: out = 24'(2856);
			38663: out = 24'(3188);
			38664: out = 24'(1128);
			38665: out = 24'(-2164);
			38666: out = 24'(-3680);
			38667: out = 24'(-3088);
			38668: out = 24'(-500);
			38669: out = 24'(-144);
			38670: out = 24'(-368);
			38671: out = 24'(224);
			38672: out = 24'(2316);
			38673: out = 24'(700);
			38674: out = 24'(-1572);
			38675: out = 24'(-2176);
			38676: out = 24'(560);
			38677: out = 24'(1480);
			38678: out = 24'(1392);
			38679: out = 24'(-300);
			38680: out = 24'(-992);
			38681: out = 24'(-3384);
			38682: out = 24'(-1628);
			38683: out = 24'(0);
			38684: out = 24'(420);
			38685: out = 24'(-332);
			38686: out = 24'(1416);
			38687: out = 24'(-16);
			38688: out = 24'(-4632);
			38689: out = 24'(-3088);
			38690: out = 24'(316);
			38691: out = 24'(2116);
			38692: out = 24'(-648);
			38693: out = 24'(-1956);
			38694: out = 24'(-2412);
			38695: out = 24'(520);
			38696: out = 24'(2068);
			38697: out = 24'(1976);
			38698: out = 24'(-1284);
			38699: out = 24'(-936);
			38700: out = 24'(84);
			38701: out = 24'(-336);
			38702: out = 24'(-4316);
			38703: out = 24'(-2760);
			38704: out = 24'(912);
			38705: out = 24'(2556);
			38706: out = 24'(68);
			38707: out = 24'(1412);
			38708: out = 24'(1732);
			38709: out = 24'(-700);
			38710: out = 24'(-5260);
			38711: out = 24'(-3992);
			38712: out = 24'(-1348);
			38713: out = 24'(776);
			38714: out = 24'(1984);
			38715: out = 24'(660);
			38716: out = 24'(-1184);
			38717: out = 24'(-444);
			38718: out = 24'(2960);
			38719: out = 24'(3844);
			38720: out = 24'(1612);
			38721: out = 24'(-800);
			38722: out = 24'(-1076);
			38723: out = 24'(-4020);
			38724: out = 24'(-2036);
			38725: out = 24'(836);
			38726: out = 24'(2824);
			38727: out = 24'(1944);
			38728: out = 24'(1876);
			38729: out = 24'(2316);
			38730: out = 24'(1684);
			38731: out = 24'(-2708);
			38732: out = 24'(-1928);
			38733: out = 24'(-740);
			38734: out = 24'(1104);
			38735: out = 24'(1752);
			38736: out = 24'(2680);
			38737: out = 24'(292);
			38738: out = 24'(-1476);
			38739: out = 24'(-1016);
			38740: out = 24'(-1864);
			38741: out = 24'(-1336);
			38742: out = 24'(-596);
			38743: out = 24'(-28);
			38744: out = 24'(-184);
			38745: out = 24'(336);
			38746: out = 24'(532);
			38747: out = 24'(620);
			38748: out = 24'(560);
			38749: out = 24'(1584);
			38750: out = 24'(1460);
			38751: out = 24'(-612);
			38752: out = 24'(-3112);
			38753: out = 24'(-884);
			38754: out = 24'(1460);
			38755: out = 24'(1076);
			38756: out = 24'(-1172);
			38757: out = 24'(-1196);
			38758: out = 24'(-228);
			38759: out = 24'(-1200);
			38760: out = 24'(-3300);
			38761: out = 24'(-1772);
			38762: out = 24'(1536);
			38763: out = 24'(1960);
			38764: out = 24'(-800);
			38765: out = 24'(-520);
			38766: out = 24'(-612);
			38767: out = 24'(564);
			38768: out = 24'(236);
			38769: out = 24'(84);
			38770: out = 24'(-1732);
			38771: out = 24'(-256);
			38772: out = 24'(316);
			38773: out = 24'(-1184);
			38774: out = 24'(-2304);
			38775: out = 24'(-956);
			38776: out = 24'(344);
			38777: out = 24'(-20);
			38778: out = 24'(696);
			38779: out = 24'(744);
			38780: out = 24'(424);
			38781: out = 24'(232);
			38782: out = 24'(1948);
			38783: out = 24'(500);
			38784: out = 24'(-972);
			38785: out = 24'(-1336);
			38786: out = 24'(488);
			38787: out = 24'(-1824);
			38788: out = 24'(-3116);
			38789: out = 24'(-1588);
			38790: out = 24'(3208);
			38791: out = 24'(3536);
			38792: out = 24'(1972);
			38793: out = 24'(-2956);
			38794: out = 24'(-5948);
			38795: out = 24'(-3672);
			38796: out = 24'(2632);
			38797: out = 24'(4424);
			38798: out = 24'(1888);
			38799: out = 24'(-756);
			38800: out = 24'(1280);
			38801: out = 24'(1408);
			38802: out = 24'(-392);
			38803: out = 24'(784);
			38804: out = 24'(-1308);
			38805: out = 24'(-2620);
			38806: out = 24'(-2548);
			38807: out = 24'(320);
			38808: out = 24'(420);
			38809: out = 24'(524);
			38810: out = 24'(-480);
			38811: out = 24'(-692);
			38812: out = 24'(-232);
			38813: out = 24'(1452);
			38814: out = 24'(2160);
			38815: out = 24'(1684);
			38816: out = 24'(4);
			38817: out = 24'(-1816);
			38818: out = 24'(-1752);
			38819: out = 24'(856);
			38820: out = 24'(1504);
			38821: out = 24'(1428);
			38822: out = 24'(-3024);
			38823: out = 24'(-4656);
			38824: out = 24'(384);
			38825: out = 24'(2296);
			38826: out = 24'(1332);
			38827: out = 24'(-248);
			38828: out = 24'(780);
			38829: out = 24'(-44);
			38830: out = 24'(-1384);
			38831: out = 24'(-2704);
			38832: out = 24'(-1912);
			38833: out = 24'(-188);
			38834: out = 24'(688);
			38835: out = 24'(460);
			38836: out = 24'(-168);
			38837: out = 24'(-760);
			38838: out = 24'(-516);
			38839: out = 24'(1108);
			38840: out = 24'(1784);
			38841: out = 24'(-92);
			38842: out = 24'(-112);
			38843: out = 24'(1108);
			38844: out = 24'(1760);
			38845: out = 24'(-472);
			38846: out = 24'(-588);
			38847: out = 24'(-1656);
			38848: out = 24'(-1156);
			38849: out = 24'(-216);
			38850: out = 24'(-804);
			38851: out = 24'(-468);
			38852: out = 24'(964);
			38853: out = 24'(1804);
			38854: out = 24'(0);
			38855: out = 24'(-764);
			38856: out = 24'(-564);
			38857: out = 24'(20);
			38858: out = 24'(-80);
			38859: out = 24'(12);
			38860: out = 24'(-216);
			38861: out = 24'(480);
			38862: out = 24'(2748);
			38863: out = 24'(1780);
			38864: out = 24'(2088);
			38865: out = 24'(596);
			38866: out = 24'(-2216);
			38867: out = 24'(-3960);
			38868: out = 24'(-3132);
			38869: out = 24'(-2312);
			38870: out = 24'(-2192);
			38871: out = 24'(-28);
			38872: out = 24'(1504);
			38873: out = 24'(2144);
			38874: out = 24'(1872);
			38875: out = 24'(1928);
			38876: out = 24'(1928);
			38877: out = 24'(520);
			38878: out = 24'(-1996);
			38879: out = 24'(-3040);
			38880: out = 24'(-880);
			38881: out = 24'(1796);
			38882: out = 24'(2108);
			38883: out = 24'(332);
			38884: out = 24'(-140);
			38885: out = 24'(-172);
			38886: out = 24'(-640);
			38887: out = 24'(-2180);
			38888: out = 24'(-3028);
			38889: out = 24'(-2540);
			38890: out = 24'(200);
			38891: out = 24'(2216);
			38892: out = 24'(2576);
			38893: out = 24'(820);
			38894: out = 24'(-336);
			38895: out = 24'(-1924);
			38896: out = 24'(-3988);
			38897: out = 24'(-4292);
			38898: out = 24'(-628);
			38899: out = 24'(3224);
			38900: out = 24'(3048);
			38901: out = 24'(-884);
			38902: out = 24'(-1020);
			38903: out = 24'(860);
			38904: out = 24'(1280);
			38905: out = 24'(516);
			38906: out = 24'(-1208);
			38907: out = 24'(-772);
			38908: out = 24'(612);
			38909: out = 24'(-300);
			38910: out = 24'(424);
			38911: out = 24'(-288);
			38912: out = 24'(-464);
			38913: out = 24'(1652);
			38914: out = 24'(1936);
			38915: out = 24'(668);
			38916: out = 24'(-2288);
			38917: out = 24'(-3992);
			38918: out = 24'(-4184);
			38919: out = 24'(-1524);
			38920: out = 24'(896);
			38921: out = 24'(1628);
			38922: out = 24'(1628);
			38923: out = 24'(504);
			38924: out = 24'(-604);
			38925: out = 24'(-528);
			38926: out = 24'(364);
			38927: out = 24'(1844);
			38928: out = 24'(880);
			38929: out = 24'(-1544);
			38930: out = 24'(-1844);
			38931: out = 24'(-568);
			38932: out = 24'(120);
			38933: out = 24'(-836);
			38934: out = 24'(-1156);
			38935: out = 24'(-484);
			38936: out = 24'(2144);
			38937: out = 24'(2836);
			38938: out = 24'(1036);
			38939: out = 24'(-1232);
			38940: out = 24'(-1640);
			38941: out = 24'(-1188);
			38942: out = 24'(-948);
			38943: out = 24'(-2032);
			38944: out = 24'(-572);
			38945: out = 24'(316);
			38946: out = 24'(152);
			38947: out = 24'(-820);
			38948: out = 24'(-64);
			38949: out = 24'(-484);
			38950: out = 24'(-524);
			38951: out = 24'(532);
			38952: out = 24'(2952);
			38953: out = 24'(1408);
			38954: out = 24'(-1156);
			38955: out = 24'(-1628);
			38956: out = 24'(1768);
			38957: out = 24'(856);
			38958: out = 24'(-968);
			38959: out = 24'(-1224);
			38960: out = 24'(-408);
			38961: out = 24'(-480);
			38962: out = 24'(-1432);
			38963: out = 24'(-1972);
			38964: out = 24'(-1244);
			38965: out = 24'(-328);
			38966: out = 24'(972);
			38967: out = 24'(1836);
			38968: out = 24'(1516);
			38969: out = 24'(152);
			38970: out = 24'(-172);
			38971: out = 24'(0);
			38972: out = 24'(-108);
			38973: out = 24'(-828);
			38974: out = 24'(-44);
			38975: out = 24'(428);
			38976: out = 24'(-252);
			38977: out = 24'(28);
			38978: out = 24'(-1064);
			38979: out = 24'(-1460);
			38980: out = 24'(-1140);
			38981: out = 24'(20);
			38982: out = 24'(-64);
			38983: out = 24'(276);
			38984: out = 24'(304);
			38985: out = 24'(0);
			38986: out = 24'(-152);
			38987: out = 24'(1140);
			38988: out = 24'(2744);
			38989: out = 24'(3528);
			38990: out = 24'(3092);
			38991: out = 24'(1028);
			38992: out = 24'(-1892);
			38993: out = 24'(-3172);
			38994: out = 24'(-1204);
			38995: out = 24'(124);
			38996: out = 24'(-52);
			38997: out = 24'(712);
			38998: out = 24'(4684);
			38999: out = 24'(4132);
			39000: out = 24'(-44);
			39001: out = 24'(-4192);
			39002: out = 24'(-3112);
			39003: out = 24'(-552);
			39004: out = 24'(436);
			39005: out = 24'(-476);
			39006: out = 24'(492);
			39007: out = 24'(-1692);
			39008: out = 24'(-616);
			39009: out = 24'(-980);
			39010: out = 24'(-2000);
			39011: out = 24'(-1632);
			39012: out = 24'(1004);
			39013: out = 24'(2300);
			39014: out = 24'(1732);
			39015: out = 24'(368);
			39016: out = 24'(1204);
			39017: out = 24'(728);
			39018: out = 24'(-644);
			39019: out = 24'(-1540);
			39020: out = 24'(-480);
			39021: out = 24'(-760);
			39022: out = 24'(-1976);
			39023: out = 24'(-2764);
			39024: out = 24'(-2728);
			39025: out = 24'(-1496);
			39026: out = 24'(1624);
			39027: out = 24'(4252);
			39028: out = 24'(960);
			39029: out = 24'(-4052);
			39030: out = 24'(-5616);
			39031: out = 24'(-1248);
			39032: out = 24'(1536);
			39033: out = 24'(3480);
			39034: out = 24'(1704);
			39035: out = 24'(228);
			39036: out = 24'(-300);
			39037: out = 24'(100);
			39038: out = 24'(-1208);
			39039: out = 24'(-1892);
			39040: out = 24'(-744);
			39041: out = 24'(0);
			39042: out = 24'(-1024);
			39043: out = 24'(-532);
			39044: out = 24'(1668);
			39045: out = 24'(700);
			39046: out = 24'(-936);
			39047: out = 24'(-372);
			39048: out = 24'(2436);
			39049: out = 24'(1896);
			39050: out = 24'(1684);
			39051: out = 24'(1372);
			39052: out = 24'(1172);
			39053: out = 24'(-296);
			39054: out = 24'(-8);
			39055: out = 24'(880);
			39056: out = 24'(1076);
			39057: out = 24'(-436);
			39058: out = 24'(-1988);
			39059: out = 24'(-1264);
			39060: out = 24'(-4);
			39061: out = 24'(-316);
			39062: out = 24'(184);
			39063: out = 24'(1076);
			39064: out = 24'(768);
			39065: out = 24'(-1408);
			39066: out = 24'(-2036);
			39067: out = 24'(-1968);
			39068: out = 24'(-888);
			39069: out = 24'(-76);
			39070: out = 24'(1520);
			39071: out = 24'(140);
			39072: out = 24'(-384);
			39073: out = 24'(-140);
			39074: out = 24'(-288);
			39075: out = 24'(-232);
			39076: out = 24'(-1108);
			39077: out = 24'(-1256);
			39078: out = 24'(0);
			39079: out = 24'(1716);
			39080: out = 24'(1172);
			39081: out = 24'(-160);
			39082: out = 24'(-128);
			39083: out = 24'(-1008);
			39084: out = 24'(-924);
			39085: out = 24'(-1036);
			39086: out = 24'(-820);
			39087: out = 24'(-976);
			39088: out = 24'(960);
			39089: out = 24'(1148);
			39090: out = 24'(152);
			39091: out = 24'(320);
			39092: out = 24'(-204);
			39093: out = 24'(-248);
			39094: out = 24'(-72);
			39095: out = 24'(360);
			39096: out = 24'(320);
			39097: out = 24'(20);
			39098: out = 24'(-352);
			39099: out = 24'(-120);
			39100: out = 24'(116);
			39101: out = 24'(492);
			39102: out = 24'(-1248);
			39103: out = 24'(-3456);
			39104: out = 24'(-908);
			39105: out = 24'(-944);
			39106: out = 24'(-568);
			39107: out = 24'(300);
			39108: out = 24'(2036);
			39109: out = 24'(2148);
			39110: out = 24'(780);
			39111: out = 24'(-160);
			39112: out = 24'(1608);
			39113: out = 24'(-148);
			39114: out = 24'(-244);
			39115: out = 24'(-420);
			39116: out = 24'(-316);
			39117: out = 24'(-3312);
			39118: out = 24'(-2312);
			39119: out = 24'(-1144);
			39120: out = 24'(-728);
			39121: out = 24'(-240);
			39122: out = 24'(1240);
			39123: out = 24'(584);
			39124: out = 24'(-1040);
			39125: out = 24'(-12);
			39126: out = 24'(1116);
			39127: out = 24'(868);
			39128: out = 24'(-828);
			39129: out = 24'(-700);
			39130: out = 24'(-112);
			39131: out = 24'(1148);
			39132: out = 24'(1556);
			39133: out = 24'(1916);
			39134: out = 24'(380);
			39135: out = 24'(-800);
			39136: out = 24'(-2544);
			39137: out = 24'(-3116);
			39138: out = 24'(-512);
			39139: out = 24'(512);
			39140: out = 24'(-716);
			39141: out = 24'(-2160);
			39142: out = 24'(-1432);
			39143: out = 24'(1208);
			39144: out = 24'(2828);
			39145: out = 24'(2688);
			39146: out = 24'(1284);
			39147: out = 24'(-428);
			39148: out = 24'(-2236);
			39149: out = 24'(-2172);
			39150: out = 24'(460);
			39151: out = 24'(1336);
			39152: out = 24'(808);
			39153: out = 24'(-88);
			39154: out = 24'(-244);
			39155: out = 24'(-280);
			39156: out = 24'(-720);
			39157: out = 24'(-808);
			39158: out = 24'(-28);
			39159: out = 24'(124);
			39160: out = 24'(-184);
			39161: out = 24'(-196);
			39162: out = 24'(704);
			39163: out = 24'(1252);
			39164: out = 24'(260);
			39165: out = 24'(-1820);
			39166: out = 24'(-2820);
			39167: out = 24'(-1924);
			39168: out = 24'(1020);
			39169: out = 24'(1140);
			39170: out = 24'(-308);
			39171: out = 24'(-808);
			39172: out = 24'(-328);
			39173: out = 24'(-96);
			39174: out = 24'(-300);
			39175: out = 24'(-116);
			39176: out = 24'(-284);
			39177: out = 24'(256);
			39178: out = 24'(-28);
			39179: out = 24'(112);
			39180: out = 24'(1376);
			39181: out = 24'(776);
			39182: out = 24'(-908);
			39183: out = 24'(-1100);
			39184: out = 24'(336);
			39185: out = 24'(1468);
			39186: out = 24'(-332);
			39187: out = 24'(-1456);
			39188: out = 24'(52);
			39189: out = 24'(1760);
			39190: out = 24'(592);
			39191: out = 24'(-388);
			39192: out = 24'(4);
			39193: out = 24'(-2836);
			39194: out = 24'(-2880);
			39195: out = 24'(-1820);
			39196: out = 24'(480);
			39197: out = 24'(1296);
			39198: out = 24'(2072);
			39199: out = 24'(888);
			39200: out = 24'(-760);
			39201: out = 24'(-1568);
			39202: out = 24'(-2688);
			39203: out = 24'(-2424);
			39204: out = 24'(-1856);
			39205: out = 24'(-1160);
			39206: out = 24'(1748);
			39207: out = 24'(3256);
			39208: out = 24'(2952);
			39209: out = 24'(1004);
			39210: out = 24'(-736);
			39211: out = 24'(-2348);
			39212: out = 24'(-2964);
			39213: out = 24'(-2300);
			39214: out = 24'(-112);
			39215: out = 24'(-660);
			39216: out = 24'(-612);
			39217: out = 24'(436);
			39218: out = 24'(1416);
			39219: out = 24'(252);
			39220: out = 24'(-436);
			39221: out = 24'(640);
			39222: out = 24'(1792);
			39223: out = 24'(-320);
			39224: out = 24'(-2388);
			39225: out = 24'(-1192);
			39226: out = 24'(2472);
			39227: out = 24'(1408);
			39228: out = 24'(548);
			39229: out = 24'(-1028);
			39230: out = 24'(-2596);
			39231: out = 24'(-5160);
			39232: out = 24'(-3812);
			39233: out = 24'(-1504);
			39234: out = 24'(496);
			39235: out = 24'(556);
			39236: out = 24'(2904);
			39237: out = 24'(2620);
			39238: out = 24'(1028);
			39239: out = 24'(536);
			39240: out = 24'(1308);
			39241: out = 24'(1764);
			39242: out = 24'(672);
			39243: out = 24'(-836);
			39244: out = 24'(64);
			39245: out = 24'(1596);
			39246: out = 24'(1616);
			39247: out = 24'(-340);
			39248: out = 24'(-3800);
			39249: out = 24'(-1464);
			39250: out = 24'(1356);
			39251: out = 24'(1576);
			39252: out = 24'(-836);
			39253: out = 24'(-1852);
			39254: out = 24'(-1664);
			39255: out = 24'(4);
			39256: out = 24'(1612);
			39257: out = 24'(2952);
			39258: out = 24'(1672);
			39259: out = 24'(-932);
			39260: out = 24'(-3516);
			39261: out = 24'(-2656);
			39262: out = 24'(-2092);
			39263: out = 24'(60);
			39264: out = 24'(2360);
			39265: out = 24'(3080);
			39266: out = 24'(336);
			39267: out = 24'(-1272);
			39268: out = 24'(-584);
			39269: out = 24'(-204);
			39270: out = 24'(-1056);
			39271: out = 24'(-1412);
			39272: out = 24'(-144);
			39273: out = 24'(1560);
			39274: out = 24'(632);
			39275: out = 24'(396);
			39276: out = 24'(132);
			39277: out = 24'(-956);
			39278: out = 24'(-1400);
			39279: out = 24'(-388);
			39280: out = 24'(1252);
			39281: out = 24'(1848);
			39282: out = 24'(-32);
			39283: out = 24'(-256);
			39284: out = 24'(-768);
			39285: out = 24'(-1624);
			39286: out = 24'(-1376);
			39287: out = 24'(-48);
			39288: out = 24'(408);
			39289: out = 24'(-576);
			39290: out = 24'(-1252);
			39291: out = 24'(-2112);
			39292: out = 24'(-888);
			39293: out = 24'(80);
			39294: out = 24'(-140);
			39295: out = 24'(-1180);
			39296: out = 24'(-1428);
			39297: out = 24'(-1100);
			39298: out = 24'(-604);
			39299: out = 24'(308);
			39300: out = 24'(1336);
			39301: out = 24'(1732);
			39302: out = 24'(1416);
			39303: out = 24'(-72);
			39304: out = 24'(-8);
			39305: out = 24'(-632);
			39306: out = 24'(-1504);
			39307: out = 24'(-620);
			39308: out = 24'(968);
			39309: out = 24'(2580);
			39310: out = 24'(2820);
			39311: out = 24'(1192);
			39312: out = 24'(176);
			39313: out = 24'(-1848);
			39314: out = 24'(-2832);
			39315: out = 24'(-1704);
			39316: out = 24'(1552);
			39317: out = 24'(1956);
			39318: out = 24'(708);
			39319: out = 24'(-272);
			39320: out = 24'(-300);
			39321: out = 24'(964);
			39322: out = 24'(1164);
			39323: out = 24'(-232);
			39324: out = 24'(-1408);
			39325: out = 24'(-2908);
			39326: out = 24'(-1336);
			39327: out = 24'(512);
			39328: out = 24'(-292);
			39329: out = 24'(280);
			39330: out = 24'(1216);
			39331: out = 24'(2212);
			39332: out = 24'(1736);
			39333: out = 24'(2092);
			39334: out = 24'(392);
			39335: out = 24'(-904);
			39336: out = 24'(-1968);
			39337: out = 24'(-3344);
			39338: out = 24'(-2888);
			39339: out = 24'(-500);
			39340: out = 24'(1720);
			39341: out = 24'(1336);
			39342: out = 24'(-284);
			39343: out = 24'(-1812);
			39344: out = 24'(-2196);
			39345: out = 24'(-2116);
			39346: out = 24'(-1160);
			39347: out = 24'(-740);
			39348: out = 24'(-1272);
			39349: out = 24'(-1880);
			39350: out = 24'(72);
			39351: out = 24'(2220);
			39352: out = 24'(3348);
			39353: out = 24'(2660);
			39354: out = 24'(488);
			39355: out = 24'(-2112);
			39356: out = 24'(-4484);
			39357: out = 24'(-3856);
			39358: out = 24'(-444);
			39359: out = 24'(1708);
			39360: out = 24'(-476);
			39361: out = 24'(-2476);
			39362: out = 24'(132);
			39363: out = 24'(3052);
			39364: out = 24'(2244);
			39365: out = 24'(-940);
			39366: out = 24'(-2496);
			39367: out = 24'(-516);
			39368: out = 24'(64);
			39369: out = 24'(0);
			39370: out = 24'(524);
			39371: out = 24'(-104);
			39372: out = 24'(-968);
			39373: out = 24'(-1152);
			39374: out = 24'(400);
			39375: out = 24'(1340);
			39376: out = 24'(884);
			39377: out = 24'(-932);
			39378: out = 24'(-2468);
			39379: out = 24'(-3208);
			39380: out = 24'(-872);
			39381: out = 24'(1044);
			39382: out = 24'(1320);
			39383: out = 24'(-224);
			39384: out = 24'(-1668);
			39385: out = 24'(-2188);
			39386: out = 24'(-1536);
			39387: out = 24'(-640);
			39388: out = 24'(-676);
			39389: out = 24'(80);
			39390: out = 24'(1176);
			39391: out = 24'(1540);
			39392: out = 24'(644);
			39393: out = 24'(84);
			39394: out = 24'(128);
			39395: out = 24'(772);
			39396: out = 24'(1604);
			39397: out = 24'(260);
			39398: out = 24'(-212);
			39399: out = 24'(-76);
			39400: out = 24'(-1004);
			39401: out = 24'(-692);
			39402: out = 24'(-1232);
			39403: out = 24'(-840);
			39404: out = 24'(864);
			39405: out = 24'(1872);
			39406: out = 24'(1328);
			39407: out = 24'(-448);
			39408: out = 24'(-1432);
			39409: out = 24'(-1456);
			39410: out = 24'(-48);
			39411: out = 24'(368);
			39412: out = 24'(-72);
			39413: out = 24'(624);
			39414: out = 24'(-64);
			39415: out = 24'(760);
			39416: out = 24'(1560);
			39417: out = 24'(260);
			39418: out = 24'(1624);
			39419: out = 24'(-396);
			39420: out = 24'(-3052);
			39421: out = 24'(-3456);
			39422: out = 24'(1420);
			39423: out = 24'(3440);
			39424: out = 24'(2904);
			39425: out = 24'(1156);
			39426: out = 24'(-4);
			39427: out = 24'(-12);
			39428: out = 24'(916);
			39429: out = 24'(1184);
			39430: out = 24'(-192);
			39431: out = 24'(-3136);
			39432: out = 24'(-4004);
			39433: out = 24'(-1516);
			39434: out = 24'(1544);
			39435: out = 24'(1688);
			39436: out = 24'(532);
			39437: out = 24'(-788);
			39438: out = 24'(-1400);
			39439: out = 24'(-308);
			39440: out = 24'(-52);
			39441: out = 24'(-384);
			39442: out = 24'(-884);
			39443: out = 24'(-844);
			39444: out = 24'(676);
			39445: out = 24'(2640);
			39446: out = 24'(3176);
			39447: out = 24'(320);
			39448: out = 24'(-76);
			39449: out = 24'(-1792);
			39450: out = 24'(-3696);
			39451: out = 24'(-2396);
			39452: out = 24'(-912);
			39453: out = 24'(1504);
			39454: out = 24'(1224);
			39455: out = 24'(-1648);
			39456: out = 24'(-3756);
			39457: out = 24'(-1916);
			39458: out = 24'(1448);
			39459: out = 24'(2932);
			39460: out = 24'(200);
			39461: out = 24'(-312);
			39462: out = 24'(0);
			39463: out = 24'(-308);
			39464: out = 24'(-812);
			39465: out = 24'(876);
			39466: out = 24'(1900);
			39467: out = 24'(1044);
			39468: out = 24'(-868);
			39469: out = 24'(-1356);
			39470: out = 24'(-1440);
			39471: out = 24'(-1724);
			39472: out = 24'(-2652);
			39473: out = 24'(-1452);
			39474: out = 24'(-636);
			39475: out = 24'(868);
			39476: out = 24'(2116);
			39477: out = 24'(1840);
			39478: out = 24'(-1552);
			39479: out = 24'(-3404);
			39480: out = 24'(-1064);
			39481: out = 24'(1740);
			39482: out = 24'(2584);
			39483: out = 24'(560);
			39484: out = 24'(-1888);
			39485: out = 24'(-2372);
			39486: out = 24'(412);
			39487: out = 24'(3584);
			39488: out = 24'(3804);
			39489: out = 24'(220);
			39490: out = 24'(404);
			39491: out = 24'(80);
			39492: out = 24'(-444);
			39493: out = 24'(-860);
			39494: out = 24'(-296);
			39495: out = 24'(-116);
			39496: out = 24'(-488);
			39497: out = 24'(-892);
			39498: out = 24'(-992);
			39499: out = 24'(88);
			39500: out = 24'(280);
			39501: out = 24'(-452);
			39502: out = 24'(-1364);
			39503: out = 24'(-460);
			39504: out = 24'(8);
			39505: out = 24'(-200);
			39506: out = 24'(36);
			39507: out = 24'(1588);
			39508: out = 24'(2340);
			39509: out = 24'(1476);
			39510: out = 24'(304);
			39511: out = 24'(-272);
			39512: out = 24'(-780);
			39513: out = 24'(-2720);
			39514: out = 24'(-4596);
			39515: out = 24'(-2832);
			39516: out = 24'(284);
			39517: out = 24'(2644);
			39518: out = 24'(2880);
			39519: out = 24'(1592);
			39520: out = 24'(-664);
			39521: out = 24'(-2368);
			39522: out = 24'(-2224);
			39523: out = 24'(-40);
			39524: out = 24'(1256);
			39525: out = 24'(1396);
			39526: out = 24'(624);
			39527: out = 24'(-212);
			39528: out = 24'(-780);
			39529: out = 24'(-608);
			39530: out = 24'(548);
			39531: out = 24'(1268);
			39532: out = 24'(-1076);
			39533: out = 24'(-2592);
			39534: out = 24'(-1652);
			39535: out = 24'(808);
			39536: out = 24'(340);
			39537: out = 24'(88);
			39538: out = 24'(-372);
			39539: out = 24'(232);
			39540: out = 24'(1492);
			39541: out = 24'(272);
			39542: out = 24'(-356);
			39543: out = 24'(-60);
			39544: out = 24'(-388);
			39545: out = 24'(456);
			39546: out = 24'(0);
			39547: out = 24'(-28);
			39548: out = 24'(432);
			39549: out = 24'(1532);
			39550: out = 24'(-92);
			39551: out = 24'(-1004);
			39552: out = 24'(316);
			39553: out = 24'(1688);
			39554: out = 24'(740);
			39555: out = 24'(-2000);
			39556: out = 24'(-3108);
			39557: out = 24'(-888);
			39558: out = 24'(-256);
			39559: out = 24'(120);
			39560: out = 24'(880);
			39561: out = 24'(1940);
			39562: out = 24'(1708);
			39563: out = 24'(40);
			39564: out = 24'(-1264);
			39565: out = 24'(-1508);
			39566: out = 24'(152);
			39567: out = 24'(-1580);
			39568: out = 24'(-2580);
			39569: out = 24'(116);
			39570: out = 24'(3692);
			39571: out = 24'(3220);
			39572: out = 24'(600);
			39573: out = 24'(-1768);
			39574: out = 24'(-2808);
			39575: out = 24'(-2416);
			39576: out = 24'(-1688);
			39577: out = 24'(-896);
			39578: out = 24'(-92);
			39579: out = 24'(-200);
			39580: out = 24'(536);
			39581: out = 24'(1432);
			39582: out = 24'(1384);
			39583: out = 24'(-48);
			39584: out = 24'(-772);
			39585: out = 24'(-540);
			39586: out = 24'(-128);
			39587: out = 24'(-264);
			39588: out = 24'(-196);
			39589: out = 24'(-24);
			39590: out = 24'(292);
			39591: out = 24'(-272);
			39592: out = 24'(156);
			39593: out = 24'(40);
			39594: out = 24'(-224);
			39595: out = 24'(-296);
			39596: out = 24'(-1764);
			39597: out = 24'(-2480);
			39598: out = 24'(-1204);
			39599: out = 24'(1312);
			39600: out = 24'(1236);
			39601: out = 24'(-244);
			39602: out = 24'(-1184);
			39603: out = 24'(272);
			39604: out = 24'(884);
			39605: out = 24'(1632);
			39606: out = 24'(820);
			39607: out = 24'(-316);
			39608: out = 24'(-348);
			39609: out = 24'(-188);
			39610: out = 24'(-452);
			39611: out = 24'(-808);
			39612: out = 24'(-740);
			39613: out = 24'(1108);
			39614: out = 24'(1476);
			39615: out = 24'(692);
			39616: out = 24'(232);
			39617: out = 24'(-200);
			39618: out = 24'(-296);
			39619: out = 24'(-572);
			39620: out = 24'(-772);
			39621: out = 24'(-216);
			39622: out = 24'(8);
			39623: out = 24'(576);
			39624: out = 24'(1068);
			39625: out = 24'(1044);
			39626: out = 24'(316);
			39627: out = 24'(-580);
			39628: out = 24'(-1620);
			39629: out = 24'(-2192);
			39630: out = 24'(-2084);
			39631: out = 24'(-524);
			39632: out = 24'(232);
			39633: out = 24'(-132);
			39634: out = 24'(-20);
			39635: out = 24'(1440);
			39636: out = 24'(2080);
			39637: out = 24'(232);
			39638: out = 24'(-976);
			39639: out = 24'(-1836);
			39640: out = 24'(-1184);
			39641: out = 24'(-20);
			39642: out = 24'(636);
			39643: out = 24'(1228);
			39644: out = 24'(1252);
			39645: out = 24'(152);
			39646: out = 24'(-1216);
			39647: out = 24'(-1496);
			39648: out = 24'(-656);
			39649: out = 24'(-132);
			39650: out = 24'(200);
			39651: out = 24'(-368);
			39652: out = 24'(624);
			39653: out = 24'(520);
			39654: out = 24'(-1452);
			39655: out = 24'(-724);
			39656: out = 24'(-516);
			39657: out = 24'(-172);
			39658: out = 24'(-352);
			39659: out = 24'(-128);
			39660: out = 24'(-292);
			39661: out = 24'(-184);
			39662: out = 24'(-288);
			39663: out = 24'(-772);
			39664: out = 24'(-128);
			39665: out = 24'(684);
			39666: out = 24'(1128);
			39667: out = 24'(996);
			39668: out = 24'(-792);
			39669: out = 24'(-2312);
			39670: out = 24'(-2360);
			39671: out = 24'(-452);
			39672: out = 24'(864);
			39673: out = 24'(1304);
			39674: out = 24'(600);
			39675: out = 24'(-176);
			39676: out = 24'(176);
			39677: out = 24'(324);
			39678: out = 24'(-4);
			39679: out = 24'(-164);
			39680: out = 24'(284);
			39681: out = 24'(-164);
			39682: out = 24'(-36);
			39683: out = 24'(268);
			39684: out = 24'(-308);
			39685: out = 24'(-556);
			39686: out = 24'(-1416);
			39687: out = 24'(-1288);
			39688: out = 24'(-48);
			39689: out = 24'(1008);
			39690: out = 24'(-84);
			39691: out = 24'(-1836);
			39692: out = 24'(-1848);
			39693: out = 24'(-400);
			39694: out = 24'(684);
			39695: out = 24'(392);
			39696: out = 24'(-36);
			39697: out = 24'(1120);
			39698: out = 24'(912);
			39699: out = 24'(264);
			39700: out = 24'(-320);
			39701: out = 24'(-108);
			39702: out = 24'(-224);
			39703: out = 24'(44);
			39704: out = 24'(92);
			39705: out = 24'(184);
			39706: out = 24'(-152);
			39707: out = 24'(-188);
			39708: out = 24'(-496);
			39709: out = 24'(-1200);
			39710: out = 24'(-844);
			39711: out = 24'(480);
			39712: out = 24'(1140);
			39713: out = 24'(452);
			39714: out = 24'(-120);
			39715: out = 24'(-404);
			39716: out = 24'(204);
			39717: out = 24'(596);
			39718: out = 24'(-232);
			39719: out = 24'(-240);
			39720: out = 24'(-236);
			39721: out = 24'(-720);
			39722: out = 24'(-2200);
			39723: out = 24'(-588);
			39724: out = 24'(128);
			39725: out = 24'(180);
			39726: out = 24'(-252);
			39727: out = 24'(-60);
			39728: out = 24'(-272);
			39729: out = 24'(304);
			39730: out = 24'(1148);
			39731: out = 24'(1156);
			39732: out = 24'(176);
			39733: out = 24'(-328);
			39734: out = 24'(-252);
			39735: out = 24'(252);
			39736: out = 24'(-148);
			39737: out = 24'(332);
			39738: out = 24'(1024);
			39739: out = 24'(596);
			39740: out = 24'(-1336);
			39741: out = 24'(-1164);
			39742: out = 24'(272);
			39743: out = 24'(448);
			39744: out = 24'(400);
			39745: out = 24'(-492);
			39746: out = 24'(-848);
			39747: out = 24'(-760);
			39748: out = 24'(-296);
			39749: out = 24'(56);
			39750: out = 24'(240);
			39751: out = 24'(200);
			39752: out = 24'(24);
			39753: out = 24'(-52);
			39754: out = 24'(-552);
			39755: out = 24'(-816);
			39756: out = 24'(-816);
			39757: out = 24'(-344);
			39758: out = 24'(-300);
			39759: out = 24'(168);
			39760: out = 24'(1424);
			39761: out = 24'(1576);
			39762: out = 24'(-128);
			39763: out = 24'(-1848);
			39764: out = 24'(-1600);
			39765: out = 24'(-652);
			39766: out = 24'(112);
			39767: out = 24'(120);
			39768: out = 24'(68);
			39769: out = 24'(-244);
			39770: out = 24'(604);
			39771: out = 24'(1220);
			39772: out = 24'(656);
			39773: out = 24'(-200);
			39774: out = 24'(-1896);
			39775: out = 24'(-2260);
			39776: out = 24'(-1316);
			39777: out = 24'(-196);
			39778: out = 24'(104);
			39779: out = 24'(608);
			39780: out = 24'(1236);
			39781: out = 24'(892);
			39782: out = 24'(-144);
			39783: out = 24'(-1064);
			39784: out = 24'(-1608);
			39785: out = 24'(-2396);
			39786: out = 24'(-2620);
			39787: out = 24'(-2164);
			39788: out = 24'(-352);
			39789: out = 24'(0);
			default: out = 0;
		endcase
	end
endmodule
