module closed_hihat_lookup(index, out);
	input logic unsigned [12:0] index;
	output logic signed [15:0] out;
	always_comb begin
		case(index)
			0: out = 16'(0);
			1: out = 16'(0);
			2: out = 16'(32);
			3: out = 16'(-119);
			4: out = 16'(58);
			5: out = 16'(-153);
			6: out = 16'(92);
			7: out = 16'(-190);
			8: out = 16'(136);
			9: out = 16'(-246);
			10: out = 16'(200);
			11: out = 16'(-319);
			12: out = 16'(297);
			13: out = 16'(-483);
			14: out = 16'(547);
			15: out = 16'(-878);
			16: out = 16'(1307);
			17: out = 16'(-3640);
			18: out = 16'(10313);
			19: out = 16'(28235);
			20: out = 16'(-7945);
			21: out = 16'(-14803);
			22: out = 16'(-10656);
			23: out = 16'(16897);
			24: out = 16'(11531);
			25: out = 16'(25476);
			26: out = 16'(18093);
			27: out = 16'(-24016);
			28: out = 16'(-32233);
			29: out = 16'(-18973);
			30: out = 16'(21890);
			31: out = 16'(32766);
			32: out = 16'(2660);
			33: out = 16'(-26774);
			34: out = 16'(2755);
			35: out = 16'(19409);
			36: out = 16'(18764);
			37: out = 16'(2127);
			38: out = 16'(-23090);
			39: out = 16'(-6566);
			40: out = 16'(25030);
			41: out = 16'(13385);
			42: out = 16'(-3886);
			43: out = 16'(-21541);
			44: out = 16'(-6370);
			45: out = 16'(-19167);
			46: out = 16'(13611);
			47: out = 16'(29083);
			48: out = 16'(10383);
			49: out = 16'(-21719);
			50: out = 16'(-26613);
			51: out = 16'(2850);
			52: out = 16'(26300);
			53: out = 16'(21752);
			54: out = 16'(-3890);
			55: out = 16'(-27220);
			56: out = 16'(-30392);
			57: out = 16'(-18168);
			58: out = 16'(10331);
			59: out = 16'(12542);
			60: out = 16'(28421);
			61: out = 16'(25950);
			62: out = 16'(-2113);
			63: out = 16'(-29121);
			64: out = 16'(-21128);
			65: out = 16'(9847);
			66: out = 16'(2457);
			67: out = 16'(-19081);
			68: out = 16'(-21331);
			69: out = 16'(20606);
			70: out = 16'(22360);
			71: out = 16'(6566);
			72: out = 16'(-19978);
			73: out = 16'(-22152);
			74: out = 16'(-2669);
			75: out = 16'(6393);
			76: out = 16'(-32767);
			77: out = 16'(10745);
			78: out = 16'(31143);
			79: out = 16'(27750);
			80: out = 16'(-21633);
			81: out = 16'(-21762);
			82: out = 16'(4059);
			83: out = 16'(29968);
			84: out = 16'(7570);
			85: out = 16'(11368);
			86: out = 16'(25175);
			87: out = 16'(2197);
			88: out = 16'(-22613);
			89: out = 16'(-29578);
			90: out = 16'(-819);
			91: out = 16'(22699);
			92: out = 16'(26716);
			93: out = 16'(15728);
			94: out = 16'(-16111);
			95: out = 16'(-27365);
			96: out = 16'(-29169);
			97: out = 16'(-27843);
			98: out = 16'(-16531);
			99: out = 16'(6147);
			100: out = 16'(18385);
			101: out = 16'(9038);
			102: out = 16'(-2680);
			103: out = 16'(-5933);
			104: out = 16'(-5193);
			105: out = 16'(20765);
			106: out = 16'(-2375);
			107: out = 16'(-31471);
			108: out = 16'(-29787);
			109: out = 16'(-10570);
			110: out = 16'(23451);
			111: out = 16'(11859);
			112: out = 16'(-16740);
			113: out = 16'(-29622);
			114: out = 16'(-11348);
			115: out = 16'(-31784);
			116: out = 16'(4696);
			117: out = 16'(3193);
			118: out = 16'(-27904);
			119: out = 16'(-30997);
			120: out = 16'(-2524);
			121: out = 16'(23725);
			122: out = 16'(-22580);
			123: out = 16'(-22543);
			124: out = 16'(-21225);
			125: out = 16'(-11261);
			126: out = 16'(-18980);
			127: out = 16'(-20967);
			128: out = 16'(-19514);
			129: out = 16'(19149);
			130: out = 16'(-15289);
			131: out = 16'(-25307);
			132: out = 16'(-2883);
			133: out = 16'(-8548);
			134: out = 16'(-18715);
			135: out = 16'(-28011);
			136: out = 16'(-24819);
			137: out = 16'(-7845);
			138: out = 16'(3022);
			139: out = 16'(-1948);
			140: out = 16'(-25456);
			141: out = 16'(-21096);
			142: out = 16'(-5243);
			143: out = 16'(-25887);
			144: out = 16'(-757);
			145: out = 16'(13870);
			146: out = 16'(10923);
			147: out = 16'(-12363);
			148: out = 16'(-23698);
			149: out = 16'(-3094);
			150: out = 16'(31576);
			151: out = 16'(29227);
			152: out = 16'(27094);
			153: out = 16'(-123);
			154: out = 16'(-26866);
			155: out = 16'(-29840);
			156: out = 16'(-24229);
			157: out = 16'(7490);
			158: out = 16'(29208);
			159: out = 16'(26027);
			160: out = 16'(12825);
			161: out = 16'(-6994);
			162: out = 16'(-2322);
			163: out = 16'(11179);
			164: out = 16'(17303);
			165: out = 16'(2396);
			166: out = 16'(-19236);
			167: out = 16'(-29909);
			168: out = 16'(-22368);
			169: out = 16'(-13192);
			170: out = 16'(121);
			171: out = 16'(16890);
			172: out = 16'(5157);
			173: out = 16'(-15963);
			174: out = 16'(-23413);
			175: out = 16'(24180);
			176: out = 16'(31981);
			177: out = 16'(25222);
			178: out = 16'(6692);
			179: out = 16'(-13205);
			180: out = 16'(-17461);
			181: out = 16'(-378);
			182: out = 16'(27364);
			183: out = 16'(30401);
			184: out = 16'(30359);
			185: out = 16'(29769);
			186: out = 16'(26778);
			187: out = 16'(7114);
			188: out = 16'(-13277);
			189: out = 16'(-29324);
			190: out = 16'(-11204);
			191: out = 16'(15276);
			192: out = 16'(29788);
			193: out = 16'(-5911);
			194: out = 16'(-15930);
			195: out = 16'(-452);
			196: out = 16'(26357);
			197: out = 16'(15611);
			198: out = 16'(-2919);
			199: out = 16'(-18125);
			200: out = 16'(4856);
			201: out = 16'(11315);
			202: out = 16'(13671);
			203: out = 16'(28373);
			204: out = 16'(30656);
			205: out = 16'(9212);
			206: out = 16'(-28914);
			207: out = 16'(-22552);
			208: out = 16'(8766);
			209: out = 16'(32766);
			210: out = 16'(28179);
			211: out = 16'(27023);
			212: out = 16'(14752);
			213: out = 16'(-2100);
			214: out = 16'(-24482);
			215: out = 16'(-31229);
			216: out = 16'(-19310);
			217: out = 16'(25686);
			218: out = 16'(32471);
			219: out = 16'(15052);
			220: out = 16'(-20949);
			221: out = 16'(11501);
			222: out = 16'(24393);
			223: out = 16'(18304);
			224: out = 16'(-25892);
			225: out = 16'(-15257);
			226: out = 16'(-9582);
			227: out = 16'(-20440);
			228: out = 16'(20486);
			229: out = 16'(15056);
			230: out = 16'(4730);
			231: out = 16'(5779);
			232: out = 16'(22830);
			233: out = 16'(21238);
			234: out = 16'(1232);
			235: out = 16'(-15494);
			236: out = 16'(-4983);
			237: out = 16'(15591);
			238: out = 16'(-2770);
			239: out = 16'(11574);
			240: out = 16'(1735);
			241: out = 16'(-7430);
			242: out = 16'(-16940);
			243: out = 16'(10551);
			244: out = 16'(25648);
			245: out = 16'(4839);
			246: out = 16'(-6407);
			247: out = 16'(-20793);
			248: out = 16'(-24023);
			249: out = 16'(24459);
			250: out = 16'(12010);
			251: out = 16'(-17913);
			252: out = 16'(-30199);
			253: out = 16'(-16960);
			254: out = 16'(4461);
			255: out = 16'(6767);
			256: out = 16'(-30566);
			257: out = 16'(-1381);
			258: out = 16'(32030);
			259: out = 16'(10007);
			260: out = 16'(-20486);
			261: out = 16'(-31854);
			262: out = 16'(-9272);
			263: out = 16'(22594);
			264: out = 16'(32444);
			265: out = 16'(18535);
			266: out = 16'(-1817);
			267: out = 16'(-2525);
			268: out = 16'(13230);
			269: out = 16'(25660);
			270: out = 16'(20524);
			271: out = 16'(13523);
			272: out = 16'(4507);
			273: out = 16'(-11142);
			274: out = 16'(20275);
			275: out = 16'(19323);
			276: out = 16'(6085);
			277: out = 16'(-2843);
			278: out = 16'(10518);
			279: out = 16'(7933);
			280: out = 16'(-28064);
			281: out = 16'(3506);
			282: out = 16'(16738);
			283: out = 16'(13564);
			284: out = 16'(-15251);
			285: out = 16'(-27896);
			286: out = 16'(-21700);
			287: out = 16'(4130);
			288: out = 16'(-18181);
			289: out = 16'(-26075);
			290: out = 16'(-20910);
			291: out = 16'(-18414);
			292: out = 16'(9407);
			293: out = 16'(12578);
			294: out = 16'(-15925);
			295: out = 16'(-6746);
			296: out = 16'(-10846);
			297: out = 16'(-19473);
			298: out = 16'(-29847);
			299: out = 16'(-27873);
			300: out = 16'(-25394);
			301: out = 16'(-13186);
			302: out = 16'(618);
			303: out = 16'(10618);
			304: out = 16'(5104);
			305: out = 16'(-8343);
			306: out = 16'(-26901);
			307: out = 16'(-21427);
			308: out = 16'(1985);
			309: out = 16'(-8295);
			310: out = 16'(-22516);
			311: out = 16'(-18475);
			312: out = 16'(28628);
			313: out = 16'(16891);
			314: out = 16'(-4064);
			315: out = 16'(-25675);
			316: out = 16'(-4314);
			317: out = 16'(16827);
			318: out = 16'(19455);
			319: out = 16'(-22561);
			320: out = 16'(-5934);
			321: out = 16'(16410);
			322: out = 16'(27761);
			323: out = 16'(-25570);
			324: out = 16'(-16181);
			325: out = 16'(20439);
			326: out = 16'(30048);
			327: out = 16'(27279);
			328: out = 16'(16992);
			329: out = 16'(4472);
			330: out = 16'(12107);
			331: out = 16'(-3678);
			332: out = 16'(-17622);
			333: out = 16'(-16105);
			334: out = 16'(15579);
			335: out = 16'(28585);
			336: out = 16'(16512);
			337: out = 16'(20042);
			338: out = 16'(3659);
			339: out = 16'(2059);
			340: out = 16'(14227);
			341: out = 16'(9301);
			342: out = 16'(-1203);
			343: out = 16'(-7583);
			344: out = 16'(-7928);
			345: out = 16'(17121);
			346: out = 16'(28800);
			347: out = 16'(15328);
			348: out = 16'(13063);
			349: out = 16'(17819);
			350: out = 16'(24164);
			351: out = 16'(-22047);
			352: out = 16'(-10250);
			353: out = 16'(8816);
			354: out = 16'(16130);
			355: out = 16'(4773);
			356: out = 16'(-8411);
			357: out = 16'(-14291);
			358: out = 16'(-1145);
			359: out = 16'(6195);
			360: out = 16'(15400);
			361: out = 16'(29084);
			362: out = 16'(-3308);
			363: out = 16'(-6547);
			364: out = 16'(7418);
			365: out = 16'(9688);
			366: out = 16'(17827);
			367: out = 16'(7374);
			368: out = 16'(-21302);
			369: out = 16'(3017);
			370: out = 16'(12675);
			371: out = 16'(12620);
			372: out = 16'(-623);
			373: out = 16'(11053);
			374: out = 16'(16109);
			375: out = 16'(2992);
			376: out = 16'(-23777);
			377: out = 16'(-30909);
			378: out = 16'(-23457);
			379: out = 16'(11711);
			380: out = 16'(20332);
			381: out = 16'(18352);
			382: out = 16'(14185);
			383: out = 16'(-11184);
			384: out = 16'(-15717);
			385: out = 16'(-4567);
			386: out = 16'(2804);
			387: out = 16'(2952);
			388: out = 16'(-6198);
			389: out = 16'(-9197);
			390: out = 16'(-21073);
			391: out = 16'(-8928);
			392: out = 16'(5307);
			393: out = 16'(25064);
			394: out = 16'(-10637);
			395: out = 16'(-16388);
			396: out = 16'(11831);
			397: out = 16'(-15765);
			398: out = 16'(-27727);
			399: out = 16'(-27583);
			400: out = 16'(-14907);
			401: out = 16'(22003);
			402: out = 16'(24287);
			403: out = 16'(3375);
			404: out = 16'(-27780);
			405: out = 16'(-13503);
			406: out = 16'(14516);
			407: out = 16'(13001);
			408: out = 16'(-6313);
			409: out = 16'(-24102);
			410: out = 16'(-28598);
			411: out = 16'(14224);
			412: out = 16'(264);
			413: out = 16'(-28344);
			414: out = 16'(-29081);
			415: out = 16'(7652);
			416: out = 16'(29519);
			417: out = 16'(11972);
			418: out = 16'(2273);
			419: out = 16'(-19840);
			420: out = 16'(-26033);
			421: out = 16'(-9151);
			422: out = 16'(-24140);
			423: out = 16'(-20022);
			424: out = 16'(8942);
			425: out = 16'(17468);
			426: out = 16'(19887);
			427: out = 16'(7694);
			428: out = 16'(-7338);
			429: out = 16'(-14157);
			430: out = 16'(-9353);
			431: out = 16'(1049);
			432: out = 16'(3709);
			433: out = 16'(12002);
			434: out = 16'(8639);
			435: out = 16'(-16621);
			436: out = 16'(-4412);
			437: out = 16'(15822);
			438: out = 16'(30162);
			439: out = 16'(-5194);
			440: out = 16'(-1628);
			441: out = 16'(3143);
			442: out = 16'(1664);
			443: out = 16'(-23770);
			444: out = 16'(-23719);
			445: out = 16'(-666);
			446: out = 16'(5058);
			447: out = 16'(974);
			448: out = 16'(2710);
			449: out = 16'(32766);
			450: out = 16'(-8029);
			451: out = 16'(-3051);
			452: out = 16'(17824);
			453: out = 16'(30077);
			454: out = 16'(-1083);
			455: out = 16'(-23216);
			456: out = 16'(-3526);
			457: out = 16'(8506);
			458: out = 16'(19768);
			459: out = 16'(17438);
			460: out = 16'(25091);
			461: out = 16'(17229);
			462: out = 16'(13445);
			463: out = 16'(260);
			464: out = 16'(20024);
			465: out = 16'(4517);
			466: out = 16'(-11559);
			467: out = 16'(-908);
			468: out = 16'(21219);
			469: out = 16'(28620);
			470: out = 16'(17271);
			471: out = 16'(2415);
			472: out = 16'(-2060);
			473: out = 16'(332);
			474: out = 16'(-9150);
			475: out = 16'(-23582);
			476: out = 16'(-28281);
			477: out = 16'(-8129);
			478: out = 16'(7363);
			479: out = 16'(17100);
			480: out = 16'(8733);
			481: out = 16'(-10473);
			482: out = 16'(-16026);
			483: out = 16'(-2913);
			484: out = 16'(12005);
			485: out = 16'(3660);
			486: out = 16'(-3130);
			487: out = 16'(-3702);
			488: out = 16'(-12917);
			489: out = 16'(6951);
			490: out = 16'(7135);
			491: out = 16'(-1084);
			492: out = 16'(-25264);
			493: out = 16'(-3377);
			494: out = 16'(24640);
			495: out = 16'(30195);
			496: out = 16'(-7991);
			497: out = 16'(-22948);
			498: out = 16'(-1049);
			499: out = 16'(-16471);
			500: out = 16'(-20898);
			501: out = 16'(-25869);
			502: out = 16'(-14664);
			503: out = 16'(-672);
			504: out = 16'(2844);
			505: out = 16'(-9734);
			506: out = 16'(-8171);
			507: out = 16'(2169);
			508: out = 16'(10660);
			509: out = 16'(-23955);
			510: out = 16'(8484);
			511: out = 16'(-1717);
			512: out = 16'(-29522);
			513: out = 16'(-21418);
			514: out = 16'(2386);
			515: out = 16'(24855);
			516: out = 16'(20245);
			517: out = 16'(11440);
			518: out = 16'(-15752);
			519: out = 16'(-28866);
			520: out = 16'(-26682);
			521: out = 16'(-2734);
			522: out = 16'(9361);
			523: out = 16'(-3122);
			524: out = 16'(3174);
			525: out = 16'(14930);
			526: out = 16'(25218);
			527: out = 16'(-12218);
			528: out = 16'(-7976);
			529: out = 16'(4826);
			530: out = 16'(25348);
			531: out = 16'(2672);
			532: out = 16'(-6230);
			533: out = 16'(-10615);
			534: out = 16'(20066);
			535: out = 16'(-9232);
			536: out = 16'(-13470);
			537: out = 16'(28608);
			538: out = 16'(20535);
			539: out = 16'(14964);
			540: out = 16'(495);
			541: out = 16'(-7010);
			542: out = 16'(-8486);
			543: out = 16'(-3988);
			544: out = 16'(-6032);
			545: out = 16'(4052);
			546: out = 16'(6201);
			547: out = 16'(8241);
			548: out = 16'(4094);
			549: out = 16'(12408);
			550: out = 16'(17129);
			551: out = 16'(17955);
			552: out = 16'(-3744);
			553: out = 16'(-5455);
			554: out = 16'(4102);
			555: out = 16'(42);
			556: out = 16'(12077);
			557: out = 16'(12665);
			558: out = 16'(6751);
			559: out = 16'(-10514);
			560: out = 16'(-8647);
			561: out = 16'(6434);
			562: out = 16'(23561);
			563: out = 16'(13176);
			564: out = 16'(4890);
			565: out = 16'(8140);
			566: out = 16'(-1031);
			567: out = 16'(6332);
			568: out = 16'(13640);
			569: out = 16'(18006);
			570: out = 16'(1575);
			571: out = 16'(-898);
			572: out = 16'(17079);
			573: out = 16'(-15635);
			574: out = 16'(-2406);
			575: out = 16'(12248);
			576: out = 16'(331);
			577: out = 16'(8295);
			578: out = 16'(4143);
			579: out = 16'(-13044);
			580: out = 16'(-4560);
			581: out = 16'(-20023);
			582: out = 16'(-22814);
			583: out = 16'(7397);
			584: out = 16'(17999);
			585: out = 16'(15026);
			586: out = 16'(5424);
			587: out = 16'(-18054);
			588: out = 16'(-7671);
			589: out = 16'(5519);
			590: out = 16'(-7330);
			591: out = 16'(-3855);
			592: out = 16'(18);
			593: out = 16'(2705);
			594: out = 16'(-650);
			595: out = 16'(-18085);
			596: out = 16'(-21929);
			597: out = 16'(11662);
			598: out = 16'(18017);
			599: out = 16'(7732);
			600: out = 16'(-17755);
			601: out = 16'(-12227);
			602: out = 16'(-20751);
			603: out = 16'(-25393);
			604: out = 16'(-23343);
			605: out = 16'(-1374);
			606: out = 16'(18831);
			607: out = 16'(21906);
			608: out = 16'(23453);
			609: out = 16'(-10789);
			610: out = 16'(-27226);
			611: out = 16'(-2452);
			612: out = 16'(19537);
			613: out = 16'(12328);
			614: out = 16'(-11044);
			615: out = 16'(279);
			616: out = 16'(11578);
			617: out = 16'(18618);
			618: out = 16'(-1923);
			619: out = 16'(13629);
			620: out = 16'(611);
			621: out = 16'(-16581);
			622: out = 16'(-2622);
			623: out = 16'(1798);
			624: out = 16'(8556);
			625: out = 16'(10551);
			626: out = 16'(11044);
			627: out = 16'(2705);
			628: out = 16'(1718);
			629: out = 16'(16656);
			630: out = 16'(18554);
			631: out = 16'(2132);
			632: out = 16'(-22761);
			633: out = 16'(-25862);
			634: out = 16'(122);
			635: out = 16'(21182);
			636: out = 16'(8110);
			637: out = 16'(-14666);
			638: out = 16'(-21967);
			639: out = 16'(2736);
			640: out = 16'(-982);
			641: out = 16'(-8192);
			642: out = 16'(-19218);
			643: out = 16'(-24204);
			644: out = 16'(-8186);
			645: out = 16'(6136);
			646: out = 16'(10913);
			647: out = 16'(-10378);
			648: out = 16'(1469);
			649: out = 16'(14109);
			650: out = 16'(-25453);
			651: out = 16'(-26219);
			652: out = 16'(-11320);
			653: out = 16'(15891);
			654: out = 16'(6678);
			655: out = 16'(-7943);
			656: out = 16'(-23581);
			657: out = 16'(-5938);
			658: out = 16'(779);
			659: out = 16'(9809);
			660: out = 16'(9692);
			661: out = 16'(-12914);
			662: out = 16'(-21523);
			663: out = 16'(-15190);
			664: out = 16'(-10762);
			665: out = 16'(7253);
			666: out = 16'(15193);
			667: out = 16'(15549);
			668: out = 16'(13935);
			669: out = 16'(5765);
			670: out = 16'(-8039);
			671: out = 16'(-25348);
			672: out = 16'(-18389);
			673: out = 16'(-1458);
			674: out = 16'(8651);
			675: out = 16'(7511);
			676: out = 16'(1353);
			677: out = 16'(-4431);
			678: out = 16'(-23508);
			679: out = 16'(9787);
			680: out = 16'(13761);
			681: out = 16'(-10646);
			682: out = 16'(-17264);
			683: out = 16'(-17625);
			684: out = 16'(-2321);
			685: out = 16'(1854);
			686: out = 16'(14822);
			687: out = 16'(4441);
			688: out = 16'(-9321);
			689: out = 16'(8321);
			690: out = 16'(13474);
			691: out = 16'(9969);
			692: out = 16'(7118);
			693: out = 16'(-20523);
			694: out = 16'(-20575);
			695: out = 16'(6276);
			696: out = 16'(19165);
			697: out = 16'(19316);
			698: out = 16'(7505);
			699: out = 16'(-546);
			700: out = 16'(-19665);
			701: out = 16'(-20120);
			702: out = 16'(-4254);
			703: out = 16'(9821);
			704: out = 16'(18910);
			705: out = 16'(12070);
			706: out = 16'(-9693);
			707: out = 16'(-24634);
			708: out = 16'(-17847);
			709: out = 16'(11329);
			710: out = 16'(6114);
			711: out = 16'(23623);
			712: out = 16'(13725);
			713: out = 16'(-13533);
			714: out = 16'(-23919);
			715: out = 16'(-9551);
			716: out = 16'(12699);
			717: out = 16'(18610);
			718: out = 16'(12876);
			719: out = 16'(8686);
			720: out = 16'(4944);
			721: out = 16'(24042);
			722: out = 16'(7229);
			723: out = 16'(-19109);
			724: out = 16'(-28435);
			725: out = 16'(-1116);
			726: out = 16'(21919);
			727: out = 16'(15881);
			728: out = 16'(-9466);
			729: out = 16'(-16760);
			730: out = 16'(28);
			731: out = 16'(12719);
			732: out = 16'(3564);
			733: out = 16'(-13620);
			734: out = 16'(-16295);
			735: out = 16'(-6185);
			736: out = 16'(14413);
			737: out = 16'(16101);
			738: out = 16'(-21519);
			739: out = 16'(-29577);
			740: out = 16'(-22364);
			741: out = 16'(1153);
			742: out = 16'(13984);
			743: out = 16'(23263);
			744: out = 16'(14259);
			745: out = 16'(-18282);
			746: out = 16'(-27107);
			747: out = 16'(-11955);
			748: out = 16'(12463);
			749: out = 16'(6018);
			750: out = 16'(-5565);
			751: out = 16'(-7775);
			752: out = 16'(20148);
			753: out = 16'(8618);
			754: out = 16'(-8104);
			755: out = 16'(-21291);
			756: out = 16'(-13534);
			757: out = 16'(8549);
			758: out = 16'(17434);
			759: out = 16'(4434);
			760: out = 16'(-13370);
			761: out = 16'(-12143);
			762: out = 16'(10499);
			763: out = 16'(17903);
			764: out = 16'(15641);
			765: out = 16'(4099);
			766: out = 16'(-15948);
			767: out = 16'(6193);
			768: out = 16'(16850);
			769: out = 16'(12467);
			770: out = 16'(-13673);
			771: out = 16'(296);
			772: out = 16'(18247);
			773: out = 16'(2532);
			774: out = 16'(732);
			775: out = 16'(-11757);
			776: out = 16'(-15997);
			777: out = 16'(-204);
			778: out = 16'(10597);
			779: out = 16'(7854);
			780: out = 16'(-15860);
			781: out = 16'(-4137);
			782: out = 16'(-11385);
			783: out = 16'(-28755);
			784: out = 16'(-9148);
			785: out = 16'(2499);
			786: out = 16'(13694);
			787: out = 16'(19061);
			788: out = 16'(14979);
			789: out = 16'(9993);
			790: out = 16'(5434);
			791: out = 16'(-7056);
			792: out = 16'(-7923);
			793: out = 16'(-7876);
			794: out = 16'(-15983);
			795: out = 16'(13077);
			796: out = 16'(18090);
			797: out = 16'(7996);
			798: out = 16'(-3335);
			799: out = 16'(-1985);
			800: out = 16'(10569);
			801: out = 16'(22871);
			802: out = 16'(5805);
			803: out = 16'(-5342);
			804: out = 16'(-5949);
			805: out = 16'(11812);
			806: out = 16'(12542);
			807: out = 16'(4623);
			808: out = 16'(-10949);
			809: out = 16'(198);
			810: out = 16'(5498);
			811: out = 16'(9807);
			812: out = 16'(13609);
			813: out = 16'(14890);
			814: out = 16'(11256);
			815: out = 16'(7420);
			816: out = 16'(1400);
			817: out = 16'(4872);
			818: out = 16'(8508);
			819: out = 16'(11919);
			820: out = 16'(-1543);
			821: out = 16'(-562);
			822: out = 16'(17953);
			823: out = 16'(12866);
			824: out = 16'(166);
			825: out = 16'(-17470);
			826: out = 16'(1047);
			827: out = 16'(-2755);
			828: out = 16'(9358);
			829: out = 16'(19427);
			830: out = 16'(7050);
			831: out = 16'(-13801);
			832: out = 16'(-26106);
			833: out = 16'(-8796);
			834: out = 16'(10249);
			835: out = 16'(18612);
			836: out = 16'(14183);
			837: out = 16'(-13174);
			838: out = 16'(-13033);
			839: out = 16'(3142);
			840: out = 16'(233);
			841: out = 16'(14082);
			842: out = 16'(8977);
			843: out = 16'(-1986);
			844: out = 16'(1282);
			845: out = 16'(8408);
			846: out = 16'(6424);
			847: out = 16'(-25946);
			848: out = 16'(-20664);
			849: out = 16'(-9139);
			850: out = 16'(5966);
			851: out = 16'(-1768);
			852: out = 16'(9110);
			853: out = 16'(13868);
			854: out = 16'(3339);
			855: out = 16'(-11559);
			856: out = 16'(-16093);
			857: out = 16'(-1043);
			858: out = 16'(-19040);
			859: out = 16'(3096);
			860: out = 16'(17848);
			861: out = 16'(-1643);
			862: out = 16'(2346);
			863: out = 16'(-6092);
			864: out = 16'(-14584);
			865: out = 16'(-15161);
			866: out = 16'(-2763);
			867: out = 16'(7805);
			868: out = 16'(3647);
			869: out = 16'(9322);
			870: out = 16'(9637);
			871: out = 16'(8196);
			872: out = 16'(-8493);
			873: out = 16'(-10647);
			874: out = 16'(-8490);
			875: out = 16'(-2671);
			876: out = 16'(-7461);
			877: out = 16'(-5000);
			878: out = 16'(2245);
			879: out = 16'(1716);
			880: out = 16'(7102);
			881: out = 16'(4303);
			882: out = 16'(-18154);
			883: out = 16'(-7313);
			884: out = 16'(-2831);
			885: out = 16'(1555);
			886: out = 16'(-15554);
			887: out = 16'(2023);
			888: out = 16'(12055);
			889: out = 16'(6496);
			890: out = 16'(-17987);
			891: out = 16'(-21016);
			892: out = 16'(-772);
			893: out = 16'(8210);
			894: out = 16'(12380);
			895: out = 16'(8046);
			896: out = 16'(5311);
			897: out = 16'(-2268);
			898: out = 16'(-3901);
			899: out = 16'(-1733);
			900: out = 16'(-3370);
			901: out = 16'(2260);
			902: out = 16'(-2886);
			903: out = 16'(-19922);
			904: out = 16'(-538);
			905: out = 16'(15206);
			906: out = 16'(16593);
			907: out = 16'(2156);
			908: out = 16'(-19063);
			909: out = 16'(-22447);
			910: out = 16'(3327);
			911: out = 16'(15346);
			912: out = 16'(11876);
			913: out = 16'(-5791);
			914: out = 16'(-18674);
			915: out = 16'(-22128);
			916: out = 16'(-14857);
			917: out = 16'(-12278);
			918: out = 16'(7787);
			919: out = 16'(5530);
			920: out = 16'(-2086);
			921: out = 16'(-8449);
			922: out = 16'(-11618);
			923: out = 16'(-12491);
			924: out = 16'(-7150);
			925: out = 16'(-12059);
			926: out = 16'(-827);
			927: out = 16'(10940);
			928: out = 16'(15626);
			929: out = 16'(-2723);
			930: out = 16'(-19459);
			931: out = 16'(-24052);
			932: out = 16'(-2161);
			933: out = 16'(8622);
			934: out = 16'(3171);
			935: out = 16'(-22877);
			936: out = 16'(-13669);
			937: out = 16'(-2353);
			938: out = 16'(1527);
			939: out = 16'(18908);
			940: out = 16'(14538);
			941: out = 16'(9101);
			942: out = 16'(14913);
			943: out = 16'(-4408);
			944: out = 16'(-19628);
			945: out = 16'(-26228);
			946: out = 16'(5374);
			947: out = 16'(14462);
			948: out = 16'(11908);
			949: out = 16'(2168);
			950: out = 16'(7380);
			951: out = 16'(4695);
			952: out = 16'(-4087);
			953: out = 16'(-8160);
			954: out = 16'(-4591);
			955: out = 16'(270);
			956: out = 16'(-8428);
			957: out = 16'(7852);
			958: out = 16'(11191);
			959: out = 16'(6624);
			960: out = 16'(-78);
			961: out = 16'(-2224);
			962: out = 16'(1563);
			963: out = 16'(10507);
			964: out = 16'(291);
			965: out = 16'(8680);
			966: out = 16'(26090);
			967: out = 16'(-16376);
			968: out = 16'(3856);
			969: out = 16'(12469);
			970: out = 16'(852);
			971: out = 16'(-4407);
			972: out = 16'(3487);
			973: out = 16'(14742);
			974: out = 16'(13798);
			975: out = 16'(720);
			976: out = 16'(-5809);
			977: out = 16'(3380);
			978: out = 16'(10034);
			979: out = 16'(5173);
			980: out = 16'(-7462);
			981: out = 16'(-21981);
			982: out = 16'(-6281);
			983: out = 16'(11294);
			984: out = 16'(10593);
			985: out = 16'(3070);
			986: out = 16'(-2963);
			987: out = 16'(-599);
			988: out = 16'(10347);
			989: out = 16'(-2279);
			990: out = 16'(-4264);
			991: out = 16'(18076);
			992: out = 16'(1636);
			993: out = 16'(-5240);
			994: out = 16'(-12279);
			995: out = 16'(28794);
			996: out = 16'(-12425);
			997: out = 16'(-22953);
			998: out = 16'(8080);
			999: out = 16'(17832);
			1000: out = 16'(17711);
			1001: out = 16'(5487);
			1002: out = 16'(-17147);
			1003: out = 16'(-10529);
			1004: out = 16'(-591);
			1005: out = 16'(-1027);
			1006: out = 16'(-10913);
			1007: out = 16'(-16845);
			1008: out = 16'(-11126);
			1009: out = 16'(4985);
			1010: out = 16'(6175);
			1011: out = 16'(15);
			1012: out = 16'(-10699);
			1013: out = 16'(-11211);
			1014: out = 16'(-11621);
			1015: out = 16'(-6243);
			1016: out = 16'(-370);
			1017: out = 16'(10063);
			1018: out = 16'(10129);
			1019: out = 16'(6631);
			1020: out = 16'(-9759);
			1021: out = 16'(1970);
			1022: out = 16'(8711);
			1023: out = 16'(-27507);
			1024: out = 16'(-17276);
			1025: out = 16'(-609);
			1026: out = 16'(17551);
			1027: out = 16'(14575);
			1028: out = 16'(7835);
			1029: out = 16'(-5310);
			1030: out = 16'(-9783);
			1031: out = 16'(-4162);
			1032: out = 16'(8501);
			1033: out = 16'(10088);
			1034: out = 16'(15394);
			1035: out = 16'(447);
			1036: out = 16'(-7818);
			1037: out = 16'(-12965);
			1038: out = 16'(12991);
			1039: out = 16'(11646);
			1040: out = 16'(-4769);
			1041: out = 16'(-17216);
			1042: out = 16'(-2760);
			1043: out = 16'(14016);
			1044: out = 16'(10754);
			1045: out = 16'(-7441);
			1046: out = 16'(-10055);
			1047: out = 16'(8654);
			1048: out = 16'(-13031);
			1049: out = 16'(-1577);
			1050: out = 16'(4120);
			1051: out = 16'(-89);
			1052: out = 16'(-3277);
			1053: out = 16'(-10125);
			1054: out = 16'(-15554);
			1055: out = 16'(-2603);
			1056: out = 16'(4601);
			1057: out = 16'(7527);
			1058: out = 16'(5001);
			1059: out = 16'(12);
			1060: out = 16'(223);
			1061: out = 16'(5330);
			1062: out = 16'(4426);
			1063: out = 16'(6099);
			1064: out = 16'(5356);
			1065: out = 16'(4943);
			1066: out = 16'(3668);
			1067: out = 16'(4869);
			1068: out = 16'(5947);
			1069: out = 16'(-3479);
			1070: out = 16'(7990);
			1071: out = 16'(15840);
			1072: out = 16'(9005);
			1073: out = 16'(2350);
			1074: out = 16'(-6043);
			1075: out = 16'(-5324);
			1076: out = 16'(-16948);
			1077: out = 16'(7190);
			1078: out = 16'(12947);
			1079: out = 16'(-5379);
			1080: out = 16'(41);
			1081: out = 16'(10039);
			1082: out = 16'(17998);
			1083: out = 16'(-8036);
			1084: out = 16'(-6585);
			1085: out = 16'(-4672);
			1086: out = 16'(2158);
			1087: out = 16'(-10612);
			1088: out = 16'(-9521);
			1089: out = 16'(-1697);
			1090: out = 16'(10088);
			1091: out = 16'(3948);
			1092: out = 16'(3658);
			1093: out = 16'(17624);
			1094: out = 16'(-11638);
			1095: out = 16'(-656);
			1096: out = 16'(16616);
			1097: out = 16'(11408);
			1098: out = 16'(4657);
			1099: out = 16'(1012);
			1100: out = 16'(12427);
			1101: out = 16'(-15722);
			1102: out = 16'(-9957);
			1103: out = 16'(5309);
			1104: out = 16'(21885);
			1105: out = 16'(543);
			1106: out = 16'(-14124);
			1107: out = 16'(-11153);
			1108: out = 16'(7812);
			1109: out = 16'(18081);
			1110: out = 16'(14257);
			1111: out = 16'(5170);
			1112: out = 16'(-9350);
			1113: out = 16'(-16437);
			1114: out = 16'(-13914);
			1115: out = 16'(1195);
			1116: out = 16'(8948);
			1117: out = 16'(8505);
			1118: out = 16'(-3104);
			1119: out = 16'(-4214);
			1120: out = 16'(-9319);
			1121: out = 16'(-12702);
			1122: out = 16'(1741);
			1123: out = 16'(8975);
			1124: out = 16'(8475);
			1125: out = 16'(6535);
			1126: out = 16'(-12425);
			1127: out = 16'(-8216);
			1128: out = 16'(15457);
			1129: out = 16'(-16410);
			1130: out = 16'(-7324);
			1131: out = 16'(-2116);
			1132: out = 16'(-12288);
			1133: out = 16'(-5028);
			1134: out = 16'(4188);
			1135: out = 16'(9002);
			1136: out = 16'(4077);
			1137: out = 16'(-11483);
			1138: out = 16'(-21604);
			1139: out = 16'(-933);
			1140: out = 16'(-12805);
			1141: out = 16'(-624);
			1142: out = 16'(16169);
			1143: out = 16'(-8049);
			1144: out = 16'(-12472);
			1145: out = 16'(-14638);
			1146: out = 16'(-7056);
			1147: out = 16'(-3438);
			1148: out = 16'(3135);
			1149: out = 16'(3382);
			1150: out = 16'(13811);
			1151: out = 16'(-1127);
			1152: out = 16'(-4139);
			1153: out = 16'(8268);
			1154: out = 16'(14558);
			1155: out = 16'(-3280);
			1156: out = 16'(-30596);
			1157: out = 16'(-13482);
			1158: out = 16'(-4306);
			1159: out = 16'(2818);
			1160: out = 16'(-4450);
			1161: out = 16'(12396);
			1162: out = 16'(17147);
			1163: out = 16'(15359);
			1164: out = 16'(-23782);
			1165: out = 16'(-10070);
			1166: out = 16'(8249);
			1167: out = 16'(12161);
			1168: out = 16'(7297);
			1169: out = 16'(-2565);
			1170: out = 16'(-7933);
			1171: out = 16'(-2160);
			1172: out = 16'(5528);
			1173: out = 16'(7434);
			1174: out = 16'(-765);
			1175: out = 16'(10999);
			1176: out = 16'(7811);
			1177: out = 16'(3966);
			1178: out = 16'(7949);
			1179: out = 16'(9425);
			1180: out = 16'(4353);
			1181: out = 16'(-10286);
			1182: out = 16'(5257);
			1183: out = 16'(-1500);
			1184: out = 16'(-13603);
			1185: out = 16'(-8474);
			1186: out = 16'(-8606);
			1187: out = 16'(1317);
			1188: out = 16'(9119);
			1189: out = 16'(6261);
			1190: out = 16'(-8252);
			1191: out = 16'(-20247);
			1192: out = 16'(-12752);
			1193: out = 16'(-2624);
			1194: out = 16'(9199);
			1195: out = 16'(17105);
			1196: out = 16'(-3826);
			1197: out = 16'(-2897);
			1198: out = 16'(4240);
			1199: out = 16'(14531);
			1200: out = 16'(-9639);
			1201: out = 16'(-15384);
			1202: out = 16'(7118);
			1203: out = 16'(-7814);
			1204: out = 16'(6325);
			1205: out = 16'(13736);
			1206: out = 16'(5798);
			1207: out = 16'(1793);
			1208: out = 16'(-6527);
			1209: out = 16'(-14285);
			1210: out = 16'(-6249);
			1211: out = 16'(2020);
			1212: out = 16'(7604);
			1213: out = 16'(3261);
			1214: out = 16'(4375);
			1215: out = 16'(-372);
			1216: out = 16'(-5032);
			1217: out = 16'(-2363);
			1218: out = 16'(258);
			1219: out = 16'(181);
			1220: out = 16'(-3687);
			1221: out = 16'(-311);
			1222: out = 16'(6884);
			1223: out = 16'(13986);
			1224: out = 16'(6999);
			1225: out = 16'(5624);
			1226: out = 16'(-355);
			1227: out = 16'(-13111);
			1228: out = 16'(2477);
			1229: out = 16'(11970);
			1230: out = 16'(10097);
			1231: out = 16'(-3527);
			1232: out = 16'(-2771);
			1233: out = 16'(7753);
			1234: out = 16'(11419);
			1235: out = 16'(10606);
			1236: out = 16'(-8846);
			1237: out = 16'(-26719);
			1238: out = 16'(-13434);
			1239: out = 16'(7148);
			1240: out = 16'(16536);
			1241: out = 16'(13235);
			1242: out = 16'(-9618);
			1243: out = 16'(-11618);
			1244: out = 16'(3661);
			1245: out = 16'(12020);
			1246: out = 16'(5426);
			1247: out = 16'(-2543);
			1248: out = 16'(2717);
			1249: out = 16'(10311);
			1250: out = 16'(8095);
			1251: out = 16'(-3914);
			1252: out = 16'(15681);
			1253: out = 16'(-10345);
			1254: out = 16'(-17756);
			1255: out = 16'(3261);
			1256: out = 16'(-1925);
			1257: out = 16'(2008);
			1258: out = 16'(4400);
			1259: out = 16'(10964);
			1260: out = 16'(-3828);
			1261: out = 16'(-11892);
			1262: out = 16'(-3031);
			1263: out = 16'(-9366);
			1264: out = 16'(-6092);
			1265: out = 16'(-2311);
			1266: out = 16'(15505);
			1267: out = 16'(-4358);
			1268: out = 16'(-14919);
			1269: out = 16'(-10748);
			1270: out = 16'(-9838);
			1271: out = 16'(-8190);
			1272: out = 16'(-3520);
			1273: out = 16'(9302);
			1274: out = 16'(12283);
			1275: out = 16'(2429);
			1276: out = 16'(-18318);
			1277: out = 16'(-19437);
			1278: out = 16'(-4470);
			1279: out = 16'(11441);
			1280: out = 16'(-18702);
			1281: out = 16'(-1820);
			1282: out = 16'(6342);
			1283: out = 16'(15664);
			1284: out = 16'(-16696);
			1285: out = 16'(-3379);
			1286: out = 16'(14828);
			1287: out = 16'(12316);
			1288: out = 16'(-4890);
			1289: out = 16'(-16681);
			1290: out = 16'(-9918);
			1291: out = 16'(4833);
			1292: out = 16'(8201);
			1293: out = 16'(2592);
			1294: out = 16'(7466);
			1295: out = 16'(-2360);
			1296: out = 16'(2033);
			1297: out = 16'(12979);
			1298: out = 16'(5861);
			1299: out = 16'(8695);
			1300: out = 16'(8878);
			1301: out = 16'(2328);
			1302: out = 16'(4061);
			1303: out = 16'(6475);
			1304: out = 16'(7785);
			1305: out = 16'(3915);
			1306: out = 16'(-3672);
			1307: out = 16'(-7677);
			1308: out = 16'(2438);
			1309: out = 16'(7707);
			1310: out = 16'(13027);
			1311: out = 16'(11038);
			1312: out = 16'(8454);
			1313: out = 16'(-705);
			1314: out = 16'(-7250);
			1315: out = 16'(-14628);
			1316: out = 16'(4787);
			1317: out = 16'(12134);
			1318: out = 16'(7372);
			1319: out = 16'(-10678);
			1320: out = 16'(-14251);
			1321: out = 16'(-7198);
			1322: out = 16'(7047);
			1323: out = 16'(-1185);
			1324: out = 16'(879);
			1325: out = 16'(8848);
			1326: out = 16'(3506);
			1327: out = 16'(3571);
			1328: out = 16'(1356);
			1329: out = 16'(775);
			1330: out = 16'(-798);
			1331: out = 16'(2397);
			1332: out = 16'(6074);
			1333: out = 16'(1426);
			1334: out = 16'(-3786);
			1335: out = 16'(-8080);
			1336: out = 16'(1530);
			1337: out = 16'(-12508);
			1338: out = 16'(-3340);
			1339: out = 16'(10459);
			1340: out = 16'(8817);
			1341: out = 16'(-1324);
			1342: out = 16'(-9959);
			1343: out = 16'(-9170);
			1344: out = 16'(-1360);
			1345: out = 16'(-773);
			1346: out = 16'(-6233);
			1347: out = 16'(-13349);
			1348: out = 16'(-2271);
			1349: out = 16'(9018);
			1350: out = 16'(9201);
			1351: out = 16'(-4234);
			1352: out = 16'(-8288);
			1353: out = 16'(-1238);
			1354: out = 16'(-4045);
			1355: out = 16'(4810);
			1356: out = 16'(5502);
			1357: out = 16'(2793);
			1358: out = 16'(-571);
			1359: out = 16'(598);
			1360: out = 16'(1857);
			1361: out = 16'(112);
			1362: out = 16'(1510);
			1363: out = 16'(3876);
			1364: out = 16'(4712);
			1365: out = 16'(9210);
			1366: out = 16'(7076);
			1367: out = 16'(860);
			1368: out = 16'(-21681);
			1369: out = 16'(-9416);
			1370: out = 16'(4355);
			1371: out = 16'(10361);
			1372: out = 16'(-320);
			1373: out = 16'(-805);
			1374: out = 16'(2639);
			1375: out = 16'(2879);
			1376: out = 16'(5516);
			1377: out = 16'(7859);
			1378: out = 16'(8313);
			1379: out = 16'(5400);
			1380: out = 16'(-1015);
			1381: out = 16'(-3563);
			1382: out = 16'(1742);
			1383: out = 16'(1139);
			1384: out = 16'(-1776);
			1385: out = 16'(-2592);
			1386: out = 16'(-24265);
			1387: out = 16'(-10760);
			1388: out = 16'(10015);
			1389: out = 16'(12066);
			1390: out = 16'(488);
			1391: out = 16'(-8067);
			1392: out = 16'(-3062);
			1393: out = 16'(-6752);
			1394: out = 16'(-4563);
			1395: out = 16'(-3230);
			1396: out = 16'(14206);
			1397: out = 16'(-13013);
			1398: out = 16'(-13926);
			1399: out = 16'(6968);
			1400: out = 16'(-2999);
			1401: out = 16'(9966);
			1402: out = 16'(8177);
			1403: out = 16'(-22105);
			1404: out = 16'(-9229);
			1405: out = 16'(-2786);
			1406: out = 16'(-2977);
			1407: out = 16'(4730);
			1408: out = 16'(3899);
			1409: out = 16'(1085);
			1410: out = 16'(-14008);
			1411: out = 16'(10600);
			1412: out = 16'(10332);
			1413: out = 16'(-3522);
			1414: out = 16'(-19195);
			1415: out = 16'(-16286);
			1416: out = 16'(-318);
			1417: out = 16'(13454);
			1418: out = 16'(4173);
			1419: out = 16'(-3253);
			1420: out = 16'(-5848);
			1421: out = 16'(-325);
			1422: out = 16'(-2991);
			1423: out = 16'(-5782);
			1424: out = 16'(-4598);
			1425: out = 16'(1899);
			1426: out = 16'(2552);
			1427: out = 16'(-1398);
			1428: out = 16'(2642);
			1429: out = 16'(359);
			1430: out = 16'(485);
			1431: out = 16'(777);
			1432: out = 16'(3870);
			1433: out = 16'(2990);
			1434: out = 16'(2368);
			1435: out = 16'(11575);
			1436: out = 16'(3045);
			1437: out = 16'(-1311);
			1438: out = 16'(4797);
			1439: out = 16'(-5186);
			1440: out = 16'(138);
			1441: out = 16'(7156);
			1442: out = 16'(2246);
			1443: out = 16'(2901);
			1444: out = 16'(-209);
			1445: out = 16'(-4776);
			1446: out = 16'(1781);
			1447: out = 16'(2391);
			1448: out = 16'(1739);
			1449: out = 16'(10903);
			1450: out = 16'(926);
			1451: out = 16'(-6095);
			1452: out = 16'(-9018);
			1453: out = 16'(3117);
			1454: out = 16'(1417);
			1455: out = 16'(-4137);
			1456: out = 16'(7469);
			1457: out = 16'(-4013);
			1458: out = 16'(-7768);
			1459: out = 16'(-5457);
			1460: out = 16'(7072);
			1461: out = 16'(7283);
			1462: out = 16'(3832);
			1463: out = 16'(3478);
			1464: out = 16'(152);
			1465: out = 16'(-4591);
			1466: out = 16'(-9077);
			1467: out = 16'(-1932);
			1468: out = 16'(3087);
			1469: out = 16'(4199);
			1470: out = 16'(1154);
			1471: out = 16'(-2346);
			1472: out = 16'(-870);
			1473: out = 16'(3679);
			1474: out = 16'(512);
			1475: out = 16'(-999);
			1476: out = 16'(-535);
			1477: out = 16'(2508);
			1478: out = 16'(4293);
			1479: out = 16'(5338);
			1480: out = 16'(7723);
			1481: out = 16'(-4446);
			1482: out = 16'(5216);
			1483: out = 16'(9480);
			1484: out = 16'(-7015);
			1485: out = 16'(-2235);
			1486: out = 16'(658);
			1487: out = 16'(2403);
			1488: out = 16'(9954);
			1489: out = 16'(-2933);
			1490: out = 16'(-13230);
			1491: out = 16'(-928);
			1492: out = 16'(3519);
			1493: out = 16'(7711);
			1494: out = 16'(2278);
			1495: out = 16'(-4687);
			1496: out = 16'(-7208);
			1497: out = 16'(-2032);
			1498: out = 16'(-4808);
			1499: out = 16'(13367);
			1500: out = 16'(10820);
			1501: out = 16'(2174);
			1502: out = 16'(-20460);
			1503: out = 16'(-13635);
			1504: out = 16'(-656);
			1505: out = 16'(9684);
			1506: out = 16'(-6196);
			1507: out = 16'(-3180);
			1508: out = 16'(8992);
			1509: out = 16'(4750);
			1510: out = 16'(-3749);
			1511: out = 16'(-11960);
			1512: out = 16'(-8841);
			1513: out = 16'(4032);
			1514: out = 16'(10549);
			1515: out = 16'(7673);
			1516: out = 16'(-7603);
			1517: out = 16'(-216);
			1518: out = 16'(2952);
			1519: out = 16'(-12703);
			1520: out = 16'(-6535);
			1521: out = 16'(-2240);
			1522: out = 16'(6455);
			1523: out = 16'(9290);
			1524: out = 16'(7074);
			1525: out = 16'(-1635);
			1526: out = 16'(-7510);
			1527: out = 16'(-8080);
			1528: out = 16'(426);
			1529: out = 16'(6165);
			1530: out = 16'(384);
			1531: out = 16'(-3482);
			1532: out = 16'(-1598);
			1533: out = 16'(8434);
			1534: out = 16'(5953);
			1535: out = 16'(1820);
			1536: out = 16'(-7801);
			1537: out = 16'(-10647);
			1538: out = 16'(-14414);
			1539: out = 16'(-5578);
			1540: out = 16'(5378);
			1541: out = 16'(8848);
			1542: out = 16'(-2051);
			1543: out = 16'(-11151);
			1544: out = 16'(-426);
			1545: out = 16'(7616);
			1546: out = 16'(6780);
			1547: out = 16'(-4801);
			1548: out = 16'(-3920);
			1549: out = 16'(-427);
			1550: out = 16'(4899);
			1551: out = 16'(1508);
			1552: out = 16'(-1465);
			1553: out = 16'(-2447);
			1554: out = 16'(3417);
			1555: out = 16'(-7605);
			1556: out = 16'(-8207);
			1557: out = 16'(-6314);
			1558: out = 16'(-1434);
			1559: out = 16'(4380);
			1560: out = 16'(5974);
			1561: out = 16'(-353);
			1562: out = 16'(6722);
			1563: out = 16'(2263);
			1564: out = 16'(1640);
			1565: out = 16'(3232);
			1566: out = 16'(8837);
			1567: out = 16'(4215);
			1568: out = 16'(-3834);
			1569: out = 16'(1427);
			1570: out = 16'(5236);
			1571: out = 16'(5497);
			1572: out = 16'(8751);
			1573: out = 16'(-6237);
			1574: out = 16'(-1798);
			1575: out = 16'(12297);
			1576: out = 16'(-491);
			1577: out = 16'(-9856);
			1578: out = 16'(-13213);
			1579: out = 16'(1580);
			1580: out = 16'(8485);
			1581: out = 16'(6847);
			1582: out = 16'(-3413);
			1583: out = 16'(-20486);
			1584: out = 16'(-9235);
			1585: out = 16'(10630);
			1586: out = 16'(6333);
			1587: out = 16'(10347);
			1588: out = 16'(-1400);
			1589: out = 16'(-9011);
			1590: out = 16'(-7748);
			1591: out = 16'(6010);
			1592: out = 16'(12383);
			1593: out = 16'(8226);
			1594: out = 16'(-5654);
			1595: out = 16'(-14201);
			1596: out = 16'(-12372);
			1597: out = 16'(6013);
			1598: out = 16'(10120);
			1599: out = 16'(9222);
			1600: out = 16'(4896);
			1601: out = 16'(3262);
			1602: out = 16'(-6358);
			1603: out = 16'(-15949);
			1604: out = 16'(-2911);
			1605: out = 16'(5667);
			1606: out = 16'(9955);
			1607: out = 16'(4274);
			1608: out = 16'(-3303);
			1609: out = 16'(-12366);
			1610: out = 16'(-13467);
			1611: out = 16'(5013);
			1612: out = 16'(1555);
			1613: out = 16'(-4542);
			1614: out = 16'(-1401);
			1615: out = 16'(-13464);
			1616: out = 16'(-8915);
			1617: out = 16'(563);
			1618: out = 16'(5615);
			1619: out = 16'(-470);
			1620: out = 16'(-5356);
			1621: out = 16'(-1822);
			1622: out = 16'(1809);
			1623: out = 16'(5151);
			1624: out = 16'(3264);
			1625: out = 16'(72);
			1626: out = 16'(-4822);
			1627: out = 16'(-315);
			1628: out = 16'(12531);
			1629: out = 16'(-9286);
			1630: out = 16'(-15094);
			1631: out = 16'(-10418);
			1632: out = 16'(5618);
			1633: out = 16'(3433);
			1634: out = 16'(-1586);
			1635: out = 16'(-5642);
			1636: out = 16'(-3237);
			1637: out = 16'(-474);
			1638: out = 16'(1036);
			1639: out = 16'(-1945);
			1640: out = 16'(2206);
			1641: out = 16'(4913);
			1642: out = 16'(5194);
			1643: out = 16'(1035);
			1644: out = 16'(-1496);
			1645: out = 16'(-3240);
			1646: out = 16'(-4610);
			1647: out = 16'(-1775);
			1648: out = 16'(4325);
			1649: out = 16'(9120);
			1650: out = 16'(-2152);
			1651: out = 16'(-8145);
			1652: out = 16'(-7661);
			1653: out = 16'(4072);
			1654: out = 16'(3447);
			1655: out = 16'(3320);
			1656: out = 16'(4849);
			1657: out = 16'(5112);
			1658: out = 16'(8040);
			1659: out = 16'(4208);
			1660: out = 16'(-14606);
			1661: out = 16'(-9043);
			1662: out = 16'(-141);
			1663: out = 16'(6924);
			1664: out = 16'(5858);
			1665: out = 16'(5547);
			1666: out = 16'(5072);
			1667: out = 16'(591);
			1668: out = 16'(3655);
			1669: out = 16'(4812);
			1670: out = 16'(7559);
			1671: out = 16'(-17787);
			1672: out = 16'(-8441);
			1673: out = 16'(4252);
			1674: out = 16'(9835);
			1675: out = 16'(-9194);
			1676: out = 16'(-16430);
			1677: out = 16'(-9473);
			1678: out = 16'(9096);
			1679: out = 16'(288);
			1680: out = 16'(-7591);
			1681: out = 16'(6763);
			1682: out = 16'(3928);
			1683: out = 16'(2968);
			1684: out = 16'(-3247);
			1685: out = 16'(-1069);
			1686: out = 16'(524);
			1687: out = 16'(5888);
			1688: out = 16'(6752);
			1689: out = 16'(3290);
			1690: out = 16'(-3442);
			1691: out = 16'(-5913);
			1692: out = 16'(-3579);
			1693: out = 16'(4611);
			1694: out = 16'(8429);
			1695: out = 16'(5179);
			1696: out = 16'(1064);
			1697: out = 16'(-4418);
			1698: out = 16'(-7393);
			1699: out = 16'(-5182);
			1700: out = 16'(594);
			1701: out = 16'(5595);
			1702: out = 16'(4702);
			1703: out = 16'(8216);
			1704: out = 16'(-384);
			1705: out = 16'(-11666);
			1706: out = 16'(-8926);
			1707: out = 16'(-5222);
			1708: out = 16'(2906);
			1709: out = 16'(6590);
			1710: out = 16'(8821);
			1711: out = 16'(3265);
			1712: out = 16'(-969);
			1713: out = 16'(-463);
			1714: out = 16'(4691);
			1715: out = 16'(4175);
			1716: out = 16'(-2982);
			1717: out = 16'(-4535);
			1718: out = 16'(-2206);
			1719: out = 16'(984);
			1720: out = 16'(-10685);
			1721: out = 16'(605);
			1722: out = 16'(9219);
			1723: out = 16'(9313);
			1724: out = 16'(6372);
			1725: out = 16'(-6074);
			1726: out = 16'(-12911);
			1727: out = 16'(9553);
			1728: out = 16'(3510);
			1729: out = 16'(-3536);
			1730: out = 16'(-12923);
			1731: out = 16'(5046);
			1732: out = 16'(8688);
			1733: out = 16'(7185);
			1734: out = 16'(1644);
			1735: out = 16'(1097);
			1736: out = 16'(1985);
			1737: out = 16'(5556);
			1738: out = 16'(-7401);
			1739: out = 16'(-5188);
			1740: out = 16'(-348);
			1741: out = 16'(3078);
			1742: out = 16'(-5203);
			1743: out = 16'(-5649);
			1744: out = 16'(4290);
			1745: out = 16'(5652);
			1746: out = 16'(6423);
			1747: out = 16'(3802);
			1748: out = 16'(9152);
			1749: out = 16'(-1474);
			1750: out = 16'(732);
			1751: out = 16'(10048);
			1752: out = 16'(-1433);
			1753: out = 16'(1072);
			1754: out = 16'(934);
			1755: out = 16'(-11351);
			1756: out = 16'(-2304);
			1757: out = 16'(1370);
			1758: out = 16'(-636);
			1759: out = 16'(-1721);
			1760: out = 16'(-5447);
			1761: out = 16'(-4862);
			1762: out = 16'(4274);
			1763: out = 16'(-259);
			1764: out = 16'(338);
			1765: out = 16'(4033);
			1766: out = 16'(-1955);
			1767: out = 16'(-791);
			1768: out = 16'(-1705);
			1769: out = 16'(-5651);
			1770: out = 16'(2161);
			1771: out = 16'(8608);
			1772: out = 16'(8416);
			1773: out = 16'(1574);
			1774: out = 16'(-8177);
			1775: out = 16'(-9613);
			1776: out = 16'(3346);
			1777: out = 16'(693);
			1778: out = 16'(-967);
			1779: out = 16'(-2262);
			1780: out = 16'(-216);
			1781: out = 16'(1942);
			1782: out = 16'(1989);
			1783: out = 16'(390);
			1784: out = 16'(-368);
			1785: out = 16'(2320);
			1786: out = 16'(4066);
			1787: out = 16'(1135);
			1788: out = 16'(-2913);
			1789: out = 16'(-2667);
			1790: out = 16'(328);
			1791: out = 16'(9451);
			1792: out = 16'(501);
			1793: out = 16'(-14184);
			1794: out = 16'(530);
			1795: out = 16'(3476);
			1796: out = 16'(2416);
			1797: out = 16'(-13718);
			1798: out = 16'(1291);
			1799: out = 16'(666);
			1800: out = 16'(-1112);
			1801: out = 16'(3090);
			1802: out = 16'(6749);
			1803: out = 16'(692);
			1804: out = 16'(-19576);
			1805: out = 16'(-5732);
			1806: out = 16'(-909);
			1807: out = 16'(2946);
			1808: out = 16'(9768);
			1809: out = 16'(6924);
			1810: out = 16'(-271);
			1811: out = 16'(-8045);
			1812: out = 16'(-8517);
			1813: out = 16'(-2216);
			1814: out = 16'(4051);
			1815: out = 16'(104);
			1816: out = 16'(-2475);
			1817: out = 16'(-6075);
			1818: out = 16'(-5221);
			1819: out = 16'(-2072);
			1820: out = 16'(1206);
			1821: out = 16'(-819);
			1822: out = 16'(-4941);
			1823: out = 16'(-7081);
			1824: out = 16'(-53);
			1825: out = 16'(9686);
			1826: out = 16'(1942);
			1827: out = 16'(496);
			1828: out = 16'(388);
			1829: out = 16'(-13916);
			1830: out = 16'(3699);
			1831: out = 16'(9627);
			1832: out = 16'(6749);
			1833: out = 16'(-7490);
			1834: out = 16'(-4636);
			1835: out = 16'(1260);
			1836: out = 16'(2931);
			1837: out = 16'(-3376);
			1838: out = 16'(515);
			1839: out = 16'(8644);
			1840: out = 16'(3246);
			1841: out = 16'(-12001);
			1842: out = 16'(-18894);
			1843: out = 16'(7371);
			1844: out = 16'(8885);
			1845: out = 16'(2683);
			1846: out = 16'(-12663);
			1847: out = 16'(-8071);
			1848: out = 16'(-3450);
			1849: out = 16'(4564);
			1850: out = 16'(8289);
			1851: out = 16'(2057);
			1852: out = 16'(410);
			1853: out = 16'(5616);
			1854: out = 16'(8356);
			1855: out = 16'(5842);
			1856: out = 16'(-31);
			1857: out = 16'(-3404);
			1858: out = 16'(-646);
			1859: out = 16'(1302);
			1860: out = 16'(130);
			1861: out = 16'(-2840);
			1862: out = 16'(-124);
			1863: out = 16'(3612);
			1864: out = 16'(4506);
			1865: out = 16'(-4141);
			1866: out = 16'(-2816);
			1867: out = 16'(6490);
			1868: out = 16'(-16685);
			1869: out = 16'(-1689);
			1870: out = 16'(8612);
			1871: out = 16'(5104);
			1872: out = 16'(-2629);
			1873: out = 16'(-6933);
			1874: out = 16'(-2710);
			1875: out = 16'(3667);
			1876: out = 16'(6364);
			1877: out = 16'(2272);
			1878: out = 16'(-3379);
			1879: out = 16'(-1915);
			1880: out = 16'(3274);
			1881: out = 16'(5631);
			1882: out = 16'(3394);
			1883: out = 16'(-2958);
			1884: out = 16'(-2428);
			1885: out = 16'(7027);
			1886: out = 16'(-576);
			1887: out = 16'(-5158);
			1888: out = 16'(-6684);
			1889: out = 16'(3677);
			1890: out = 16'(5119);
			1891: out = 16'(4672);
			1892: out = 16'(1701);
			1893: out = 16'(2457);
			1894: out = 16'(-999);
			1895: out = 16'(-4352);
			1896: out = 16'(4350);
			1897: out = 16'(121);
			1898: out = 16'(1903);
			1899: out = 16'(5200);
			1900: out = 16'(4097);
			1901: out = 16'(-8024);
			1902: out = 16'(-17752);
			1903: out = 16'(396);
			1904: out = 16'(6745);
			1905: out = 16'(11160);
			1906: out = 16'(7738);
			1907: out = 16'(3252);
			1908: out = 16'(-2693);
			1909: out = 16'(-4556);
			1910: out = 16'(-4901);
			1911: out = 16'(901);
			1912: out = 16'(3451);
			1913: out = 16'(2523);
			1914: out = 16'(2130);
			1915: out = 16'(1077);
			1916: out = 16'(565);
			1917: out = 16'(-606);
			1918: out = 16'(-865);
			1919: out = 16'(-554);
			1920: out = 16'(1888);
			1921: out = 16'(1982);
			1922: out = 16'(4794);
			1923: out = 16'(5292);
			1924: out = 16'(5935);
			1925: out = 16'(-1447);
			1926: out = 16'(-778);
			1927: out = 16'(5850);
			1928: out = 16'(4593);
			1929: out = 16'(2970);
			1930: out = 16'(1126);
			1931: out = 16'(4154);
			1932: out = 16'(3951);
			1933: out = 16'(2789);
			1934: out = 16'(-681);
			1935: out = 16'(118);
			1936: out = 16'(1304);
			1937: out = 16'(2087);
			1938: out = 16'(-5101);
			1939: out = 16'(-2608);
			1940: out = 16'(-3788);
			1941: out = 16'(-2310);
			1942: out = 16'(115);
			1943: out = 16'(7431);
			1944: out = 16'(5333);
			1945: out = 16'(-10126);
			1946: out = 16'(-13862);
			1947: out = 16'(-8008);
			1948: out = 16'(5650);
			1949: out = 16'(4659);
			1950: out = 16'(6916);
			1951: out = 16'(4309);
			1952: out = 16'(3326);
			1953: out = 16'(-4828);
			1954: out = 16'(-6612);
			1955: out = 16'(-5071);
			1956: out = 16'(-578);
			1957: out = 16'(1716);
			1958: out = 16'(3769);
			1959: out = 16'(2775);
			1960: out = 16'(2711);
			1961: out = 16'(-1625);
			1962: out = 16'(-4397);
			1963: out = 16'(-5655);
			1964: out = 16'(375);
			1965: out = 16'(1482);
			1966: out = 16'(-3269);
			1967: out = 16'(-8585);
			1968: out = 16'(-4118);
			1969: out = 16'(4459);
			1970: out = 16'(1103);
			1971: out = 16'(-1462);
			1972: out = 16'(-3001);
			1973: out = 16'(2256);
			1974: out = 16'(2197);
			1975: out = 16'(2399);
			1976: out = 16'(221);
			1977: out = 16'(608);
			1978: out = 16'(-3058);
			1979: out = 16'(-6044);
			1980: out = 16'(-7564);
			1981: out = 16'(-1772);
			1982: out = 16'(2247);
			1983: out = 16'(3142);
			1984: out = 16'(8118);
			1985: out = 16'(554);
			1986: out = 16'(117);
			1987: out = 16'(7009);
			1988: out = 16'(4734);
			1989: out = 16'(367);
			1990: out = 16'(-5363);
			1991: out = 16'(-12022);
			1992: out = 16'(-1876);
			1993: out = 16'(5461);
			1994: out = 16'(2471);
			1995: out = 16'(3275);
			1996: out = 16'(-588);
			1997: out = 16'(-2355);
			1998: out = 16'(356);
			1999: out = 16'(-2545);
			2000: out = 16'(-2437);
			2001: out = 16'(2051);
			2002: out = 16'(-560);
			2003: out = 16'(2697);
			2004: out = 16'(6066);
			2005: out = 16'(3929);
			2006: out = 16'(2033);
			2007: out = 16'(-5644);
			2008: out = 16'(-13372);
			2009: out = 16'(-8951);
			2010: out = 16'(1960);
			2011: out = 16'(8159);
			2012: out = 16'(1015);
			2013: out = 16'(-1701);
			2014: out = 16'(-981);
			2015: out = 16'(4299);
			2016: out = 16'(-4910);
			2017: out = 16'(-7598);
			2018: out = 16'(-5895);
			2019: out = 16'(6166);
			2020: out = 16'(2057);
			2021: out = 16'(-2216);
			2022: out = 16'(-7147);
			2023: out = 16'(-2775);
			2024: out = 16'(-1120);
			2025: out = 16'(243);
			2026: out = 16'(-3010);
			2027: out = 16'(4224);
			2028: out = 16'(1728);
			2029: out = 16'(-7362);
			2030: out = 16'(6749);
			2031: out = 16'(469);
			2032: out = 16'(-5878);
			2033: out = 16'(-8021);
			2034: out = 16'(2);
			2035: out = 16'(3217);
			2036: out = 16'(253);
			2037: out = 16'(6756);
			2038: out = 16'(1641);
			2039: out = 16'(-3265);
			2040: out = 16'(-8260);
			2041: out = 16'(1119);
			2042: out = 16'(5841);
			2043: out = 16'(4401);
			2044: out = 16'(-4039);
			2045: out = 16'(-8474);
			2046: out = 16'(-8149);
			2047: out = 16'(-2232);
			2048: out = 16'(728);
			2049: out = 16'(4);
			2050: out = 16'(-4779);
			2051: out = 16'(6100);
			2052: out = 16'(-3528);
			2053: out = 16'(-6048);
			2054: out = 16'(3437);
			2055: out = 16'(8144);
			2056: out = 16'(4996);
			2057: out = 16'(-4104);
			2058: out = 16'(-3824);
			2059: out = 16'(-5909);
			2060: out = 16'(-1632);
			2061: out = 16'(5656);
			2062: out = 16'(4306);
			2063: out = 16'(362);
			2064: out = 16'(-4902);
			2065: out = 16'(2663);
			2066: out = 16'(-5204);
			2067: out = 16'(-4360);
			2068: out = 16'(7394);
			2069: out = 16'(4823);
			2070: out = 16'(401);
			2071: out = 16'(-6056);
			2072: out = 16'(-5609);
			2073: out = 16'(1649);
			2074: out = 16'(8152);
			2075: out = 16'(3914);
			2076: out = 16'(6594);
			2077: out = 16'(-3305);
			2078: out = 16'(-11479);
			2079: out = 16'(-11377);
			2080: out = 16'(632);
			2081: out = 16'(8719);
			2082: out = 16'(6209);
			2083: out = 16'(2564);
			2084: out = 16'(-2397);
			2085: out = 16'(-1122);
			2086: out = 16'(6486);
			2087: out = 16'(6771);
			2088: out = 16'(866);
			2089: out = 16'(-7900);
			2090: out = 16'(-3852);
			2091: out = 16'(-1364);
			2092: out = 16'(1194);
			2093: out = 16'(8006);
			2094: out = 16'(-262);
			2095: out = 16'(-2861);
			2096: out = 16'(1740);
			2097: out = 16'(-1449);
			2098: out = 16'(155);
			2099: out = 16'(1140);
			2100: out = 16'(1901);
			2101: out = 16'(1263);
			2102: out = 16'(3104);
			2103: out = 16'(6820);
			2104: out = 16'(-2420);
			2105: out = 16'(-1283);
			2106: out = 16'(1336);
			2107: out = 16'(2835);
			2108: out = 16'(1746);
			2109: out = 16'(1830);
			2110: out = 16'(2039);
			2111: out = 16'(420);
			2112: out = 16'(-1733);
			2113: out = 16'(-3168);
			2114: out = 16'(-8147);
			2115: out = 16'(3505);
			2116: out = 16'(3952);
			2117: out = 16'(-3655);
			2118: out = 16'(-4067);
			2119: out = 16'(796);
			2120: out = 16'(5147);
			2121: out = 16'(-5919);
			2122: out = 16'(2965);
			2123: out = 16'(3990);
			2124: out = 16'(4959);
			2125: out = 16'(744);
			2126: out = 16'(5726);
			2127: out = 16'(5563);
			2128: out = 16'(-1336);
			2129: out = 16'(-4536);
			2130: out = 16'(-376);
			2131: out = 16'(7287);
			2132: out = 16'(1596);
			2133: out = 16'(1884);
			2134: out = 16'(-1227);
			2135: out = 16'(-9085);
			2136: out = 16'(-311);
			2137: out = 16'(4335);
			2138: out = 16'(5630);
			2139: out = 16'(2504);
			2140: out = 16'(3521);
			2141: out = 16'(451);
			2142: out = 16'(-8615);
			2143: out = 16'(-6907);
			2144: out = 16'(-1738);
			2145: out = 16'(3953);
			2146: out = 16'(4226);
			2147: out = 16'(-1955);
			2148: out = 16'(-5766);
			2149: out = 16'(1569);
			2150: out = 16'(-4614);
			2151: out = 16'(-3074);
			2152: out = 16'(-781);
			2153: out = 16'(4882);
			2154: out = 16'(540);
			2155: out = 16'(-1046);
			2156: out = 16'(2813);
			2157: out = 16'(-4281);
			2158: out = 16'(-7147);
			2159: out = 16'(-5729);
			2160: out = 16'(7846);
			2161: out = 16'(4882);
			2162: out = 16'(3327);
			2163: out = 16'(5961);
			2164: out = 16'(-2094);
			2165: out = 16'(-2124);
			2166: out = 16'(-473);
			2167: out = 16'(-7048);
			2168: out = 16'(-3892);
			2169: out = 16'(-813);
			2170: out = 16'(2617);
			2171: out = 16'(255);
			2172: out = 16'(3653);
			2173: out = 16'(4804);
			2174: out = 16'(-9714);
			2175: out = 16'(-3149);
			2176: out = 16'(3306);
			2177: out = 16'(4785);
			2178: out = 16'(6593);
			2179: out = 16'(1388);
			2180: out = 16'(-3382);
			2181: out = 16'(-3984);
			2182: out = 16'(1186);
			2183: out = 16'(3289);
			2184: out = 16'(-307);
			2185: out = 16'(2958);
			2186: out = 16'(148);
			2187: out = 16'(-2363);
			2188: out = 16'(111);
			2189: out = 16'(236);
			2190: out = 16'(2858);
			2191: out = 16'(4213);
			2192: out = 16'(4832);
			2193: out = 16'(-4027);
			2194: out = 16'(-11456);
			2195: out = 16'(-3208);
			2196: out = 16'(2121);
			2197: out = 16'(7096);
			2198: out = 16'(4562);
			2199: out = 16'(4207);
			2200: out = 16'(-5269);
			2201: out = 16'(-12231);
			2202: out = 16'(-14154);
			2203: out = 16'(-4000);
			2204: out = 16'(1754);
			2205: out = 16'(433);
			2206: out = 16'(7817);
			2207: out = 16'(2973);
			2208: out = 16'(-1861);
			2209: out = 16'(655);
			2210: out = 16'(-7581);
			2211: out = 16'(-9206);
			2212: out = 16'(-5320);
			2213: out = 16'(-4372);
			2214: out = 16'(-2279);
			2215: out = 16'(366);
			2216: out = 16'(6641);
			2217: out = 16'(299);
			2218: out = 16'(-4274);
			2219: out = 16'(-6192);
			2220: out = 16'(-3239);
			2221: out = 16'(2281);
			2222: out = 16'(7068);
			2223: out = 16'(7222);
			2224: out = 16'(-1218);
			2225: out = 16'(-11367);
			2226: out = 16'(-15974);
			2227: out = 16'(-5367);
			2228: out = 16'(5401);
			2229: out = 16'(8596);
			2230: out = 16'(1782);
			2231: out = 16'(1546);
			2232: out = 16'(1318);
			2233: out = 16'(2117);
			2234: out = 16'(-2882);
			2235: out = 16'(-3228);
			2236: out = 16'(-2176);
			2237: out = 16'(987);
			2238: out = 16'(-1821);
			2239: out = 16'(-2599);
			2240: out = 16'(-1527);
			2241: out = 16'(-1025);
			2242: out = 16'(2479);
			2243: out = 16'(1637);
			2244: out = 16'(-6861);
			2245: out = 16'(-5908);
			2246: out = 16'(-3323);
			2247: out = 16'(2257);
			2248: out = 16'(-5782);
			2249: out = 16'(2844);
			2250: out = 16'(3986);
			2251: out = 16'(-4203);
			2252: out = 16'(1292);
			2253: out = 16'(2620);
			2254: out = 16'(854);
			2255: out = 16'(6624);
			2256: out = 16'(-6638);
			2257: out = 16'(-8500);
			2258: out = 16'(8429);
			2259: out = 16'(3301);
			2260: out = 16'(2551);
			2261: out = 16'(-1162);
			2262: out = 16'(-1222);
			2263: out = 16'(-2563);
			2264: out = 16'(-2480);
			2265: out = 16'(-4983);
			2266: out = 16'(4434);
			2267: out = 16'(4294);
			2268: out = 16'(2517);
			2269: out = 16'(5099);
			2270: out = 16'(1774);
			2271: out = 16'(-308);
			2272: out = 16'(581);
			2273: out = 16'(-2504);
			2274: out = 16'(254);
			2275: out = 16'(3358);
			2276: out = 16'(3229);
			2277: out = 16'(2787);
			2278: out = 16'(1083);
			2279: out = 16'(-1545);
			2280: out = 16'(-1766);
			2281: out = 16'(-1007);
			2282: out = 16'(2591);
			2283: out = 16'(4750);
			2284: out = 16'(6403);
			2285: out = 16'(1354);
			2286: out = 16'(-4830);
			2287: out = 16'(-5800);
			2288: out = 16'(506);
			2289: out = 16'(5866);
			2290: out = 16'(8057);
			2291: out = 16'(-3767);
			2292: out = 16'(-6999);
			2293: out = 16'(-5);
			2294: out = 16'(755);
			2295: out = 16'(-708);
			2296: out = 16'(-2512);
			2297: out = 16'(4460);
			2298: out = 16'(6820);
			2299: out = 16'(7039);
			2300: out = 16'(1875);
			2301: out = 16'(1036);
			2302: out = 16'(-434);
			2303: out = 16'(-589);
			2304: out = 16'(-8854);
			2305: out = 16'(19);
			2306: out = 16'(3421);
			2307: out = 16'(5199);
			2308: out = 16'(-5812);
			2309: out = 16'(-1158);
			2310: out = 16'(3788);
			2311: out = 16'(7764);
			2312: out = 16'(-3424);
			2313: out = 16'(-3897);
			2314: out = 16'(3054);
			2315: out = 16'(8219);
			2316: out = 16'(3300);
			2317: out = 16'(-4327);
			2318: out = 16'(-8839);
			2319: out = 16'(-2062);
			2320: out = 16'(2528);
			2321: out = 16'(2652);
			2322: out = 16'(328);
			2323: out = 16'(1351);
			2324: out = 16'(1075);
			2325: out = 16'(-2659);
			2326: out = 16'(-2533);
			2327: out = 16'(1905);
			2328: out = 16'(6547);
			2329: out = 16'(-320);
			2330: out = 16'(-2878);
			2331: out = 16'(-1792);
			2332: out = 16'(6585);
			2333: out = 16'(-2934);
			2334: out = 16'(-8408);
			2335: out = 16'(-9730);
			2336: out = 16'(6623);
			2337: out = 16'(7502);
			2338: out = 16'(6498);
			2339: out = 16'(2473);
			2340: out = 16'(1980);
			2341: out = 16'(-1190);
			2342: out = 16'(-3931);
			2343: out = 16'(-11464);
			2344: out = 16'(-3040);
			2345: out = 16'(4013);
			2346: out = 16'(3672);
			2347: out = 16'(745);
			2348: out = 16'(-3135);
			2349: out = 16'(-3502);
			2350: out = 16'(-1038);
			2351: out = 16'(2560);
			2352: out = 16'(3509);
			2353: out = 16'(2388);
			2354: out = 16'(-1344);
			2355: out = 16'(-1243);
			2356: out = 16'(673);
			2357: out = 16'(260);
			2358: out = 16'(-254);
			2359: out = 16'(-2172);
			2360: out = 16'(-3018);
			2361: out = 16'(-4352);
			2362: out = 16'(-964);
			2363: out = 16'(1536);
			2364: out = 16'(-4775);
			2365: out = 16'(389);
			2366: out = 16'(4163);
			2367: out = 16'(4987);
			2368: out = 16'(141);
			2369: out = 16'(-4084);
			2370: out = 16'(-5204);
			2371: out = 16'(1363);
			2372: out = 16'(-879);
			2373: out = 16'(-2215);
			2374: out = 16'(-1977);
			2375: out = 16'(4595);
			2376: out = 16'(5082);
			2377: out = 16'(851);
			2378: out = 16'(-7531);
			2379: out = 16'(-7693);
			2380: out = 16'(-3092);
			2381: out = 16'(3448);
			2382: out = 16'(4600);
			2383: out = 16'(1922);
			2384: out = 16'(-3592);
			2385: out = 16'(-5176);
			2386: out = 16'(-5389);
			2387: out = 16'(665);
			2388: out = 16'(5100);
			2389: out = 16'(2171);
			2390: out = 16'(-5575);
			2391: out = 16'(-8374);
			2392: out = 16'(1959);
			2393: out = 16'(4604);
			2394: out = 16'(2134);
			2395: out = 16'(-6166);
			2396: out = 16'(-765);
			2397: out = 16'(-3195);
			2398: out = 16'(-2917);
			2399: out = 16'(825);
			2400: out = 16'(-2874);
			2401: out = 16'(-4227);
			2402: out = 16'(-1325);
			2403: out = 16'(-1172);
			2404: out = 16'(4555);
			2405: out = 16'(5442);
			2406: out = 16'(-1186);
			2407: out = 16'(228);
			2408: out = 16'(461);
			2409: out = 16'(393);
			2410: out = 16'(2421);
			2411: out = 16'(-1564);
			2412: out = 16'(-4552);
			2413: out = 16'(-1267);
			2414: out = 16'(-1207);
			2415: out = 16'(1722);
			2416: out = 16'(2975);
			2417: out = 16'(1183);
			2418: out = 16'(-2119);
			2419: out = 16'(-4065);
			2420: out = 16'(-3855);
			2421: out = 16'(3403);
			2422: out = 16'(5473);
			2423: out = 16'(3024);
			2424: out = 16'(4695);
			2425: out = 16'(-726);
			2426: out = 16'(-3129);
			2427: out = 16'(-1383);
			2428: out = 16'(1697);
			2429: out = 16'(1824);
			2430: out = 16'(-960);
			2431: out = 16'(-1924);
			2432: out = 16'(-2312);
			2433: out = 16'(1214);
			2434: out = 16'(5631);
			2435: out = 16'(3839);
			2436: out = 16'(252);
			2437: out = 16'(-1826);
			2438: out = 16'(2490);
			2439: out = 16'(2786);
			2440: out = 16'(51);
			2441: out = 16'(-5521);
			2442: out = 16'(1302);
			2443: out = 16'(3863);
			2444: out = 16'(3967);
			2445: out = 16'(6930);
			2446: out = 16'(1173);
			2447: out = 16'(-755);
			2448: out = 16'(1156);
			2449: out = 16'(-91);
			2450: out = 16'(-3132);
			2451: out = 16'(-5395);
			2452: out = 16'(-2002);
			2453: out = 16'(2640);
			2454: out = 16'(3275);
			2455: out = 16'(-2397);
			2456: out = 16'(-115);
			2457: out = 16'(570);
			2458: out = 16'(1962);
			2459: out = 16'(-4722);
			2460: out = 16'(1815);
			2461: out = 16'(2961);
			2462: out = 16'(189);
			2463: out = 16'(4131);
			2464: out = 16'(1015);
			2465: out = 16'(-4093);
			2466: out = 16'(-1248);
			2467: out = 16'(-5974);
			2468: out = 16'(-1162);
			2469: out = 16'(6485);
			2470: out = 16'(5181);
			2471: out = 16'(-2055);
			2472: out = 16'(-9384);
			2473: out = 16'(-10714);
			2474: out = 16'(1128);
			2475: out = 16'(8476);
			2476: out = 16'(5832);
			2477: out = 16'(-3322);
			2478: out = 16'(-5704);
			2479: out = 16'(-1470);
			2480: out = 16'(-324);
			2481: out = 16'(6163);
			2482: out = 16'(4391);
			2483: out = 16'(-543);
			2484: out = 16'(-5981);
			2485: out = 16'(-3453);
			2486: out = 16'(2265);
			2487: out = 16'(4247);
			2488: out = 16'(5119);
			2489: out = 16'(-728);
			2490: out = 16'(-7520);
			2491: out = 16'(4343);
			2492: out = 16'(4857);
			2493: out = 16'(3002);
			2494: out = 16'(-651);
			2495: out = 16'(-1198);
			2496: out = 16'(-2684);
			2497: out = 16'(-3399);
			2498: out = 16'(3529);
			2499: out = 16'(4200);
			2500: out = 16'(2531);
			2501: out = 16'(-2352);
			2502: out = 16'(2673);
			2503: out = 16'(1958);
			2504: out = 16'(-1588);
			2505: out = 16'(4808);
			2506: out = 16'(1523);
			2507: out = 16'(-186);
			2508: out = 16'(87);
			2509: out = 16'(621);
			2510: out = 16'(-1263);
			2511: out = 16'(-2940);
			2512: out = 16'(3774);
			2513: out = 16'(3217);
			2514: out = 16'(1535);
			2515: out = 16'(-403);
			2516: out = 16'(1086);
			2517: out = 16'(2323);
			2518: out = 16'(1009);
			2519: out = 16'(-9417);
			2520: out = 16'(-5810);
			2521: out = 16'(1991);
			2522: out = 16'(5241);
			2523: out = 16'(5250);
			2524: out = 16'(-3738);
			2525: out = 16'(-11044);
			2526: out = 16'(-3513);
			2527: out = 16'(2211);
			2528: out = 16'(4321);
			2529: out = 16'(1738);
			2530: out = 16'(-23);
			2531: out = 16'(1529);
			2532: out = 16'(3716);
			2533: out = 16'(2567);
			2534: out = 16'(-1619);
			2535: out = 16'(-2266);
			2536: out = 16'(2936);
			2537: out = 16'(3654);
			2538: out = 16'(3177);
			2539: out = 16'(346);
			2540: out = 16'(-3802);
			2541: out = 16'(755);
			2542: out = 16'(3722);
			2543: out = 16'(1816);
			2544: out = 16'(-2144);
			2545: out = 16'(-1494);
			2546: out = 16'(2190);
			2547: out = 16'(-1372);
			2548: out = 16'(370);
			2549: out = 16'(-1180);
			2550: out = 16'(-697);
			2551: out = 16'(-3629);
			2552: out = 16'(547);
			2553: out = 16'(2811);
			2554: out = 16'(2620);
			2555: out = 16'(-3407);
			2556: out = 16'(-4094);
			2557: out = 16'(-354);
			2558: out = 16'(1273);
			2559: out = 16'(-1701);
			2560: out = 16'(-3623);
			2561: out = 16'(1452);
			2562: out = 16'(3484);
			2563: out = 16'(1302);
			2564: out = 16'(-5092);
			2565: out = 16'(-7075);
			2566: out = 16'(-3757);
			2567: out = 16'(2020);
			2568: out = 16'(608);
			2569: out = 16'(4703);
			2570: out = 16'(835);
			2571: out = 16'(-7037);
			2572: out = 16'(-2862);
			2573: out = 16'(-6698);
			2574: out = 16'(-5308);
			2575: out = 16'(7480);
			2576: out = 16'(2597);
			2577: out = 16'(-3243);
			2578: out = 16'(-9989);
			2579: out = 16'(-1239);
			2580: out = 16'(602);
			2581: out = 16'(2843);
			2582: out = 16'(4251);
			2583: out = 16'(2294);
			2584: out = 16'(-1456);
			2585: out = 16'(-4005);
			2586: out = 16'(-2770);
			2587: out = 16'(1316);
			2588: out = 16'(2237);
			2589: out = 16'(-5515);
			2590: out = 16'(3021);
			2591: out = 16'(3973);
			2592: out = 16'(1292);
			2593: out = 16'(1023);
			2594: out = 16'(-787);
			2595: out = 16'(-1840);
			2596: out = 16'(-3245);
			2597: out = 16'(1225);
			2598: out = 16'(2752);
			2599: out = 16'(1941);
			2600: out = 16'(-725);
			2601: out = 16'(-1013);
			2602: out = 16'(98);
			2603: out = 16'(1601);
			2604: out = 16'(1006);
			2605: out = 16'(-663);
			2606: out = 16'(-2598);
			2607: out = 16'(-767);
			2608: out = 16'(-408);
			2609: out = 16'(1312);
			2610: out = 16'(2229);
			2611: out = 16'(3548);
			2612: out = 16'(1696);
			2613: out = 16'(111);
			2614: out = 16'(192);
			2615: out = 16'(804);
			2616: out = 16'(1590);
			2617: out = 16'(5037);
			2618: out = 16'(-7286);
			2619: out = 16'(-6275);
			2620: out = 16'(195);
			2621: out = 16'(6424);
			2622: out = 16'(-980);
			2623: out = 16'(-5631);
			2624: out = 16'(-847);
			2625: out = 16'(1059);
			2626: out = 16'(3124);
			2627: out = 16'(1393);
			2628: out = 16'(4);
			2629: out = 16'(1048);
			2630: out = 16'(3561);
			2631: out = 16'(3109);
			2632: out = 16'(-1911);
			2633: out = 16'(-2488);
			2634: out = 16'(689);
			2635: out = 16'(-10133);
			2636: out = 16'(2524);
			2637: out = 16'(4460);
			2638: out = 16'(-127);
			2639: out = 16'(-6855);
			2640: out = 16'(-1228);
			2641: out = 16'(4323);
			2642: out = 16'(-4572);
			2643: out = 16'(-6094);
			2644: out = 16'(-3538);
			2645: out = 16'(4455);
			2646: out = 16'(4874);
			2647: out = 16'(1096);
			2648: out = 16'(-4014);
			2649: out = 16'(1278);
			2650: out = 16'(1696);
			2651: out = 16'(4294);
			2652: out = 16'(3530);
			2653: out = 16'(-1088);
			2654: out = 16'(-4476);
			2655: out = 16'(-2884);
			2656: out = 16'(3323);
			2657: out = 16'(1823);
			2658: out = 16'(-2076);
			2659: out = 16'(-5447);
			2660: out = 16'(1463);
			2661: out = 16'(3656);
			2662: out = 16'(2200);
			2663: out = 16'(-3897);
			2664: out = 16'(-2538);
			2665: out = 16'(-826);
			2666: out = 16'(623);
			2667: out = 16'(970);
			2668: out = 16'(857);
			2669: out = 16'(495);
			2670: out = 16'(487);
			2671: out = 16'(486);
			2672: out = 16'(651);
			2673: out = 16'(475);
			2674: out = 16'(676);
			2675: out = 16'(58);
			2676: out = 16'(720);
			2677: out = 16'(3624);
			2678: out = 16'(1394);
			2679: out = 16'(-1492);
			2680: out = 16'(-3938);
			2681: out = 16'(4274);
			2682: out = 16'(1627);
			2683: out = 16'(-2213);
			2684: out = 16'(-4474);
			2685: out = 16'(-1764);
			2686: out = 16'(-605);
			2687: out = 16'(-1927);
			2688: out = 16'(5561);
			2689: out = 16'(-937);
			2690: out = 16'(-5601);
			2691: out = 16'(-3074);
			2692: out = 16'(453);
			2693: out = 16'(3460);
			2694: out = 16'(2257);
			2695: out = 16'(-399);
			2696: out = 16'(-4908);
			2697: out = 16'(-3726);
			2698: out = 16'(4765);
			2699: out = 16'(1549);
			2700: out = 16'(-1210);
			2701: out = 16'(-3661);
			2702: out = 16'(6336);
			2703: out = 16'(1404);
			2704: out = 16'(-3610);
			2705: out = 16'(-8833);
			2706: out = 16'(1445);
			2707: out = 16'(5259);
			2708: out = 16'(4563);
			2709: out = 16'(-5171);
			2710: out = 16'(-139);
			2711: out = 16'(2707);
			2712: out = 16'(37);
			2713: out = 16'(1134);
			2714: out = 16'(3026);
			2715: out = 16'(4097);
			2716: out = 16'(-4201);
			2717: out = 16'(-2901);
			2718: out = 16'(-628);
			2719: out = 16'(1206);
			2720: out = 16'(3016);
			2721: out = 16'(46);
			2722: out = 16'(-3540);
			2723: out = 16'(-3214);
			2724: out = 16'(1128);
			2725: out = 16'(2646);
			2726: out = 16'(-1968);
			2727: out = 16'(1628);
			2728: out = 16'(1374);
			2729: out = 16'(1392);
			2730: out = 16'(-2918);
			2731: out = 16'(-1235);
			2732: out = 16'(-63);
			2733: out = 16'(3170);
			2734: out = 16'(3121);
			2735: out = 16'(4334);
			2736: out = 16'(1546);
			2737: out = 16'(587);
			2738: out = 16'(-7929);
			2739: out = 16'(-4499);
			2740: out = 16'(6246);
			2741: out = 16'(4609);
			2742: out = 16'(-354);
			2743: out = 16'(-5873);
			2744: out = 16'(-5259);
			2745: out = 16'(1417);
			2746: out = 16'(5036);
			2747: out = 16'(3044);
			2748: out = 16'(139);
			2749: out = 16'(122);
			2750: out = 16'(350);
			2751: out = 16'(-4768);
			2752: out = 16'(-1163);
			2753: out = 16'(1454);
			2754: out = 16'(1503);
			2755: out = 16'(5752);
			2756: out = 16'(-4479);
			2757: out = 16'(-11715);
			2758: out = 16'(-1345);
			2759: out = 16'(1483);
			2760: out = 16'(4395);
			2761: out = 16'(1898);
			2762: out = 16'(-243);
			2763: out = 16'(-2707);
			2764: out = 16'(-1759);
			2765: out = 16'(-1546);
			2766: out = 16'(2455);
			2767: out = 16'(1141);
			2768: out = 16'(-1458);
			2769: out = 16'(3305);
			2770: out = 16'(2971);
			2771: out = 16'(2344);
			2772: out = 16'(2997);
			2773: out = 16'(-143);
			2774: out = 16'(-1114);
			2775: out = 16'(-682);
			2776: out = 16'(3139);
			2777: out = 16'(1387);
			2778: out = 16'(-1041);
			2779: out = 16'(-3009);
			2780: out = 16'(735);
			2781: out = 16'(2169);
			2782: out = 16'(1146);
			2783: out = 16'(-4275);
			2784: out = 16'(-634);
			2785: out = 16'(2996);
			2786: out = 16'(563);
			2787: out = 16'(2123);
			2788: out = 16'(-2941);
			2789: out = 16'(-6364);
			2790: out = 16'(2309);
			2791: out = 16'(4093);
			2792: out = 16'(2028);
			2793: out = 16'(-6067);
			2794: out = 16'(1453);
			2795: out = 16'(-214);
			2796: out = 16'(-3637);
			2797: out = 16'(2556);
			2798: out = 16'(-488);
			2799: out = 16'(-1829);
			2800: out = 16'(-1770);
			2801: out = 16'(1223);
			2802: out = 16'(-602);
			2803: out = 16'(-3447);
			2804: out = 16'(2599);
			2805: out = 16'(1741);
			2806: out = 16'(-137);
			2807: out = 16'(-7699);
			2808: out = 16'(3352);
			2809: out = 16'(-785);
			2810: out = 16'(-5820);
			2811: out = 16'(-3732);
			2812: out = 16'(1676);
			2813: out = 16'(2460);
			2814: out = 16'(-2475);
			2815: out = 16'(-2750);
			2816: out = 16'(-213);
			2817: out = 16'(2100);
			2818: out = 16'(-4296);
			2819: out = 16'(-3248);
			2820: out = 16'(-1436);
			2821: out = 16'(543);
			2822: out = 16'(315);
			2823: out = 16'(-3751);
			2824: out = 16'(-5427);
			2825: out = 16'(4618);
			2826: out = 16'(1438);
			2827: out = 16'(-2723);
			2828: out = 16'(-6592);
			2829: out = 16'(-6968);
			2830: out = 16'(-422);
			2831: out = 16'(5765);
			2832: out = 16'(3599);
			2833: out = 16'(935);
			2834: out = 16'(-1520);
			2835: out = 16'(380);
			2836: out = 16'(207);
			2837: out = 16'(2091);
			2838: out = 16'(1751);
			2839: out = 16'(1030);
			2840: out = 16'(-1014);
			2841: out = 16'(-211);
			2842: out = 16'(1984);
			2843: out = 16'(1181);
			2844: out = 16'(763);
			2845: out = 16'(-715);
			2846: out = 16'(-3158);
			2847: out = 16'(-1954);
			2848: out = 16'(171);
			2849: out = 16'(1761);
			2850: out = 16'(680);
			2851: out = 16'(-1348);
			2852: out = 16'(-1622);
			2853: out = 16'(3872);
			2854: out = 16'(-564);
			2855: out = 16'(-1859);
			2856: out = 16'(-1567);
			2857: out = 16'(1692);
			2858: out = 16'(-402);
			2859: out = 16'(-2011);
			2860: out = 16'(1299);
			2861: out = 16'(1203);
			2862: out = 16'(2348);
			2863: out = 16'(2044);
			2864: out = 16'(2201);
			2865: out = 16'(530);
			2866: out = 16'(9);
			2867: out = 16'(-702);
			2868: out = 16'(1788);
			2869: out = 16'(1390);
			2870: out = 16'(581);
			2871: out = 16'(-237);
			2872: out = 16'(1060);
			2873: out = 16'(1082);
			2874: out = 16'(1866);
			2875: out = 16'(-3315);
			2876: out = 16'(-659);
			2877: out = 16'(3253);
			2878: out = 16'(-2254);
			2879: out = 16'(-5956);
			2880: out = 16'(-5292);
			2881: out = 16'(2514);
			2882: out = 16'(4775);
			2883: out = 16'(1343);
			2884: out = 16'(-5064);
			2885: out = 16'(3418);
			2886: out = 16'(1276);
			2887: out = 16'(207);
			2888: out = 16'(-2943);
			2889: out = 16'(3156);
			2890: out = 16'(1778);
			2891: out = 16'(-1622);
			2892: out = 16'(626);
			2893: out = 16'(-307);
			2894: out = 16'(1169);
			2895: out = 16'(3204);
			2896: out = 16'(2414);
			2897: out = 16'(-403);
			2898: out = 16'(-1831);
			2899: out = 16'(3567);
			2900: out = 16'(3849);
			2901: out = 16'(1845);
			2902: out = 16'(-2497);
			2903: out = 16'(-290);
			2904: out = 16'(1215);
			2905: out = 16'(2243);
			2906: out = 16'(-180);
			2907: out = 16'(382);
			2908: out = 16'(-775);
			2909: out = 16'(-3502);
			2910: out = 16'(3037);
			2911: out = 16'(3895);
			2912: out = 16'(2477);
			2913: out = 16'(-1493);
			2914: out = 16'(795);
			2915: out = 16'(1926);
			2916: out = 16'(1135);
			2917: out = 16'(1567);
			2918: out = 16'(837);
			2919: out = 16'(-301);
			2920: out = 16'(-470);
			2921: out = 16'(-1852);
			2922: out = 16'(-124);
			2923: out = 16'(2983);
			2924: out = 16'(2642);
			2925: out = 16'(-503);
			2926: out = 16'(-3096);
			2927: out = 16'(395);
			2928: out = 16'(2009);
			2929: out = 16'(2460);
			2930: out = 16'(-332);
			2931: out = 16'(3135);
			2932: out = 16'(786);
			2933: out = 16'(-1427);
			2934: out = 16'(-4812);
			2935: out = 16'(1133);
			2936: out = 16'(3222);
			2937: out = 16'(965);
			2938: out = 16'(-394);
			2939: out = 16'(-3300);
			2940: out = 16'(-3040);
			2941: out = 16'(3250);
			2942: out = 16'(611);
			2943: out = 16'(887);
			2944: out = 16'(2555);
			2945: out = 16'(-109);
			2946: out = 16'(239);
			2947: out = 16'(780);
			2948: out = 16'(670);
			2949: out = 16'(-829);
			2950: out = 16'(-3419);
			2951: out = 16'(-4731);
			2952: out = 16'(2011);
			2953: out = 16'(3404);
			2954: out = 16'(1421);
			2955: out = 16'(-3795);
			2956: out = 16'(-1726);
			2957: out = 16'(994);
			2958: out = 16'(2711);
			2959: out = 16'(31);
			2960: out = 16'(246);
			2961: out = 16'(29);
			2962: out = 16'(-4231);
			2963: out = 16'(843);
			2964: out = 16'(-21);
			2965: out = 16'(-1541);
			2966: out = 16'(1456);
			2967: out = 16'(4000);
			2968: out = 16'(1873);
			2969: out = 16'(-5884);
			2970: out = 16'(-5661);
			2971: out = 16'(-1319);
			2972: out = 16'(3856);
			2973: out = 16'(1686);
			2974: out = 16'(-1827);
			2975: out = 16'(-3480);
			2976: out = 16'(2472);
			2977: out = 16'(-1082);
			2978: out = 16'(-141);
			2979: out = 16'(84);
			2980: out = 16'(-1043);
			2981: out = 16'(70);
			2982: out = 16'(2131);
			2983: out = 16'(2422);
			2984: out = 16'(-223);
			2985: out = 16'(-2296);
			2986: out = 16'(-1215);
			2987: out = 16'(191);
			2988: out = 16'(1897);
			2989: out = 16'(561);
			2990: out = 16'(369);
			2991: out = 16'(-5690);
			2992: out = 16'(-1821);
			2993: out = 16'(2067);
			2994: out = 16'(239);
			2995: out = 16'(-6923);
			2996: out = 16'(-6699);
			2997: out = 16'(4682);
			2998: out = 16'(4213);
			2999: out = 16'(2970);
			3000: out = 16'(-2687);
			3001: out = 16'(-6617);
			3002: out = 16'(-6510);
			3003: out = 16'(-1736);
			3004: out = 16'(2102);
			3005: out = 16'(2397);
			3006: out = 16'(65);
			3007: out = 16'(-2055);
			3008: out = 16'(-2050);
			3009: out = 16'(-1720);
			3010: out = 16'(-678);
			3011: out = 16'(-31);
			3012: out = 16'(1626);
			3013: out = 16'(-214);
			3014: out = 16'(-1715);
			3015: out = 16'(1404);
			3016: out = 16'(-255);
			3017: out = 16'(-1441);
			3018: out = 16'(-2289);
			3019: out = 16'(-33);
			3020: out = 16'(704);
			3021: out = 16'(340);
			3022: out = 16'(-1809);
			3023: out = 16'(49);
			3024: out = 16'(558);
			3025: out = 16'(-995);
			3026: out = 16'(2254);
			3027: out = 16'(-642);
			3028: out = 16'(-3053);
			3029: out = 16'(-3320);
			3030: out = 16'(1800);
			3031: out = 16'(3043);
			3032: out = 16'(18);
			3033: out = 16'(3259);
			3034: out = 16'(63);
			3035: out = 16'(-2220);
			3036: out = 16'(-1865);
			3037: out = 16'(-2541);
			3038: out = 16'(-1827);
			3039: out = 16'(-61);
			3040: out = 16'(3141);
			3041: out = 16'(2111);
			3042: out = 16'(642);
			3043: out = 16'(3145);
			3044: out = 16'(-2657);
			3045: out = 16'(-2985);
			3046: out = 16'(-160);
			3047: out = 16'(2855);
			3048: out = 16'(2015);
			3049: out = 16'(-378);
			3050: out = 16'(-2379);
			3051: out = 16'(1346);
			3052: out = 16'(3541);
			3053: out = 16'(2775);
			3054: out = 16'(1364);
			3055: out = 16'(-2235);
			3056: out = 16'(-3146);
			3057: out = 16'(603);
			3058: out = 16'(-79);
			3059: out = 16'(955);
			3060: out = 16'(1819);
			3061: out = 16'(2934);
			3062: out = 16'(2271);
			3063: out = 16'(1103);
			3064: out = 16'(-1397);
			3065: out = 16'(1453);
			3066: out = 16'(470);
			3067: out = 16'(-1382);
			3068: out = 16'(-619);
			3069: out = 16'(325);
			3070: out = 16'(1223);
			3071: out = 16'(1437);
			3072: out = 16'(370);
			3073: out = 16'(329);
			3074: out = 16'(988);
			3075: out = 16'(3339);
			3076: out = 16'(609);
			3077: out = 16'(171);
			3078: out = 16'(3994);
			3079: out = 16'(-157);
			3080: out = 16'(-263);
			3081: out = 16'(59);
			3082: out = 16'(508);
			3083: out = 16'(260);
			3084: out = 16'(148);
			3085: out = 16'(119);
			3086: out = 16'(1376);
			3087: out = 16'(2860);
			3088: out = 16'(2900);
			3089: out = 16'(-4227);
			3090: out = 16'(-1277);
			3091: out = 16'(1433);
			3092: out = 16'(3229);
			3093: out = 16'(-4192);
			3094: out = 16'(-4286);
			3095: out = 16'(-1298);
			3096: out = 16'(-1959);
			3097: out = 16'(820);
			3098: out = 16'(1686);
			3099: out = 16'(1898);
			3100: out = 16'(331);
			3101: out = 16'(78);
			3102: out = 16'(-106);
			3103: out = 16'(163);
			3104: out = 16'(-1370);
			3105: out = 16'(-1390);
			3106: out = 16'(330);
			3107: out = 16'(965);
			3108: out = 16'(1228);
			3109: out = 16'(362);
			3110: out = 16'(-810);
			3111: out = 16'(-953);
			3112: out = 16'(-1366);
			3113: out = 16'(-2912);
			3114: out = 16'(1978);
			3115: out = 16'(598);
			3116: out = 16'(-631);
			3117: out = 16'(194);
			3118: out = 16'(702);
			3119: out = 16'(-1354);
			3120: out = 16'(-4673);
			3121: out = 16'(1109);
			3122: out = 16'(2748);
			3123: out = 16'(2900);
			3124: out = 16'(1857);
			3125: out = 16'(-557);
			3126: out = 16'(-1506);
			3127: out = 16'(-948);
			3128: out = 16'(-1163);
			3129: out = 16'(77);
			3130: out = 16'(1346);
			3131: out = 16'(67);
			3132: out = 16'(2119);
			3133: out = 16'(203);
			3134: out = 16'(-2610);
			3135: out = 16'(-4336);
			3136: out = 16'(-557);
			3137: out = 16'(2391);
			3138: out = 16'(1259);
			3139: out = 16'(-2425);
			3140: out = 16'(-2515);
			3141: out = 16'(1190);
			3142: out = 16'(2393);
			3143: out = 16'(91);
			3144: out = 16'(-2207);
			3145: out = 16'(3337);
			3146: out = 16'(-4433);
			3147: out = 16'(-3529);
			3148: out = 16'(826);
			3149: out = 16'(2808);
			3150: out = 16'(1940);
			3151: out = 16'(-73);
			3152: out = 16'(-617);
			3153: out = 16'(-77);
			3154: out = 16'(287);
			3155: out = 16'(-977);
			3156: out = 16'(505);
			3157: out = 16'(-1957);
			3158: out = 16'(-1412);
			3159: out = 16'(1322);
			3160: out = 16'(3286);
			3161: out = 16'(-206);
			3162: out = 16'(-5375);
			3163: out = 16'(-3163);
			3164: out = 16'(-1097);
			3165: out = 16'(1765);
			3166: out = 16'(1950);
			3167: out = 16'(-23);
			3168: out = 16'(-1873);
			3169: out = 16'(-1273);
			3170: out = 16'(-228);
			3171: out = 16'(1643);
			3172: out = 16'(349);
			3173: out = 16'(-2999);
			3174: out = 16'(-2107);
			3175: out = 16'(-57);
			3176: out = 16'(1817);
			3177: out = 16'(537);
			3178: out = 16'(561);
			3179: out = 16'(-868);
			3180: out = 16'(-3296);
			3181: out = 16'(1576);
			3182: out = 16'(2325);
			3183: out = 16'(1465);
			3184: out = 16'(43);
			3185: out = 16'(326);
			3186: out = 16'(1293);
			3187: out = 16'(2592);
			3188: out = 16'(-5075);
			3189: out = 16'(-4601);
			3190: out = 16'(-129);
			3191: out = 16'(2418);
			3192: out = 16'(3835);
			3193: out = 16'(2358);
			3194: out = 16'(280);
			3195: out = 16'(-4003);
			3196: out = 16'(-2627);
			3197: out = 16'(549);
			3198: out = 16'(-714);
			3199: out = 16'(2735);
			3200: out = 16'(2554);
			3201: out = 16'(1270);
			3202: out = 16'(-2216);
			3203: out = 16'(83);
			3204: out = 16'(2339);
			3205: out = 16'(-94);
			3206: out = 16'(-1387);
			3207: out = 16'(-1558);
			3208: out = 16'(1239);
			3209: out = 16'(1219);
			3210: out = 16'(2046);
			3211: out = 16'(240);
			3212: out = 16'(-2102);
			3213: out = 16'(-3961);
			3214: out = 16'(-1964);
			3215: out = 16'(1192);
			3216: out = 16'(3098);
			3217: out = 16'(-1393);
			3218: out = 16'(-5381);
			3219: out = 16'(-365);
			3220: out = 16'(-3112);
			3221: out = 16'(-129);
			3222: out = 16'(3008);
			3223: out = 16'(2089);
			3224: out = 16'(-551);
			3225: out = 16'(-1396);
			3226: out = 16'(2493);
			3227: out = 16'(-654);
			3228: out = 16'(-1229);
			3229: out = 16'(-123);
			3230: out = 16'(1490);
			3231: out = 16'(1885);
			3232: out = 16'(69);
			3233: out = 16'(-2600);
			3234: out = 16'(-3354);
			3235: out = 16'(-600);
			3236: out = 16'(3014);
			3237: out = 16'(3558);
			3238: out = 16'(1534);
			3239: out = 16'(-1922);
			3240: out = 16'(-5315);
			3241: out = 16'(-2257);
			3242: out = 16'(-93);
			3243: out = 16'(1285);
			3244: out = 16'(2539);
			3245: out = 16'(2783);
			3246: out = 16'(838);
			3247: out = 16'(-2678);
			3248: out = 16'(-2032);
			3249: out = 16'(52);
			3250: out = 16'(1980);
			3251: out = 16'(3725);
			3252: out = 16'(-219);
			3253: out = 16'(-2068);
			3254: out = 16'(544);
			3255: out = 16'(300);
			3256: out = 16'(-546);
			3257: out = 16'(-1620);
			3258: out = 16'(3020);
			3259: out = 16'(1491);
			3260: out = 16'(-491);
			3261: out = 16'(-3093);
			3262: out = 16'(394);
			3263: out = 16'(2313);
			3264: out = 16'(2205);
			3265: out = 16'(-2838);
			3266: out = 16'(-2513);
			3267: out = 16'(-1656);
			3268: out = 16'(-1172);
			3269: out = 16'(374);
			3270: out = 16'(-483);
			3271: out = 16'(-938);
			3272: out = 16'(2502);
			3273: out = 16'(2219);
			3274: out = 16'(791);
			3275: out = 16'(-2105);
			3276: out = 16'(763);
			3277: out = 16'(590);
			3278: out = 16'(88);
			3279: out = 16'(266);
			3280: out = 16'(-243);
			3281: out = 16'(-392);
			3282: out = 16'(-15);
			3283: out = 16'(2142);
			3284: out = 16'(1933);
			3285: out = 16'(373);
			3286: out = 16'(-437);
			3287: out = 16'(-1372);
			3288: out = 16'(-361);
			3289: out = 16'(1035);
			3290: out = 16'(647);
			3291: out = 16'(-140);
			3292: out = 16'(-283);
			3293: out = 16'(427);
			3294: out = 16'(883);
			3295: out = 16'(292);
			3296: out = 16'(-201);
			3297: out = 16'(-264);
			3298: out = 16'(1993);
			3299: out = 16'(1813);
			3300: out = 16'(-4570);
			3301: out = 16'(-3428);
			3302: out = 16'(-1116);
			3303: out = 16'(1530);
			3304: out = 16'(459);
			3305: out = 16'(-1782);
			3306: out = 16'(-3172);
			3307: out = 16'(814);
			3308: out = 16'(1);
			3309: out = 16'(394);
			3310: out = 16'(-576);
			3311: out = 16'(-29);
			3312: out = 16'(-3252);
			3313: out = 16'(-3458);
			3314: out = 16'(3075);
			3315: out = 16'(1001);
			3316: out = 16'(1218);
			3317: out = 16'(1518);
			3318: out = 16'(-3022);
			3319: out = 16'(-2681);
			3320: out = 16'(-975);
			3321: out = 16'(2);
			3322: out = 16'(1981);
			3323: out = 16'(850);
			3324: out = 16'(-1769);
			3325: out = 16'(1850);
			3326: out = 16'(-399);
			3327: out = 16'(-1570);
			3328: out = 16'(-944);
			3329: out = 16'(2082);
			3330: out = 16'(1651);
			3331: out = 16'(-1415);
			3332: out = 16'(-1217);
			3333: out = 16'(-2543);
			3334: out = 16'(-1050);
			3335: out = 16'(2167);
			3336: out = 16'(1664);
			3337: out = 16'(777);
			3338: out = 16'(-141);
			3339: out = 16'(-1665);
			3340: out = 16'(-401);
			3341: out = 16'(1039);
			3342: out = 16'(1647);
			3343: out = 16'(1194);
			3344: out = 16'(-67);
			3345: out = 16'(-1379);
			3346: out = 16'(862);
			3347: out = 16'(-1044);
			3348: out = 16'(-1276);
			3349: out = 16'(421);
			3350: out = 16'(996);
			3351: out = 16'(808);
			3352: out = 16'(439);
			3353: out = 16'(835);
			3354: out = 16'(1008);
			3355: out = 16'(-341);
			3356: out = 16'(-2751);
			3357: out = 16'(-4533);
			3358: out = 16'(-1045);
			3359: out = 16'(3594);
			3360: out = 16'(-1707);
			3361: out = 16'(2092);
			3362: out = 16'(1422);
			3363: out = 16'(-1652);
			3364: out = 16'(-2693);
			3365: out = 16'(-259);
			3366: out = 16'(2283);
			3367: out = 16'(-2704);
			3368: out = 16'(501);
			3369: out = 16'(1167);
			3370: out = 16'(77);
			3371: out = 16'(-2108);
			3372: out = 16'(-2114);
			3373: out = 16'(-753);
			3374: out = 16'(675);
			3375: out = 16'(459);
			3376: out = 16'(177);
			3377: out = 16'(663);
			3378: out = 16'(607);
			3379: out = 16'(745);
			3380: out = 16'(550);
			3381: out = 16'(1781);
			3382: out = 16'(-1363);
			3383: out = 16'(-1362);
			3384: out = 16'(1945);
			3385: out = 16'(2938);
			3386: out = 16'(2209);
			3387: out = 16'(-121);
			3388: out = 16'(3017);
			3389: out = 16'(-4848);
			3390: out = 16'(-4444);
			3391: out = 16'(1684);
			3392: out = 16'(1692);
			3393: out = 16'(597);
			3394: out = 16'(-1362);
			3395: out = 16'(245);
			3396: out = 16'(1046);
			3397: out = 16'(1687);
			3398: out = 16'(-219);
			3399: out = 16'(-420);
			3400: out = 16'(-2604);
			3401: out = 16'(-1666);
			3402: out = 16'(2263);
			3403: out = 16'(2335);
			3404: out = 16'(1304);
			3405: out = 16'(519);
			3406: out = 16'(-1081);
			3407: out = 16'(940);
			3408: out = 16'(1449);
			3409: out = 16'(-1021);
			3410: out = 16'(-2488);
			3411: out = 16'(-848);
			3412: out = 16'(2867);
			3413: out = 16'(1763);
			3414: out = 16'(536);
			3415: out = 16'(-1485);
			3416: out = 16'(-87);
			3417: out = 16'(-2474);
			3418: out = 16'(-507);
			3419: out = 16'(1903);
			3420: out = 16'(1510);
			3421: out = 16'(360);
			3422: out = 16'(-750);
			3423: out = 16'(-1074);
			3424: out = 16'(-962);
			3425: out = 16'(-466);
			3426: out = 16'(317);
			3427: out = 16'(-1654);
			3428: out = 16'(1078);
			3429: out = 16'(1924);
			3430: out = 16'(-490);
			3431: out = 16'(-1305);
			3432: out = 16'(-1058);
			3433: out = 16'(569);
			3434: out = 16'(-986);
			3435: out = 16'(1079);
			3436: out = 16'(998);
			3437: out = 16'(-1640);
			3438: out = 16'(1886);
			3439: out = 16'(1528);
			3440: out = 16'(-449);
			3441: out = 16'(-2083);
			3442: out = 16'(-869);
			3443: out = 16'(639);
			3444: out = 16'(-530);
			3445: out = 16'(2546);
			3446: out = 16'(-184);
			3447: out = 16'(-3019);
			3448: out = 16'(-604);
			3449: out = 16'(1279);
			3450: out = 16'(1872);
			3451: out = 16'(-834);
			3452: out = 16'(245);
			3453: out = 16'(-192);
			3454: out = 16'(185);
			3455: out = 16'(-2417);
			3456: out = 16'(1062);
			3457: out = 16'(1845);
			3458: out = 16'(1274);
			3459: out = 16'(-1706);
			3460: out = 16'(-140);
			3461: out = 16'(1340);
			3462: out = 16'(-897);
			3463: out = 16'(-1723);
			3464: out = 16'(-777);
			3465: out = 16'(1315);
			3466: out = 16'(1203);
			3467: out = 16'(-1655);
			3468: out = 16'(-4445);
			3469: out = 16'(-4110);
			3470: out = 16'(1122);
			3471: out = 16'(3557);
			3472: out = 16'(1287);
			3473: out = 16'(1909);
			3474: out = 16'(1065);
			3475: out = 16'(957);
			3476: out = 16'(-1903);
			3477: out = 16'(-90);
			3478: out = 16'(221);
			3479: out = 16'(326);
			3480: out = 16'(-1233);
			3481: out = 16'(30);
			3482: out = 16'(1679);
			3483: out = 16'(3120);
			3484: out = 16'(-123);
			3485: out = 16'(-1448);
			3486: out = 16'(79);
			3487: out = 16'(-500);
			3488: out = 16'(1691);
			3489: out = 16'(2010);
			3490: out = 16'(247);
			3491: out = 16'(-586);
			3492: out = 16'(403);
			3493: out = 16'(2050);
			3494: out = 16'(-214);
			3495: out = 16'(-608);
			3496: out = 16'(-610);
			3497: out = 16'(-675);
			3498: out = 16'(1304);
			3499: out = 16'(1403);
			3500: out = 16'(251);
			3501: out = 16'(-1727);
			3502: out = 16'(-255);
			3503: out = 16'(1611);
			3504: out = 16'(1037);
			3505: out = 16'(-30);
			3506: out = 16'(-682);
			3507: out = 16'(644);
			3508: out = 16'(-1739);
			3509: out = 16'(1013);
			3510: out = 16'(1568);
			3511: out = 16'(269);
			3512: out = 16'(-3068);
			3513: out = 16'(-2753);
			3514: out = 16'(-94);
			3515: out = 16'(1777);
			3516: out = 16'(982);
			3517: out = 16'(-67);
			3518: out = 16'(241);
			3519: out = 16'(256);
			3520: out = 16'(-31);
			3521: out = 16'(-404);
			3522: out = 16'(484);
			3523: out = 16'(1389);
			3524: out = 16'(1584);
			3525: out = 16'(1018);
			3526: out = 16'(-2859);
			3527: out = 16'(-3221);
			3528: out = 16'(-738);
			3529: out = 16'(1903);
			3530: out = 16'(2039);
			3531: out = 16'(282);
			3532: out = 16'(-2770);
			3533: out = 16'(184);
			3534: out = 16'(-983);
			3535: out = 16'(-2872);
			3536: out = 16'(1291);
			3537: out = 16'(803);
			3538: out = 16'(361);
			3539: out = 16'(-1106);
			3540: out = 16'(891);
			3541: out = 16'(306);
			3542: out = 16'(-337);
			3543: out = 16'(1734);
			3544: out = 16'(587);
			3545: out = 16'(-244);
			3546: out = 16'(-1008);
			3547: out = 16'(1131);
			3548: out = 16'(-46);
			3549: out = 16'(-1727);
			3550: out = 16'(1100);
			3551: out = 16'(-92);
			3552: out = 16'(407);
			3553: out = 16'(1569);
			3554: out = 16'(176);
			3555: out = 16'(-399);
			3556: out = 16'(-2);
			3557: out = 16'(1321);
			3558: out = 16'(142);
			3559: out = 16'(-2778);
			3560: out = 16'(-6070);
			3561: out = 16'(-2816);
			3562: out = 16'(665);
			3563: out = 16'(2797);
			3564: out = 16'(620);
			3565: out = 16'(-292);
			3566: out = 16'(-2311);
			3567: out = 16'(-3142);
			3568: out = 16'(-961);
			3569: out = 16'(1518);
			3570: out = 16'(1883);
			3571: out = 16'(-634);
			3572: out = 16'(-2074);
			3573: out = 16'(-2236);
			3574: out = 16'(-881);
			3575: out = 16'(801);
			3576: out = 16'(1267);
			3577: out = 16'(344);
			3578: out = 16'(-2174);
			3579: out = 16'(-815);
			3580: out = 16'(137);
			3581: out = 16'(215);
			3582: out = 16'(1192);
			3583: out = 16'(-368);
			3584: out = 16'(-2252);
			3585: out = 16'(-1230);
			3586: out = 16'(-2478);
			3587: out = 16'(-928);
			3588: out = 16'(844);
			3589: out = 16'(1642);
			3590: out = 16'(-554);
			3591: out = 16'(-2079);
			3592: out = 16'(-1693);
			3593: out = 16'(951);
			3594: out = 16'(610);
			3595: out = 16'(-1518);
			3596: out = 16'(-493);
			3597: out = 16'(749);
			3598: out = 16'(1585);
			3599: out = 16'(1239);
			3600: out = 16'(-1320);
			3601: out = 16'(-710);
			3602: out = 16'(1891);
			3603: out = 16'(-622);
			3604: out = 16'(25);
			3605: out = 16'(170);
			3606: out = 16'(-784);
			3607: out = 16'(1469);
			3608: out = 16'(1263);
			3609: out = 16'(-147);
			3610: out = 16'(-5644);
			3611: out = 16'(-2183);
			3612: out = 16'(1078);
			3613: out = 16'(127);
			3614: out = 16'(1123);
			3615: out = 16'(1887);
			3616: out = 16'(2180);
			3617: out = 16'(-3882);
			3618: out = 16'(-4056);
			3619: out = 16'(-1854);
			3620: out = 16'(1795);
			3621: out = 16'(2576);
			3622: out = 16'(1848);
			3623: out = 16'(-91);
			3624: out = 16'(-4195);
			3625: out = 16'(-1863);
			3626: out = 16'(728);
			3627: out = 16'(1055);
			3628: out = 16'(-143);
			3629: out = 16'(-100);
			3630: out = 16'(1189);
			3631: out = 16'(980);
			3632: out = 16'(1246);
			3633: out = 16'(-241);
			3634: out = 16'(-2974);
			3635: out = 16'(1469);
			3636: out = 16'(1789);
			3637: out = 16'(499);
			3638: out = 16'(-1320);
			3639: out = 16'(-130);
			3640: out = 16'(1239);
			3641: out = 16'(1574);
			3642: out = 16'(786);
			3643: out = 16'(274);
			3644: out = 16'(277);
			3645: out = 16'(1600);
			3646: out = 16'(1092);
			3647: out = 16'(1631);
			3648: out = 16'(2246);
			3649: out = 16'(1995);
			3650: out = 16'(-515);
			3651: out = 16'(-2137);
			3652: out = 16'(970);
			3653: out = 16'(993);
			3654: out = 16'(110);
			3655: out = 16'(-2170);
			3656: out = 16'(524);
			3657: out = 16'(1193);
			3658: out = 16'(1391);
			3659: out = 16'(-379);
			3660: out = 16'(994);
			3661: out = 16'(1404);
			3662: out = 16'(1238);
			3663: out = 16'(-519);
			3664: out = 16'(-537);
			3665: out = 16'(275);
			3666: out = 16'(1200);
			3667: out = 16'(1295);
			3668: out = 16'(860);
			3669: out = 16'(337);
			3670: out = 16'(237);
			3671: out = 16'(636);
			3672: out = 16'(778);
			3673: out = 16'(-469);
			3674: out = 16'(895);
			3675: out = 16'(1395);
			3676: out = 16'(1204);
			3677: out = 16'(-727);
			3678: out = 16'(-232);
			3679: out = 16'(655);
			3680: out = 16'(371);
			3681: out = 16'(240);
			3682: out = 16'(-426);
			3683: out = 16'(-400);
			3684: out = 16'(-528);
			3685: out = 16'(1572);
			3686: out = 16'(2220);
			3687: out = 16'(304);
			3688: out = 16'(-2216);
			3689: out = 16'(-3678);
			3690: out = 16'(-2362);
			3691: out = 16'(1104);
			3692: out = 16'(1983);
			3693: out = 16'(893);
			3694: out = 16'(160);
			3695: out = 16'(-1947);
			3696: out = 16'(-1100);
			3697: out = 16'(499);
			3698: out = 16'(1675);
			3699: out = 16'(626);
			3700: out = 16'(-686);
			3701: out = 16'(-2660);
			3702: out = 16'(1736);
			3703: out = 16'(1514);
			3704: out = 16'(-529);
			3705: out = 16'(-3031);
			3706: out = 16'(-26);
			3707: out = 16'(1945);
			3708: out = 16'(-158);
			3709: out = 16'(-92);
			3710: out = 16'(-1060);
			3711: out = 16'(-893);
			3712: out = 16'(905);
			3713: out = 16'(-96);
			3714: out = 16'(-804);
			3715: out = 16'(96);
			3716: out = 16'(-956);
			3717: out = 16'(-933);
			3718: out = 16'(-449);
			3719: out = 16'(1027);
			3720: out = 16'(781);
			3721: out = 16'(-166);
			3722: out = 16'(-1159);
			3723: out = 16'(-1321);
			3724: out = 16'(-65);
			3725: out = 16'(579);
			3726: out = 16'(-1516);
			3727: out = 16'(-2297);
			3728: out = 16'(-1232);
			3729: out = 16'(1750);
			3730: out = 16'(823);
			3731: out = 16'(419);
			3732: out = 16'(-286);
			3733: out = 16'(-67);
			3734: out = 16'(-210);
			3735: out = 16'(-49);
			3736: out = 16'(-70);
			3737: out = 16'(-935);
			3738: out = 16'(-1040);
			3739: out = 16'(-343);
			3740: out = 16'(1663);
			3741: out = 16'(-451);
			3742: out = 16'(-1704);
			3743: out = 16'(-1084);
			3744: out = 16'(-768);
			3745: out = 16'(437);
			3746: out = 16'(735);
			3747: out = 16'(-343);
			3748: out = 16'(-511);
			3749: out = 16'(-625);
			3750: out = 16'(-568);
			3751: out = 16'(-986);
			3752: out = 16'(-395);
			3753: out = 16'(316);
			3754: out = 16'(29);
			3755: out = 16'(392);
			3756: out = 16'(387);
			3757: out = 16'(593);
			3758: out = 16'(-1085);
			3759: out = 16'(-700);
			3760: out = 16'(-674);
			3761: out = 16'(-2186);
			3762: out = 16'(-2005);
			3763: out = 16'(-1165);
			3764: out = 16'(303);
			3765: out = 16'(1961);
			3766: out = 16'(1895);
			3767: out = 16'(532);
			3768: out = 16'(-2028);
			3769: out = 16'(-827);
			3770: out = 16'(-126);
			3771: out = 16'(-400);
			3772: out = 16'(-1225);
			3773: out = 16'(-594);
			3774: out = 16'(916);
			3775: out = 16'(1062);
			3776: out = 16'(1612);
			3777: out = 16'(-145);
			3778: out = 16'(-2030);
			3779: out = 16'(-2734);
			3780: out = 16'(-652);
			3781: out = 16'(546);
			3782: out = 16'(-1686);
			3783: out = 16'(-119);
			3784: out = 16'(595);
			3785: out = 16'(960);
			3786: out = 16'(-1026);
			3787: out = 16'(-1078);
			3788: out = 16'(-504);
			3789: out = 16'(881);
			3790: out = 16'(344);
			3791: out = 16'(339);
			3792: out = 16'(261);
			3793: out = 16'(-924);
			3794: out = 16'(-458);
			3795: out = 16'(-95);
			3796: out = 16'(-718);
			3797: out = 16'(588);
			3798: out = 16'(674);
			3799: out = 16'(419);
			3800: out = 16'(1082);
			3801: out = 16'(856);
			3802: out = 16'(1156);
			3803: out = 16'(2139);
			3804: out = 16'(-1137);
			3805: out = 16'(-2964);
			3806: out = 16'(-3118);
			3807: out = 16'(320);
			3808: out = 16'(382);
			3809: out = 16'(833);
			3810: out = 16'(2201);
			3811: out = 16'(-376);
			3812: out = 16'(-1390);
			3813: out = 16'(-1417);
			3814: out = 16'(1296);
			3815: out = 16'(104);
			3816: out = 16'(-115);
			3817: out = 16'(1303);
			3818: out = 16'(206);
			3819: out = 16'(415);
			3820: out = 16'(628);
			3821: out = 16'(1001);
			3822: out = 16'(711);
			3823: out = 16'(521);
			3824: out = 16'(100);
			3825: out = 16'(1099);
			3826: out = 16'(451);
			3827: out = 16'(-76);
			3828: out = 16'(1018);
			3829: out = 16'(942);
			3830: out = 16'(724);
			3831: out = 16'(92);
			3832: out = 16'(-84);
			3833: out = 16'(-407);
			3834: out = 16'(-108);
			3835: out = 16'(1580);
			3836: out = 16'(1525);
			3837: out = 16'(875);
			3838: out = 16'(-953);
			3839: out = 16'(-117);
			3840: out = 16'(-1245);
			3841: out = 16'(-1317);
			3842: out = 16'(-757);
			3843: out = 16'(1596);
			3844: out = 16'(1371);
			3845: out = 16'(-79);
			3846: out = 16'(-2438);
			3847: out = 16'(-328);
			3848: out = 16'(1889);
			3849: out = 16'(1291);
			3850: out = 16'(-1245);
			3851: out = 16'(-1295);
			3852: out = 16'(1901);
			3853: out = 16'(648);
			3854: out = 16'(879);
			3855: out = 16'(-25);
			3856: out = 16'(168);
			3857: out = 16'(-74);
			3858: out = 16'(684);
			3859: out = 16'(513);
			3860: out = 16'(-441);
			3861: out = 16'(-1764);
			3862: out = 16'(-1130);
			3863: out = 16'(1487);
			3864: out = 16'(1271);
			3865: out = 16'(664);
			3866: out = 16'(328);
			3867: out = 16'(-1857);
			3868: out = 16'(3);
			3869: out = 16'(1397);
			3870: out = 16'(1067);
			3871: out = 16'(-472);
			3872: out = 16'(-80);
			3873: out = 16'(1562);
			3874: out = 16'(-224);
			3875: out = 16'(19);
			3876: out = 16'(-685);
			3877: out = 16'(-2817);
			3878: out = 16'(870);
			3879: out = 16'(2229);
			3880: out = 16'(1535);
			3881: out = 16'(-3408);
			3882: out = 16'(-1453);
			3883: out = 16'(1390);
			3884: out = 16'(1495);
			3885: out = 16'(615);
			3886: out = 16'(-1345);
			3887: out = 16'(-2177);
			3888: out = 16'(-2518);
			3889: out = 16'(-408);
			3890: out = 16'(788);
			3891: out = 16'(414);
			3892: out = 16'(48);
			3893: out = 16'(-395);
			3894: out = 16'(-415);
			3895: out = 16'(-6);
			3896: out = 16'(-5);
			3897: out = 16'(133);
			3898: out = 16'(670);
			3899: out = 16'(-469);
			3900: out = 16'(-513);
			3901: out = 16'(-124);
			3902: out = 16'(67);
			3903: out = 16'(255);
			3904: out = 16'(-60);
			3905: out = 16'(-776);
			3906: out = 16'(-36);
			3907: out = 16'(397);
			3908: out = 16'(658);
			3909: out = 16'(490);
			3910: out = 16'(187);
			3911: out = 16'(-321);
			3912: out = 16'(-601);
			3913: out = 16'(-583);
			3914: out = 16'(-137);
			3915: out = 16'(131);
			3916: out = 16'(137);
			3917: out = 16'(-553);
			3918: out = 16'(-945);
			3919: out = 16'(-734);
			3920: out = 16'(93);
			3921: out = 16'(352);
			3922: out = 16'(53);
			3923: out = 16'(-695);
			3924: out = 16'(-168);
			3925: out = 16'(304);
			3926: out = 16'(262);
			3927: out = 16'(-198);
			3928: out = 16'(-604);
			3929: out = 16'(-632);
			3930: out = 16'(-442);
			3931: out = 16'(372);
			3932: out = 16'(693);
			3933: out = 16'(391);
			3934: out = 16'(1016);
			3935: out = 16'(393);
			3936: out = 16'(-529);
			3937: out = 16'(-1636);
			3938: out = 16'(-1263);
			3939: out = 16'(-602);
			3940: out = 16'(164);
			3941: out = 16'(-724);
			3942: out = 16'(440);
			3943: out = 16'(1026);
			3944: out = 16'(-854);
			3945: out = 16'(-930);
			3946: out = 16'(-1098);
			3947: out = 16'(-354);
			3948: out = 16'(-2262);
			3949: out = 16'(-477);
			3950: out = 16'(908);
			3951: out = 16'(1335);
			3952: out = 16'(-1300);
			3953: out = 16'(-2026);
			3954: out = 16'(-544);
			3955: out = 16'(1477);
			3956: out = 16'(993);
			3957: out = 16'(-871);
			3958: out = 16'(-2264);
			3959: out = 16'(-1759);
			3960: out = 16'(32);
			3961: out = 16'(1324);
			3962: out = 16'(561);
			3963: out = 16'(-291);
			3964: out = 16'(-1155);
			3965: out = 16'(-1485);
			3966: out = 16'(167);
			3967: out = 16'(1290);
			3968: out = 16'(1152);
			3969: out = 16'(427);
			3970: out = 16'(-1059);
			3971: out = 16'(-1280);
			3972: out = 16'(217);
			3973: out = 16'(363);
			3974: out = 16'(-19);
			3975: out = 16'(-688);
			3976: out = 16'(928);
			3977: out = 16'(796);
			3978: out = 16'(924);
			3979: out = 16'(823);
			3980: out = 16'(417);
			3981: out = 16'(54);
			3982: out = 16'(-248);
			3983: out = 16'(-3580);
			3984: out = 16'(-881);
			3985: out = 16'(1334);
			3986: out = 16'(1065);
			3987: out = 16'(908);
			3988: out = 16'(-305);
			3989: out = 16'(-970);
			3990: out = 16'(-644);
			3991: out = 16'(381);
			3992: out = 16'(835);
			3993: out = 16'(85);
			3994: out = 16'(406);
			3995: out = 16'(-52);
			3996: out = 16'(-95);
			3997: out = 16'(-303);
			3998: out = 16'(555);
			3999: out = 16'(598);
			4000: out = 16'(597);
			4001: out = 16'(-998);
			4002: out = 16'(341);
			4003: out = 16'(1706);
			4004: out = 16'(965);
			4005: out = 16'(-356);
			4006: out = 16'(-576);
			4007: out = 16'(933);
			4008: out = 16'(812);
			4009: out = 16'(205);
			4010: out = 16'(-767);
			4011: out = 16'(-268);
			4012: out = 16'(421);
			4013: out = 16'(984);
			4014: out = 16'(518);
			4015: out = 16'(278);
			4016: out = 16'(-74);
			4017: out = 16'(211);
			4018: out = 16'(765);
			4019: out = 16'(305);
			4020: out = 16'(-302);
			4021: out = 16'(-376);
			4022: out = 16'(-757);
			4023: out = 16'(-601);
			4024: out = 16'(-179);
			4025: out = 16'(1751);
			4026: out = 16'(-308);
			4027: out = 16'(-1226);
			4028: out = 16'(-1004);
			4029: out = 16'(1079);
			4030: out = 16'(889);
			4031: out = 16'(100);
			4032: out = 16'(416);
			4033: out = 16'(-238);
			4034: out = 16'(-205);
			4035: out = 16'(11);
			4036: out = 16'(285);
			4037: out = 16'(18);
			4038: out = 16'(-233);
			4039: out = 16'(170);
			4040: out = 16'(670);
			4041: out = 16'(1030);
			4042: out = 16'(384);
			4043: out = 16'(93);
			4044: out = 16'(-1985);
			4045: out = 16'(-2140);
			4046: out = 16'(1532);
			4047: out = 16'(1341);
			4048: out = 16'(999);
			4049: out = 16'(-163);
			4050: out = 16'(-1592);
			4051: out = 16'(-1091);
			4052: out = 16'(193);
			4053: out = 16'(-132);
			4054: out = 16'(1273);
			4055: out = 16'(355);
			4056: out = 16'(-885);
			4057: out = 16'(-412);
			4058: out = 16'(230);
			4059: out = 16'(558);
			4060: out = 16'(345);
			4061: out = 16'(-642);
			4062: out = 16'(-265);
			4063: out = 16'(625);
			4064: out = 16'(-1714);
			4065: out = 16'(-785);
			4066: out = 16'(372);
			4067: out = 16'(1072);
			4068: out = 16'(490);
			4069: out = 16'(-63);
			4070: out = 16'(-316);
			4071: out = 16'(-1333);
			4072: out = 16'(15);
			4073: out = 16'(849);
			4074: out = 16'(442);
			4075: out = 16'(153);
			4076: out = 16'(277);
			4077: out = 16'(607);
			4078: out = 16'(-965);
			4079: out = 16'(-661);
			4080: out = 16'(-593);
			4081: out = 16'(-635);
			4082: out = 16'(117);
			4083: out = 16'(444);
			4084: out = 16'(386);
			4085: out = 16'(103);
			4086: out = 16'(32);
			4087: out = 16'(-341);
			4088: out = 16'(-1330);
			4089: out = 16'(-74);
			4090: out = 16'(341);
			4091: out = 16'(423);
			4092: out = 16'(-1208);
			4093: out = 16'(-287);
			4094: out = 16'(87);
			4095: out = 16'(110);
			4096: out = 16'(-1237);
			4097: out = 16'(-638);
			4098: out = 16'(177);
			4099: out = 16'(-408);
			4100: out = 16'(-673);
			4101: out = 16'(-67);
			4102: out = 16'(1363);
			4103: out = 16'(-219);
			4104: out = 16'(-986);
			4105: out = 16'(-1225);
			4106: out = 16'(651);
			4107: out = 16'(192);
			4108: out = 16'(292);
			4109: out = 16'(480);
			4110: out = 16'(-171);
			4111: out = 16'(-483);
			4112: out = 16'(-640);
			4113: out = 16'(-772);
			4114: out = 16'(-445);
			4115: out = 16'(160);
			4116: out = 16'(621);
			4117: out = 16'(-1361);
			4118: out = 16'(-1421);
			4119: out = 16'(-597);
			4120: out = 16'(-108);
			4121: out = 16'(1055);
			4122: out = 16'(608);
			4123: out = 16'(-578);
			4124: out = 16'(-579);
			4125: out = 16'(-338);
			4126: out = 16'(-108);
			4127: out = 16'(-538);
			4128: out = 16'(31);
			4129: out = 16'(421);
			4130: out = 16'(539);
			4131: out = 16'(727);
			4132: out = 16'(-319);
			4133: out = 16'(-1022);
			4134: out = 16'(-265);
			4135: out = 16'(728);
			4136: out = 16'(1367);
			4137: out = 16'(1052);
			4138: out = 16'(1509);
			4139: out = 16'(509);
			4140: out = 16'(-264);
			4141: out = 16'(-1041);
			4142: out = 16'(281);
			4143: out = 16'(444);
			4144: out = 16'(58);
			4145: out = 16'(211);
			4146: out = 16'(524);
			4147: out = 16'(675);
			4148: out = 16'(162);
			4149: out = 16'(126);
			4150: out = 16'(-341);
			4151: out = 16'(-647);
			4152: out = 16'(-11);
			4153: out = 16'(375);
			4154: out = 16'(402);
			4155: out = 16'(-621);
			4156: out = 16'(783);
			4157: out = 16'(560);
			4158: out = 16'(73);
			4159: out = 16'(-473);
			4160: out = 16'(802);
			4161: out = 16'(1165);
			4162: out = 16'(-126);
			4163: out = 16'(369);
			4164: out = 16'(366);
			4165: out = 16'(425);
			4166: out = 16'(534);
			4167: out = 16'(113);
			4168: out = 16'(-223);
			4169: out = 16'(-273);
			4170: out = 16'(356);
			4171: out = 16'(441);
			4172: out = 16'(375);
			4173: out = 16'(247);
			4174: out = 16'(445);
			4175: out = 16'(302);
			4176: out = 16'(169);
			4177: out = 16'(-2010);
			4178: out = 16'(-1527);
			4179: out = 16'(163);
			4180: out = 16'(1336);
			4181: out = 16'(959);
			4182: out = 16'(302);
			4183: out = 16'(-208);
			4184: out = 16'(133);
			4185: out = 16'(-1173);
			4186: out = 16'(-2256);
			4187: out = 16'(484);
			4188: out = 16'(663);
			4189: out = 16'(1245);
			4190: out = 16'(936);
			4191: out = 16'(571);
			4192: out = 16'(-777);
			4193: out = 16'(-1302);
			4194: out = 16'(-172);
			4195: out = 16'(343);
			4196: out = 16'(-54);
			4197: out = 16'(-1278);
			4198: out = 16'(-186);
			4199: out = 16'(319);
			4200: out = 16'(496);
			4201: out = 16'(-1208);
			4202: out = 16'(105);
			4203: out = 16'(554);
			4204: out = 16'(519);
			4205: out = 16'(-775);
			4206: out = 16'(-472);
			4207: out = 16'(-64);
			4208: out = 16'(-375);
			4209: out = 16'(-632);
			4210: out = 16'(-188);
			4211: out = 16'(703);
			4212: out = 16'(-838);
			4213: out = 16'(-782);
			4214: out = 16'(-292);
			4215: out = 16'(223);
			4216: out = 16'(153);
			4217: out = 16'(-378);
			4218: out = 16'(-747);
			4219: out = 16'(-366);
			4220: out = 16'(227);
			4221: out = 16'(44);
			4222: out = 16'(-939);
			4223: out = 16'(-1113);
			4224: out = 16'(-292);
			4225: out = 16'(574);
			4226: out = 16'(844);
			4227: out = 16'(-492);
			4228: out = 16'(-1052);
			4229: out = 16'(214);
			4230: out = 16'(607);
			4231: out = 16'(-351);
			4232: out = 16'(-1969);
			4233: out = 16'(-338);
			4234: out = 16'(472);
			4235: out = 16'(755);
			4236: out = 16'(-305);
			4237: out = 16'(-692);
			4238: out = 16'(-587);
			4239: out = 16'(147);
			4240: out = 16'(28);
			4241: out = 16'(-130);
			4242: out = 16'(-47);
			4243: out = 16'(892);
			4244: out = 16'(412);
			4245: out = 16'(-109);
			4246: out = 16'(-654);
			4247: out = 16'(246);
			4248: out = 16'(445);
			4249: out = 16'(422);
			4250: out = 16'(-55);
			4251: out = 16'(230);
			4252: out = 16'(589);
			4253: out = 16'(701);
			4254: out = 16'(-1249);
			4255: out = 16'(-1243);
			4256: out = 16'(-603);
			4257: out = 16'(634);
			4258: out = 16'(12);
			4259: out = 16'(-21);
			4260: out = 16'(105);
			4261: out = 16'(1147);
			4262: out = 16'(160);
			4263: out = 16'(-352);
			4264: out = 16'(217);
			4265: out = 16'(-1147);
			4266: out = 16'(-968);
			4267: out = 16'(-255);
			4268: out = 16'(6);
			4269: out = 16'(675);
			4270: out = 16'(882);
			4271: out = 16'(515);
			4272: out = 16'(296);
			4273: out = 16'(-684);
			4274: out = 16'(-1511);
			4275: out = 16'(-485);
			4276: out = 16'(-683);
			4277: out = 16'(-328);
			4278: out = 16'(208);
			4279: out = 16'(532);
			4280: out = 16'(111);
			4281: out = 16'(-509);
			4282: out = 16'(-486);
			4283: out = 16'(-222);
			4284: out = 16'(177);
			4285: out = 16'(226);
			4286: out = 16'(682);
			4287: out = 16'(170);
			4288: out = 16'(-104);
			4289: out = 16'(806);
			4290: out = 16'(417);
			4291: out = 16'(-20);
			4292: out = 16'(-571);
			4293: out = 16'(753);
			4294: out = 16'(766);
			4295: out = 16'(325);
			4296: out = 16'(-796);
			4297: out = 16'(70);
			4298: out = 16'(605);
			4299: out = 16'(584);
			4300: out = 16'(-797);
			4301: out = 16'(-871);
			4302: out = 16'(-440);
			4303: out = 16'(-452);
			4304: out = 16'(399);
			4305: out = 16'(443);
			4306: out = 16'(-119);
			4307: out = 16'(636);
			4308: out = 16'(55);
			4309: out = 16'(-496);
			4310: out = 16'(-878);
			4311: out = 16'(72);
			4312: out = 16'(285);
			4313: out = 16'(-137);
			4314: out = 16'(-376);
			4315: out = 16'(139);
			4316: out = 16'(634);
			4317: out = 16'(-222);
			4318: out = 16'(505);
			4319: out = 16'(293);
			4320: out = 16'(-194);
			4321: out = 16'(-2419);
			4322: out = 16'(-1447);
			4323: out = 16'(343);
			4324: out = 16'(1100);
			4325: out = 16'(940);
			4326: out = 16'(-9);
			4327: out = 16'(-651);
			4328: out = 16'(-369);
			4329: out = 16'(191);
			4330: out = 16'(376);
			4331: out = 16'(202);
			4332: out = 16'(-408);
			4333: out = 16'(-152);
			4334: out = 16'(259);
			4335: out = 16'(-1327);
			4336: out = 16'(-1431);
			4337: out = 16'(-874);
			4338: out = 16'(319);
			4339: out = 16'(552);
			4340: out = 16'(607);
			4341: out = 16'(362);
			4342: out = 16'(-589);
			4343: out = 16'(-219);
			4344: out = 16'(-124);
			4345: out = 16'(-865);
			4346: out = 16'(-588);
			4347: out = 16'(-333);
			4348: out = 16'(247);
			4349: out = 16'(292);
			4350: out = 16'(718);
			4351: out = 16'(550);
			4352: out = 16'(19);
			4353: out = 16'(-187);
			4354: out = 16'(-439);
			4355: out = 16'(-560);
			4356: out = 16'(32);
			4357: out = 16'(-279);
			4358: out = 16'(-378);
			4359: out = 16'(-119);
			4360: out = 16'(26);
			4361: out = 16'(61);
			4362: out = 16'(-19);
			4363: out = 16'(91);
			4364: out = 16'(-10);
			4365: out = 16'(20);
			4366: out = 16'(59);
			4367: out = 16'(6);
			4368: out = 16'(-131);
			4369: out = 16'(-209);
			4370: out = 16'(271);
			4371: out = 16'(-116);
			4372: out = 16'(-216);
			4373: out = 16'(47);
			4374: out = 16'(179);
			4375: out = 16'(127);
			4376: out = 16'(64);
			4377: out = 16'(1031);
			4378: out = 16'(-268);
			4379: out = 16'(-668);
			4380: out = 16'(-146);
			4381: out = 16'(-105);
			4382: out = 16'(179);
			4383: out = 16'(138);
			4384: out = 16'(-190);
			4385: out = 16'(60);
			4386: out = 16'(-155);
			4387: out = 16'(-1024);
			4388: out = 16'(723);
			4389: out = 16'(-136);
			4390: out = 16'(-895);
			4391: out = 16'(-154);
			4392: out = 16'(388);
			4393: out = 16'(718);
			4394: out = 16'(276);
			4395: out = 16'(738);
			4396: out = 16'(-352);
			4397: out = 16'(-942);
			4398: out = 16'(63);
			4399: out = 16'(294);
			4400: out = 16'(639);
			4401: out = 16'(636);
			4402: out = 16'(370);
			4403: out = 16'(98);
			4404: out = 16'(-227);
			4405: out = 16'(-1377);
			4406: out = 16'(91);
			4407: out = 16'(473);
			4408: out = 16'(209);
			4409: out = 16'(-233);
			4410: out = 16'(30);
			4411: out = 16'(355);
			4412: out = 16'(245);
			4413: out = 16'(-212);
			4414: out = 16'(-171);
			4415: out = 16'(374);
			4416: out = 16'(-72);
			4417: out = 16'(-105);
			4418: out = 16'(-306);
			4419: out = 16'(224);
			4420: out = 16'(-170);
			4421: out = 16'(510);
			4422: out = 16'(871);
			4423: out = 16'(-233);
			4424: out = 16'(-1087);
			4425: out = 16'(-1200);
			4426: out = 16'(-463);
			4427: out = 16'(171);
			4428: out = 16'(286);
			4429: out = 16'(163);
			4430: out = 16'(-967);
			4431: out = 16'(234);
			4432: out = 16'(657);
			4433: out = 16'(-306);
			4434: out = 16'(-995);
			4435: out = 16'(-668);
			4436: out = 16'(411);
			4437: out = 16'(336);
			4438: out = 16'(-106);
			4439: out = 16'(-676);
			4440: out = 16'(-265);
			4441: out = 16'(-128);
			4442: out = 16'(279);
			4443: out = 16'(327);
			4444: out = 16'(269);
			4445: out = 16'(-72);
			4446: out = 16'(-61);
			4447: out = 16'(404);
			4448: out = 16'(-413);
			4449: out = 16'(-123);
			4450: out = 16'(433);
			4451: out = 16'(56);
			4452: out = 16'(23);
			4453: out = 16'(87);
			4454: out = 16'(722);
			4455: out = 16'(-177);
			4456: out = 16'(-494);
			4457: out = 16'(-668);
			4458: out = 16'(566);
			4459: out = 16'(-201);
			4460: out = 16'(-88);
			4461: out = 16'(459);
			4462: out = 16'(1051);
			4463: out = 16'(-204);
			4464: out = 16'(-1426);
			4465: out = 16'(513);
			4466: out = 16'(56);
			4467: out = 16'(-237);
			4468: out = 16'(-944);
			4469: out = 16'(552);
			4470: out = 16'(457);
			4471: out = 16'(49);
			4472: out = 16'(-326);
			4473: out = 16'(-187);
			4474: out = 16'(69);
			4475: out = 16'(178);
			4476: out = 16'(62);
			4477: out = 16'(-161);
			4478: out = 16'(-268);
			4479: out = 16'(-214);
			4480: out = 16'(92);
			4481: out = 16'(229);
			4482: out = 16'(140);
			4483: out = 16'(-711);
			4484: out = 16'(-379);
			4485: out = 16'(71);
			4486: out = 16'(-1185);
			4487: out = 16'(-83);
			4488: out = 16'(-244);
			4489: out = 16'(-1083);
			4490: out = 16'(159);
			4491: out = 16'(612);
			4492: out = 16'(621);
			4493: out = 16'(-650);
			4494: out = 16'(38);
			4495: out = 16'(169);
			4496: out = 16'(-49);
			4497: out = 16'(-1342);
			4498: out = 16'(-873);
			4499: out = 16'(128);
			4500: out = 16'(422);
			4501: out = 16'(626);
			4502: out = 16'(37);
			4503: out = 16'(-543);
			4504: out = 16'(-22);
			4505: out = 16'(336);
			4506: out = 16'(327);
			4507: out = 16'(-202);
			4508: out = 16'(-21);
			4509: out = 16'(196);
			4510: out = 16'(346);
			4511: out = 16'(41);
			4512: out = 16'(-726);
			4513: out = 16'(-1021);
			4514: out = 16'(476);
			4515: out = 16'(-874);
			4516: out = 16'(-335);
			4517: out = 16'(640);
			4518: out = 16'(-309);
			4519: out = 16'(-253);
			4520: out = 16'(-62);
			4521: out = 16'(541);
			4522: out = 16'(-650);
			4523: out = 16'(-1160);
			4524: out = 16'(-881);
			4525: out = 16'(544);
			4526: out = 16'(748);
			4527: out = 16'(262);
			4528: out = 16'(-725);
			4529: out = 16'(-682);
			4530: out = 16'(-565);
			4531: out = 16'(-265);
			4532: out = 16'(579);
			4533: out = 16'(285);
			4534: out = 16'(-265);
			4535: out = 16'(-935);
			4536: out = 16'(-492);
			4537: out = 16'(-363);
			4538: out = 16'(-414);
			4539: out = 16'(-719);
			4540: out = 16'(-98);
			4541: out = 16'(414);
			4542: out = 16'(488);
			4543: out = 16'(220);
			4544: out = 16'(-110);
			4545: out = 16'(-340);
			4546: out = 16'(-191);
			4547: out = 16'(-453);
			4548: out = 16'(-394);
			4549: out = 16'(-6);
			4550: out = 16'(440);
			4551: out = 16'(468);
			4552: out = 16'(318);
			4553: out = 16'(447);
			4554: out = 16'(293);
			4555: out = 16'(-142);
			4556: out = 16'(-916);
			4557: out = 16'(-58);
			4558: out = 16'(362);
			4559: out = 16'(624);
			4560: out = 16'(238);
			4561: out = 16'(522);
			4562: out = 16'(369);
			4563: out = 16'(123);
			4564: out = 16'(-456);
			4565: out = 16'(-97);
			4566: out = 16'(391);
			4567: out = 16'(414);
			4568: out = 16'(151);
			4569: out = 16'(-139);
			4570: out = 16'(-205);
			4571: out = 16'(-228);
			4572: out = 16'(-55);
			4573: out = 16'(159);
			4574: out = 16'(170);
			4575: out = 16'(171);
			4576: out = 16'(-176);
			4577: out = 16'(-377);
			4578: out = 16'(47);
			4579: out = 16'(451);
			4580: out = 16'(444);
			4581: out = 16'(368);
			4582: out = 16'(-646);
			4583: out = 16'(-335);
			4584: out = 16'(777);
			4585: out = 16'(351);
			4586: out = 16'(163);
			4587: out = 16'(-227);
			4588: out = 16'(-183);
			4589: out = 16'(-4);
			4590: out = 16'(188);
			4591: out = 16'(104);
			4592: out = 16'(-68);
			4593: out = 16'(-87);
			4594: out = 16'(-63);
			4595: out = 16'(-319);
			4596: out = 16'(-24);
			4597: out = 16'(200);
			4598: out = 16'(384);
			4599: out = 16'(-489);
			4600: out = 16'(-80);
			4601: out = 16'(309);
			4602: out = 16'(324);
			4603: out = 16'(100);
			4604: out = 16'(-62);
			4605: out = 16'(-36);
			4606: out = 16'(-472);
			4607: out = 16'(39);
			4608: out = 16'(296);
			4609: out = 16'(-84);
			4610: out = 16'(258);
			4611: out = 16'(246);
			4612: out = 16'(157);
			4613: out = 16'(69);
			4614: out = 16'(-59);
			4615: out = 16'(-166);
			4616: out = 16'(-96);
			4617: out = 16'(-180);
			4618: out = 16'(157);
			4619: out = 16'(501);
			4620: out = 16'(203);
			4621: out = 16'(34);
			4622: out = 16'(-108);
			4623: out = 16'(105);
			4624: out = 16'(125);
			4625: out = 16'(220);
			4626: out = 16'(25);
			4627: out = 16'(501);
			4628: out = 16'(-545);
			4629: out = 16'(-741);
			4630: out = 16'(57);
			4631: out = 16'(420);
			4632: out = 16'(-34);
			4633: out = 16'(-788);
			4634: out = 16'(474);
			4635: out = 16'(-308);
			4636: out = 16'(-547);
			4637: out = 16'(-433);
			4638: out = 16'(-56);
			4639: out = 16'(-120);
			4640: out = 16'(-206);
			4641: out = 16'(360);
			4642: out = 16'(116);
			4643: out = 16'(55);
			4644: out = 16'(84);
			4645: out = 16'(-184);
			4646: out = 16'(-392);
			4647: out = 16'(-385);
			4648: out = 16'(4);
			4649: out = 16'(177);
			4650: out = 16'(143);
			4651: out = 16'(-96);
			4652: out = 16'(-215);
			4653: out = 16'(-183);
			4654: out = 16'(46);
			4655: out = 16'(233);
			4656: out = 16'(294);
			4657: out = 16'(55);
			4658: out = 16'(-292);
			4659: out = 16'(-316);
			4660: out = 16'(-265);
			4661: out = 16'(-149);
			4662: out = 16'(-30);
			4663: out = 16'(190);
			4664: out = 16'(302);
			4665: out = 16'(276);
			4666: out = 16'(182);
			4667: out = 16'(-149);
			4668: out = 16'(-235);
			4669: out = 16'(485);
			4670: out = 16'(-158);
			4671: out = 16'(-375);
			4672: out = 16'(-220);
			4673: out = 16'(-133);
			4674: out = 16'(66);
			4675: out = 16'(219);
			4676: out = 16'(506);
			4677: out = 16'(-182);
			4678: out = 16'(-603);
			4679: out = 16'(-602);
			4680: out = 16'(127);
			4681: out = 16'(246);
			4682: out = 16'(6);
			4683: out = 16'(-322);
			4684: out = 16'(-371);
			4685: out = 16'(-174);
			4686: out = 16'(-7);
			4687: out = 16'(-36);
			4688: out = 16'(-187);
			4689: out = 16'(-237);
			4690: out = 16'(-123);
			4691: out = 16'(115);
			4692: out = 16'(63);
			4693: out = 16'(-230);
			4694: out = 16'(-796);
			4695: out = 16'(-380);
			4696: out = 16'(421);
			4697: out = 16'(730);
			4698: out = 16'(316);
			4699: out = 16'(-622);
			4700: out = 16'(-1239);
			4701: out = 16'(-120);
			4702: out = 16'(514);
			4703: out = 16'(463);
			4704: out = 16'(-606);
			4705: out = 16'(-476);
			4706: out = 16'(-660);
			4707: out = 16'(-480);
			4708: out = 16'(657);
			4709: out = 16'(622);
			4710: out = 16'(206);
			4711: out = 16'(-228);
			4712: out = 16'(-267);
			4713: out = 16'(-62);
			4714: out = 16'(168);
			4715: out = 16'(110);
			4716: out = 16'(14);
			4717: out = 16'(-43);
			4718: out = 16'(154);
			4719: out = 16'(-44);
			4720: out = 16'(-7);
			4721: out = 16'(-4);
			4722: out = 16'(304);
			4723: out = 16'(-176);
			4724: out = 16'(-321);
			4725: out = 16'(65);
			4726: out = 16'(80);
			4727: out = 16'(-50);
			4728: out = 16'(-366);
			4729: out = 16'(13);
			4730: out = 16'(-393);
			4731: out = 16'(-170);
			4732: out = 16'(389);
			4733: out = 16'(235);
			4734: out = 16'(57);
			4735: out = 16'(-131);
			4736: out = 16'(-447);
			4737: out = 16'(-227);
			4738: out = 16'(-340);
			4739: out = 16'(-755);
			4740: out = 16'(-125);
			4741: out = 16'(300);
			4742: out = 16'(501);
			4743: out = 16'(301);
			4744: out = 16'(-227);
			4745: out = 16'(-669);
			4746: out = 16'(-804);
			4747: out = 16'(333);
			4748: out = 16'(343);
			4749: out = 16'(-92);
			4750: out = 16'(-278);
			4751: out = 16'(-302);
			4752: out = 16'(-5);
			4753: out = 16'(229);
			4754: out = 16'(71);
			4755: out = 16'(-184);
			4756: out = 16'(-262);
			4757: out = 16'(445);
			4758: out = 16'(-275);
			4759: out = 16'(-436);
			4760: out = 16'(-125);
			4761: out = 16'(287);
			4762: out = 16'(184);
			4763: out = 16'(66);
			4764: out = 16'(560);
			4765: out = 16'(-121);
			4766: out = 16'(-376);
			4767: out = 16'(-344);
			4768: out = 16'(351);
			4769: out = 16'(216);
			4770: out = 16'(-83);
			4771: out = 16'(-66);
			4772: out = 16'(-422);
			4773: out = 16'(-377);
			4774: out = 16'(-137);
			4775: out = 16'(553);
			4776: out = 16'(279);
			4777: out = 16'(75);
			4778: out = 16'(530);
			4779: out = 16'(-261);
			4780: out = 16'(-354);
			4781: out = 16'(-119);
			4782: out = 16'(-871);
			4783: out = 16'(-398);
			4784: out = 16'(179);
			4785: out = 16'(507);
			4786: out = 16'(85);
			4787: out = 16'(-154);
			4788: out = 16'(-141);
			4789: out = 16'(-138);
			4790: out = 16'(19);
			4791: out = 16'(55);
			4792: out = 16'(-46);
			4793: out = 16'(58);
			4794: out = 16'(-7);
			4795: out = 16'(-157);
			4796: out = 16'(-385);
			4797: out = 16'(-108);
			4798: out = 16'(294);
			4799: out = 16'(378);
			4800: out = 16'(163);
			4801: out = 16'(-214);
			4802: out = 16'(-469);
			4803: out = 16'(-494);
			4804: out = 16'(64);
			4805: out = 16'(274);
			4806: out = 16'(-186);
			4807: out = 16'(-190);
			4808: out = 16'(-387);
			4809: out = 16'(-275);
			4810: out = 16'(111);
			4811: out = 16'(429);
			4812: out = 16'(109);
			4813: out = 16'(-760);
			4814: out = 16'(-153);
			4815: out = 16'(-172);
			4816: out = 16'(-247);
			4817: out = 16'(569);
			4818: out = 16'(100);
			4819: out = 16'(46);
			4820: out = 16'(269);
			4821: out = 16'(346);
			4822: out = 16'(63);
			4823: out = 16'(-160);
			4824: out = 16'(156);
			4825: out = 16'(257);
			4826: out = 16'(153);
			4827: out = 16'(-108);
			4828: out = 16'(-776);
			4829: out = 16'(-510);
			4830: out = 16'(160);
			4831: out = 16'(591);
			4832: out = 16'(189);
			4833: out = 16'(-355);
			4834: out = 16'(-690);
			4835: out = 16'(110);
			4836: out = 16'(0);
			4837: out = 16'(-302);
			4838: out = 16'(191);
			4839: out = 16'(-333);
			4840: out = 16'(-483);
			4841: out = 16'(-442);
			4842: out = 16'(53);
			4843: out = 16'(137);
			4844: out = 16'(24);
			4845: out = 16'(41);
			4846: out = 16'(-348);
			4847: out = 16'(-207);
			4848: out = 16'(314);
			4849: out = 16'(-42);
			4850: out = 16'(-70);
			4851: out = 16'(-12);
			4852: out = 16'(457);
			4853: out = 16'(-214);
			4854: out = 16'(-205);
			4855: out = 16'(342);
			4856: out = 16'(-124);
			4857: out = 16'(343);
			4858: out = 16'(409);
			4859: out = 16'(-61);
			4860: out = 16'(-522);
			4861: out = 16'(-469);
			4862: out = 16'(95);
			4863: out = 16'(-96);
			4864: out = 16'(84);
			4865: out = 16'(63);
			4866: out = 16'(118);
			4867: out = 16'(-33);
			4868: out = 16'(-1);
			4869: out = 16'(8);
			4870: out = 16'(-22);
			4871: out = 16'(-246);
			4872: out = 16'(-217);
			4873: out = 16'(162);
			4874: out = 16'(147);
			4875: out = 16'(102);
			4876: out = 16'(-17);
			4877: out = 16'(295);
			4878: out = 16'(141);
			4879: out = 16'(-35);
			4880: out = 16'(-391);
			4881: out = 16'(35);
			4882: out = 16'(-2);
			4883: out = 16'(-226);
			4884: out = 16'(75);
			4885: out = 16'(27);
			4886: out = 16'(-14);
			4887: out = 16'(85);
			4888: out = 16'(-57);
			4889: out = 16'(52);
			4890: out = 16'(200);
			4891: out = 16'(214);
			4892: out = 16'(63);
			4893: out = 16'(-123);
			4894: out = 16'(-278);
			4895: out = 16'(-45);
			4896: out = 16'(71);
			4897: out = 16'(102);
			4898: out = 16'(44);
			4899: out = 16'(137);
			4900: out = 16'(51);
			4901: out = 16'(-356);
			4902: out = 16'(109);
			4903: out = 16'(78);
			4904: out = 16'(-109);
			4905: out = 16'(26);
			4906: out = 16'(-218);
			4907: out = 16'(-279);
			4908: out = 16'(-274);
			4909: out = 16'(161);
			4910: out = 16'(124);
			4911: out = 16'(-48);
			4912: out = 16'(-333);
			4913: out = 16'(27);
			4914: out = 16'(162);
			4915: out = 16'(-52);
			4916: out = 16'(-185);
			4917: out = 16'(-24);
			4918: out = 16'(268);
			4919: out = 16'(-306);
			4920: out = 16'(30);
			4921: out = 16'(84);
			4922: out = 16'(113);
			4923: out = 16'(77);
			4924: out = 16'(191);
			4925: out = 16'(100);
			4926: out = 16'(-254);
			4927: out = 16'(-217);
			4928: out = 16'(118);
			4929: out = 16'(414);
			4930: out = 16'(-25);
			4931: out = 16'(-256);
			4932: out = 16'(-211);
			4933: out = 16'(-392);
			4934: out = 16'(269);
			4935: out = 16'(359);
			4936: out = 16'(181);
			4937: out = 16'(-782);
			4938: out = 16'(-528);
			4939: out = 16'(85);
			4940: out = 16'(440);
			4941: out = 16'(-380);
			4942: out = 16'(-645);
			4943: out = 16'(-69);
			4944: out = 16'(156);
			4945: out = 16'(-65);
			4946: out = 16'(-586);
			4947: out = 16'(-298);
			4948: out = 16'(-201);
			4949: out = 16'(168);
			4950: out = 16'(144);
			4951: out = 16'(248);
			4952: out = 16'(-335);
			4953: out = 16'(-631);
			4954: out = 16'(-489);
			4955: out = 16'(116);
			4956: out = 16'(343);
			4957: out = 16'(174);
			4958: out = 16'(-334);
			4959: out = 16'(-218);
			4960: out = 16'(93);
			4961: out = 16'(115);
			4962: out = 16'(102);
			4963: out = 16'(-119);
			4964: out = 16'(-245);
			4965: out = 16'(100);
			4966: out = 16'(-60);
			4967: out = 16'(-378);
			4968: out = 16'(-631);
			4969: out = 16'(-648);
			4970: out = 16'(-328);
			4971: out = 16'(90);
			4972: out = 16'(310);
			4973: out = 16'(380);
			4974: out = 16'(250);
			4975: out = 16'(86);
			4976: out = 16'(-317);
			4977: out = 16'(-326);
			4978: out = 16'(8);
			4979: out = 16'(-297);
			4980: out = 16'(102);
			4981: out = 16'(285);
			4982: out = 16'(233);
			4983: out = 16'(-297);
			4984: out = 16'(-321);
			4985: out = 16'(31);
			4986: out = 16'(177);
			4987: out = 16'(146);
			4988: out = 16'(-47);
			4989: out = 16'(-44);
			4990: out = 16'(-571);
			4991: out = 16'(-471);
			4992: out = 16'(-96);
			4993: out = 16'(0);
			default: out = 0;
		endcase
	end
endmodule
