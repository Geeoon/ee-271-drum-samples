module crash1_lookup(index, out);
	input logic unsigned [15:0] index;
	output logic signed [15:0] out;
	always_comb begin
		case(index)
			0: out = 16'(0);
			1: out = 16'(0);
			2: out = 16'(5);
			3: out = 16'(-85);
			4: out = 16'(2);
			5: out = 16'(-81);
			6: out = 16'(26);
			7: out = 16'(-116);
			8: out = 16'(51);
			9: out = 16'(-155);
			10: out = 16'(108);
			11: out = 16'(-214);
			12: out = 16'(221);
			13: out = 16'(-355);
			14: out = 16'(-24);
			15: out = 16'(-394);
			16: out = 16'(7393);
			17: out = 16'(3989);
			18: out = 16'(-2028);
			19: out = 16'(3994);
			20: out = 16'(-7947);
			21: out = 16'(-7500);
			22: out = 16'(-932);
			23: out = 16'(2320);
			24: out = 16'(-17672);
			25: out = 16'(-16391);
			26: out = 16'(5131);
			27: out = 16'(19256);
			28: out = 16'(1158);
			29: out = 16'(-11713);
			30: out = 16'(-11705);
			31: out = 16'(-2208);
			32: out = 16'(-3561);
			33: out = 16'(-2903);
			34: out = 16'(-2243);
			35: out = 16'(531);
			36: out = 16'(4337);
			37: out = 16'(554);
			38: out = 16'(-5370);
			39: out = 16'(-6750);
			40: out = 16'(5764);
			41: out = 16'(-991);
			42: out = 16'(3305);
			43: out = 16'(1223);
			44: out = 16'(-6430);
			45: out = 16'(-9847);
			46: out = 16'(8458);
			47: out = 16'(14656);
			48: out = 16'(1002);
			49: out = 16'(4918);
			50: out = 16'(1138);
			51: out = 16'(-8092);
			52: out = 16'(-17884);
			53: out = 16'(326);
			54: out = 16'(10806);
			55: out = 16'(12850);
			56: out = 16'(4223);
			57: out = 16'(-2535);
			58: out = 16'(-8663);
			59: out = 16'(-5332);
			60: out = 16'(1278);
			61: out = 16'(3697);
			62: out = 16'(-967);
			63: out = 16'(-7813);
			64: out = 16'(-3472);
			65: out = 16'(9585);
			66: out = 16'(2421);
			67: out = 16'(-11468);
			68: out = 16'(-15365);
			69: out = 16'(2250);
			70: out = 16'(-4540);
			71: out = 16'(7663);
			72: out = 16'(7238);
			73: out = 16'(1222);
			74: out = 16'(-12657);
			75: out = 16'(3466);
			76: out = 16'(4586);
			77: out = 16'(-4136);
			78: out = 16'(-2000);
			79: out = 16'(11168);
			80: out = 16'(8160);
			81: out = 16'(-5380);
			82: out = 16'(-7293);
			83: out = 16'(-5069);
			84: out = 16'(2571);
			85: out = 16'(4488);
			86: out = 16'(2210);
			87: out = 16'(-5395);
			88: out = 16'(-4257);
			89: out = 16'(4895);
			90: out = 16'(12416);
			91: out = 16'(4907);
			92: out = 16'(1746);
			93: out = 16'(-54);
			94: out = 16'(-1907);
			95: out = 16'(-358);
			96: out = 16'(-2157);
			97: out = 16'(6729);
			98: out = 16'(12609);
			99: out = 16'(1815);
			100: out = 16'(-1052);
			101: out = 16'(6369);
			102: out = 16'(11850);
			103: out = 16'(-4194);
			104: out = 16'(1123);
			105: out = 16'(-4039);
			106: out = 16'(-647);
			107: out = 16'(2964);
			108: out = 16'(5095);
			109: out = 16'(-8906);
			110: out = 16'(-9033);
			111: out = 16'(2941);
			112: out = 16'(-1967);
			113: out = 16'(-7771);
			114: out = 16'(-4322);
			115: out = 16'(3973);
			116: out = 16'(-7995);
			117: out = 16'(-4264);
			118: out = 16'(582);
			119: out = 16'(898);
			120: out = 16'(-19886);
			121: out = 16'(1450);
			122: out = 16'(2156);
			123: out = 16'(-1779);
			124: out = 16'(-774);
			125: out = 16'(4418);
			126: out = 16'(-2307);
			127: out = 16'(-6184);
			128: out = 16'(1002);
			129: out = 16'(3681);
			130: out = 16'(1924);
			131: out = 16'(-1972);
			132: out = 16'(328);
			133: out = 16'(-1635);
			134: out = 16'(6873);
			135: out = 16'(4138);
			136: out = 16'(-2747);
			137: out = 16'(-8818);
			138: out = 16'(2507);
			139: out = 16'(-1404);
			140: out = 16'(-8747);
			141: out = 16'(1155);
			142: out = 16'(2874);
			143: out = 16'(8082);
			144: out = 16'(5024);
			145: out = 16'(-1340);
			146: out = 16'(-6642);
			147: out = 16'(-2874);
			148: out = 16'(-2132);
			149: out = 16'(-6922);
			150: out = 16'(-274);
			151: out = 16'(-868);
			152: out = 16'(-93);
			153: out = 16'(615);
			154: out = 16'(10371);
			155: out = 16'(-3392);
			156: out = 16'(-4889);
			157: out = 16'(514);
			158: out = 16'(3124);
			159: out = 16'(-641);
			160: out = 16'(2324);
			161: out = 16'(5029);
			162: out = 16'(4735);
			163: out = 16'(-1217);
			164: out = 16'(3380);
			165: out = 16'(-2421);
			166: out = 16'(-20005);
			167: out = 16'(-14994);
			168: out = 16'(-6473);
			169: out = 16'(-2756);
			170: out = 16'(-6239);
			171: out = 16'(-2078);
			172: out = 16'(-15);
			173: out = 16'(-2387);
			174: out = 16'(-4160);
			175: out = 16'(5979);
			176: out = 16'(10069);
			177: out = 16'(4681);
			178: out = 16'(-3455);
			179: out = 16'(309);
			180: out = 16'(-4101);
			181: out = 16'(-3233);
			182: out = 16'(1544);
			183: out = 16'(11215);
			184: out = 16'(5284);
			185: out = 16'(2252);
			186: out = 16'(-2298);
			187: out = 16'(-3089);
			188: out = 16'(-18236);
			189: out = 16'(-2871);
			190: out = 16'(4099);
			191: out = 16'(-291);
			192: out = 16'(4678);
			193: out = 16'(11890);
			194: out = 16'(17760);
			195: out = 16'(15518);
			196: out = 16'(9490);
			197: out = 16'(-742);
			198: out = 16'(-4026);
			199: out = 16'(-1851);
			200: out = 16'(1824);
			201: out = 16'(19102);
			202: out = 16'(14598);
			203: out = 16'(-2368);
			204: out = 16'(-19023);
			205: out = 16'(-4833);
			206: out = 16'(-5151);
			207: out = 16'(-8287);
			208: out = 16'(-7128);
			209: out = 16'(4354);
			210: out = 16'(-4405);
			211: out = 16'(-9249);
			212: out = 16'(-3696);
			213: out = 16'(4484);
			214: out = 16'(-375);
			215: out = 16'(-2605);
			216: out = 16'(3813);
			217: out = 16'(14260);
			218: out = 16'(1918);
			219: out = 16'(3941);
			220: out = 16'(12465);
			221: out = 16'(10904);
			222: out = 16'(9430);
			223: out = 16'(-572);
			224: out = 16'(277);
			225: out = 16'(9536);
			226: out = 16'(3752);
			227: out = 16'(-3190);
			228: out = 16'(-11942);
			229: out = 16'(-14937);
			230: out = 16'(-13663);
			231: out = 16'(-9859);
			232: out = 16'(-6189);
			233: out = 16'(-3731);
			234: out = 16'(-14845);
			235: out = 16'(762);
			236: out = 16'(952);
			237: out = 16'(-2209);
			238: out = 16'(820);
			239: out = 16'(17103);
			240: out = 16'(11610);
			241: out = 16'(1640);
			242: out = 16'(-542);
			243: out = 16'(-428);
			244: out = 16'(-1676);
			245: out = 16'(6740);
			246: out = 16'(18101);
			247: out = 16'(4595);
			248: out = 16'(-5131);
			249: out = 16'(-9772);
			250: out = 16'(-5436);
			251: out = 16'(-250);
			252: out = 16'(-18131);
			253: out = 16'(-26100);
			254: out = 16'(-10556);
			255: out = 16'(8970);
			256: out = 16'(-1421);
			257: out = 16'(-12343);
			258: out = 16'(-9417);
			259: out = 16'(1759);
			260: out = 16'(-9221);
			261: out = 16'(-12792);
			262: out = 16'(-7804);
			263: out = 16'(-969);
			264: out = 16'(-1311);
			265: out = 16'(628);
			266: out = 16'(-1375);
			267: out = 16'(-6875);
			268: out = 16'(1662);
			269: out = 16'(734);
			270: out = 16'(1879);
			271: out = 16'(1820);
			272: out = 16'(10664);
			273: out = 16'(-8969);
			274: out = 16'(-3112);
			275: out = 16'(14710);
			276: out = 16'(17930);
			277: out = 16'(16237);
			278: out = 16'(19640);
			279: out = 16'(23235);
			280: out = 16'(14586);
			281: out = 16'(2030);
			282: out = 16'(-1272);
			283: out = 16'(10908);
			284: out = 16'(19457);
			285: out = 16'(3533);
			286: out = 16'(7740);
			287: out = 16'(13771);
			288: out = 16'(7105);
			289: out = 16'(-6195);
			290: out = 16'(-19068);
			291: out = 16'(-12803);
			292: out = 16'(-5882);
			293: out = 16'(-21986);
			294: out = 16'(-22013);
			295: out = 16'(-15125);
			296: out = 16'(-6544);
			297: out = 16'(-6590);
			298: out = 16'(-3981);
			299: out = 16'(-5886);
			300: out = 16'(-10904);
			301: out = 16'(-17920);
			302: out = 16'(-15649);
			303: out = 16'(-9992);
			304: out = 16'(-5890);
			305: out = 16'(-6987);
			306: out = 16'(-6044);
			307: out = 16'(1482);
			308: out = 16'(7079);
			309: out = 16'(3452);
			310: out = 16'(2673);
			311: out = 16'(-8832);
			312: out = 16'(-3427);
			313: out = 16'(8424);
			314: out = 16'(11434);
			315: out = 16'(10763);
			316: out = 16'(7874);
			317: out = 16'(7220);
			318: out = 16'(12724);
			319: out = 16'(16714);
			320: out = 16'(26215);
			321: out = 16'(23518);
			322: out = 16'(14274);
			323: out = 16'(20683);
			324: out = 16'(23310);
			325: out = 16'(13030);
			326: out = 16'(-2278);
			327: out = 16'(13843);
			328: out = 16'(13998);
			329: out = 16'(14505);
			330: out = 16'(8707);
			331: out = 16'(11415);
			332: out = 16'(-8432);
			333: out = 16'(-6588);
			334: out = 16'(-4054);
			335: out = 16'(-15117);
			336: out = 16'(-12070);
			337: out = 16'(-4805);
			338: out = 16'(-6856);
			339: out = 16'(-20500);
			340: out = 16'(-11037);
			341: out = 16'(-2887);
			342: out = 16'(260);
			343: out = 16'(-7544);
			344: out = 16'(-26753);
			345: out = 16'(-28955);
			346: out = 16'(-22755);
			347: out = 16'(-15592);
			348: out = 16'(-32767);
			349: out = 16'(-8010);
			350: out = 16'(-2501);
			351: out = 16'(-13308);
			352: out = 16'(-18141);
			353: out = 16'(8020);
			354: out = 16'(-1928);
			355: out = 16'(-23078);
			356: out = 16'(-21127);
			357: out = 16'(-11644);
			358: out = 16'(-16310);
			359: out = 16'(-16828);
			360: out = 16'(3286);
			361: out = 16'(-3376);
			362: out = 16'(514);
			363: out = 16'(235);
			364: out = 16'(-3470);
			365: out = 16'(-1499);
			366: out = 16'(-17009);
			367: out = 16'(-14315);
			368: out = 16'(799);
			369: out = 16'(4225);
			370: out = 16'(3141);
			371: out = 16'(17180);
			372: out = 16'(25093);
			373: out = 16'(6615);
			374: out = 16'(-5663);
			375: out = 16'(409);
			376: out = 16'(11789);
			377: out = 16'(2846);
			378: out = 16'(14168);
			379: out = 16'(10910);
			380: out = 16'(13533);
			381: out = 16'(16469);
			382: out = 16'(25656);
			383: out = 16'(17277);
			384: out = 16'(14706);
			385: out = 16'(14979);
			386: out = 16'(9237);
			387: out = 16'(6237);
			388: out = 16'(10960);
			389: out = 16'(20177);
			390: out = 16'(17709);
			391: out = 16'(25465);
			392: out = 16'(14511);
			393: out = 16'(6433);
			394: out = 16'(9271);
			395: out = 16'(15517);
			396: out = 16'(8254);
			397: out = 16'(3139);
			398: out = 16'(9354);
			399: out = 16'(11421);
			400: out = 16'(12531);
			401: out = 16'(12582);
			402: out = 16'(16394);
			403: out = 16'(22741);
			404: out = 16'(11216);
			405: out = 16'(3260);
			406: out = 16'(8041);
			407: out = 16'(18299);
			408: out = 16'(15009);
			409: out = 16'(5838);
			410: out = 16'(-881);
			411: out = 16'(815);
			412: out = 16'(3977);
			413: out = 16'(2382);
			414: out = 16'(-5823);
			415: out = 16'(-10762);
			416: out = 16'(-14221);
			417: out = 16'(-5859);
			418: out = 16'(-8003);
			419: out = 16'(-19665);
			420: out = 16'(-22545);
			421: out = 16'(-9754);
			422: out = 16'(-8712);
			423: out = 16'(-24411);
			424: out = 16'(-19618);
			425: out = 16'(-24123);
			426: out = 16'(-18816);
			427: out = 16'(-17198);
			428: out = 16'(-21414);
			429: out = 16'(-25655);
			430: out = 16'(-27430);
			431: out = 16'(-29691);
			432: out = 16'(-27693);
			433: out = 16'(-28502);
			434: out = 16'(-19172);
			435: out = 16'(-19292);
			436: out = 16'(-24426);
			437: out = 16'(-29479);
			438: out = 16'(-12307);
			439: out = 16'(-5071);
			440: out = 16'(-11647);
			441: out = 16'(-23035);
			442: out = 16'(-7143);
			443: out = 16'(-7725);
			444: out = 16'(-20014);
			445: out = 16'(-6644);
			446: out = 16'(3109);
			447: out = 16'(538);
			448: out = 16'(-9526);
			449: out = 16'(-14828);
			450: out = 16'(-3716);
			451: out = 16'(-11462);
			452: out = 16'(-14599);
			453: out = 16'(5346);
			454: out = 16'(5942);
			455: out = 16'(-3268);
			456: out = 16'(3090);
			457: out = 16'(31340);
			458: out = 16'(22972);
			459: out = 16'(17738);
			460: out = 16'(6749);
			461: out = 16'(4258);
			462: out = 16'(-3808);
			463: out = 16'(14197);
			464: out = 16'(24628);
			465: out = 16'(27016);
			466: out = 16'(22365);
			467: out = 16'(27890);
			468: out = 16'(24224);
			469: out = 16'(15948);
			470: out = 16'(7482);
			471: out = 16'(17782);
			472: out = 16'(17326);
			473: out = 16'(9033);
			474: out = 16'(-2224);
			475: out = 16'(1200);
			476: out = 16'(-221);
			477: out = 16'(6545);
			478: out = 16'(15437);
			479: out = 16'(7366);
			480: out = 16'(-2707);
			481: out = 16'(-11192);
			482: out = 16'(-9207);
			483: out = 16'(-20);
			484: out = 16'(3994);
			485: out = 16'(4550);
			486: out = 16'(10691);
			487: out = 16'(26013);
			488: out = 16'(14931);
			489: out = 16'(10897);
			490: out = 16'(9408);
			491: out = 16'(8879);
			492: out = 16'(-5093);
			493: out = 16'(-5286);
			494: out = 16'(-2080);
			495: out = 16'(928);
			496: out = 16'(12536);
			497: out = 16'(17154);
			498: out = 16'(10193);
			499: out = 16'(-1322);
			500: out = 16'(137);
			501: out = 16'(-2673);
			502: out = 16'(-5901);
			503: out = 16'(-5742);
			504: out = 16'(2192);
			505: out = 16'(4194);
			506: out = 16'(1817);
			507: out = 16'(3345);
			508: out = 16'(13298);
			509: out = 16'(5462);
			510: out = 16'(-2956);
			511: out = 16'(-10526);
			512: out = 16'(-15771);
			513: out = 16'(-13256);
			514: out = 16'(-11866);
			515: out = 16'(-758);
			516: out = 16'(12724);
			517: out = 16'(4979);
			518: out = 16'(-1369);
			519: out = 16'(-423);
			520: out = 16'(1337);
			521: out = 16'(-24577);
			522: out = 16'(-18935);
			523: out = 16'(-7937);
			524: out = 16'(-1993);
			525: out = 16'(-2150);
			526: out = 16'(-7050);
			527: out = 16'(-5089);
			528: out = 16'(-1422);
			529: out = 16'(-1993);
			530: out = 16'(-5338);
			531: out = 16'(-2835);
			532: out = 16'(-6330);
			533: out = 16'(-20060);
			534: out = 16'(-13681);
			535: out = 16'(-5083);
			536: out = 16'(-1587);
			537: out = 16'(-6119);
			538: out = 16'(6928);
			539: out = 16'(3311);
			540: out = 16'(-4005);
			541: out = 16'(-12504);
			542: out = 16'(2587);
			543: out = 16'(-18162);
			544: out = 16'(-13910);
			545: out = 16'(6592);
			546: out = 16'(8798);
			547: out = 16'(-146);
			548: out = 16'(-6615);
			549: out = 16'(-981);
			550: out = 16'(2572);
			551: out = 16'(7963);
			552: out = 16'(4931);
			553: out = 16'(8200);
			554: out = 16'(12472);
			555: out = 16'(23875);
			556: out = 16'(10872);
			557: out = 16'(6812);
			558: out = 16'(7870);
			559: out = 16'(957);
			560: out = 16'(-15854);
			561: out = 16'(-10163);
			562: out = 16'(9148);
			563: out = 16'(4470);
			564: out = 16'(2671);
			565: out = 16'(-469);
			566: out = 16'(-614);
			567: out = 16'(-5735);
			568: out = 16'(-148);
			569: out = 16'(6535);
			570: out = 16'(13103);
			571: out = 16'(12530);
			572: out = 16'(5009);
			573: out = 16'(4055);
			574: out = 16'(4778);
			575: out = 16'(-52);
			576: out = 16'(-5199);
			577: out = 16'(-4659);
			578: out = 16'(336);
			579: out = 16'(1127);
			580: out = 16'(673);
			581: out = 16'(5901);
			582: out = 16'(10901);
			583: out = 16'(7918);
			584: out = 16'(5693);
			585: out = 16'(-986);
			586: out = 16'(3403);
			587: out = 16'(772);
			588: out = 16'(-7553);
			589: out = 16'(104);
			590: out = 16'(16586);
			591: out = 16'(16577);
			592: out = 16'(2574);
			593: out = 16'(-3206);
			594: out = 16'(5651);
			595: out = 16'(3283);
			596: out = 16'(-11750);
			597: out = 16'(-12375);
			598: out = 16'(6305);
			599: out = 16'(14875);
			600: out = 16'(5113);
			601: out = 16'(104);
			602: out = 16'(1612);
			603: out = 16'(9009);
			604: out = 16'(12496);
			605: out = 16'(12037);
			606: out = 16'(-969);
			607: out = 16'(-14619);
			608: out = 16'(-16871);
			609: out = 16'(-2734);
			610: out = 16'(-9620);
			611: out = 16'(-5669);
			612: out = 16'(271);
			613: out = 16'(5431);
			614: out = 16'(-8958);
			615: out = 16'(-2919);
			616: out = 16'(-3622);
			617: out = 16'(-8979);
			618: out = 16'(-2535);
			619: out = 16'(-1574);
			620: out = 16'(77);
			621: out = 16'(-4232);
			622: out = 16'(-14085);
			623: out = 16'(-10278);
			624: out = 16'(-2983);
			625: out = 16'(-2370);
			626: out = 16'(-13719);
			627: out = 16'(-22194);
			628: out = 16'(-26303);
			629: out = 16'(-19455);
			630: out = 16'(-10341);
			631: out = 16'(-6203);
			632: out = 16'(-9408);
			633: out = 16'(-5898);
			634: out = 16'(5856);
			635: out = 16'(19382);
			636: out = 16'(6907);
			637: out = 16'(2838);
			638: out = 16'(11388);
			639: out = 16'(10105);
			640: out = 16'(12018);
			641: out = 16'(891);
			642: out = 16'(-3124);
			643: out = 16'(7803);
			644: out = 16'(22072);
			645: out = 16'(17561);
			646: out = 16'(5306);
			647: out = 16'(1028);
			648: out = 16'(4045);
			649: out = 16'(12051);
			650: out = 16'(16064);
			651: out = 16'(17144);
			652: out = 16'(13512);
			653: out = 16'(11401);
			654: out = 16'(576);
			655: out = 16'(-7143);
			656: out = 16'(13765);
			657: out = 16'(-4035);
			658: out = 16'(-13937);
			659: out = 16'(-13038);
			660: out = 16'(-3408);
			661: out = 16'(-12808);
			662: out = 16'(-9885);
			663: out = 16'(4779);
			664: out = 16'(18258);
			665: out = 16'(1227);
			666: out = 16'(-1105);
			667: out = 16'(-4154);
			668: out = 16'(-13912);
			669: out = 16'(-12167);
			670: out = 16'(-10455);
			671: out = 16'(-5412);
			672: out = 16'(-2011);
			673: out = 16'(74);
			674: out = 16'(-5726);
			675: out = 16'(-8622);
			676: out = 16'(-7978);
			677: out = 16'(-12957);
			678: out = 16'(-26099);
			679: out = 16'(-27658);
			680: out = 16'(-13154);
			681: out = 16'(-2912);
			682: out = 16'(10642);
			683: out = 16'(769);
			684: out = 16'(-5501);
			685: out = 16'(-144);
			686: out = 16'(431);
			687: out = 16'(-10645);
			688: out = 16'(-11745);
			689: out = 16'(1133);
			690: out = 16'(-5715);
			691: out = 16'(-6702);
			692: out = 16'(-5953);
			693: out = 16'(-2966);
			694: out = 16'(-3071);
			695: out = 16'(-5070);
			696: out = 16'(422);
			697: out = 16'(8465);
			698: out = 16'(11086);
			699: out = 16'(3930);
			700: out = 16'(7514);
			701: out = 16'(14470);
			702: out = 16'(14222);
			703: out = 16'(3487);
			704: out = 16'(6878);
			705: out = 16'(16680);
			706: out = 16'(22595);
			707: out = 16'(10993);
			708: out = 16'(21627);
			709: out = 16'(22129);
			710: out = 16'(13772);
			711: out = 16'(18428);
			712: out = 16'(14613);
			713: out = 16'(2031);
			714: out = 16'(-6684);
			715: out = 16'(14338);
			716: out = 16'(13065);
			717: out = 16'(8918);
			718: out = 16'(1225);
			719: out = 16'(897);
			720: out = 16'(6047);
			721: out = 16'(12554);
			722: out = 16'(5339);
			723: out = 16'(-14340);
			724: out = 16'(2245);
			725: out = 16'(5823);
			726: out = 16'(12334);
			727: out = 16'(16443);
			728: out = 16'(19977);
			729: out = 16'(-7012);
			730: out = 16'(-21073);
			731: out = 16'(-14297);
			732: out = 16'(-11133);
			733: out = 16'(-12755);
			734: out = 16'(-10074);
			735: out = 16'(-2663);
			736: out = 16'(-4249);
			737: out = 16'(-1836);
			738: out = 16'(3976);
			739: out = 16'(7654);
			740: out = 16'(-3572);
			741: out = 16'(-7015);
			742: out = 16'(-22052);
			743: out = 16'(-29858);
			744: out = 16'(-25717);
			745: out = 16'(2491);
			746: out = 16'(16417);
			747: out = 16'(11132);
			748: out = 16'(-2156);
			749: out = 16'(-66);
			750: out = 16'(-17594);
			751: out = 16'(-29400);
			752: out = 16'(-27933);
			753: out = 16'(-24731);
			754: out = 16'(-9789);
			755: out = 16'(-5947);
			756: out = 16'(-2498);
			757: out = 16'(10775);
			758: out = 16'(6232);
			759: out = 16'(-3637);
			760: out = 16'(-16482);
			761: out = 16'(-18483);
			762: out = 16'(-8938);
			763: out = 16'(5323);
			764: out = 16'(9109);
			765: out = 16'(7800);
			766: out = 16'(8286);
			767: out = 16'(10958);
			768: out = 16'(3692);
			769: out = 16'(-8259);
			770: out = 16'(-11606);
			771: out = 16'(-3864);
			772: out = 16'(1722);
			773: out = 16'(2051);
			774: out = 16'(3784);
			775: out = 16'(12812);
			776: out = 16'(14163);
			777: out = 16'(9176);
			778: out = 16'(4813);
			779: out = 16'(6006);
			780: out = 16'(6236);
			781: out = 16'(5179);
			782: out = 16'(980);
			783: out = 16'(-392);
			784: out = 16'(-8821);
			785: out = 16'(-7141);
			786: out = 16'(1570);
			787: out = 16'(-1068);
			788: out = 16'(-1973);
			789: out = 16'(6292);
			790: out = 16'(16890);
			791: out = 16'(12803);
			792: out = 16'(3884);
			793: out = 16'(-1059);
			794: out = 16'(1063);
			795: out = 16'(148);
			796: out = 16'(7636);
			797: out = 16'(14643);
			798: out = 16'(19876);
			799: out = 16'(15226);
			800: out = 16'(9802);
			801: out = 16'(1069);
			802: out = 16'(-860);
			803: out = 16'(-1282);
			804: out = 16'(4994);
			805: out = 16'(-11769);
			806: out = 16'(-15294);
			807: out = 16'(2737);
			808: out = 16'(16544);
			809: out = 16'(5519);
			810: out = 16'(-9958);
			811: out = 16'(-11699);
			812: out = 16'(-1286);
			813: out = 16'(-1461);
			814: out = 16'(-5725);
			815: out = 16'(-3324);
			816: out = 16'(4287);
			817: out = 16'(-3943);
			818: out = 16'(-17528);
			819: out = 16'(-23121);
			820: out = 16'(-9631);
			821: out = 16'(-9305);
			822: out = 16'(2598);
			823: out = 16'(5156);
			824: out = 16'(1387);
			825: out = 16'(-7155);
			826: out = 16'(-1083);
			827: out = 16'(-2212);
			828: out = 16'(-6432);
			829: out = 16'(969);
			830: out = 16'(3986);
			831: out = 16'(2234);
			832: out = 16'(3138);
			833: out = 16'(13785);
			834: out = 16'(4107);
			835: out = 16'(-3228);
			836: out = 16'(-3794);
			837: out = 16'(1462);
			838: out = 16'(-6045);
			839: out = 16'(-5347);
			840: out = 16'(5442);
			841: out = 16'(15581);
			842: out = 16'(15324);
			843: out = 16'(3092);
			844: out = 16'(-4987);
			845: out = 16'(-4565);
			846: out = 16'(5643);
			847: out = 16'(-1062);
			848: out = 16'(2964);
			849: out = 16'(8116);
			850: out = 16'(3784);
			851: out = 16'(319);
			852: out = 16'(13205);
			853: out = 16'(17062);
			854: out = 16'(-3641);
			855: out = 16'(7902);
			856: out = 16'(21212);
			857: out = 16'(25963);
			858: out = 16'(13275);
			859: out = 16'(14227);
			860: out = 16'(1927);
			861: out = 16'(-3114);
			862: out = 16'(-3914);
			863: out = 16'(-19363);
			864: out = 16'(-8510);
			865: out = 16'(5852);
			866: out = 16'(12568);
			867: out = 16'(2257);
			868: out = 16'(14594);
			869: out = 16'(1700);
			870: out = 16'(-19429);
			871: out = 16'(-21788);
			872: out = 16'(8113);
			873: out = 16'(22099);
			874: out = 16'(16453);
			875: out = 16'(6196);
			876: out = 16'(-2632);
			877: out = 16'(-19042);
			878: out = 16'(-23954);
			879: out = 16'(-8595);
			880: out = 16'(-20192);
			881: out = 16'(-16123);
			882: out = 16'(-12439);
			883: out = 16'(-5359);
			884: out = 16'(-9895);
			885: out = 16'(-403);
			886: out = 16'(-12864);
			887: out = 16'(-30324);
			888: out = 16'(-27961);
			889: out = 16'(-29449);
			890: out = 16'(-25274);
			891: out = 16'(-17584);
			892: out = 16'(-8170);
			893: out = 16'(9672);
			894: out = 16'(9210);
			895: out = 16'(-9562);
			896: out = 16'(-29960);
			897: out = 16'(-22583);
			898: out = 16'(-25809);
			899: out = 16'(-28426);
			900: out = 16'(-21383);
			901: out = 16'(2903);
			902: out = 16'(800);
			903: out = 16'(4455);
			904: out = 16'(14054);
			905: out = 16'(2980);
			906: out = 16'(-2895);
			907: out = 16'(-15434);
			908: out = 16'(-17361);
			909: out = 16'(-6627);
			910: out = 16'(10857);
			911: out = 16'(14713);
			912: out = 16'(19201);
			913: out = 16'(30143);
			914: out = 16'(30228);
			915: out = 16'(17717);
			916: out = 16'(-2415);
			917: out = 16'(-8153);
			918: out = 16'(639);
			919: out = 16'(22078);
			920: out = 16'(28022);
			921: out = 16'(23563);
			922: out = 16'(16163);
			923: out = 16'(26584);
			924: out = 16'(22157);
			925: out = 16'(12450);
			926: out = 16'(18424);
			927: out = 16'(13168);
			928: out = 16'(11160);
			929: out = 16'(9639);
			930: out = 16'(13533);
			931: out = 16'(21956);
			932: out = 16'(25390);
			933: out = 16'(19948);
			934: out = 16'(9643);
			935: out = 16'(11104);
			936: out = 16'(566);
			937: out = 16'(-8290);
			938: out = 16'(-9229);
			939: out = 16'(508);
			940: out = 16'(-2854);
			941: out = 16'(-2277);
			942: out = 16'(4522);
			943: out = 16'(5155);
			944: out = 16'(-1266);
			945: out = 16'(-8826);
			946: out = 16'(-8534);
			947: out = 16'(-3308);
			948: out = 16'(-12704);
			949: out = 16'(-14352);
			950: out = 16'(-6240);
			951: out = 16'(-5182);
			952: out = 16'(-1768);
			953: out = 16'(-15184);
			954: out = 16'(-18367);
			955: out = 16'(-8113);
			956: out = 16'(-8200);
			957: out = 16'(-11489);
			958: out = 16'(-8009);
			959: out = 16'(1534);
			960: out = 16'(9948);
			961: out = 16'(-1571);
			962: out = 16'(-5576);
			963: out = 16'(-1663);
			964: out = 16'(-2295);
			965: out = 16'(-11416);
			966: out = 16'(-5983);
			967: out = 16'(6476);
			968: out = 16'(4576);
			969: out = 16'(6059);
			970: out = 16'(4350);
			971: out = 16'(1168);
			972: out = 16'(-7556);
			973: out = 16'(-23441);
			974: out = 16'(-20515);
			975: out = 16'(-6279);
			976: out = 16'(369);
			977: out = 16'(-4017);
			978: out = 16'(-8843);
			979: out = 16'(-13166);
			980: out = 16'(-15972);
			981: out = 16'(-10127);
			982: out = 16'(-3004);
			983: out = 16'(1990);
			984: out = 16'(-162);
			985: out = 16'(-9274);
			986: out = 16'(-962);
			987: out = 16'(3645);
			988: out = 16'(2925);
			989: out = 16'(1487);
			990: out = 16'(-2827);
			991: out = 16'(-8452);
			992: out = 16'(-10333);
			993: out = 16'(-751);
			994: out = 16'(12898);
			995: out = 16'(22695);
			996: out = 16'(19447);
			997: out = 16'(10608);
			998: out = 16'(11634);
			999: out = 16'(5200);
			1000: out = 16'(978);
			1001: out = 16'(1934);
			1002: out = 16'(5355);
			1003: out = 16'(1055);
			1004: out = 16'(-5885);
			1005: out = 16'(-1696);
			1006: out = 16'(19210);
			1007: out = 16'(22460);
			1008: out = 16'(18576);
			1009: out = 16'(6765);
			1010: out = 16'(-4442);
			1011: out = 16'(-3530);
			1012: out = 16'(-2129);
			1013: out = 16'(-3539);
			1014: out = 16'(789);
			1015: out = 16'(20578);
			1016: out = 16'(25613);
			1017: out = 16'(16780);
			1018: out = 16'(6233);
			1019: out = 16'(8555);
			1020: out = 16'(2284);
			1021: out = 16'(-4726);
			1022: out = 16'(-7243);
			1023: out = 16'(-3608);
			1024: out = 16'(9917);
			1025: out = 16'(16198);
			1026: out = 16'(16007);
			1027: out = 16'(9245);
			1028: out = 16'(816);
			1029: out = 16'(-11256);
			1030: out = 16'(-8333);
			1031: out = 16'(7315);
			1032: out = 16'(6528);
			1033: out = 16'(2349);
			1034: out = 16'(4827);
			1035: out = 16'(8626);
			1036: out = 16'(-9055);
			1037: out = 16'(-23152);
			1038: out = 16'(-18438);
			1039: out = 16'(1561);
			1040: out = 16'(-1910);
			1041: out = 16'(7795);
			1042: out = 16'(8114);
			1043: out = 16'(6719);
			1044: out = 16'(-2983);
			1045: out = 16'(7877);
			1046: out = 16'(-6411);
			1047: out = 16'(-25881);
			1048: out = 16'(-27792);
			1049: out = 16'(-22278);
			1050: out = 16'(-10197);
			1051: out = 16'(-7937);
			1052: out = 16'(-12221);
			1053: out = 16'(-8409);
			1054: out = 16'(-6097);
			1055: out = 16'(-9723);
			1056: out = 16'(-20419);
			1057: out = 16'(-27533);
			1058: out = 16'(-20537);
			1059: out = 16'(-5231);
			1060: out = 16'(2770);
			1061: out = 16'(5170);
			1062: out = 16'(-16645);
			1063: out = 16'(-25623);
			1064: out = 16'(-23466);
			1065: out = 16'(-18794);
			1066: out = 16'(-7689);
			1067: out = 16'(4657);
			1068: out = 16'(7132);
			1069: out = 16'(1248);
			1070: out = 16'(7743);
			1071: out = 16'(6280);
			1072: out = 16'(-6367);
			1073: out = 16'(-19895);
			1074: out = 16'(2565);
			1075: out = 16'(15067);
			1076: out = 16'(23171);
			1077: out = 16'(23932);
			1078: out = 16'(22900);
			1079: out = 16'(25707);
			1080: out = 16'(23630);
			1081: out = 16'(12634);
			1082: out = 16'(-1110);
			1083: out = 16'(4059);
			1084: out = 16'(8211);
			1085: out = 16'(9845);
			1086: out = 16'(13707);
			1087: out = 16'(8094);
			1088: out = 16'(10043);
			1089: out = 16'(6043);
			1090: out = 16'(-3120);
			1091: out = 16'(-23190);
			1092: out = 16'(-5970);
			1093: out = 16'(11000);
			1094: out = 16'(5340);
			1095: out = 16'(-10199);
			1096: out = 16'(-18143);
			1097: out = 16'(-13121);
			1098: out = 16'(-6888);
			1099: out = 16'(-7232);
			1100: out = 16'(-5625);
			1101: out = 16'(-1977);
			1102: out = 16'(4098);
			1103: out = 16'(12035);
			1104: out = 16'(17191);
			1105: out = 16'(17855);
			1106: out = 16'(13326);
			1107: out = 16'(7710);
			1108: out = 16'(5233);
			1109: out = 16'(-3469);
			1110: out = 16'(-9436);
			1111: out = 16'(-6240);
			1112: out = 16'(-20997);
			1113: out = 16'(-4538);
			1114: out = 16'(-2463);
			1115: out = 16'(-5804);
			1116: out = 16'(5609);
			1117: out = 16'(15234);
			1118: out = 16'(6155);
			1119: out = 16'(-9635);
			1120: out = 16'(-10415);
			1121: out = 16'(-2701);
			1122: out = 16'(1197);
			1123: out = 16'(1321);
			1124: out = 16'(6630);
			1125: out = 16'(9705);
			1126: out = 16'(10381);
			1127: out = 16'(11147);
			1128: out = 16'(11709);
			1129: out = 16'(3960);
			1130: out = 16'(-4411);
			1131: out = 16'(-1345);
			1132: out = 16'(8179);
			1133: out = 16'(-3537);
			1134: out = 16'(2008);
			1135: out = 16'(1419);
			1136: out = 16'(-1174);
			1137: out = 16'(-670);
			1138: out = 16'(-7179);
			1139: out = 16'(-8129);
			1140: out = 16'(-4527);
			1141: out = 16'(1946);
			1142: out = 16'(8116);
			1143: out = 16'(7634);
			1144: out = 16'(-5854);
			1145: out = 16'(-23358);
			1146: out = 16'(-29272);
			1147: out = 16'(-17902);
			1148: out = 16'(-10680);
			1149: out = 16'(-12804);
			1150: out = 16'(-10694);
			1151: out = 16'(13882);
			1152: out = 16'(24704);
			1153: out = 16'(11546);
			1154: out = 16'(-9432);
			1155: out = 16'(-10895);
			1156: out = 16'(-9359);
			1157: out = 16'(-16929);
			1158: out = 16'(-26426);
			1159: out = 16'(-19842);
			1160: out = 16'(-5960);
			1161: out = 16'(-436);
			1162: out = 16'(-4774);
			1163: out = 16'(11119);
			1164: out = 16'(6126);
			1165: out = 16'(-4834);
			1166: out = 16'(-6954);
			1167: out = 16'(10770);
			1168: out = 16'(13411);
			1169: out = 16'(11396);
			1170: out = 16'(13374);
			1171: out = 16'(16692);
			1172: out = 16'(9150);
			1173: out = 16'(-3871);
			1174: out = 16'(-9204);
			1175: out = 16'(1154);
			1176: out = 16'(-362);
			1177: out = 16'(-391);
			1178: out = 16'(3131);
			1179: out = 16'(6356);
			1180: out = 16'(12437);
			1181: out = 16'(6997);
			1182: out = 16'(-2925);
			1183: out = 16'(-13391);
			1184: out = 16'(-5198);
			1185: out = 16'(-9435);
			1186: out = 16'(-6012);
			1187: out = 16'(9736);
			1188: out = 16'(29368);
			1189: out = 16'(21453);
			1190: out = 16'(16545);
			1191: out = 16'(14871);
			1192: out = 16'(11433);
			1193: out = 16'(-11888);
			1194: out = 16'(-12571);
			1195: out = 16'(5788);
			1196: out = 16'(13264);
			1197: out = 16'(10858);
			1198: out = 16'(12834);
			1199: out = 16'(16831);
			1200: out = 16'(9859);
			1201: out = 16'(4050);
			1202: out = 16'(-2301);
			1203: out = 16'(-7109);
			1204: out = 16'(-16045);
			1205: out = 16'(-8622);
			1206: out = 16'(-7517);
			1207: out = 16'(-1411);
			1208: out = 16'(-1901);
			1209: out = 16'(-11175);
			1210: out = 16'(-21229);
			1211: out = 16'(-20423);
			1212: out = 16'(-19354);
			1213: out = 16'(-22675);
			1214: out = 16'(-15988);
			1215: out = 16'(8253);
			1216: out = 16'(24059);
			1217: out = 16'(21704);
			1218: out = 16'(11564);
			1219: out = 16'(8780);
			1220: out = 16'(-7037);
			1221: out = 16'(-29514);
			1222: out = 16'(-28519);
			1223: out = 16'(-11774);
			1224: out = 16'(2463);
			1225: out = 16'(2181);
			1226: out = 16'(14452);
			1227: out = 16'(19981);
			1228: out = 16'(13727);
			1229: out = 16'(-3483);
			1230: out = 16'(-5777);
			1231: out = 16'(-17699);
			1232: out = 16'(-16273);
			1233: out = 16'(-6305);
			1234: out = 16'(6947);
			1235: out = 16'(10885);
			1236: out = 16'(8613);
			1237: out = 16'(8805);
			1238: out = 16'(18541);
			1239: out = 16'(-564);
			1240: out = 16'(-195);
			1241: out = 16'(-2586);
			1242: out = 16'(-11737);
			1243: out = 16'(-27165);
			1244: out = 16'(-7581);
			1245: out = 16'(18719);
			1246: out = 16'(20791);
			1247: out = 16'(2227);
			1248: out = 16'(-2303);
			1249: out = 16'(873);
			1250: out = 16'(105);
			1251: out = 16'(-4349);
			1252: out = 16'(-853);
			1253: out = 16'(12283);
			1254: out = 16'(15501);
			1255: out = 16'(2787);
			1256: out = 16'(816);
			1257: out = 16'(906);
			1258: out = 16'(1489);
			1259: out = 16'(-105);
			1260: out = 16'(-469);
			1261: out = 16'(2337);
			1262: out = 16'(3164);
			1263: out = 16'(632);
			1264: out = 16'(-7604);
			1265: out = 16'(269);
			1266: out = 16'(3675);
			1267: out = 16'(1045);
			1268: out = 16'(1666);
			1269: out = 16'(-740);
			1270: out = 16'(-11100);
			1271: out = 16'(-19830);
			1272: out = 16'(-7854);
			1273: out = 16'(2563);
			1274: out = 16'(5864);
			1275: out = 16'(-1867);
			1276: out = 16'(-3010);
			1277: out = 16'(5977);
			1278: out = 16'(19972);
			1279: out = 16'(14345);
			1280: out = 16'(-5735);
			1281: out = 16'(-19890);
			1282: out = 16'(-5711);
			1283: out = 16'(17313);
			1284: out = 16'(19474);
			1285: out = 16'(-4561);
			1286: out = 16'(-3311);
			1287: out = 16'(9434);
			1288: out = 16'(14989);
			1289: out = 16'(-3685);
			1290: out = 16'(4314);
			1291: out = 16'(-1596);
			1292: out = 16'(-14437);
			1293: out = 16'(-28399);
			1294: out = 16'(-3247);
			1295: out = 16'(2544);
			1296: out = 16'(-1812);
			1297: out = 16'(-5988);
			1298: out = 16'(-2974);
			1299: out = 16'(-14326);
			1300: out = 16'(-15772);
			1301: out = 16'(-2625);
			1302: out = 16'(445);
			1303: out = 16'(-2651);
			1304: out = 16'(-2851);
			1305: out = 16'(1939);
			1306: out = 16'(-1277);
			1307: out = 16'(-1101);
			1308: out = 16'(5182);
			1309: out = 16'(10808);
			1310: out = 16'(87);
			1311: out = 16'(9137);
			1312: out = 16'(7556);
			1313: out = 16'(3215);
			1314: out = 16'(-5783);
			1315: out = 16'(4288);
			1316: out = 16'(-8330);
			1317: out = 16'(-22715);
			1318: out = 16'(-25883);
			1319: out = 16'(-6391);
			1320: out = 16'(3907);
			1321: out = 16'(10221);
			1322: out = 16'(10611);
			1323: out = 16'(7326);
			1324: out = 16'(-8149);
			1325: out = 16'(-8625);
			1326: out = 16'(2016);
			1327: out = 16'(4168);
			1328: out = 16'(-2058);
			1329: out = 16'(-6271);
			1330: out = 16'(-6604);
			1331: out = 16'(-8308);
			1332: out = 16'(-8266);
			1333: out = 16'(-2103);
			1334: out = 16'(3020);
			1335: out = 16'(3050);
			1336: out = 16'(17227);
			1337: out = 16'(8160);
			1338: out = 16'(-6457);
			1339: out = 16'(-11719);
			1340: out = 16'(3799);
			1341: out = 16'(2837);
			1342: out = 16'(-6517);
			1343: out = 16'(-4494);
			1344: out = 16'(18826);
			1345: out = 16'(16846);
			1346: out = 16'(5853);
			1347: out = 16'(-53);
			1348: out = 16'(6393);
			1349: out = 16'(3771);
			1350: out = 16'(-2283);
			1351: out = 16'(6760);
			1352: out = 16'(31091);
			1353: out = 16'(26752);
			1354: out = 16'(26052);
			1355: out = 16'(17223);
			1356: out = 16'(3455);
			1357: out = 16'(-19888);
			1358: out = 16'(-14743);
			1359: out = 16'(9385);
			1360: out = 16'(26760);
			1361: out = 16'(21648);
			1362: out = 16'(19638);
			1363: out = 16'(14755);
			1364: out = 16'(7279);
			1365: out = 16'(-2559);
			1366: out = 16'(-20136);
			1367: out = 16'(-15339);
			1368: out = 16'(6783);
			1369: out = 16'(16817);
			1370: out = 16'(10379);
			1371: out = 16'(6847);
			1372: out = 16'(13749);
			1373: out = 16'(14448);
			1374: out = 16'(-1719);
			1375: out = 16'(-15929);
			1376: out = 16'(-11542);
			1377: out = 16'(-1163);
			1378: out = 16'(-11021);
			1379: out = 16'(-19892);
			1380: out = 16'(-13204);
			1381: out = 16'(1906);
			1382: out = 16'(-2859);
			1383: out = 16'(732);
			1384: out = 16'(-1612);
			1385: out = 16'(-4987);
			1386: out = 16'(-9528);
			1387: out = 16'(-20304);
			1388: out = 16'(-19702);
			1389: out = 16'(-8751);
			1390: out = 16'(-1057);
			1391: out = 16'(-11494);
			1392: out = 16'(-15479);
			1393: out = 16'(-14952);
			1394: out = 16'(-14728);
			1395: out = 16'(-10716);
			1396: out = 16'(-8223);
			1397: out = 16'(-2639);
			1398: out = 16'(-916);
			1399: out = 16'(-21329);
			1400: out = 16'(-5439);
			1401: out = 16'(9836);
			1402: out = 16'(9335);
			1403: out = 16'(-11731);
			1404: out = 16'(-2046);
			1405: out = 16'(-6977);
			1406: out = 16'(-20004);
			1407: out = 16'(-26172);
			1408: out = 16'(-12692);
			1409: out = 16'(-2737);
			1410: out = 16'(-1682);
			1411: out = 16'(-4281);
			1412: out = 16'(917);
			1413: out = 16'(7443);
			1414: out = 16'(15133);
			1415: out = 16'(12340);
			1416: out = 16'(-444);
			1417: out = 16'(-7640);
			1418: out = 16'(11087);
			1419: out = 16'(26438);
			1420: out = 16'(5225);
			1421: out = 16'(2102);
			1422: out = 16'(7817);
			1423: out = 16'(9876);
			1424: out = 16'(-8713);
			1425: out = 16'(-8285);
			1426: out = 16'(-3675);
			1427: out = 16'(-2645);
			1428: out = 16'(-11264);
			1429: out = 16'(-2116);
			1430: out = 16'(16440);
			1431: out = 16'(25368);
			1432: out = 16'(13522);
			1433: out = 16'(5079);
			1434: out = 16'(-2794);
			1435: out = 16'(-1007);
			1436: out = 16'(2353);
			1437: out = 16'(12741);
			1438: out = 16'(10677);
			1439: out = 16'(10401);
			1440: out = 16'(7055);
			1441: out = 16'(4178);
			1442: out = 16'(-8825);
			1443: out = 16'(-6630);
			1444: out = 16'(5541);
			1445: out = 16'(16159);
			1446: out = 16'(9127);
			1447: out = 16'(13573);
			1448: out = 16'(14327);
			1449: out = 16'(4344);
			1450: out = 16'(18679);
			1451: out = 16'(10267);
			1452: out = 16'(-4301);
			1453: out = 16'(-15274);
			1454: out = 16'(3123);
			1455: out = 16'(1095);
			1456: out = 16'(-2273);
			1457: out = 16'(4684);
			1458: out = 16'(28753);
			1459: out = 16'(10410);
			1460: out = 16'(-6596);
			1461: out = 16'(-10345);
			1462: out = 16'(7318);
			1463: out = 16'(-5435);
			1464: out = 16'(-5132);
			1465: out = 16'(2355);
			1466: out = 16'(11363);
			1467: out = 16'(-2860);
			1468: out = 16'(-1048);
			1469: out = 16'(-5544);
			1470: out = 16'(-20395);
			1471: out = 16'(-19137);
			1472: out = 16'(-11244);
			1473: out = 16'(-4500);
			1474: out = 16'(-1151);
			1475: out = 16'(7282);
			1476: out = 16'(14546);
			1477: out = 16'(5733);
			1478: out = 16'(-6757);
			1479: out = 16'(8793);
			1480: out = 16'(3906);
			1481: out = 16'(1846);
			1482: out = 16'(-994);
			1483: out = 16'(7771);
			1484: out = 16'(-19413);
			1485: out = 16'(-17380);
			1486: out = 16'(-7136);
			1487: out = 16'(-3652);
			1488: out = 16'(-20609);
			1489: out = 16'(-10200);
			1490: out = 16'(-4894);
			1491: out = 16'(-25191);
			1492: out = 16'(-28061);
			1493: out = 16'(-28195);
			1494: out = 16'(-10684);
			1495: out = 16'(6611);
			1496: out = 16'(14451);
			1497: out = 16'(5170);
			1498: out = 16'(-2161);
			1499: out = 16'(-3186);
			1500: out = 16'(1539);
			1501: out = 16'(-7890);
			1502: out = 16'(-9013);
			1503: out = 16'(-2913);
			1504: out = 16'(841);
			1505: out = 16'(-12640);
			1506: out = 16'(-14138);
			1507: out = 16'(-705);
			1508: out = 16'(12664);
			1509: out = 16'(6336);
			1510: out = 16'(2929);
			1511: out = 16'(4211);
			1512: out = 16'(4469);
			1513: out = 16'(-18941);
			1514: out = 16'(-6141);
			1515: out = 16'(5445);
			1516: out = 16'(6388);
			1517: out = 16'(2208);
			1518: out = 16'(4737);
			1519: out = 16'(8457);
			1520: out = 16'(10826);
			1521: out = 16'(9385);
			1522: out = 16'(3202);
			1523: out = 16'(-524);
			1524: out = 16'(554);
			1525: out = 16'(3738);
			1526: out = 16'(13783);
			1527: out = 16'(13834);
			1528: out = 16'(15374);
			1529: out = 16'(14601);
			1530: out = 16'(4782);
			1531: out = 16'(-1376);
			1532: out = 16'(934);
			1533: out = 16'(-108);
			1534: out = 16'(-20304);
			1535: out = 16'(-8375);
			1536: out = 16'(16537);
			1537: out = 16'(29531);
			1538: out = 16'(22276);
			1539: out = 16'(20140);
			1540: out = 16'(17814);
			1541: out = 16'(9597);
			1542: out = 16'(-8440);
			1543: out = 16'(-3590);
			1544: out = 16'(-445);
			1545: out = 16'(5563);
			1546: out = 16'(11805);
			1547: out = 16'(20407);
			1548: out = 16'(17720);
			1549: out = 16'(7577);
			1550: out = 16'(-3965);
			1551: out = 16'(-1685);
			1552: out = 16'(-3074);
			1553: out = 16'(311);
			1554: out = 16'(4479);
			1555: out = 16'(11247);
			1556: out = 16'(14372);
			1557: out = 16'(16182);
			1558: out = 16'(2375);
			1559: out = 16'(-26679);
			1560: out = 16'(-17036);
			1561: out = 16'(-6148);
			1562: out = 16'(-5639);
			1563: out = 16'(-19224);
			1564: out = 16'(-16407);
			1565: out = 16'(-19079);
			1566: out = 16'(-19632);
			1567: out = 16'(-22515);
			1568: out = 16'(-9386);
			1569: out = 16'(-12585);
			1570: out = 16'(-5549);
			1571: out = 16'(-1894);
			1572: out = 16'(-8155);
			1573: out = 16'(-22044);
			1574: out = 16'(-7620);
			1575: out = 16'(11635);
			1576: out = 16'(2575);
			1577: out = 16'(-2591);
			1578: out = 16'(-7366);
			1579: out = 16'(-14139);
			1580: out = 16'(-29284);
			1581: out = 16'(-21650);
			1582: out = 16'(-12074);
			1583: out = 16'(-7617);
			1584: out = 16'(-8502);
			1585: out = 16'(17140);
			1586: out = 16'(9103);
			1587: out = 16'(-10340);
			1588: out = 16'(-26305);
			1589: out = 16'(-7259);
			1590: out = 16'(-7895);
			1591: out = 16'(-9003);
			1592: out = 16'(-2927);
			1593: out = 16'(20011);
			1594: out = 16'(12372);
			1595: out = 16'(10045);
			1596: out = 16'(5757);
			1597: out = 16'(2215);
			1598: out = 16'(-18531);
			1599: out = 16'(-10116);
			1600: out = 16'(5363);
			1601: out = 16'(5180);
			1602: out = 16'(4104);
			1603: out = 16'(7035);
			1604: out = 16'(16618);
			1605: out = 16'(18960);
			1606: out = 16'(6340);
			1607: out = 16'(1057);
			1608: out = 16'(-3316);
			1609: out = 16'(-9950);
			1610: out = 16'(-14297);
			1611: out = 16'(-7983);
			1612: out = 16'(12422);
			1613: out = 16'(30349);
			1614: out = 16'(29382);
			1615: out = 16'(27011);
			1616: out = 16'(10184);
			1617: out = 16'(-3004);
			1618: out = 16'(-5293);
			1619: out = 16'(-12533);
			1620: out = 16'(-437);
			1621: out = 16'(19380);
			1622: out = 16'(29766);
			1623: out = 16'(29856);
			1624: out = 16'(23168);
			1625: out = 16'(9557);
			1626: out = 16'(-7513);
			1627: out = 16'(-17207);
			1628: out = 16'(-27639);
			1629: out = 16'(-20404);
			1630: out = 16'(2072);
			1631: out = 16'(22909);
			1632: out = 16'(29054);
			1633: out = 16'(30592);
			1634: out = 16'(23079);
			1635: out = 16'(-4155);
			1636: out = 16'(-24524);
			1637: out = 16'(-27794);
			1638: out = 16'(-8146);
			1639: out = 16'(6734);
			1640: out = 16'(6092);
			1641: out = 16'(-1759);
			1642: out = 16'(10035);
			1643: out = 16'(22251);
			1644: out = 16'(-4616);
			1645: out = 16'(-25375);
			1646: out = 16'(-24244);
			1647: out = 16'(-6703);
			1648: out = 16'(-11861);
			1649: out = 16'(-25712);
			1650: out = 16'(-24997);
			1651: out = 16'(-3648);
			1652: out = 16'(7062);
			1653: out = 16'(-8443);
			1654: out = 16'(-25979);
			1655: out = 16'(-22990);
			1656: out = 16'(-1514);
			1657: out = 16'(-608);
			1658: out = 16'(-5353);
			1659: out = 16'(-13729);
			1660: out = 16'(-15227);
			1661: out = 16'(143);
			1662: out = 16'(3237);
			1663: out = 16'(-9845);
			1664: out = 16'(-22157);
			1665: out = 16'(-3287);
			1666: out = 16'(11538);
			1667: out = 16'(14565);
			1668: out = 16'(586);
			1669: out = 16'(-21671);
			1670: out = 16'(-12135);
			1671: out = 16'(-86);
			1672: out = 16'(-3645);
			1673: out = 16'(-15686);
			1674: out = 16'(-13917);
			1675: out = 16'(2973);
			1676: out = 16'(13052);
			1677: out = 16'(5015);
			1678: out = 16'(1380);
			1679: out = 16'(3747);
			1680: out = 16'(13772);
			1681: out = 16'(13216);
			1682: out = 16'(5022);
			1683: out = 16'(-1241);
			1684: out = 16'(11196);
			1685: out = 16'(19325);
			1686: out = 16'(6143);
			1687: out = 16'(2542);
			1688: out = 16'(13161);
			1689: out = 16'(16276);
			1690: out = 16'(-5506);
			1691: out = 16'(-10802);
			1692: out = 16'(-742);
			1693: out = 16'(14355);
			1694: out = 16'(13183);
			1695: out = 16'(17907);
			1696: out = 16'(9810);
			1697: out = 16'(1703);
			1698: out = 16'(-4446);
			1699: out = 16'(8698);
			1700: out = 16'(3686);
			1701: out = 16'(-2696);
			1702: out = 16'(-2178);
			1703: out = 16'(16315);
			1704: out = 16'(13918);
			1705: out = 16'(10977);
			1706: out = 16'(7217);
			1707: out = 16'(7166);
			1708: out = 16'(6942);
			1709: out = 16'(8162);
			1710: out = 16'(2004);
			1711: out = 16'(-5855);
			1712: out = 16'(-6164);
			1713: out = 16'(1326);
			1714: out = 16'(-1310);
			1715: out = 16'(-9325);
			1716: out = 16'(-2202);
			1717: out = 16'(12662);
			1718: out = 16'(12327);
			1719: out = 16'(1768);
			1720: out = 16'(4071);
			1721: out = 16'(422);
			1722: out = 16'(-16152);
			1723: out = 16'(-25990);
			1724: out = 16'(4424);
			1725: out = 16'(11171);
			1726: out = 16'(1674);
			1727: out = 16'(-6624);
			1728: out = 16'(9898);
			1729: out = 16'(12376);
			1730: out = 16'(6090);
			1731: out = 16'(-7875);
			1732: out = 16'(-9330);
			1733: out = 16'(-18781);
			1734: out = 16'(-17847);
			1735: out = 16'(-23660);
			1736: out = 16'(-21883);
			1737: out = 16'(-2703);
			1738: out = 16'(17402);
			1739: out = 16'(8648);
			1740: out = 16'(-11117);
			1741: out = 16'(-8367);
			1742: out = 16'(-8568);
			1743: out = 16'(-11559);
			1744: out = 16'(-11492);
			1745: out = 16'(854);
			1746: out = 16'(-3768);
			1747: out = 16'(-9964);
			1748: out = 16'(-1352);
			1749: out = 16'(21511);
			1750: out = 16'(20559);
			1751: out = 16'(7435);
			1752: out = 16'(-2471);
			1753: out = 16'(1283);
			1754: out = 16'(-8177);
			1755: out = 16'(-10507);
			1756: out = 16'(-3497);
			1757: out = 16'(12475);
			1758: out = 16'(11320);
			1759: out = 16'(15690);
			1760: out = 16'(12287);
			1761: out = 16'(4850);
			1762: out = 16'(-15126);
			1763: out = 16'(-12100);
			1764: out = 16'(-6746);
			1765: out = 16'(831);
			1766: out = 16'(-622);
			1767: out = 16'(7047);
			1768: out = 16'(463);
			1769: out = 16'(3320);
			1770: out = 16'(11452);
			1771: out = 16'(7892);
			1772: out = 16'(-18660);
			1773: out = 16'(-24247);
			1774: out = 16'(3391);
			1775: out = 16'(12405);
			1776: out = 16'(11441);
			1777: out = 16'(10109);
			1778: out = 16'(8676);
			1779: out = 16'(-16821);
			1780: out = 16'(-26954);
			1781: out = 16'(-25120);
			1782: out = 16'(-15833);
			1783: out = 16'(-24911);
			1784: out = 16'(-7289);
			1785: out = 16'(7211);
			1786: out = 16'(19357);
			1787: out = 16'(19057);
			1788: out = 16'(17035);
			1789: out = 16'(5732);
			1790: out = 16'(6179);
			1791: out = 16'(11865);
			1792: out = 16'(3870);
			1793: out = 16'(-703);
			1794: out = 16'(9314);
			1795: out = 16'(20607);
			1796: out = 16'(11913);
			1797: out = 16'(83);
			1798: out = 16'(-40);
			1799: out = 16'(13122);
			1800: out = 16'(21502);
			1801: out = 16'(14705);
			1802: out = 16'(9135);
			1803: out = 16'(4883);
			1804: out = 16'(-3368);
			1805: out = 16'(-659);
			1806: out = 16'(9143);
			1807: out = 16'(12784);
			1808: out = 16'(351);
			1809: out = 16'(6362);
			1810: out = 16'(-5096);
			1811: out = 16'(-18424);
			1812: out = 16'(-26189);
			1813: out = 16'(9390);
			1814: out = 16'(2826);
			1815: out = 16'(-518);
			1816: out = 16'(6527);
			1817: out = 16'(23361);
			1818: out = 16'(-9819);
			1819: out = 16'(-30688);
			1820: out = 16'(-27999);
			1821: out = 16'(-28396);
			1822: out = 16'(-2820);
			1823: out = 16'(22045);
			1824: out = 16'(25757);
			1825: out = 16'(13229);
			1826: out = 16'(-8430);
			1827: out = 16'(-11558);
			1828: out = 16'(-14539);
			1829: out = 16'(-29313);
			1830: out = 16'(-28804);
			1831: out = 16'(-18812);
			1832: out = 16'(597);
			1833: out = 16'(6372);
			1834: out = 16'(9170);
			1835: out = 16'(2366);
			1836: out = 16'(2798);
			1837: out = 16'(6023);
			1838: out = 16'(12238);
			1839: out = 16'(-11400);
			1840: out = 16'(-23380);
			1841: out = 16'(-16985);
			1842: out = 16'(1602);
			1843: out = 16'(-14621);
			1844: out = 16'(-9950);
			1845: out = 16'(8062);
			1846: out = 16'(15357);
			1847: out = 16'(-8889);
			1848: out = 16'(-24961);
			1849: out = 16'(-25227);
			1850: out = 16'(-7837);
			1851: out = 16'(15270);
			1852: out = 16'(29692);
			1853: out = 16'(27384);
			1854: out = 16'(19897);
			1855: out = 16'(12251);
			1856: out = 16'(13742);
			1857: out = 16'(1251);
			1858: out = 16'(-10704);
			1859: out = 16'(2010);
			1860: out = 16'(15591);
			1861: out = 16'(17112);
			1862: out = 16'(9563);
			1863: out = 16'(12902);
			1864: out = 16'(6914);
			1865: out = 16'(9766);
			1866: out = 16'(808);
			1867: out = 16'(-12540);
			1868: out = 16'(-16246);
			1869: out = 16'(2696);
			1870: out = 16'(19240);
			1871: out = 16'(19088);
			1872: out = 16'(110);
			1873: out = 16'(11744);
			1874: out = 16'(22593);
			1875: out = 16'(17795);
			1876: out = 16'(-7322);
			1877: out = 16'(-2856);
			1878: out = 16'(-4770);
			1879: out = 16'(-12395);
			1880: out = 16'(-20276);
			1881: out = 16'(11);
			1882: out = 16'(2734);
			1883: out = 16'(-1893);
			1884: out = 16'(-685);
			1885: out = 16'(-802);
			1886: out = 16'(-12797);
			1887: out = 16'(-18941);
			1888: out = 16'(-5284);
			1889: out = 16'(-1976);
			1890: out = 16'(-6004);
			1891: out = 16'(-16204);
			1892: out = 16'(-16091);
			1893: out = 16'(-20522);
			1894: out = 16'(-3290);
			1895: out = 16'(-2548);
			1896: out = 16'(-11409);
			1897: out = 16'(-21909);
			1898: out = 16'(857);
			1899: out = 16'(6962);
			1900: out = 16'(1100);
			1901: out = 16'(260);
			1902: out = 16'(8660);
			1903: out = 16'(-152);
			1904: out = 16'(-17523);
			1905: out = 16'(-24567);
			1906: out = 16'(-2272);
			1907: out = 16'(1274);
			1908: out = 16'(-4188);
			1909: out = 16'(-684);
			1910: out = 16'(12199);
			1911: out = 16'(5484);
			1912: out = 16'(-7498);
			1913: out = 16'(-14960);
			1914: out = 16'(-23865);
			1915: out = 16'(-122);
			1916: out = 16'(15637);
			1917: out = 16'(16919);
			1918: out = 16'(10217);
			1919: out = 16'(9388);
			1920: out = 16'(4620);
			1921: out = 16'(-768);
			1922: out = 16'(-3415);
			1923: out = 16'(8781);
			1924: out = 16'(7382);
			1925: out = 16'(5592);
			1926: out = 16'(12503);
			1927: out = 16'(24304);
			1928: out = 16'(20376);
			1929: out = 16'(8602);
			1930: out = 16'(-2721);
			1931: out = 16'(-11039);
			1932: out = 16'(-9280);
			1933: out = 16'(-4568);
			1934: out = 16'(-1124);
			1935: out = 16'(1930);
			1936: out = 16'(23570);
			1937: out = 16'(31196);
			1938: out = 16'(19028);
			1939: out = 16'(-3607);
			1940: out = 16'(-1739);
			1941: out = 16'(-5590);
			1942: out = 16'(-16971);
			1943: out = 16'(-23737);
			1944: out = 16'(4277);
			1945: out = 16'(26264);
			1946: out = 16'(25579);
			1947: out = 16'(11989);
			1948: out = 16'(5058);
			1949: out = 16'(10072);
			1950: out = 16'(11818);
			1951: out = 16'(3629);
			1952: out = 16'(-607);
			1953: out = 16'(-3073);
			1954: out = 16'(3235);
			1955: out = 16'(6434);
			1956: out = 16'(4304);
			1957: out = 16'(-9145);
			1958: out = 16'(-8785);
			1959: out = 16'(-307);
			1960: out = 16'(959);
			1961: out = 16'(-22453);
			1962: out = 16'(-31143);
			1963: out = 16'(-20926);
			1964: out = 16'(-2176);
			1965: out = 16'(-15556);
			1966: out = 16'(-8824);
			1967: out = 16'(-4613);
			1968: out = 16'(-1071);
			1969: out = 16'(11168);
			1970: out = 16'(125);
			1971: out = 16'(-20341);
			1972: out = 16'(-27377);
			1973: out = 16'(-1785);
			1974: out = 16'(-3437);
			1975: out = 16'(-8481);
			1976: out = 16'(-6908);
			1977: out = 16'(5051);
			1978: out = 16'(-8392);
			1979: out = 16'(-12143);
			1980: out = 16'(-6988);
			1981: out = 16'(8442);
			1982: out = 16'(15518);
			1983: out = 16'(12688);
			1984: out = 16'(-4462);
			1985: out = 16'(-13482);
			1986: out = 16'(3463);
			1987: out = 16'(21541);
			1988: out = 16'(21647);
			1989: out = 16'(15224);
			1990: out = 16'(11111);
			1991: out = 16'(3943);
			1992: out = 16'(-9548);
			1993: out = 16'(-12719);
			1994: out = 16'(-4555);
			1995: out = 16'(-1327);
			1996: out = 16'(-19029);
			1997: out = 16'(-18371);
			1998: out = 16'(12028);
			1999: out = 16'(12632);
			2000: out = 16'(-3824);
			2001: out = 16'(-3782);
			2002: out = 16'(23990);
			2003: out = 16'(13684);
			2004: out = 16'(11136);
			2005: out = 16'(113);
			2006: out = 16'(1934);
			2007: out = 16'(-2155);
			2008: out = 16'(2846);
			2009: out = 16'(-13314);
			2010: out = 16'(-19881);
			2011: out = 16'(-1266);
			2012: out = 16'(11172);
			2013: out = 16'(5711);
			2014: out = 16'(1337);
			2015: out = 16'(4859);
			2016: out = 16'(-2869);
			2017: out = 16'(-17859);
			2018: out = 16'(-15938);
			2019: out = 16'(7034);
			2020: out = 16'(6701);
			2021: out = 16'(3506);
			2022: out = 16'(2350);
			2023: out = 16'(8241);
			2024: out = 16'(3534);
			2025: out = 16'(9971);
			2026: out = 16'(14024);
			2027: out = 16'(9659);
			2028: out = 16'(-12478);
			2029: out = 16'(-27598);
			2030: out = 16'(-23760);
			2031: out = 16'(-4396);
			2032: out = 16'(3820);
			2033: out = 16'(5273);
			2034: out = 16'(5716);
			2035: out = 16'(7284);
			2036: out = 16'(528);
			2037: out = 16'(2499);
			2038: out = 16'(-6839);
			2039: out = 16'(-3892);
			2040: out = 16'(4423);
			2041: out = 16'(1005);
			2042: out = 16'(-6546);
			2043: out = 16'(-3399);
			2044: out = 16'(11248);
			2045: out = 16'(25347);
			2046: out = 16'(9211);
			2047: out = 16'(-2259);
			2048: out = 16'(-5585);
			2049: out = 16'(-3250);
			2050: out = 16'(-6028);
			2051: out = 16'(9485);
			2052: out = 16'(25514);
			2053: out = 16'(22789);
			2054: out = 16'(13118);
			2055: out = 16'(2614);
			2056: out = 16'(-4264);
			2057: out = 16'(-11918);
			2058: out = 16'(-18899);
			2059: out = 16'(-10826);
			2060: out = 16'(-156);
			2061: out = 16'(-1354);
			2062: out = 16'(1272);
			2063: out = 16'(3890);
			2064: out = 16'(19073);
			2065: out = 16'(23918);
			2066: out = 16'(12578);
			2067: out = 16'(-7471);
			2068: out = 16'(-14865);
			2069: out = 16'(-12527);
			2070: out = 16'(-5230);
			2071: out = 16'(-2542);
			2072: out = 16'(14289);
			2073: out = 16'(24202);
			2074: out = 16'(21421);
			2075: out = 16'(5932);
			2076: out = 16'(754);
			2077: out = 16'(-17435);
			2078: out = 16'(-29281);
			2079: out = 16'(-30090);
			2080: out = 16'(-2894);
			2081: out = 16'(15179);
			2082: out = 16'(9527);
			2083: out = 16'(14662);
			2084: out = 16'(20287);
			2085: out = 16'(9601);
			2086: out = 16'(-10543);
			2087: out = 16'(1673);
			2088: out = 16'(1339);
			2089: out = 16'(7409);
			2090: out = 16'(-9233);
			2091: out = 16'(-26145);
			2092: out = 16'(-30297);
			2093: out = 16'(234);
			2094: out = 16'(12915);
			2095: out = 16'(537);
			2096: out = 16'(-9101);
			2097: out = 16'(-5461);
			2098: out = 16'(-15580);
			2099: out = 16'(-30952);
			2100: out = 16'(-19274);
			2101: out = 16'(8565);
			2102: out = 16'(22473);
			2103: out = 16'(15846);
			2104: out = 16'(3380);
			2105: out = 16'(-8977);
			2106: out = 16'(-22545);
			2107: out = 16'(-25031);
			2108: out = 16'(-8430);
			2109: out = 16'(-10761);
			2110: out = 16'(-15804);
			2111: out = 16'(-4003);
			2112: out = 16'(26137);
			2113: out = 16'(26566);
			2114: out = 16'(10647);
			2115: out = 16'(-8625);
			2116: out = 16'(-9917);
			2117: out = 16'(-23906);
			2118: out = 16'(-13767);
			2119: out = 16'(-11156);
			2120: out = 16'(-2676);
			2121: out = 16'(8156);
			2122: out = 16'(15926);
			2123: out = 16'(-10518);
			2124: out = 16'(-29676);
			2125: out = 16'(-11966);
			2126: out = 16'(16747);
			2127: out = 16'(7423);
			2128: out = 16'(-11215);
			2129: out = 16'(-3511);
			2130: out = 16'(12722);
			2131: out = 16'(10156);
			2132: out = 16'(-4748);
			2133: out = 16'(-3167);
			2134: out = 16'(13084);
			2135: out = 16'(21540);
			2136: out = 16'(12546);
			2137: out = 16'(6078);
			2138: out = 16'(14415);
			2139: out = 16'(10667);
			2140: out = 16'(-3202);
			2141: out = 16'(-17964);
			2142: out = 16'(-23693);
			2143: out = 16'(-2307);
			2144: out = 16'(15266);
			2145: out = 16'(17128);
			2146: out = 16'(6330);
			2147: out = 16'(5340);
			2148: out = 16'(6123);
			2149: out = 16'(17528);
			2150: out = 16'(25892);
			2151: out = 16'(21881);
			2152: out = 16'(0);
			2153: out = 16'(-14588);
			2154: out = 16'(-15157);
			2155: out = 16'(-9704);
			2156: out = 16'(-10997);
			2157: out = 16'(4402);
			2158: out = 16'(23001);
			2159: out = 16'(13447);
			2160: out = 16'(907);
			2161: out = 16'(-5263);
			2162: out = 16'(1289);
			2163: out = 16'(-2038);
			2164: out = 16'(1036);
			2165: out = 16'(-3030);
			2166: out = 16'(-461);
			2167: out = 16'(-340);
			2168: out = 16'(1089);
			2169: out = 16'(-8382);
			2170: out = 16'(-1591);
			2171: out = 16'(16133);
			2172: out = 16'(19887);
			2173: out = 16'(13346);
			2174: out = 16'(7385);
			2175: out = 16'(215);
			2176: out = 16'(-12990);
			2177: out = 16'(-18252);
			2178: out = 16'(-1080);
			2179: out = 16'(17376);
			2180: out = 16'(13250);
			2181: out = 16'(2653);
			2182: out = 16'(6845);
			2183: out = 16'(10821);
			2184: out = 16'(-17002);
			2185: out = 16'(-27622);
			2186: out = 16'(-27295);
			2187: out = 16'(-2360);
			2188: out = 16'(17223);
			2189: out = 16'(18141);
			2190: out = 16'(11210);
			2191: out = 16'(6371);
			2192: out = 16'(-653);
			2193: out = 16'(-9167);
			2194: out = 16'(-22266);
			2195: out = 16'(-15867);
			2196: out = 16'(5659);
			2197: out = 16'(19725);
			2198: out = 16'(18538);
			2199: out = 16'(13277);
			2200: out = 16'(8794);
			2201: out = 16'(6814);
			2202: out = 16'(-22502);
			2203: out = 16'(-29653);
			2204: out = 16'(-29173);
			2205: out = 16'(-25789);
			2206: out = 16'(-4362);
			2207: out = 16'(9759);
			2208: out = 16'(385);
			2209: out = 16'(-16848);
			2210: out = 16'(-6530);
			2211: out = 16'(7392);
			2212: out = 16'(1498);
			2213: out = 16'(-18318);
			2214: out = 16'(-21736);
			2215: out = 16'(-9452);
			2216: out = 16'(-12309);
			2217: out = 16'(-31590);
			2218: out = 16'(-25747);
			2219: out = 16'(693);
			2220: out = 16'(29407);
			2221: out = 16'(20808);
			2222: out = 16'(1732);
			2223: out = 16'(-24457);
			2224: out = 16'(-10276);
			2225: out = 16'(-2522);
			2226: out = 16'(-16804);
			2227: out = 16'(-25726);
			2228: out = 16'(1685);
			2229: out = 16'(24917);
			2230: out = 16'(19519);
			2231: out = 16'(7404);
			2232: out = 16'(6012);
			2233: out = 16'(5937);
			2234: out = 16'(-624);
			2235: out = 16'(-6493);
			2236: out = 16'(5025);
			2237: out = 16'(10764);
			2238: out = 16'(10863);
			2239: out = 16'(16640);
			2240: out = 16'(18653);
			2241: out = 16'(15732);
			2242: out = 16'(10600);
			2243: out = 16'(12786);
			2244: out = 16'(13314);
			2245: out = 16'(8298);
			2246: out = 16'(-1922);
			2247: out = 16'(-5248);
			2248: out = 16'(-6792);
			2249: out = 16'(10136);
			2250: out = 16'(15555);
			2251: out = 16'(3378);
			2252: out = 16'(-28151);
			2253: out = 16'(-13364);
			2254: out = 16'(2368);
			2255: out = 16'(6882);
			2256: out = 16'(3211);
			2257: out = 16'(13422);
			2258: out = 16'(7786);
			2259: out = 16'(3555);
			2260: out = 16'(8164);
			2261: out = 16'(10759);
			2262: out = 16'(3999);
			2263: out = 16'(744);
			2264: out = 16'(1842);
			2265: out = 16'(235);
			2266: out = 16'(-14004);
			2267: out = 16'(-7028);
			2268: out = 16'(17481);
			2269: out = 16'(14036);
			2270: out = 16'(-1541);
			2271: out = 16'(-18104);
			2272: out = 16'(-17872);
			2273: out = 16'(-14970);
			2274: out = 16'(-17031);
			2275: out = 16'(-13237);
			2276: out = 16'(7967);
			2277: out = 16'(19414);
			2278: out = 16'(23829);
			2279: out = 16'(-6320);
			2280: out = 16'(-30415);
			2281: out = 16'(-26656);
			2282: out = 16'(13842);
			2283: out = 16'(13265);
			2284: out = 16'(-4518);
			2285: out = 16'(-3313);
			2286: out = 16'(24344);
			2287: out = 16'(21713);
			2288: out = 16'(4611);
			2289: out = 16'(-15326);
			2290: out = 16'(-28961);
			2291: out = 16'(-28028);
			2292: out = 16'(-23344);
			2293: out = 16'(-11141);
			2294: out = 16'(1612);
			2295: out = 16'(16383);
			2296: out = 16'(10390);
			2297: out = 16'(-5472);
			2298: out = 16'(-15438);
			2299: out = 16'(-20768);
			2300: out = 16'(-3253);
			2301: out = 16'(13819);
			2302: out = 16'(14287);
			2303: out = 16'(13712);
			2304: out = 16'(11127);
			2305: out = 16'(14214);
			2306: out = 16'(12674);
			2307: out = 16'(7954);
			2308: out = 16'(-11029);
			2309: out = 16'(-15475);
			2310: out = 16'(-5551);
			2311: out = 16'(3246);
			2312: out = 16'(-14452);
			2313: out = 16'(-18083);
			2314: out = 16'(638);
			2315: out = 16'(16465);
			2316: out = 16'(211);
			2317: out = 16'(-13267);
			2318: out = 16'(-13940);
			2319: out = 16'(-8464);
			2320: out = 16'(-10776);
			2321: out = 16'(-12048);
			2322: out = 16'(-9101);
			2323: out = 16'(-3163);
			2324: out = 16'(12820);
			2325: out = 16'(11724);
			2326: out = 16'(4995);
			2327: out = 16'(-6106);
			2328: out = 16'(-3797);
			2329: out = 16'(-6769);
			2330: out = 16'(11719);
			2331: out = 16'(25111);
			2332: out = 16'(17099);
			2333: out = 16'(-1914);
			2334: out = 16'(-3906);
			2335: out = 16'(2368);
			2336: out = 16'(-139);
			2337: out = 16'(-15350);
			2338: out = 16'(-4592);
			2339: out = 16'(15001);
			2340: out = 16'(15360);
			2341: out = 16'(3100);
			2342: out = 16'(1446);
			2343: out = 16'(6890);
			2344: out = 16'(6541);
			2345: out = 16'(8136);
			2346: out = 16'(9344);
			2347: out = 16'(15405);
			2348: out = 16'(14074);
			2349: out = 16'(3294);
			2350: out = 16'(-14455);
			2351: out = 16'(-15051);
			2352: out = 16'(4282);
			2353: out = 16'(18246);
			2354: out = 16'(15003);
			2355: out = 16'(1253);
			2356: out = 16'(-2367);
			2357: out = 16'(6125);
			2358: out = 16'(3546);
			2359: out = 16'(-13436);
			2360: out = 16'(-24766);
			2361: out = 16'(-7471);
			2362: out = 16'(13117);
			2363: out = 16'(20906);
			2364: out = 16'(8291);
			2365: out = 16'(513);
			2366: out = 16'(7859);
			2367: out = 16'(17479);
			2368: out = 16'(1515);
			2369: out = 16'(-24333);
			2370: out = 16'(-28444);
			2371: out = 16'(-15699);
			2372: out = 16'(-8864);
			2373: out = 16'(-17411);
			2374: out = 16'(-21636);
			2375: out = 16'(-17413);
			2376: out = 16'(98);
			2377: out = 16'(8655);
			2378: out = 16'(3129);
			2379: out = 16'(160);
			2380: out = 16'(6482);
			2381: out = 16'(16239);
			2382: out = 16'(9304);
			2383: out = 16'(-9183);
			2384: out = 16'(-26963);
			2385: out = 16'(-8832);
			2386: out = 16'(18106);
			2387: out = 16'(9155);
			2388: out = 16'(110);
			2389: out = 16'(4202);
			2390: out = 16'(17511);
			2391: out = 16'(8348);
			2392: out = 16'(-259);
			2393: out = 16'(-15369);
			2394: out = 16'(-10292);
			2395: out = 16'(3975);
			2396: out = 16'(6676);
			2397: out = 16'(-4680);
			2398: out = 16'(-3384);
			2399: out = 16'(14394);
			2400: out = 16'(24137);
			2401: out = 16'(15780);
			2402: out = 16'(-2036);
			2403: out = 16'(-18677);
			2404: out = 16'(-24786);
			2405: out = 16'(-15303);
			2406: out = 16'(1968);
			2407: out = 16'(6874);
			2408: out = 16'(-3279);
			2409: out = 16'(-5700);
			2410: out = 16'(2221);
			2411: out = 16'(6402);
			2412: out = 16'(-330);
			2413: out = 16'(-1683);
			2414: out = 16'(10239);
			2415: out = 16'(17819);
			2416: out = 16'(8130);
			2417: out = 16'(-1662);
			2418: out = 16'(-11358);
			2419: out = 16'(-14699);
			2420: out = 16'(-18824);
			2421: out = 16'(-24053);
			2422: out = 16'(-5381);
			2423: out = 16'(17326);
			2424: out = 16'(19549);
			2425: out = 16'(3987);
			2426: out = 16'(-9482);
			2427: out = 16'(-11891);
			2428: out = 16'(-6383);
			2429: out = 16'(-1396);
			2430: out = 16'(-7550);
			2431: out = 16'(-1352);
			2432: out = 16'(6580);
			2433: out = 16'(2380);
			2434: out = 16'(-5943);
			2435: out = 16'(-10307);
			2436: out = 16'(-2331);
			2437: out = 16'(4406);
			2438: out = 16'(1758);
			2439: out = 16'(-11671);
			2440: out = 16'(-10380);
			2441: out = 16'(5939);
			2442: out = 16'(9904);
			2443: out = 16'(15080);
			2444: out = 16'(4818);
			2445: out = 16'(-9427);
			2446: out = 16'(-19125);
			2447: out = 16'(-1904);
			2448: out = 16'(10232);
			2449: out = 16'(13300);
			2450: out = 16'(14721);
			2451: out = 16'(19517);
			2452: out = 16'(22005);
			2453: out = 16'(14625);
			2454: out = 16'(-1019);
			2455: out = 16'(-755);
			2456: out = 16'(-10772);
			2457: out = 16'(-10180);
			2458: out = 16'(-688);
			2459: out = 16'(11504);
			2460: out = 16'(7412);
			2461: out = 16'(13817);
			2462: out = 16'(22560);
			2463: out = 16'(11400);
			2464: out = 16'(-19188);
			2465: out = 16'(-32679);
			2466: out = 16'(-15876);
			2467: out = 16'(14400);
			2468: out = 16'(11188);
			2469: out = 16'(2922);
			2470: out = 16'(265);
			2471: out = 16'(2508);
			2472: out = 16'(-6403);
			2473: out = 16'(-12476);
			2474: out = 16'(-6381);
			2475: out = 16'(8529);
			2476: out = 16'(2311);
			2477: out = 16'(2269);
			2478: out = 16'(-3655);
			2479: out = 16'(-5224);
			2480: out = 16'(-8332);
			2481: out = 16'(8166);
			2482: out = 16'(-3642);
			2483: out = 16'(-25549);
			2484: out = 16'(-22438);
			2485: out = 16'(-4076);
			2486: out = 16'(10390);
			2487: out = 16'(9021);
			2488: out = 16'(8270);
			2489: out = 16'(-15);
			2490: out = 16'(6913);
			2491: out = 16'(5774);
			2492: out = 16'(-4197);
			2493: out = 16'(-25344);
			2494: out = 16'(-7071);
			2495: out = 16'(9640);
			2496: out = 16'(4357);
			2497: out = 16'(-2546);
			2498: out = 16'(10533);
			2499: out = 16'(23381);
			2500: out = 16'(8545);
			2501: out = 16'(-25486);
			2502: out = 16'(-25526);
			2503: out = 16'(-1479);
			2504: out = 16'(12132);
			2505: out = 16'(-881);
			2506: out = 16'(-8062);
			2507: out = 16'(-5334);
			2508: out = 16'(2611);
			2509: out = 16'(-2662);
			2510: out = 16'(2457);
			2511: out = 16'(4116);
			2512: out = 16'(19199);
			2513: out = 16'(25102);
			2514: out = 16'(17489);
			2515: out = 16'(-3087);
			2516: out = 16'(623);
			2517: out = 16'(12673);
			2518: out = 16'(2395);
			2519: out = 16'(-18781);
			2520: out = 16'(-22790);
			2521: out = 16'(-8876);
			2522: out = 16'(-5996);
			2523: out = 16'(515);
			2524: out = 16'(2674);
			2525: out = 16'(2730);
			2526: out = 16'(-3592);
			2527: out = 16'(1739);
			2528: out = 16'(-1555);
			2529: out = 16'(-10303);
			2530: out = 16'(-17106);
			2531: out = 16'(-4204);
			2532: out = 16'(8734);
			2533: out = 16'(13357);
			2534: out = 16'(12471);
			2535: out = 16'(14545);
			2536: out = 16'(9523);
			2537: out = 16'(1799);
			2538: out = 16'(-1568);
			2539: out = 16'(-771);
			2540: out = 16'(-4419);
			2541: out = 16'(-18484);
			2542: out = 16'(-20240);
			2543: out = 16'(1215);
			2544: out = 16'(906);
			2545: out = 16'(-5291);
			2546: out = 16'(-4075);
			2547: out = 16'(9063);
			2548: out = 16'(7427);
			2549: out = 16'(-2550);
			2550: out = 16'(-7618);
			2551: out = 16'(6997);
			2552: out = 16'(25343);
			2553: out = 16'(25790);
			2554: out = 16'(8198);
			2555: out = 16'(-15984);
			2556: out = 16'(-27201);
			2557: out = 16'(-22609);
			2558: out = 16'(1021);
			2559: out = 16'(18183);
			2560: out = 16'(18152);
			2561: out = 16'(12705);
			2562: out = 16'(5791);
			2563: out = 16'(-8512);
			2564: out = 16'(-23305);
			2565: out = 16'(1759);
			2566: out = 16'(20092);
			2567: out = 16'(5544);
			2568: out = 16'(-29418);
			2569: out = 16'(-29140);
			2570: out = 16'(-14243);
			2571: out = 16'(11460);
			2572: out = 16'(7836);
			2573: out = 16'(114);
			2574: out = 16'(-3481);
			2575: out = 16'(11381);
			2576: out = 16'(12848);
			2577: out = 16'(5236);
			2578: out = 16'(-20474);
			2579: out = 16'(2362);
			2580: out = 16'(29887);
			2581: out = 16'(16270);
			2582: out = 16'(-22184);
			2583: out = 16'(-19064);
			2584: out = 16'(15881);
			2585: out = 16'(24647);
			2586: out = 16'(-1288);
			2587: out = 16'(-24430);
			2588: out = 16'(-24373);
			2589: out = 16'(-5079);
			2590: out = 16'(2752);
			2591: out = 16'(8300);
			2592: out = 16'(1630);
			2593: out = 16'(-6259);
			2594: out = 16'(-10816);
			2595: out = 16'(-991);
			2596: out = 16'(633);
			2597: out = 16'(10277);
			2598: out = 16'(28648);
			2599: out = 16'(30811);
			2600: out = 16'(-744);
			2601: out = 16'(-32079);
			2602: out = 16'(-24425);
			2603: out = 16'(-1875);
			2604: out = 16'(7789);
			2605: out = 16'(-1805);
			2606: out = 16'(-5697);
			2607: out = 16'(-8114);
			2608: out = 16'(15634);
			2609: out = 16'(24262);
			2610: out = 16'(13370);
			2611: out = 16'(-15772);
			2612: out = 16'(-11049);
			2613: out = 16'(-1109);
			2614: out = 16'(4086);
			2615: out = 16'(275);
			2616: out = 16'(15370);
			2617: out = 16'(12128);
			2618: out = 16'(3712);
			2619: out = 16'(-272);
			2620: out = 16'(134);
			2621: out = 16'(-2289);
			2622: out = 16'(2277);
			2623: out = 16'(10942);
			2624: out = 16'(3681);
			2625: out = 16'(-3889);
			2626: out = 16'(-1105);
			2627: out = 16'(12335);
			2628: out = 16'(14913);
			2629: out = 16'(7454);
			2630: out = 16'(-7739);
			2631: out = 16'(-21300);
			2632: out = 16'(-27812);
			2633: out = 16'(-25972);
			2634: out = 16'(-16040);
			2635: out = 16'(-7387);
			2636: out = 16'(-5927);
			2637: out = 16'(9636);
			2638: out = 16'(9797);
			2639: out = 16'(-4701);
			2640: out = 16'(-17779);
			2641: out = 16'(9440);
			2642: out = 16'(23010);
			2643: out = 16'(11568);
			2644: out = 16'(-12281);
			2645: out = 16'(-15624);
			2646: out = 16'(-10881);
			2647: out = 16'(-4480);
			2648: out = 16'(-5674);
			2649: out = 16'(-5530);
			2650: out = 16'(1318);
			2651: out = 16'(8335);
			2652: out = 16'(2428);
			2653: out = 16'(-16150);
			2654: out = 16'(-23636);
			2655: out = 16'(-13023);
			2656: out = 16'(7395);
			2657: out = 16'(12915);
			2658: out = 16'(10923);
			2659: out = 16'(-381);
			2660: out = 16'(3597);
			2661: out = 16'(14153);
			2662: out = 16'(11932);
			2663: out = 16'(-934);
			2664: out = 16'(1707);
			2665: out = 16'(15758);
			2666: out = 16'(15361);
			2667: out = 16'(-4780);
			2668: out = 16'(-10544);
			2669: out = 16'(6282);
			2670: out = 16'(12198);
			2671: out = 16'(2214);
			2672: out = 16'(-11885);
			2673: out = 16'(-4303);
			2674: out = 16'(18065);
			2675: out = 16'(20066);
			2676: out = 16'(8104);
			2677: out = 16'(-3686);
			2678: out = 16'(-2571);
			2679: out = 16'(1485);
			2680: out = 16'(2729);
			2681: out = 16'(-7832);
			2682: out = 16'(-14797);
			2683: out = 16'(5203);
			2684: out = 16'(16656);
			2685: out = 16'(10598);
			2686: out = 16'(-2475);
			2687: out = 16'(4309);
			2688: out = 16'(4296);
			2689: out = 16'(5983);
			2690: out = 16'(-1327);
			2691: out = 16'(-7285);
			2692: out = 16'(-11664);
			2693: out = 16'(291);
			2694: out = 16'(5132);
			2695: out = 16'(-1148);
			2696: out = 16'(-9509);
			2697: out = 16'(1531);
			2698: out = 16'(5783);
			2699: out = 16'(-7180);
			2700: out = 16'(-13403);
			2701: out = 16'(-4251);
			2702: out = 16'(11285);
			2703: out = 16'(12320);
			2704: out = 16'(494);
			2705: out = 16'(-8010);
			2706: out = 16'(-7687);
			2707: out = 16'(-2388);
			2708: out = 16'(-637);
			2709: out = 16'(-4012);
			2710: out = 16'(-4573);
			2711: out = 16'(7255);
			2712: out = 16'(21103);
			2713: out = 16'(8677);
			2714: out = 16'(-2528);
			2715: out = 16'(-4882);
			2716: out = 16'(-2184);
			2717: out = 16'(-15081);
			2718: out = 16'(-21799);
			2719: out = 16'(-9224);
			2720: out = 16'(12894);
			2721: out = 16'(8812);
			2722: out = 16'(8486);
			2723: out = 16'(4791);
			2724: out = 16'(-108);
			2725: out = 16'(-20855);
			2726: out = 16'(-8609);
			2727: out = 16'(-4866);
			2728: out = 16'(-9309);
			2729: out = 16'(-15532);
			2730: out = 16'(-5121);
			2731: out = 16'(34);
			2732: out = 16'(1995);
			2733: out = 16'(4701);
			2734: out = 16'(1416);
			2735: out = 16'(2985);
			2736: out = 16'(7010);
			2737: out = 16'(9518);
			2738: out = 16'(-2495);
			2739: out = 16'(-955);
			2740: out = 16'(1143);
			2741: out = 16'(-931);
			2742: out = 16'(-9954);
			2743: out = 16'(-4041);
			2744: out = 16'(2433);
			2745: out = 16'(3471);
			2746: out = 16'(-1332);
			2747: out = 16'(-2656);
			2748: out = 16'(398);
			2749: out = 16'(6434);
			2750: out = 16'(6196);
			2751: out = 16'(5781);
			2752: out = 16'(-5577);
			2753: out = 16'(-8364);
			2754: out = 16'(3588);
			2755: out = 16'(22727);
			2756: out = 16'(11943);
			2757: out = 16'(-3597);
			2758: out = 16'(-6859);
			2759: out = 16'(5648);
			2760: out = 16'(-4285);
			2761: out = 16'(-19910);
			2762: out = 16'(-23072);
			2763: out = 16'(1643);
			2764: out = 16'(20560);
			2765: out = 16'(26768);
			2766: out = 16'(10019);
			2767: out = 16'(-18003);
			2768: out = 16'(-30932);
			2769: out = 16'(-11688);
			2770: out = 16'(7449);
			2771: out = 16'(3438);
			2772: out = 16'(1104);
			2773: out = 16'(17231);
			2774: out = 16'(28128);
			2775: out = 16'(14223);
			2776: out = 16'(-15931);
			2777: out = 16'(-15540);
			2778: out = 16'(2074);
			2779: out = 16'(2889);
			2780: out = 16'(-11894);
			2781: out = 16'(-7931);
			2782: out = 16'(13695);
			2783: out = 16'(22358);
			2784: out = 16'(11008);
			2785: out = 16'(6456);
			2786: out = 16'(9826);
			2787: out = 16'(9059);
			2788: out = 16'(-2208);
			2789: out = 16'(-21664);
			2790: out = 16'(-24385);
			2791: out = 16'(-12504);
			2792: out = 16'(2586);
			2793: out = 16'(10918);
			2794: out = 16'(19747);
			2795: out = 16'(13425);
			2796: out = 16'(-550);
			2797: out = 16'(-490);
			2798: out = 16'(8610);
			2799: out = 16'(8002);
			2800: out = 16'(-4094);
			2801: out = 16'(-9003);
			2802: out = 16'(-6699);
			2803: out = 16'(-5024);
			2804: out = 16'(-10215);
			2805: out = 16'(-11867);
			2806: out = 16'(2368);
			2807: out = 16'(8095);
			2808: out = 16'(-836);
			2809: out = 16'(-10367);
			2810: out = 16'(-2508);
			2811: out = 16'(4290);
			2812: out = 16'(4113);
			2813: out = 16'(4211);
			2814: out = 16'(5447);
			2815: out = 16'(3446);
			2816: out = 16'(-8944);
			2817: out = 16'(-17965);
			2818: out = 16'(-6425);
			2819: out = 16'(-5573);
			2820: out = 16'(-11862);
			2821: out = 16'(-9488);
			2822: out = 16'(10304);
			2823: out = 16'(11216);
			2824: out = 16'(2315);
			2825: out = 16'(-1833);
			2826: out = 16'(6769);
			2827: out = 16'(-3118);
			2828: out = 16'(-17742);
			2829: out = 16'(-19856);
			2830: out = 16'(4436);
			2831: out = 16'(7999);
			2832: out = 16'(10714);
			2833: out = 16'(1996);
			2834: out = 16'(-42);
			2835: out = 16'(-1139);
			2836: out = 16'(9984);
			2837: out = 16'(-1469);
			2838: out = 16'(-18108);
			2839: out = 16'(-13678);
			2840: out = 16'(3025);
			2841: out = 16'(5655);
			2842: out = 16'(-536);
			2843: out = 16'(2894);
			2844: out = 16'(414);
			2845: out = 16'(-1586);
			2846: out = 16'(-598);
			2847: out = 16'(8460);
			2848: out = 16'(5160);
			2849: out = 16'(10647);
			2850: out = 16'(13679);
			2851: out = 16'(10561);
			2852: out = 16'(1139);
			2853: out = 16'(-14933);
			2854: out = 16'(-19701);
			2855: out = 16'(-5470);
			2856: out = 16'(8859);
			2857: out = 16'(11361);
			2858: out = 16'(8812);
			2859: out = 16'(12039);
			2860: out = 16'(13722);
			2861: out = 16'(3743);
			2862: out = 16'(-8621);
			2863: out = 16'(-8241);
			2864: out = 16'(-628);
			2865: out = 16'(1291);
			2866: out = 16'(-13662);
			2867: out = 16'(-16423);
			2868: out = 16'(4670);
			2869: out = 16'(16224);
			2870: out = 16'(19507);
			2871: out = 16'(11907);
			2872: out = 16'(-1470);
			2873: out = 16'(-17701);
			2874: out = 16'(-24413);
			2875: out = 16'(-14452);
			2876: out = 16'(-2388);
			2877: out = 16'(-4757);
			2878: out = 16'(9341);
			2879: out = 16'(15386);
			2880: out = 16'(5337);
			2881: out = 16'(-11700);
			2882: out = 16'(-5292);
			2883: out = 16'(9710);
			2884: out = 16'(3524);
			2885: out = 16'(-18292);
			2886: out = 16'(-949);
			2887: out = 16'(18071);
			2888: out = 16'(15138);
			2889: out = 16'(-5880);
			2890: out = 16'(-9695);
			2891: out = 16'(2672);
			2892: out = 16'(13605);
			2893: out = 16'(9624);
			2894: out = 16'(3575);
			2895: out = 16'(-95);
			2896: out = 16'(-5971);
			2897: out = 16'(-12652);
			2898: out = 16'(-8049);
			2899: out = 16'(3312);
			2900: out = 16'(11422);
			2901: out = 16'(10631);
			2902: out = 16'(5355);
			2903: out = 16'(778);
			2904: out = 16'(-7801);
			2905: out = 16'(-10438);
			2906: out = 16'(-733);
			2907: out = 16'(13569);
			2908: out = 16'(1152);
			2909: out = 16'(-15040);
			2910: out = 16'(-11404);
			2911: out = 16'(10428);
			2912: out = 16'(2638);
			2913: out = 16'(-15655);
			2914: out = 16'(-17886);
			2915: out = 16'(3468);
			2916: out = 16'(7557);
			2917: out = 16'(2425);
			2918: out = 16'(1973);
			2919: out = 16'(5490);
			2920: out = 16'(-3797);
			2921: out = 16'(-22281);
			2922: out = 16'(-21976);
			2923: out = 16'(4486);
			2924: out = 16'(14446);
			2925: out = 16'(11387);
			2926: out = 16'(1123);
			2927: out = 16'(-8742);
			2928: out = 16'(-11244);
			2929: out = 16'(-17946);
			2930: out = 16'(-9883);
			2931: out = 16'(4847);
			2932: out = 16'(13809);
			2933: out = 16'(5488);
			2934: out = 16'(9535);
			2935: out = 16'(9494);
			2936: out = 16'(-5930);
			2937: out = 16'(-26051);
			2938: out = 16'(-9023);
			2939: out = 16'(18496);
			2940: out = 16'(15824);
			2941: out = 16'(7059);
			2942: out = 16'(2252);
			2943: out = 16'(5140);
			2944: out = 16'(2448);
			2945: out = 16'(1353);
			2946: out = 16'(-6362);
			2947: out = 16'(-9819);
			2948: out = 16'(-5948);
			2949: out = 16'(6968);
			2950: out = 16'(17445);
			2951: out = 16'(16720);
			2952: out = 16'(7532);
			2953: out = 16'(-227);
			2954: out = 16'(-117);
			2955: out = 16'(-8161);
			2956: out = 16'(-20077);
			2957: out = 16'(-15729);
			2958: out = 16'(1889);
			2959: out = 16'(18028);
			2960: out = 16'(14045);
			2961: out = 16'(2809);
			2962: out = 16'(-676);
			2963: out = 16'(3211);
			2964: out = 16'(-4064);
			2965: out = 16'(-17613);
			2966: out = 16'(-10858);
			2967: out = 16'(8532);
			2968: out = 16'(14353);
			2969: out = 16'(-2394);
			2970: out = 16'(-19953);
			2971: out = 16'(-7804);
			2972: out = 16'(12689);
			2973: out = 16'(9462);
			2974: out = 16'(-7014);
			2975: out = 16'(-27652);
			2976: out = 16'(-6853);
			2977: out = 16'(21416);
			2978: out = 16'(18384);
			2979: out = 16'(-15670);
			2980: out = 16'(-18009);
			2981: out = 16'(9904);
			2982: out = 16'(25683);
			2983: out = 16'(6965);
			2984: out = 16'(-5844);
			2985: out = 16'(-5078);
			2986: out = 16'(5926);
			2987: out = 16'(5328);
			2988: out = 16'(5673);
			2989: out = 16'(-3823);
			2990: out = 16'(-7774);
			2991: out = 16'(-461);
			2992: out = 16'(-4618);
			2993: out = 16'(-18764);
			2994: out = 16'(-23025);
			2995: out = 16'(-764);
			2996: out = 16'(2708);
			2997: out = 16'(3735);
			2998: out = 16'(-1376);
			2999: out = 16'(-2425);
			3000: out = 16'(-6999);
			3001: out = 16'(-3321);
			3002: out = 16'(-2654);
			3003: out = 16'(1719);
			3004: out = 16'(9525);
			3005: out = 16'(10246);
			3006: out = 16'(-2774);
			3007: out = 16'(-15794);
			3008: out = 16'(-17515);
			3009: out = 16'(230);
			3010: out = 16'(4598);
			3011: out = 16'(673);
			3012: out = 16'(1724);
			3013: out = 16'(8614);
			3014: out = 16'(5574);
			3015: out = 16'(5055);
			3016: out = 16'(14070);
			3017: out = 16'(7483);
			3018: out = 16'(-3292);
			3019: out = 16'(-15388);
			3020: out = 16'(-17306);
			3021: out = 16'(-16547);
			3022: out = 16'(-1411);
			3023: out = 16'(13702);
			3024: out = 16'(24754);
			3025: out = 16'(29255);
			3026: out = 16'(19483);
			3027: out = 16'(6739);
			3028: out = 16'(-1169);
			3029: out = 16'(-131);
			3030: out = 16'(-11022);
			3031: out = 16'(-11123);
			3032: out = 16'(-4215);
			3033: out = 16'(2542);
			3034: out = 16'(11437);
			3035: out = 16'(18162);
			3036: out = 16'(19404);
			3037: out = 16'(12062);
			3038: out = 16'(620);
			3039: out = 16'(-4746);
			3040: out = 16'(-3057);
			3041: out = 16'(-1031);
			3042: out = 16'(1020);
			3043: out = 16'(9347);
			3044: out = 16'(13544);
			3045: out = 16'(12);
			3046: out = 16'(-25098);
			3047: out = 16'(-15871);
			3048: out = 16'(11679);
			3049: out = 16'(17523);
			3050: out = 16'(-1848);
			3051: out = 16'(-8044);
			3052: out = 16'(5331);
			3053: out = 16'(11448);
			3054: out = 16'(-8488);
			3055: out = 16'(-9757);
			3056: out = 16'(-20917);
			3057: out = 16'(-24391);
			3058: out = 16'(-21029);
			3059: out = 16'(-884);
			3060: out = 16'(5242);
			3061: out = 16'(9210);
			3062: out = 16'(8766);
			3063: out = 16'(3280);
			3064: out = 16'(-12795);
			3065: out = 16'(-25571);
			3066: out = 16'(-24190);
			3067: out = 16'(-4998);
			3068: out = 16'(12835);
			3069: out = 16'(16439);
			3070: out = 16'(4639);
			3071: out = 16'(-10041);
			3072: out = 16'(-4491);
			3073: out = 16'(2429);
			3074: out = 16'(3806);
			3075: out = 16'(4145);
			3076: out = 16'(14880);
			3077: out = 16'(6785);
			3078: out = 16'(-12329);
			3079: out = 16'(-25463);
			3080: out = 16'(-7349);
			3081: out = 16'(-555);
			3082: out = 16'(905);
			3083: out = 16'(4991);
			3084: out = 16'(19339);
			3085: out = 16'(16675);
			3086: out = 16'(8000);
			3087: out = 16'(-3390);
			3088: out = 16'(-6531);
			3089: out = 16'(-11309);
			3090: out = 16'(-3405);
			3091: out = 16'(6439);
			3092: out = 16'(13184);
			3093: out = 16'(6730);
			3094: out = 16'(5481);
			3095: out = 16'(-2342);
			3096: out = 16'(-12681);
			3097: out = 16'(-18120);
			3098: out = 16'(-4202);
			3099: out = 16'(9189);
			3100: out = 16'(12455);
			3101: out = 16'(6673);
			3102: out = 16'(7608);
			3103: out = 16'(-1612);
			3104: out = 16'(-15727);
			3105: out = 16'(-23807);
			3106: out = 16'(-12199);
			3107: out = 16'(-1031);
			3108: out = 16'(5361);
			3109: out = 16'(10374);
			3110: out = 16'(20641);
			3111: out = 16'(10869);
			3112: out = 16'(-832);
			3113: out = 16'(-2213);
			3114: out = 16'(2788);
			3115: out = 16'(1873);
			3116: out = 16'(-1825);
			3117: out = 16'(-437);
			3118: out = 16'(3227);
			3119: out = 16'(6413);
			3120: out = 16'(7326);
			3121: out = 16'(7313);
			3122: out = 16'(169);
			3123: out = 16'(-2192);
			3124: out = 16'(-9068);
			3125: out = 16'(-10431);
			3126: out = 16'(-6384);
			3127: out = 16'(10872);
			3128: out = 16'(15193);
			3129: out = 16'(17264);
			3130: out = 16'(10860);
			3131: out = 16'(-7743);
			3132: out = 16'(-20607);
			3133: out = 16'(-5705);
			3134: out = 16'(15956);
			3135: out = 16'(19110);
			3136: out = 16'(-1949);
			3137: out = 16'(-3274);
			3138: out = 16'(6797);
			3139: out = 16'(2022);
			3140: out = 16'(-17045);
			3141: out = 16'(-11195);
			3142: out = 16'(6369);
			3143: out = 16'(749);
			3144: out = 16'(-11471);
			3145: out = 16'(-8905);
			3146: out = 16'(5276);
			3147: out = 16'(6205);
			3148: out = 16'(1641);
			3149: out = 16'(-7827);
			3150: out = 16'(-13085);
			3151: out = 16'(-10491);
			3152: out = 16'(2028);
			3153: out = 16'(11932);
			3154: out = 16'(2659);
			3155: out = 16'(-15855);
			3156: out = 16'(-15928);
			3157: out = 16'(-12670);
			3158: out = 16'(-11814);
			3159: out = 16'(-11508);
			3160: out = 16'(4938);
			3161: out = 16'(21062);
			3162: out = 16'(16720);
			3163: out = 16'(-10240);
			3164: out = 16'(-28171);
			3165: out = 16'(-20748);
			3166: out = 16'(4274);
			3167: out = 16'(10704);
			3168: out = 16'(-176);
			3169: out = 16'(-1427);
			3170: out = 16'(-375);
			3171: out = 16'(3016);
			3172: out = 16'(874);
			3173: out = 16'(-10628);
			3174: out = 16'(-14917);
			3175: out = 16'(-10235);
			3176: out = 16'(2823);
			3177: out = 16'(12459);
			3178: out = 16'(20571);
			3179: out = 16'(14768);
			3180: out = 16'(6535);
			3181: out = 16'(443);
			3182: out = 16'(-1618);
			3183: out = 16'(-4490);
			3184: out = 16'(4383);
			3185: out = 16'(16865);
			3186: out = 16'(5899);
			3187: out = 16'(-8623);
			3188: out = 16'(-10608);
			3189: out = 16'(4585);
			3190: out = 16'(16029);
			3191: out = 16'(6496);
			3192: out = 16'(-3194);
			3193: out = 16'(-959);
			3194: out = 16'(6291);
			3195: out = 16'(-3076);
			3196: out = 16'(-5776);
			3197: out = 16'(5709);
			3198: out = 16'(15766);
			3199: out = 16'(4031);
			3200: out = 16'(-1996);
			3201: out = 16'(4038);
			3202: out = 16'(8590);
			3203: out = 16'(6464);
			3204: out = 16'(1063);
			3205: out = 16'(4582);
			3206: out = 16'(7203);
			3207: out = 16'(-5261);
			3208: out = 16'(-18779);
			3209: out = 16'(-9982);
			3210: out = 16'(16361);
			3211: out = 16'(22748);
			3212: out = 16'(12324);
			3213: out = 16'(-1323);
			3214: out = 16'(-3309);
			3215: out = 16'(-2247);
			3216: out = 16'(-15101);
			3217: out = 16'(-28922);
			3218: out = 16'(-19551);
			3219: out = 16'(9257);
			3220: out = 16'(22883);
			3221: out = 16'(14853);
			3222: out = 16'(4872);
			3223: out = 16'(2497);
			3224: out = 16'(-3375);
			3225: out = 16'(-5595);
			3226: out = 16'(3369);
			3227: out = 16'(16436);
			3228: out = 16'(5663);
			3229: out = 16'(1066);
			3230: out = 16'(-1804);
			3231: out = 16'(-4376);
			3232: out = 16'(-27780);
			3233: out = 16'(-8671);
			3234: out = 16'(4315);
			3235: out = 16'(-2147);
			3236: out = 16'(-19660);
			3237: out = 16'(-8572);
			3238: out = 16'(6810);
			3239: out = 16'(7895);
			3240: out = 16'(-6666);
			3241: out = 16'(-13009);
			3242: out = 16'(-9227);
			3243: out = 16'(553);
			3244: out = 16'(929);
			3245: out = 16'(-3088);
			3246: out = 16'(1075);
			3247: out = 16'(15315);
			3248: out = 16'(14156);
			3249: out = 16'(-13079);
			3250: out = 16'(-26099);
			3251: out = 16'(-9458);
			3252: out = 16'(9252);
			3253: out = 16'(-3051);
			3254: out = 16'(1935);
			3255: out = 16'(8870);
			3256: out = 16'(-1223);
			3257: out = 16'(-28521);
			3258: out = 16'(-29926);
			3259: out = 16'(-14983);
			3260: out = 16'(12599);
			3261: out = 16'(16552);
			3262: out = 16'(11893);
			3263: out = 16'(-20);
			3264: out = 16'(-5269);
			3265: out = 16'(-3047);
			3266: out = 16'(2210);
			3267: out = 16'(1667);
			3268: out = 16'(-6303);
			3269: out = 16'(-8907);
			3270: out = 16'(6346);
			3271: out = 16'(23851);
			3272: out = 16'(22893);
			3273: out = 16'(8953);
			3274: out = 16'(-2606);
			3275: out = 16'(-889);
			3276: out = 16'(5928);
			3277: out = 16'(10944);
			3278: out = 16'(6479);
			3279: out = 16'(4357);
			3280: out = 16'(-16456);
			3281: out = 16'(-26545);
			3282: out = 16'(-12647);
			3283: out = 16'(9960);
			3284: out = 16'(8460);
			3285: out = 16'(7404);
			3286: out = 16'(11412);
			3287: out = 16'(3610);
			3288: out = 16'(-8170);
			3289: out = 16'(-11162);
			3290: out = 16'(-3186);
			3291: out = 16'(-3912);
			3292: out = 16'(3210);
			3293: out = 16'(3060);
			3294: out = 16'(-3716);
			3295: out = 16'(-14831);
			3296: out = 16'(4485);
			3297: out = 16'(22958);
			3298: out = 16'(21057);
			3299: out = 16'(-4026);
			3300: out = 16'(-13215);
			3301: out = 16'(-15053);
			3302: out = 16'(47);
			3303: out = 16'(9149);
			3304: out = 16'(18236);
			3305: out = 16'(804);
			3306: out = 16'(-2613);
			3307: out = 16'(-1841);
			3308: out = 16'(-6215);
			3309: out = 16'(-18249);
			3310: out = 16'(-920);
			3311: out = 16'(20223);
			3312: out = 16'(11837);
			3313: out = 16'(-1423);
			3314: out = 16'(-4496);
			3315: out = 16'(1540);
			3316: out = 16'(-2074);
			3317: out = 16'(-19414);
			3318: out = 16'(-11379);
			3319: out = 16'(11533);
			3320: out = 16'(17317);
			3321: out = 16'(5605);
			3322: out = 16'(-9953);
			3323: out = 16'(-13523);
			3324: out = 16'(-2532);
			3325: out = 16'(13116);
			3326: out = 16'(6467);
			3327: out = 16'(-8127);
			3328: out = 16'(-15896);
			3329: out = 16'(-6811);
			3330: out = 16'(-6675);
			3331: out = 16'(-4730);
			3332: out = 16'(5257);
			3333: out = 16'(17806);
			3334: out = 16'(-1183);
			3335: out = 16'(-14063);
			3336: out = 16'(-6317);
			3337: out = 16'(21294);
			3338: out = 16'(20145);
			3339: out = 16'(17146);
			3340: out = 16'(-65);
			3341: out = 16'(-15596);
			3342: out = 16'(-29614);
			3343: out = 16'(-16148);
			3344: out = 16'(-8583);
			3345: out = 16'(-2283);
			3346: out = 16'(12203);
			3347: out = 16'(26765);
			3348: out = 16'(17562);
			3349: out = 16'(2472);
			3350: out = 16'(-3844);
			3351: out = 16'(-4370);
			3352: out = 16'(-16891);
			3353: out = 16'(-21331);
			3354: out = 16'(-1862);
			3355: out = 16'(5855);
			3356: out = 16'(4025);
			3357: out = 16'(1977);
			3358: out = 16'(12263);
			3359: out = 16'(19517);
			3360: out = 16'(12335);
			3361: out = 16'(-402);
			3362: out = 16'(-5872);
			3363: out = 16'(-9719);
			3364: out = 16'(-3092);
			3365: out = 16'(-2620);
			3366: out = 16'(-2953);
			3367: out = 16'(117);
			3368: out = 16'(-65);
			3369: out = 16'(5789);
			3370: out = 16'(14922);
			3371: out = 16'(15091);
			3372: out = 16'(-4628);
			3373: out = 16'(-18833);
			3374: out = 16'(-14204);
			3375: out = 16'(1062);
			3376: out = 16'(436);
			3377: out = 16'(2140);
			3378: out = 16'(7418);
			3379: out = 16'(10467);
			3380: out = 16'(6822);
			3381: out = 16'(-13535);
			3382: out = 16'(-17144);
			3383: out = 16'(1801);
			3384: out = 16'(13412);
			3385: out = 16'(3485);
			3386: out = 16'(-9327);
			3387: out = 16'(-5025);
			3388: out = 16'(9567);
			3389: out = 16'(6493);
			3390: out = 16'(1139);
			3391: out = 16'(256);
			3392: out = 16'(-2304);
			3393: out = 16'(-13292);
			3394: out = 16'(-24174);
			3395: out = 16'(-10636);
			3396: out = 16'(19526);
			3397: out = 16'(24450);
			3398: out = 16'(16930);
			3399: out = 16'(1034);
			3400: out = 16'(-12558);
			3401: out = 16'(-25901);
			3402: out = 16'(-7416);
			3403: out = 16'(7332);
			3404: out = 16'(5726);
			3405: out = 16'(-870);
			3406: out = 16'(-7131);
			3407: out = 16'(3684);
			3408: out = 16'(13084);
			3409: out = 16'(9956);
			3410: out = 16'(1227);
			3411: out = 16'(-233);
			3412: out = 16'(-2607);
			3413: out = 16'(-8885);
			3414: out = 16'(-216);
			3415: out = 16'(1816);
			3416: out = 16'(-612);
			3417: out = 16'(-6425);
			3418: out = 16'(-8312);
			3419: out = 16'(-2380);
			3420: out = 16'(6167);
			3421: out = 16'(13590);
			3422: out = 16'(15218);
			3423: out = 16'(4642);
			3424: out = 16'(-16965);
			3425: out = 16'(-25332);
			3426: out = 16'(-1011);
			3427: out = 16'(10084);
			3428: out = 16'(8611);
			3429: out = 16'(-3402);
			3430: out = 16'(-7099);
			3431: out = 16'(-5194);
			3432: out = 16'(13808);
			3433: out = 16'(22402);
			3434: out = 16'(17015);
			3435: out = 16'(157);
			3436: out = 16'(-13067);
			3437: out = 16'(-24090);
			3438: out = 16'(-19744);
			3439: out = 16'(1059);
			3440: out = 16'(18866);
			3441: out = 16'(8965);
			3442: out = 16'(-10611);
			3443: out = 16'(-14309);
			3444: out = 16'(3137);
			3445: out = 16'(16074);
			3446: out = 16'(17494);
			3447: out = 16'(14816);
			3448: out = 16'(-1849);
			3449: out = 16'(-7621);
			3450: out = 16'(-5167);
			3451: out = 16'(-1100);
			3452: out = 16'(-6755);
			3453: out = 16'(-1442);
			3454: out = 16'(12997);
			3455: out = 16'(19572);
			3456: out = 16'(-389);
			3457: out = 16'(-1227);
			3458: out = 16'(-332);
			3459: out = 16'(-5736);
			3460: out = 16'(-24467);
			3461: out = 16'(-11282);
			3462: out = 16'(12890);
			3463: out = 16'(24798);
			3464: out = 16'(10502);
			3465: out = 16'(-12046);
			3466: out = 16'(-28812);
			3467: out = 16'(-18641);
			3468: out = 16'(3865);
			3469: out = 16'(10937);
			3470: out = 16'(9033);
			3471: out = 16'(7501);
			3472: out = 16'(799);
			3473: out = 16'(-18338);
			3474: out = 16'(-30418);
			3475: out = 16'(-14400);
			3476: out = 16'(13289);
			3477: out = 16'(9494);
			3478: out = 16'(-2239);
			3479: out = 16'(-13537);
			3480: out = 16'(-5645);
			3481: out = 16'(8932);
			3482: out = 16'(20677);
			3483: out = 16'(10495);
			3484: out = 16'(-2932);
			3485: out = 16'(-12663);
			3486: out = 16'(-27682);
			3487: out = 16'(-25071);
			3488: out = 16'(-5582);
			3489: out = 16'(14763);
			3490: out = 16'(15720);
			3491: out = 16'(13798);
			3492: out = 16'(10027);
			3493: out = 16'(7777);
			3494: out = 16'(1482);
			3495: out = 16'(-4225);
			3496: out = 16'(-9139);
			3497: out = 16'(-5362);
			3498: out = 16'(3767);
			3499: out = 16'(6096);
			3500: out = 16'(-1833);
			3501: out = 16'(-11392);
			3502: out = 16'(-12591);
			3503: out = 16'(-1464);
			3504: out = 16'(9375);
			3505: out = 16'(14613);
			3506: out = 16'(13269);
			3507: out = 16'(9277);
			3508: out = 16'(2106);
			3509: out = 16'(376);
			3510: out = 16'(-1707);
			3511: out = 16'(-25120);
			3512: out = 16'(-13069);
			3513: out = 16'(9673);
			3514: out = 16'(20731);
			3515: out = 16'(10445);
			3516: out = 16'(11694);
			3517: out = 16'(7588);
			3518: out = 16'(3099);
			3519: out = 16'(-881);
			3520: out = 16'(-3590);
			3521: out = 16'(-2056);
			3522: out = 16'(57);
			3523: out = 16'(-3307);
			3524: out = 16'(-6334);
			3525: out = 16'(2945);
			3526: out = 16'(17334);
			3527: out = 16'(14937);
			3528: out = 16'(7158);
			3529: out = 16'(-20663);
			3530: out = 16'(-18878);
			3531: out = 16'(5433);
			3532: out = 16'(15300);
			3533: out = 16'(3495);
			3534: out = 16'(-1802);
			3535: out = 16'(-7530);
			3536: out = 16'(-26833);
			3537: out = 16'(-30511);
			3538: out = 16'(-6027);
			3539: out = 16'(26126);
			3540: out = 16'(26803);
			3541: out = 16'(12235);
			3542: out = 16'(-7832);
			3543: out = 16'(-16395);
			3544: out = 16'(-12746);
			3545: out = 16'(58);
			3546: out = 16'(10031);
			3547: out = 16'(10438);
			3548: out = 16'(2762);
			3549: out = 16'(-1599);
			3550: out = 16'(-19904);
			3551: out = 16'(-30471);
			3552: out = 16'(-20501);
			3553: out = 16'(5817);
			3554: out = 16'(16619);
			3555: out = 16'(10685);
			3556: out = 16'(2362);
			3557: out = 16'(2321);
			3558: out = 16'(-3700);
			3559: out = 16'(-10933);
			3560: out = 16'(-9165);
			3561: out = 16'(8822);
			3562: out = 16'(11086);
			3563: out = 16'(10272);
			3564: out = 16'(-2900);
			3565: out = 16'(-11171);
			3566: out = 16'(-6112);
			3567: out = 16'(3205);
			3568: out = 16'(-529);
			3569: out = 16'(-6824);
			3570: out = 16'(-7066);
			3571: out = 16'(-6216);
			3572: out = 16'(-18356);
			3573: out = 16'(-22421);
			3574: out = 16'(3929);
			3575: out = 16'(23763);
			3576: out = 16'(23158);
			3577: out = 16'(7969);
			3578: out = 16'(-7183);
			3579: out = 16'(-10912);
			3580: out = 16'(-11780);
			3581: out = 16'(-1659);
			3582: out = 16'(14793);
			3583: out = 16'(19249);
			3584: out = 16'(2785);
			3585: out = 16'(-13956);
			3586: out = 16'(-15881);
			3587: out = 16'(-8558);
			3588: out = 16'(5594);
			3589: out = 16'(12705);
			3590: out = 16'(11665);
			3591: out = 16'(5665);
			3592: out = 16'(-1504);
			3593: out = 16'(-3448);
			3594: out = 16'(-2177);
			3595: out = 16'(794);
			3596: out = 16'(-4785);
			3597: out = 16'(10320);
			3598: out = 16'(23456);
			3599: out = 16'(18472);
			3600: out = 16'(3825);
			3601: out = 16'(-12611);
			3602: out = 16'(-19842);
			3603: out = 16'(-12550);
			3604: out = 16'(2527);
			3605: out = 16'(14159);
			3606: out = 16'(10608);
			3607: out = 16'(2146);
			3608: out = 16'(2635);
			3609: out = 16'(10159);
			3610: out = 16'(11765);
			3611: out = 16'(7083);
			3612: out = 16'(1839);
			3613: out = 16'(-14989);
			3614: out = 16'(-25720);
			3615: out = 16'(-21605);
			3616: out = 16'(-2212);
			3617: out = 16'(10819);
			3618: out = 16'(17564);
			3619: out = 16'(13928);
			3620: out = 16'(582);
			3621: out = 16'(-15816);
			3622: out = 16'(-27449);
			3623: out = 16'(-15307);
			3624: out = 16'(10010);
			3625: out = 16'(17042);
			3626: out = 16'(13028);
			3627: out = 16'(5598);
			3628: out = 16'(3234);
			3629: out = 16'(-807);
			3630: out = 16'(-7719);
			3631: out = 16'(-15399);
			3632: out = 16'(-11492);
			3633: out = 16'(561);
			3634: out = 16'(-3702);
			3635: out = 16'(-6293);
			3636: out = 16'(-3287);
			3637: out = 16'(2820);
			3638: out = 16'(1266);
			3639: out = 16'(-2452);
			3640: out = 16'(-4935);
			3641: out = 16'(-3575);
			3642: out = 16'(-992);
			3643: out = 16'(-4584);
			3644: out = 16'(-952);
			3645: out = 16'(12668);
			3646: out = 16'(18083);
			3647: out = 16'(13215);
			3648: out = 16'(-8451);
			3649: out = 16'(-19501);
			3650: out = 16'(650);
			3651: out = 16'(2927);
			3652: out = 16'(3457);
			3653: out = 16'(-90);
			3654: out = 16'(1287);
			3655: out = 16'(-9805);
			3656: out = 16'(4049);
			3657: out = 16'(16227);
			3658: out = 16'(13939);
			3659: out = 16'(-5059);
			3660: out = 16'(-4047);
			3661: out = 16'(1390);
			3662: out = 16'(-211);
			3663: out = 16'(-12984);
			3664: out = 16'(148);
			3665: out = 16'(11730);
			3666: out = 16'(7578);
			3667: out = 16'(-12114);
			3668: out = 16'(-14189);
			3669: out = 16'(-184);
			3670: out = 16'(19784);
			3671: out = 16'(18208);
			3672: out = 16'(5601);
			3673: out = 16'(-13100);
			3674: out = 16'(-348);
			3675: out = 16'(23339);
			3676: out = 16'(11250);
			3677: out = 16'(-15535);
			3678: out = 16'(-21927);
			3679: out = 16'(-1835);
			3680: out = 16'(-938);
			3681: out = 16'(586);
			3682: out = 16'(7757);
			3683: out = 16'(18168);
			3684: out = 16'(13659);
			3685: out = 16'(-1964);
			3686: out = 16'(-11115);
			3687: out = 16'(-10177);
			3688: out = 16'(-8410);
			3689: out = 16'(-1957);
			3690: out = 16'(9350);
			3691: out = 16'(11268);
			3692: out = 16'(1171);
			3693: out = 16'(4619);
			3694: out = 16'(8412);
			3695: out = 16'(4431);
			3696: out = 16'(-7269);
			3697: out = 16'(-9032);
			3698: out = 16'(-4154);
			3699: out = 16'(-5626);
			3700: out = 16'(-12994);
			3701: out = 16'(-6429);
			3702: out = 16'(2373);
			3703: out = 16'(4237);
			3704: out = 16'(233);
			3705: out = 16'(6050);
			3706: out = 16'(666);
			3707: out = 16'(-2261);
			3708: out = 16'(-7271);
			3709: out = 16'(-7755);
			3710: out = 16'(-1418);
			3711: out = 16'(6256);
			3712: out = 16'(7810);
			3713: out = 16'(4232);
			3714: out = 16'(547);
			3715: out = 16'(-12184);
			3716: out = 16'(-18457);
			3717: out = 16'(-4601);
			3718: out = 16'(13213);
			3719: out = 16'(13168);
			3720: out = 16'(-3317);
			3721: out = 16'(-8140);
			3722: out = 16'(10551);
			3723: out = 16'(12167);
			3724: out = 16'(-7967);
			3725: out = 16'(-25539);
			3726: out = 16'(-12232);
			3727: out = 16'(-2412);
			3728: out = 16'(1991);
			3729: out = 16'(2701);
			3730: out = 16'(9560);
			3731: out = 16'(2417);
			3732: out = 16'(4437);
			3733: out = 16'(8364);
			3734: out = 16'(12484);
			3735: out = 16'(4896);
			3736: out = 16'(-4003);
			3737: out = 16'(-15328);
			3738: out = 16'(-20607);
			3739: out = 16'(-19808);
			3740: out = 16'(1932);
			3741: out = 16'(19937);
			3742: out = 16'(23804);
			3743: out = 16'(11932);
			3744: out = 16'(-3787);
			3745: out = 16'(-16938);
			3746: out = 16'(-12933);
			3747: out = 16'(353);
			3748: out = 16'(-4952);
			3749: out = 16'(-13626);
			3750: out = 16'(-9141);
			3751: out = 16'(8385);
			3752: out = 16'(8153);
			3753: out = 16'(7442);
			3754: out = 16'(6253);
			3755: out = 16'(8812);
			3756: out = 16'(1618);
			3757: out = 16'(5444);
			3758: out = 16'(3694);
			3759: out = 16'(356);
			3760: out = 16'(-9291);
			3761: out = 16'(-697);
			3762: out = 16'(-3657);
			3763: out = 16'(-5489);
			3764: out = 16'(1800);
			3765: out = 16'(17710);
			3766: out = 16'(14319);
			3767: out = 16'(8130);
			3768: out = 16'(11216);
			3769: out = 16'(20746);
			3770: out = 16'(4850);
			3771: out = 16'(-18194);
			3772: out = 16'(-27578);
			3773: out = 16'(-16324);
			3774: out = 16'(-2414);
			3775: out = 16'(8390);
			3776: out = 16'(14522);
			3777: out = 16'(11307);
			3778: out = 16'(1448);
			3779: out = 16'(-6657);
			3780: out = 16'(-6003);
			3781: out = 16'(-2246);
			3782: out = 16'(4414);
			3783: out = 16'(-601);
			3784: out = 16'(-10307);
			3785: out = 16'(-18186);
			3786: out = 16'(-6459);
			3787: out = 16'(-1854);
			3788: out = 16'(4935);
			3789: out = 16'(11461);
			3790: out = 16'(5225);
			3791: out = 16'(-5382);
			3792: out = 16'(-15727);
			3793: out = 16'(-15779);
			3794: out = 16'(-3302);
			3795: out = 16'(4120);
			3796: out = 16'(6678);
			3797: out = 16'(3582);
			3798: out = 16'(-3175);
			3799: out = 16'(-10687);
			3800: out = 16'(-8461);
			3801: out = 16'(-4339);
			3802: out = 16'(-7889);
			3803: out = 16'(5214);
			3804: out = 16'(7423);
			3805: out = 16'(6384);
			3806: out = 16'(2888);
			3807: out = 16'(17619);
			3808: out = 16'(-6918);
			3809: out = 16'(-29075);
			3810: out = 16'(-26753);
			3811: out = 16'(2872);
			3812: out = 16'(21216);
			3813: out = 16'(12591);
			3814: out = 16'(-2836);
			3815: out = 16'(-6252);
			3816: out = 16'(-815);
			3817: out = 16'(12362);
			3818: out = 16'(17409);
			3819: out = 16'(13526);
			3820: out = 16'(-938);
			3821: out = 16'(-4402);
			3822: out = 16'(-7794);
			3823: out = 16'(-13179);
			3824: out = 16'(-5995);
			3825: out = 16'(13419);
			3826: out = 16'(21513);
			3827: out = 16'(12543);
			3828: out = 16'(6556);
			3829: out = 16'(7498);
			3830: out = 16'(7025);
			3831: out = 16'(-4109);
			3832: out = 16'(-9233);
			3833: out = 16'(-17373);
			3834: out = 16'(-3990);
			3835: out = 16'(13333);
			3836: out = 16'(19038);
			3837: out = 16'(-6713);
			3838: out = 16'(-10848);
			3839: out = 16'(4573);
			3840: out = 16'(14767);
			3841: out = 16'(-3929);
			3842: out = 16'(-5411);
			3843: out = 16'(7238);
			3844: out = 16'(11959);
			3845: out = 16'(-10000);
			3846: out = 16'(-18856);
			3847: out = 16'(-10651);
			3848: out = 16'(5915);
			3849: out = 16'(15719);
			3850: out = 16'(7397);
			3851: out = 16'(-2109);
			3852: out = 16'(-4444);
			3853: out = 16'(1913);
			3854: out = 16'(-92);
			3855: out = 16'(653);
			3856: out = 16'(2979);
			3857: out = 16'(5568);
			3858: out = 16'(-13459);
			3859: out = 16'(-12176);
			3860: out = 16'(2838);
			3861: out = 16'(15891);
			3862: out = 16'(13253);
			3863: out = 16'(8445);
			3864: out = 16'(-1271);
			3865: out = 16'(-7694);
			3866: out = 16'(-8216);
			3867: out = 16'(5348);
			3868: out = 16'(8111);
			3869: out = 16'(3716);
			3870: out = 16'(2569);
			3871: out = 16'(947);
			3872: out = 16'(-10426);
			3873: out = 16'(-17260);
			3874: out = 16'(-3000);
			3875: out = 16'(-996);
			3876: out = 16'(-2139);
			3877: out = 16'(-1616);
			3878: out = 16'(5637);
			3879: out = 16'(5001);
			3880: out = 16'(-3653);
			3881: out = 16'(-8081);
			3882: out = 16'(1804);
			3883: out = 16'(313);
			3884: out = 16'(-5866);
			3885: out = 16'(-21902);
			3886: out = 16'(-24964);
			3887: out = 16'(-2812);
			3888: out = 16'(17742);
			3889: out = 16'(17040);
			3890: out = 16'(6143);
			3891: out = 16'(-3245);
			3892: out = 16'(-7658);
			3893: out = 16'(-9660);
			3894: out = 16'(-4957);
			3895: out = 16'(4398);
			3896: out = 16'(8644);
			3897: out = 16'(2360);
			3898: out = 16'(-243);
			3899: out = 16'(5642);
			3900: out = 16'(-1314);
			3901: out = 16'(-3328);
			3902: out = 16'(1352);
			3903: out = 16'(10822);
			3904: out = 16'(4288);
			3905: out = 16'(3730);
			3906: out = 16'(-2813);
			3907: out = 16'(-7462);
			3908: out = 16'(-6840);
			3909: out = 16'(3888);
			3910: out = 16'(8094);
			3911: out = 16'(3195);
			3912: out = 16'(-7091);
			3913: out = 16'(-2738);
			3914: out = 16'(-209);
			3915: out = 16'(349);
			3916: out = 16'(708);
			3917: out = 16'(10316);
			3918: out = 16'(5836);
			3919: out = 16'(-1573);
			3920: out = 16'(-1553);
			3921: out = 16'(12492);
			3922: out = 16'(9261);
			3923: out = 16'(2197);
			3924: out = 16'(1258);
			3925: out = 16'(8497);
			3926: out = 16'(6127);
			3927: out = 16'(-2764);
			3928: out = 16'(-10468);
			3929: out = 16'(-5183);
			3930: out = 16'(-5319);
			3931: out = 16'(-414);
			3932: out = 16'(1307);
			3933: out = 16'(2285);
			3934: out = 16'(6101);
			3935: out = 16'(9241);
			3936: out = 16'(-1407);
			3937: out = 16'(-20154);
			3938: out = 16'(-15312);
			3939: out = 16'(-6828);
			3940: out = 16'(4990);
			3941: out = 16'(16640);
			3942: out = 16'(21585);
			3943: out = 16'(13526);
			3944: out = 16'(-9854);
			3945: out = 16'(-25943);
			3946: out = 16'(-7208);
			3947: out = 16'(9803);
			3948: out = 16'(4985);
			3949: out = 16'(-14467);
			3950: out = 16'(-20882);
			3951: out = 16'(-17889);
			3952: out = 16'(-1797);
			3953: out = 16'(11231);
			3954: out = 16'(21725);
			3955: out = 16'(16771);
			3956: out = 16'(7808);
			3957: out = 16'(-11621);
			3958: out = 16'(-20564);
			3959: out = 16'(-10204);
			3960: out = 16'(9979);
			3961: out = 16'(1460);
			3962: out = 16'(-14347);
			3963: out = 16'(-1243);
			3964: out = 16'(17742);
			3965: out = 16'(12903);
			3966: out = 16'(-6012);
			3967: out = 16'(-10565);
			3968: out = 16'(6378);
			3969: out = 16'(5162);
			3970: out = 16'(-13954);
			3971: out = 16'(-21146);
			3972: out = 16'(1179);
			3973: out = 16'(12914);
			3974: out = 16'(-1807);
			3975: out = 16'(-22033);
			3976: out = 16'(-11756);
			3977: out = 16'(1556);
			3978: out = 16'(5428);
			3979: out = 16'(-933);
			3980: out = 16'(-3376);
			3981: out = 16'(-3319);
			3982: out = 16'(8471);
			3983: out = 16'(18503);
			3984: out = 16'(14336);
			3985: out = 16'(3743);
			3986: out = 16'(-6718);
			3987: out = 16'(-13222);
			3988: out = 16'(-20258);
			3989: out = 16'(-11530);
			3990: out = 16'(-3820);
			3991: out = 16'(5887);
			3992: out = 16'(9209);
			3993: out = 16'(2706);
			3994: out = 16'(-8093);
			3995: out = 16'(-1728);
			3996: out = 16'(15956);
			3997: out = 16'(15936);
			3998: out = 16'(1420);
			3999: out = 16'(-13883);
			4000: out = 16'(-10928);
			4001: out = 16'(7880);
			4002: out = 16'(4614);
			4003: out = 16'(479);
			4004: out = 16'(7924);
			4005: out = 16'(20185);
			4006: out = 16'(14289);
			4007: out = 16'(859);
			4008: out = 16'(-11151);
			4009: out = 16'(-13958);
			4010: out = 16'(-10092);
			4011: out = 16'(212);
			4012: out = 16'(9108);
			4013: out = 16'(9535);
			4014: out = 16'(-529);
			4015: out = 16'(-4092);
			4016: out = 16'(334);
			4017: out = 16'(6302);
			4018: out = 16'(9709);
			4019: out = 16'(12262);
			4020: out = 16'(12182);
			4021: out = 16'(131);
			4022: out = 16'(-22116);
			4023: out = 16'(-26746);
			4024: out = 16'(-8751);
			4025: out = 16'(10415);
			4026: out = 16'(12851);
			4027: out = 16'(3297);
			4028: out = 16'(8473);
			4029: out = 16'(12635);
			4030: out = 16'(1830);
			4031: out = 16'(-2095);
			4032: out = 16'(-8098);
			4033: out = 16'(-3886);
			4034: out = 16'(2465);
			4035: out = 16'(9268);
			4036: out = 16'(2019);
			4037: out = 16'(-2973);
			4038: out = 16'(-3547);
			4039: out = 16'(-136);
			4040: out = 16'(-297);
			4041: out = 16'(-2576);
			4042: out = 16'(-6757);
			4043: out = 16'(-4405);
			4044: out = 16'(-2290);
			4045: out = 16'(2738);
			4046: out = 16'(-4343);
			4047: out = 16'(-15528);
			4048: out = 16'(-10718);
			4049: out = 16'(7627);
			4050: out = 16'(10069);
			4051: out = 16'(-5109);
			4052: out = 16'(-14411);
			4053: out = 16'(-5390);
			4054: out = 16'(3969);
			4055: out = 16'(4698);
			4056: out = 16'(14446);
			4057: out = 16'(4185);
			4058: out = 16'(-1781);
			4059: out = 16'(-6698);
			4060: out = 16'(-8601);
			4061: out = 16'(-13226);
			4062: out = 16'(-14272);
			4063: out = 16'(-11362);
			4064: out = 16'(-2903);
			4065: out = 16'(4572);
			4066: out = 16'(9520);
			4067: out = 16'(10389);
			4068: out = 16'(9266);
			4069: out = 16'(693);
			4070: out = 16'(557);
			4071: out = 16'(421);
			4072: out = 16'(664);
			4073: out = 16'(1768);
			4074: out = 16'(-9948);
			4075: out = 16'(-19601);
			4076: out = 16'(-8266);
			4077: out = 16'(20523);
			4078: out = 16'(22187);
			4079: out = 16'(5092);
			4080: out = 16'(-10224);
			4081: out = 16'(-672);
			4082: out = 16'(5552);
			4083: out = 16'(11044);
			4084: out = 16'(6943);
			4085: out = 16'(6332);
			4086: out = 16'(7722);
			4087: out = 16'(8320);
			4088: out = 16'(-3560);
			4089: out = 16'(-9207);
			4090: out = 16'(9862);
			4091: out = 16'(20751);
			4092: out = 16'(8886);
			4093: out = 16'(-8008);
			4094: out = 16'(-5466);
			4095: out = 16'(2220);
			4096: out = 16'(2182);
			4097: out = 16'(1354);
			4098: out = 16'(9526);
			4099: out = 16'(-3831);
			4100: out = 16'(-18223);
			4101: out = 16'(-15052);
			4102: out = 16'(11288);
			4103: out = 16'(13375);
			4104: out = 16'(6599);
			4105: out = 16'(680);
			4106: out = 16'(5907);
			4107: out = 16'(-6457);
			4108: out = 16'(-6913);
			4109: out = 16'(-8593);
			4110: out = 16'(-7513);
			4111: out = 16'(-11719);
			4112: out = 16'(-9187);
			4113: out = 16'(-6789);
			4114: out = 16'(2172);
			4115: out = 16'(10159);
			4116: out = 16'(19529);
			4117: out = 16'(9978);
			4118: out = 16'(-4018);
			4119: out = 16'(-12166);
			4120: out = 16'(3586);
			4121: out = 16'(-3054);
			4122: out = 16'(-19521);
			4123: out = 16'(-25687);
			4124: out = 16'(-9714);
			4125: out = 16'(1347);
			4126: out = 16'(6693);
			4127: out = 16'(9202);
			4128: out = 16'(571);
			4129: out = 16'(-3788);
			4130: out = 16'(-1141);
			4131: out = 16'(5903);
			4132: out = 16'(-2542);
			4133: out = 16'(3750);
			4134: out = 16'(-2770);
			4135: out = 16'(-14441);
			4136: out = 16'(-24682);
			4137: out = 16'(-2948);
			4138: out = 16'(7531);
			4139: out = 16'(5639);
			4140: out = 16'(3353);
			4141: out = 16'(9026);
			4142: out = 16'(8220);
			4143: out = 16'(1321);
			4144: out = 16'(-4348);
			4145: out = 16'(1763);
			4146: out = 16'(1413);
			4147: out = 16'(-1360);
			4148: out = 16'(-3370);
			4149: out = 16'(-4642);
			4150: out = 16'(-4727);
			4151: out = 16'(-1199);
			4152: out = 16'(8307);
			4153: out = 16'(18792);
			4154: out = 16'(18406);
			4155: out = 16'(9409);
			4156: out = 16'(-6921);
			4157: out = 16'(-26731);
			4158: out = 16'(-6647);
			4159: out = 16'(2241);
			4160: out = 16'(-1554);
			4161: out = 16'(-4681);
			4162: out = 16'(15642);
			4163: out = 16'(18838);
			4164: out = 16'(12368);
			4165: out = 16'(2458);
			4166: out = 16'(-3201);
			4167: out = 16'(-2664);
			4168: out = 16'(1166);
			4169: out = 16'(167);
			4170: out = 16'(-76);
			4171: out = 16'(-12519);
			4172: out = 16'(-11720);
			4173: out = 16'(-6817);
			4174: out = 16'(-6039);
			4175: out = 16'(5870);
			4176: out = 16'(21348);
			4177: out = 16'(23161);
			4178: out = 16'(9792);
			4179: out = 16'(-16838);
			4180: out = 16'(-14274);
			4181: out = 16'(-21);
			4182: out = 16'(4477);
			4183: out = 16'(6141);
			4184: out = 16'(11076);
			4185: out = 16'(8620);
			4186: out = 16'(-6073);
			4187: out = 16'(-20888);
			4188: out = 16'(-11432);
			4189: out = 16'(10519);
			4190: out = 16'(21531);
			4191: out = 16'(14882);
			4192: out = 16'(-1943);
			4193: out = 16'(-20661);
			4194: out = 16'(-23201);
			4195: out = 16'(-4254);
			4196: out = 16'(3467);
			4197: out = 16'(-1218);
			4198: out = 16'(-10820);
			4199: out = 16'(-9471);
			4200: out = 16'(8672);
			4201: out = 16'(11564);
			4202: out = 16'(5866);
			4203: out = 16'(4124);
			4204: out = 16'(6723);
			4205: out = 16'(6532);
			4206: out = 16'(-5225);
			4207: out = 16'(-18703);
			4208: out = 16'(-15708);
			4209: out = 16'(-8541);
			4210: out = 16'(-2753);
			4211: out = 16'(-4381);
			4212: out = 16'(-897);
			4213: out = 16'(12369);
			4214: out = 16'(22726);
			4215: out = 16'(9505);
			4216: out = 16'(-19158);
			4217: out = 16'(-29703);
			4218: out = 16'(-17077);
			4219: out = 16'(-1493);
			4220: out = 16'(1098);
			4221: out = 16'(4089);
			4222: out = 16'(5950);
			4223: out = 16'(-662);
			4224: out = 16'(-11294);
			4225: out = 16'(-7013);
			4226: out = 16'(7779);
			4227: out = 16'(16268);
			4228: out = 16'(9385);
			4229: out = 16'(-3184);
			4230: out = 16'(-10899);
			4231: out = 16'(-8014);
			4232: out = 16'(979);
			4233: out = 16'(4968);
			4234: out = 16'(5439);
			4235: out = 16'(-9843);
			4236: out = 16'(-13504);
			4237: out = 16'(8420);
			4238: out = 16'(23184);
			4239: out = 16'(15832);
			4240: out = 16'(-9151);
			4241: out = 16'(-24704);
			4242: out = 16'(-11236);
			4243: out = 16'(7627);
			4244: out = 16'(9486);
			4245: out = 16'(1690);
			4246: out = 16'(-2346);
			4247: out = 16'(3988);
			4248: out = 16'(3722);
			4249: out = 16'(-336);
			4250: out = 16'(1495);
			4251: out = 16'(8244);
			4252: out = 16'(10980);
			4253: out = 16'(4727);
			4254: out = 16'(-5593);
			4255: out = 16'(1966);
			4256: out = 16'(-4915);
			4257: out = 16'(-10294);
			4258: out = 16'(-9322);
			4259: out = 16'(-3050);
			4260: out = 16'(3835);
			4261: out = 16'(13465);
			4262: out = 16'(15808);
			4263: out = 16'(4769);
			4264: out = 16'(-8739);
			4265: out = 16'(-9460);
			4266: out = 16'(-393);
			4267: out = 16'(1202);
			4268: out = 16'(-3295);
			4269: out = 16'(-3130);
			4270: out = 16'(1750);
			4271: out = 16'(-351);
			4272: out = 16'(3130);
			4273: out = 16'(-163);
			4274: out = 16'(5770);
			4275: out = 16'(14990);
			4276: out = 16'(19631);
			4277: out = 16'(5715);
			4278: out = 16'(-4861);
			4279: out = 16'(-2654);
			4280: out = 16'(11381);
			4281: out = 16'(7171);
			4282: out = 16'(5629);
			4283: out = 16'(3346);
			4284: out = 16'(-6495);
			4285: out = 16'(-10676);
			4286: out = 16'(-7175);
			4287: out = 16'(-1522);
			4288: out = 16'(-4034);
			4289: out = 16'(8343);
			4290: out = 16'(3793);
			4291: out = 16'(-2613);
			4292: out = 16'(-2136);
			4293: out = 16'(10237);
			4294: out = 16'(5011);
			4295: out = 16'(-8479);
			4296: out = 16'(-14386);
			4297: out = 16'(2018);
			4298: out = 16'(11492);
			4299: out = 16'(5982);
			4300: out = 16'(-12495);
			4301: out = 16'(-26797);
			4302: out = 16'(-25801);
			4303: out = 16'(-10990);
			4304: out = 16'(2236);
			4305: out = 16'(6987);
			4306: out = 16'(2876);
			4307: out = 16'(1778);
			4308: out = 16'(1584);
			4309: out = 16'(-209);
			4310: out = 16'(-4229);
			4311: out = 16'(-1722);
			4312: out = 16'(3218);
			4313: out = 16'(4925);
			4314: out = 16'(614);
			4315: out = 16'(-1235);
			4316: out = 16'(-754);
			4317: out = 16'(-494);
			4318: out = 16'(-6578);
			4319: out = 16'(2917);
			4320: out = 16'(4114);
			4321: out = 16'(-1877);
			4322: out = 16'(-3918);
			4323: out = 16'(202);
			4324: out = 16'(4760);
			4325: out = 16'(6249);
			4326: out = 16'(11447);
			4327: out = 16'(19331);
			4328: out = 16'(14175);
			4329: out = 16'(-5608);
			4330: out = 16'(-21848);
			4331: out = 16'(-18446);
			4332: out = 16'(2870);
			4333: out = 16'(7125);
			4334: out = 16'(-5058);
			4335: out = 16'(-16589);
			4336: out = 16'(3059);
			4337: out = 16'(13795);
			4338: out = 16'(5846);
			4339: out = 16'(-28);
			4340: out = 16'(10592);
			4341: out = 16'(18478);
			4342: out = 16'(11736);
			4343: out = 16'(-1058);
			4344: out = 16'(-2807);
			4345: out = 16'(1279);
			4346: out = 16'(5501);
			4347: out = 16'(4493);
			4348: out = 16'(221);
			4349: out = 16'(-7708);
			4350: out = 16'(-6330);
			4351: out = 16'(437);
			4352: out = 16'(-9121);
			4353: out = 16'(-7579);
			4354: out = 16'(2053);
			4355: out = 16'(13859);
			4356: out = 16'(11547);
			4357: out = 16'(4965);
			4358: out = 16'(-7396);
			4359: out = 16'(-12874);
			4360: out = 16'(-8844);
			4361: out = 16'(6362);
			4362: out = 16'(5937);
			4363: out = 16'(-1588);
			4364: out = 16'(-3629);
			4365: out = 16'(-4671);
			4366: out = 16'(-6510);
			4367: out = 16'(-10848);
			4368: out = 16'(-5007);
			4369: out = 16'(13414);
			4370: out = 16'(19743);
			4371: out = 16'(1010);
			4372: out = 16'(-25837);
			4373: out = 16'(-21324);
			4374: out = 16'(-3298);
			4375: out = 16'(10949);
			4376: out = 16'(5220);
			4377: out = 16'(-2059);
			4378: out = 16'(-11431);
			4379: out = 16'(2471);
			4380: out = 16'(12375);
			4381: out = 16'(2209);
			4382: out = 16'(-22816);
			4383: out = 16'(-21485);
			4384: out = 16'(-1249);
			4385: out = 16'(5370);
			4386: out = 16'(-602);
			4387: out = 16'(-10391);
			4388: out = 16'(-6363);
			4389: out = 16'(4615);
			4390: out = 16'(10142);
			4391: out = 16'(9828);
			4392: out = 16'(13312);
			4393: out = 16'(15769);
			4394: out = 16'(7937);
			4395: out = 16'(-19993);
			4396: out = 16'(-30504);
			4397: out = 16'(-14350);
			4398: out = 16'(10757);
			4399: out = 16'(17874);
			4400: out = 16'(8188);
			4401: out = 16'(-11089);
			4402: out = 16'(-26820);
			4403: out = 16'(-6446);
			4404: out = 16'(9115);
			4405: out = 16'(14137);
			4406: out = 16'(11367);
			4407: out = 16'(2671);
			4408: out = 16'(-5063);
			4409: out = 16'(-12377);
			4410: out = 16'(-13646);
			4411: out = 16'(-685);
			4412: out = 16'(16989);
			4413: out = 16'(22858);
			4414: out = 16'(9596);
			4415: out = 16'(-13109);
			4416: out = 16'(-15620);
			4417: out = 16'(-2599);
			4418: out = 16'(6046);
			4419: out = 16'(29);
			4420: out = 16'(2716);
			4421: out = 16'(2113);
			4422: out = 16'(2464);
			4423: out = 16'(3173);
			4424: out = 16'(11999);
			4425: out = 16'(5996);
			4426: out = 16'(-2742);
			4427: out = 16'(-5422);
			4428: out = 16'(4721);
			4429: out = 16'(3116);
			4430: out = 16'(546);
			4431: out = 16'(787);
			4432: out = 16'(1397);
			4433: out = 16'(1210);
			4434: out = 16'(-4961);
			4435: out = 16'(-7095);
			4436: out = 16'(3515);
			4437: out = 16'(11533);
			4438: out = 16'(14819);
			4439: out = 16'(8972);
			4440: out = 16'(279);
			4441: out = 16'(-562);
			4442: out = 16'(-4008);
			4443: out = 16'(-6502);
			4444: out = 16'(-5220);
			4445: out = 16'(-6151);
			4446: out = 16'(-2400);
			4447: out = 16'(-4941);
			4448: out = 16'(-8813);
			4449: out = 16'(-4236);
			4450: out = 16'(19120);
			4451: out = 16'(23598);
			4452: out = 16'(3627);
			4453: out = 16'(-20966);
			4454: out = 16'(-23637);
			4455: out = 16'(-3024);
			4456: out = 16'(8114);
			4457: out = 16'(-769);
			4458: out = 16'(663);
			4459: out = 16'(3187);
			4460: out = 16'(4154);
			4461: out = 16'(-2041);
			4462: out = 16'(-9414);
			4463: out = 16'(-905);
			4464: out = 16'(9152);
			4465: out = 16'(2578);
			4466: out = 16'(-19656);
			4467: out = 16'(-23106);
			4468: out = 16'(-5569);
			4469: out = 16'(11541);
			4470: out = 16'(8924);
			4471: out = 16'(3322);
			4472: out = 16'(-6325);
			4473: out = 16'(-8576);
			4474: out = 16'(519);
			4475: out = 16'(11957);
			4476: out = 16'(11141);
			4477: out = 16'(-4812);
			4478: out = 16'(-24656);
			4479: out = 16'(-25954);
			4480: out = 16'(-8669);
			4481: out = 16'(9672);
			4482: out = 16'(14640);
			4483: out = 16'(15104);
			4484: out = 16'(2980);
			4485: out = 16'(-2375);
			4486: out = 16'(192);
			4487: out = 16'(2153);
			4488: out = 16'(2967);
			4489: out = 16'(557);
			4490: out = 16'(-2915);
			4491: out = 16'(-7529);
			4492: out = 16'(10190);
			4493: out = 16'(8414);
			4494: out = 16'(-3772);
			4495: out = 16'(-12554);
			4496: out = 16'(181);
			4497: out = 16'(10588);
			4498: out = 16'(15839);
			4499: out = 16'(12829);
			4500: out = 16'(3106);
			4501: out = 16'(-14985);
			4502: out = 16'(-23825);
			4503: out = 16'(-15262);
			4504: out = 16'(2038);
			4505: out = 16'(14465);
			4506: out = 16'(16305);
			4507: out = 16'(8384);
			4508: out = 16'(-783);
			4509: out = 16'(-337);
			4510: out = 16'(11252);
			4511: out = 16'(12040);
			4512: out = 16'(-5443);
			4513: out = 16'(-6328);
			4514: out = 16'(-3733);
			4515: out = 16'(1476);
			4516: out = 16'(3521);
			4517: out = 16'(22315);
			4518: out = 16'(8176);
			4519: out = 16'(-12276);
			4520: out = 16'(-25140);
			4521: out = 16'(-3747);
			4522: out = 16'(1551);
			4523: out = 16'(7264);
			4524: out = 16'(10145);
			4525: out = 16'(13520);
			4526: out = 16'(-3676);
			4527: out = 16'(-4625);
			4528: out = 16'(1470);
			4529: out = 16'(1068);
			4530: out = 16'(-2905);
			4531: out = 16'(111);
			4532: out = 16'(2291);
			4533: out = 16'(-4694);
			4534: out = 16'(-3065);
			4535: out = 16'(6462);
			4536: out = 16'(16921);
			4537: out = 16'(7992);
			4538: out = 16'(-21345);
			4539: out = 16'(-32505);
			4540: out = 16'(-18916);
			4541: out = 16'(2872);
			4542: out = 16'(7379);
			4543: out = 16'(-4035);
			4544: out = 16'(1087);
			4545: out = 16'(11746);
			4546: out = 16'(8977);
			4547: out = 16'(1799);
			4548: out = 16'(4672);
			4549: out = 16'(9910);
			4550: out = 16'(1786);
			4551: out = 16'(-22502);
			4552: out = 16'(-25696);
			4553: out = 16'(-6925);
			4554: out = 16'(9588);
			4555: out = 16'(10125);
			4556: out = 16'(8156);
			4557: out = 16'(4339);
			4558: out = 16'(-639);
			4559: out = 16'(-4591);
			4560: out = 16'(-3788);
			4561: out = 16'(-3116);
			4562: out = 16'(-1469);
			4563: out = 16'(5217);
			4564: out = 16'(-739);
			4565: out = 16'(-9115);
			4566: out = 16'(-12504);
			4567: out = 16'(-3084);
			4568: out = 16'(3606);
			4569: out = 16'(13394);
			4570: out = 16'(14952);
			4571: out = 16'(3603);
			4572: out = 16'(-15320);
			4573: out = 16'(-18460);
			4574: out = 16'(2457);
			4575: out = 16'(20887);
			4576: out = 16'(14304);
			4577: out = 16'(-3064);
			4578: out = 16'(-12584);
			4579: out = 16'(-7268);
			4580: out = 16'(3693);
			4581: out = 16'(9545);
			4582: out = 16'(13631);
			4583: out = 16'(10297);
			4584: out = 16'(-198);
			4585: out = 16'(-12451);
			4586: out = 16'(-6180);
			4587: out = 16'(3493);
			4588: out = 16'(-915);
			4589: out = 16'(-6882);
			4590: out = 16'(-3279);
			4591: out = 16'(6269);
			4592: out = 16'(9699);
			4593: out = 16'(12269);
			4594: out = 16'(10382);
			4595: out = 16'(4959);
			4596: out = 16'(-4387);
			4597: out = 16'(-10257);
			4598: out = 16'(-10017);
			4599: out = 16'(-9276);
			4600: out = 16'(-9521);
			4601: out = 16'(-902);
			4602: out = 16'(3695);
			4603: out = 16'(4413);
			4604: out = 16'(1803);
			4605: out = 16'(9845);
			4606: out = 16'(8697);
			4607: out = 16'(14446);
			4608: out = 16'(5099);
			4609: out = 16'(-12191);
			4610: out = 16'(-24433);
			4611: out = 16'(-6391);
			4612: out = 16'(7904);
			4613: out = 16'(2794);
			4614: out = 16'(-2604);
			4615: out = 16'(-4120);
			4616: out = 16'(-2504);
			4617: out = 16'(2624);
			4618: out = 16'(11291);
			4619: out = 16'(14622);
			4620: out = 16'(2066);
			4621: out = 16'(-10972);
			4622: out = 16'(-8986);
			4623: out = 16'(-5554);
			4624: out = 16'(-11583);
			4625: out = 16'(-12817);
			4626: out = 16'(2365);
			4627: out = 16'(11315);
			4628: out = 16'(8175);
			4629: out = 16'(6831);
			4630: out = 16'(11478);
			4631: out = 16'(510);
			4632: out = 16'(-13163);
			4633: out = 16'(-12732);
			4634: out = 16'(6037);
			4635: out = 16'(7360);
			4636: out = 16'(-436);
			4637: out = 16'(-16609);
			4638: out = 16'(-18828);
			4639: out = 16'(-4710);
			4640: out = 16'(12246);
			4641: out = 16'(19824);
			4642: out = 16'(19096);
			4643: out = 16'(6343);
			4644: out = 16'(-10929);
			4645: out = 16'(-24820);
			4646: out = 16'(-14106);
			4647: out = 16'(7187);
			4648: out = 16'(1768);
			4649: out = 16'(-10920);
			4650: out = 16'(-10618);
			4651: out = 16'(5233);
			4652: out = 16'(6022);
			4653: out = 16'(7548);
			4654: out = 16'(7980);
			4655: out = 16'(7608);
			4656: out = 16'(-7583);
			4657: out = 16'(-12095);
			4658: out = 16'(-11398);
			4659: out = 16'(862);
			4660: out = 16'(9384);
			4661: out = 16'(18662);
			4662: out = 16'(918);
			4663: out = 16'(-15033);
			4664: out = 16'(-7661);
			4665: out = 16'(2595);
			4666: out = 16'(7325);
			4667: out = 16'(1747);
			4668: out = 16'(-1281);
			4669: out = 16'(-5732);
			4670: out = 16'(3248);
			4671: out = 16'(3458);
			4672: out = 16'(718);
			4673: out = 16'(1263);
			4674: out = 16'(6629);
			4675: out = 16'(80);
			4676: out = 16'(-6920);
			4677: out = 16'(-533);
			4678: out = 16'(17053);
			4679: out = 16'(12073);
			4680: out = 16'(-6173);
			4681: out = 16'(-16374);
			4682: out = 16'(-1611);
			4683: out = 16'(8385);
			4684: out = 16'(7210);
			4685: out = 16'(-336);
			4686: out = 16'(-12426);
			4687: out = 16'(-12427);
			4688: out = 16'(87);
			4689: out = 16'(9126);
			4690: out = 16'(-895);
			4691: out = 16'(7735);
			4692: out = 16'(20084);
			4693: out = 16'(16021);
			4694: out = 16'(-12908);
			4695: out = 16'(-27011);
			4696: out = 16'(-16333);
			4697: out = 16'(5386);
			4698: out = 16'(2604);
			4699: out = 16'(-4436);
			4700: out = 16'(-12594);
			4701: out = 16'(-1586);
			4702: out = 16'(13689);
			4703: out = 16'(18134);
			4704: out = 16'(10961);
			4705: out = 16'(5580);
			4706: out = 16'(247);
			4707: out = 16'(996);
			4708: out = 16'(-15784);
			4709: out = 16'(-12509);
			4710: out = 16'(6037);
			4711: out = 16'(11071);
			4712: out = 16'(4377);
			4713: out = 16'(3079);
			4714: out = 16'(4944);
			4715: out = 16'(-6332);
			4716: out = 16'(14);
			4717: out = 16'(-328);
			4718: out = 16'(950);
			4719: out = 16'(1779);
			4720: out = 16'(7517);
			4721: out = 16'(-4769);
			4722: out = 16'(-22289);
			4723: out = 16'(-25752);
			4724: out = 16'(1906);
			4725: out = 16'(19838);
			4726: out = 16'(13865);
			4727: out = 16'(-2661);
			4728: out = 16'(-3643);
			4729: out = 16'(-1794);
			4730: out = 16'(-308);
			4731: out = 16'(-8399);
			4732: out = 16'(-11551);
			4733: out = 16'(-5947);
			4734: out = 16'(13227);
			4735: out = 16'(16878);
			4736: out = 16'(3541);
			4737: out = 16'(-14992);
			4738: out = 16'(-5300);
			4739: out = 16'(7502);
			4740: out = 16'(-1173);
			4741: out = 16'(-10617);
			4742: out = 16'(-6855);
			4743: out = 16'(10157);
			4744: out = 16'(13470);
			4745: out = 16'(2326);
			4746: out = 16'(-11522);
			4747: out = 16'(-3524);
			4748: out = 16'(16177);
			4749: out = 16'(20663);
			4750: out = 16'(-4050);
			4751: out = 16'(-25090);
			4752: out = 16'(-16355);
			4753: out = 16'(17089);
			4754: out = 16'(15509);
			4755: out = 16'(3879);
			4756: out = 16'(-9017);
			4757: out = 16'(-8745);
			4758: out = 16'(-6908);
			4759: out = 16'(3166);
			4760: out = 16'(1857);
			4761: out = 16'(-5152);
			4762: out = 16'(-5059);
			4763: out = 16'(8688);
			4764: out = 16'(12773);
			4765: out = 16'(6853);
			4766: out = 16'(9760);
			4767: out = 16'(8757);
			4768: out = 16'(3738);
			4769: out = 16'(-8357);
			4770: out = 16'(-14596);
			4771: out = 16'(-4860);
			4772: out = 16'(5905);
			4773: out = 16'(1254);
			4774: out = 16'(-11729);
			4775: out = 16'(-29404);
			4776: out = 16'(-9336);
			4777: out = 16'(23021);
			4778: out = 16'(27068);
			4779: out = 16'(4678);
			4780: out = 16'(-19928);
			4781: out = 16'(-29333);
			4782: out = 16'(-18361);
			4783: out = 16'(4119);
			4784: out = 16'(16230);
			4785: out = 16'(16394);
			4786: out = 16'(12080);
			4787: out = 16'(5668);
			4788: out = 16'(-8373);
			4789: out = 16'(-18451);
			4790: out = 16'(-4568);
			4791: out = 16'(22688);
			4792: out = 16'(13899);
			4793: out = 16'(-9824);
			4794: out = 16'(-22668);
			4795: out = 16'(-3252);
			4796: out = 16'(1341);
			4797: out = 16'(10769);
			4798: out = 16'(12745);
			4799: out = 16'(11048);
			4800: out = 16'(-11353);
			4801: out = 16'(-5427);
			4802: out = 16'(1356);
			4803: out = 16'(3225);
			4804: out = 16'(17);
			4805: out = 16'(1872);
			4806: out = 16'(-755);
			4807: out = 16'(-3894);
			4808: out = 16'(-3225);
			4809: out = 16'(-479);
			4810: out = 16'(-1670);
			4811: out = 16'(-2887);
			4812: out = 16'(667);
			4813: out = 16'(109);
			4814: out = 16'(5931);
			4815: out = 16'(12495);
			4816: out = 16'(11114);
			4817: out = 16'(-16838);
			4818: out = 16'(-17307);
			4819: out = 16'(-1650);
			4820: out = 16'(8766);
			4821: out = 16'(-3189);
			4822: out = 16'(-15301);
			4823: out = 16'(-14576);
			4824: out = 16'(3548);
			4825: out = 16'(10616);
			4826: out = 16'(14857);
			4827: out = 16'(2786);
			4828: out = 16'(3241);
			4829: out = 16'(14865);
			4830: out = 16'(5118);
			4831: out = 16'(-18466);
			4832: out = 16'(-23210);
			4833: out = 16'(3233);
			4834: out = 16'(6817);
			4835: out = 16'(3947);
			4836: out = 16'(-222);
			4837: out = 16'(3039);
			4838: out = 16'(3042);
			4839: out = 16'(1301);
			4840: out = 16'(3523);
			4841: out = 16'(11530);
			4842: out = 16'(12124);
			4843: out = 16'(10669);
			4844: out = 16'(698);
			4845: out = 16'(-12583);
			4846: out = 16'(-23260);
			4847: out = 16'(-14419);
			4848: out = 16'(6054);
			4849: out = 16'(17871);
			4850: out = 16'(9828);
			4851: out = 16'(-8217);
			4852: out = 16'(-16230);
			4853: out = 16'(-6998);
			4854: out = 16'(3702);
			4855: out = 16'(514);
			4856: out = 16'(3841);
			4857: out = 16'(9911);
			4858: out = 16'(5551);
			4859: out = 16'(-19954);
			4860: out = 16'(-8923);
			4861: out = 16'(10722);
			4862: out = 16'(14970);
			4863: out = 16'(4792);
			4864: out = 16'(-2935);
			4865: out = 16'(1257);
			4866: out = 16'(2016);
			4867: out = 16'(-10382);
			4868: out = 16'(-21722);
			4869: out = 16'(-13660);
			4870: out = 16'(6282);
			4871: out = 16'(16644);
			4872: out = 16'(17476);
			4873: out = 16'(3941);
			4874: out = 16'(-10861);
			4875: out = 16'(-13238);
			4876: out = 16'(531);
			4877: out = 16'(15016);
			4878: out = 16'(10821);
			4879: out = 16'(-2329);
			4880: out = 16'(-8259);
			4881: out = 16'(-1965);
			4882: out = 16'(-350);
			4883: out = 16'(-1349);
			4884: out = 16'(2088);
			4885: out = 16'(7597);
			4886: out = 16'(-7996);
			4887: out = 16'(-26173);
			4888: out = 16'(-16387);
			4889: out = 16'(8551);
			4890: out = 16'(26136);
			4891: out = 16'(15691);
			4892: out = 16'(-5834);
			4893: out = 16'(-20145);
			4894: out = 16'(-10334);
			4895: out = 16'(2815);
			4896: out = 16'(4689);
			4897: out = 16'(5964);
			4898: out = 16'(325);
			4899: out = 16'(4135);
			4900: out = 16'(8573);
			4901: out = 16'(7501);
			4902: out = 16'(2171);
			4903: out = 16'(3742);
			4904: out = 16'(5688);
			4905: out = 16'(-1515);
			4906: out = 16'(-22586);
			4907: out = 16'(-24951);
			4908: out = 16'(-6301);
			4909: out = 16'(11348);
			4910: out = 16'(16402);
			4911: out = 16'(6273);
			4912: out = 16'(1787);
			4913: out = 16'(6542);
			4914: out = 16'(8111);
			4915: out = 16'(-177);
			4916: out = 16'(-16911);
			4917: out = 16'(-24917);
			4918: out = 16'(-3516);
			4919: out = 16'(6096);
			4920: out = 16'(16151);
			4921: out = 16'(12719);
			4922: out = 16'(-1492);
			4923: out = 16'(-23088);
			4924: out = 16'(-21881);
			4925: out = 16'(-5769);
			4926: out = 16'(7619);
			4927: out = 16'(17985);
			4928: out = 16'(16691);
			4929: out = 16'(4158);
			4930: out = 16'(-13281);
			4931: out = 16'(-20373);
			4932: out = 16'(-5517);
			4933: out = 16'(6925);
			4934: out = 16'(3072);
			4935: out = 16'(2055);
			4936: out = 16'(-13149);
			4937: out = 16'(-8002);
			4938: out = 16'(5824);
			4939: out = 16'(13877);
			4940: out = 16'(7783);
			4941: out = 16'(8386);
			4942: out = 16'(7842);
			4943: out = 16'(87);
			4944: out = 16'(-11851);
			4945: out = 16'(-10761);
			4946: out = 16'(-2969);
			4947: out = 16'(1129);
			4948: out = 16'(9905);
			4949: out = 16'(7435);
			4950: out = 16'(5026);
			4951: out = 16'(320);
			4952: out = 16'(-2619);
			4953: out = 16'(-9444);
			4954: out = 16'(-4926);
			4955: out = 16'(7480);
			4956: out = 16'(19673);
			4957: out = 16'(11102);
			4958: out = 16'(1350);
			4959: out = 16'(-8416);
			4960: out = 16'(-7048);
			4961: out = 16'(-6196);
			4962: out = 16'(12900);
			4963: out = 16'(16807);
			4964: out = 16'(4945);
			4965: out = 16'(-8078);
			4966: out = 16'(-3306);
			4967: out = 16'(-4511);
			4968: out = 16'(-12136);
			4969: out = 16'(-2014);
			4970: out = 16'(12123);
			4971: out = 16'(9489);
			4972: out = 16'(-6745);
			4973: out = 16'(-10929);
			4974: out = 16'(-10727);
			4975: out = 16'(-2884);
			4976: out = 16'(7068);
			4977: out = 16'(18157);
			4978: out = 16'(5475);
			4979: out = 16'(-8169);
			4980: out = 16'(-17537);
			4981: out = 16'(-11897);
			4982: out = 16'(-6570);
			4983: out = 16'(897);
			4984: out = 16'(3385);
			4985: out = 16'(5453);
			4986: out = 16'(178);
			4987: out = 16'(-1300);
			4988: out = 16'(-3796);
			4989: out = 16'(1910);
			4990: out = 16'(8099);
			4991: out = 16'(11856);
			4992: out = 16'(-6869);
			4993: out = 16'(-25144);
			4994: out = 16'(-15133);
			4995: out = 16'(10838);
			4996: out = 16'(11159);
			4997: out = 16'(-8203);
			4998: out = 16'(-16177);
			4999: out = 16'(-5283);
			5000: out = 16'(13729);
			5001: out = 16'(14861);
			5002: out = 16'(3943);
			5003: out = 16'(-18748);
			5004: out = 16'(-5733);
			5005: out = 16'(12041);
			5006: out = 16'(12644);
			5007: out = 16'(1557);
			5008: out = 16'(-11043);
			5009: out = 16'(-18903);
			5010: out = 16'(-19623);
			5011: out = 16'(-11871);
			5012: out = 16'(4521);
			5013: out = 16'(18487);
			5014: out = 16'(20748);
			5015: out = 16'(9263);
			5016: out = 16'(-5318);
			5017: out = 16'(-17212);
			5018: out = 16'(-13598);
			5019: out = 16'(748);
			5020: out = 16'(5663);
			5021: out = 16'(7779);
			5022: out = 16'(11545);
			5023: out = 16'(12347);
			5024: out = 16'(1600);
			5025: out = 16'(-4525);
			5026: out = 16'(4886);
			5027: out = 16'(19311);
			5028: out = 16'(11384);
			5029: out = 16'(-6801);
			5030: out = 16'(-23140);
			5031: out = 16'(-11432);
			5032: out = 16'(15723);
			5033: out = 16'(16918);
			5034: out = 16'(1977);
			5035: out = 16'(-6528);
			5036: out = 16'(1297);
			5037: out = 16'(8225);
			5038: out = 16'(10172);
			5039: out = 16'(12104);
			5040: out = 16'(13308);
			5041: out = 16'(9427);
			5042: out = 16'(-10584);
			5043: out = 16'(-22835);
			5044: out = 16'(-13969);
			5045: out = 16'(162);
			5046: out = 16'(5220);
			5047: out = 16'(2742);
			5048: out = 16'(-2742);
			5049: out = 16'(-15365);
			5050: out = 16'(-3256);
			5051: out = 16'(4404);
			5052: out = 16'(3024);
			5053: out = 16'(-3038);
			5054: out = 16'(-765);
			5055: out = 16'(5788);
			5056: out = 16'(11090);
			5057: out = 16'(10417);
			5058: out = 16'(-3559);
			5059: out = 16'(-2993);
			5060: out = 16'(1203);
			5061: out = 16'(2128);
			5062: out = 16'(8868);
			5063: out = 16'(6143);
			5064: out = 16'(-3022);
			5065: out = 16'(-17747);
			5066: out = 16'(-18492);
			5067: out = 16'(-25073);
			5068: out = 16'(-11075);
			5069: out = 16'(5709);
			5070: out = 16'(5932);
			5071: out = 16'(-6393);
			5072: out = 16'(-8686);
			5073: out = 16'(-1071);
			5074: out = 16'(2961);
			5075: out = 16'(12076);
			5076: out = 16'(14553);
			5077: out = 16'(11571);
			5078: out = 16'(-1221);
			5079: out = 16'(-7753);
			5080: out = 16'(-19954);
			5081: out = 16'(-13241);
			5082: out = 16'(4117);
			5083: out = 16'(9305);
			5084: out = 16'(3367);
			5085: out = 16'(-1379);
			5086: out = 16'(-663);
			5087: out = 16'(159);
			5088: out = 16'(-2377);
			5089: out = 16'(1108);
			5090: out = 16'(7085);
			5091: out = 16'(5318);
			5092: out = 16'(-5500);
			5093: out = 16'(-8128);
			5094: out = 16'(-56);
			5095: out = 16'(5290);
			5096: out = 16'(8940);
			5097: out = 16'(5327);
			5098: out = 16'(7486);
			5099: out = 16'(7753);
			5100: out = 16'(787);
			5101: out = 16'(-15026);
			5102: out = 16'(-17374);
			5103: out = 16'(-7032);
			5104: out = 16'(284);
			5105: out = 16'(6877);
			5106: out = 16'(10907);
			5107: out = 16'(8322);
			5108: out = 16'(114);
			5109: out = 16'(-9160);
			5110: out = 16'(-3644);
			5111: out = 16'(5122);
			5112: out = 16'(8478);
			5113: out = 16'(8814);
			5114: out = 16'(5178);
			5115: out = 16'(-11238);
			5116: out = 16'(-26897);
			5117: out = 16'(-10454);
			5118: out = 16'(6518);
			5119: out = 16'(6596);
			5120: out = 16'(1807);
			5121: out = 16'(9433);
			5122: out = 16'(15356);
			5123: out = 16'(1771);
			5124: out = 16'(-11668);
			5125: out = 16'(4048);
			5126: out = 16'(17840);
			5127: out = 16'(11402);
			5128: out = 16'(-8385);
			5129: out = 16'(-17419);
			5130: out = 16'(-27259);
			5131: out = 16'(-11767);
			5132: out = 16'(12592);
			5133: out = 16'(24299);
			5134: out = 16'(10631);
			5135: out = 16'(-165);
			5136: out = 16'(-2105);
			5137: out = 16'(1365);
			5138: out = 16'(-5100);
			5139: out = 16'(-7266);
			5140: out = 16'(1925);
			5141: out = 16'(12910);
			5142: out = 16'(2992);
			5143: out = 16'(-2003);
			5144: out = 16'(-7575);
			5145: out = 16'(-109);
			5146: out = 16'(9446);
			5147: out = 16'(19404);
			5148: out = 16'(8614);
			5149: out = 16'(-3427);
			5150: out = 16'(-9383);
			5151: out = 16'(-5699);
			5152: out = 16'(-6190);
			5153: out = 16'(-1304);
			5154: out = 16'(5226);
			5155: out = 16'(4798);
			5156: out = 16'(5022);
			5157: out = 16'(8347);
			5158: out = 16'(4199);
			5159: out = 16'(-13962);
			5160: out = 16'(-26129);
			5161: out = 16'(-14416);
			5162: out = 16'(8984);
			5163: out = 16'(13837);
			5164: out = 16'(-2010);
			5165: out = 16'(-12270);
			5166: out = 16'(-7531);
			5167: out = 16'(2121);
			5168: out = 16'(2074);
			5169: out = 16'(6780);
			5170: out = 16'(9050);
			5171: out = 16'(2637);
			5172: out = 16'(-3653);
			5173: out = 16'(-8796);
			5174: out = 16'(-4598);
			5175: out = 16'(1640);
			5176: out = 16'(4751);
			5177: out = 16'(-11296);
			5178: out = 16'(-20943);
			5179: out = 16'(-14587);
			5180: out = 16'(-1153);
			5181: out = 16'(3030);
			5182: out = 16'(732);
			5183: out = 16'(-425);
			5184: out = 16'(1892);
			5185: out = 16'(15419);
			5186: out = 16'(9096);
			5187: out = 16'(-2851);
			5188: out = 16'(-6727);
			5189: out = 16'(1094);
			5190: out = 16'(6359);
			5191: out = 16'(4669);
			5192: out = 16'(-551);
			5193: out = 16'(-4197);
			5194: out = 16'(-1368);
			5195: out = 16'(1315);
			5196: out = 16'(156);
			5197: out = 16'(1258);
			5198: out = 16'(6993);
			5199: out = 16'(12363);
			5200: out = 16'(3826);
			5201: out = 16'(-15669);
			5202: out = 16'(-20217);
			5203: out = 16'(-1179);
			5204: out = 16'(17007);
			5205: out = 16'(12498);
			5206: out = 16'(8712);
			5207: out = 16'(3841);
			5208: out = 16'(6229);
			5209: out = 16'(1620);
			5210: out = 16'(-8033);
			5211: out = 16'(-10041);
			5212: out = 16'(10342);
			5213: out = 16'(23199);
			5214: out = 16'(6878);
			5215: out = 16'(-17947);
			5216: out = 16'(-22146);
			5217: out = 16'(-381);
			5218: out = 16'(11715);
			5219: out = 16'(11576);
			5220: out = 16'(747);
			5221: out = 16'(-3211);
			5222: out = 16'(232);
			5223: out = 16'(4276);
			5224: out = 16'(-2063);
			5225: out = 16'(-11012);
			5226: out = 16'(-12193);
			5227: out = 16'(1593);
			5228: out = 16'(2563);
			5229: out = 16'(-6946);
			5230: out = 16'(-15760);
			5231: out = 16'(-10020);
			5232: out = 16'(-2107);
			5233: out = 16'(3937);
			5234: out = 16'(5637);
			5235: out = 16'(5596);
			5236: out = 16'(8970);
			5237: out = 16'(5763);
			5238: out = 16'(-3808);
			5239: out = 16'(-10857);
			5240: out = 16'(-5361);
			5241: out = 16'(6392);
			5242: out = 16'(10591);
			5243: out = 16'(1764);
			5244: out = 16'(-22118);
			5245: out = 16'(-27532);
			5246: out = 16'(-13077);
			5247: out = 16'(4794);
			5248: out = 16'(8583);
			5249: out = 16'(14161);
			5250: out = 16'(12381);
			5251: out = 16'(989);
			5252: out = 16'(-9702);
			5253: out = 16'(-4219);
			5254: out = 16'(14092);
			5255: out = 16'(20538);
			5256: out = 16'(10448);
			5257: out = 16'(-19646);
			5258: out = 16'(-22149);
			5259: out = 16'(-4493);
			5260: out = 16'(3505);
			5261: out = 16'(6192);
			5262: out = 16'(5049);
			5263: out = 16'(3868);
			5264: out = 16'(-2493);
			5265: out = 16'(1679);
			5266: out = 16'(-7624);
			5267: out = 16'(-5236);
			5268: out = 16'(7520);
			5269: out = 16'(15227);
			5270: out = 16'(4210);
			5271: out = 16'(-10157);
			5272: out = 16'(-12737);
			5273: out = 16'(1487);
			5274: out = 16'(13930);
			5275: out = 16'(11994);
			5276: out = 16'(-458);
			5277: out = 16'(-7063);
			5278: out = 16'(-2075);
			5279: out = 16'(3460);
			5280: out = 16'(-3077);
			5281: out = 16'(-8319);
			5282: out = 16'(-188);
			5283: out = 16'(22107);
			5284: out = 16'(23762);
			5285: out = 16'(8630);
			5286: out = 16'(-6476);
			5287: out = 16'(-8347);
			5288: out = 16'(-15935);
			5289: out = 16'(-21991);
			5290: out = 16'(-4098);
			5291: out = 16'(19049);
			5292: out = 16'(17220);
			5293: out = 16'(-5750);
			5294: out = 16'(-26508);
			5295: out = 16'(-30075);
			5296: out = 16'(-21803);
			5297: out = 16'(7823);
			5298: out = 16'(29720);
			5299: out = 16'(28873);
			5300: out = 16'(5662);
			5301: out = 16'(-17612);
			5302: out = 16'(-20280);
			5303: out = 16'(-1303);
			5304: out = 16'(6073);
			5305: out = 16'(10103);
			5306: out = 16'(12272);
			5307: out = 16'(-2713);
			5308: out = 16'(-22711);
			5309: out = 16'(-27551);
			5310: out = 16'(-4388);
			5311: out = 16'(17065);
			5312: out = 16'(19156);
			5313: out = 16'(3082);
			5314: out = 16'(-7674);
			5315: out = 16'(-5133);
			5316: out = 16'(7260);
			5317: out = 16'(7723);
			5318: out = 16'(7671);
			5319: out = 16'(6809);
			5320: out = 16'(8);
			5321: out = 16'(-9961);
			5322: out = 16'(-6971);
			5323: out = 16'(-116);
			5324: out = 16'(-8991);
			5325: out = 16'(-7674);
			5326: out = 16'(7233);
			5327: out = 16'(13762);
			5328: out = 16'(-5005);
			5329: out = 16'(-18404);
			5330: out = 16'(-11038);
			5331: out = 16'(4425);
			5332: out = 16'(1580);
			5333: out = 16'(1647);
			5334: out = 16'(7295);
			5335: out = 16'(13986);
			5336: out = 16'(7344);
			5337: out = 16'(882);
			5338: out = 16'(-13518);
			5339: out = 16'(-20991);
			5340: out = 16'(-15320);
			5341: out = 16'(2916);
			5342: out = 16'(13281);
			5343: out = 16'(8567);
			5344: out = 16'(-5254);
			5345: out = 16'(-17365);
			5346: out = 16'(-561);
			5347: out = 16'(14739);
			5348: out = 16'(17519);
			5349: out = 16'(13173);
			5350: out = 16'(7281);
			5351: out = 16'(-5478);
			5352: out = 16'(-15302);
			5353: out = 16'(-8306);
			5354: out = 16'(12973);
			5355: out = 16'(16496);
			5356: out = 16'(3810);
			5357: out = 16'(-9040);
			5358: out = 16'(-10355);
			5359: out = 16'(-1644);
			5360: out = 16'(2400);
			5361: out = 16'(-972);
			5362: out = 16'(-3552);
			5363: out = 16'(13710);
			5364: out = 16'(24109);
			5365: out = 16'(14909);
			5366: out = 16'(-1761);
			5367: out = 16'(-21156);
			5368: out = 16'(-12183);
			5369: out = 16'(9220);
			5370: out = 16'(14117);
			5371: out = 16'(3019);
			5372: out = 16'(-3707);
			5373: out = 16'(-2467);
			5374: out = 16'(-2146);
			5375: out = 16'(3892);
			5376: out = 16'(-954);
			5377: out = 16'(1386);
			5378: out = 16'(6772);
			5379: out = 16'(7560);
			5380: out = 16'(-12000);
			5381: out = 16'(-19264);
			5382: out = 16'(-2656);
			5383: out = 16'(14725);
			5384: out = 16'(21271);
			5385: out = 16'(8063);
			5386: out = 16'(-11044);
			5387: out = 16'(-24941);
			5388: out = 16'(-13822);
			5389: out = 16'(-4039);
			5390: out = 16'(-658);
			5391: out = 16'(1677);
			5392: out = 16'(8395);
			5393: out = 16'(4864);
			5394: out = 16'(-7870);
			5395: out = 16'(-13367);
			5396: out = 16'(16987);
			5397: out = 16'(15101);
			5398: out = 16'(3742);
			5399: out = 16'(-5903);
			5400: out = 16'(-1331);
			5401: out = 16'(-2457);
			5402: out = 16'(1882);
			5403: out = 16'(3412);
			5404: out = 16'(-5883);
			5405: out = 16'(-3070);
			5406: out = 16'(-8094);
			5407: out = 16'(-12219);
			5408: out = 16'(-8456);
			5409: out = 16'(1905);
			5410: out = 16'(13909);
			5411: out = 16'(19350);
			5412: out = 16'(11148);
			5413: out = 16'(-13994);
			5414: out = 16'(-19147);
			5415: out = 16'(-7390);
			5416: out = 16'(-270);
			5417: out = 16'(-4871);
			5418: out = 16'(569);
			5419: out = 16'(16065);
			5420: out = 16'(18115);
			5421: out = 16'(6434);
			5422: out = 16'(-19013);
			5423: out = 16'(-12750);
			5424: out = 16'(2031);
			5425: out = 16'(-4102);
			5426: out = 16'(-7278);
			5427: out = 16'(2557);
			5428: out = 16'(9147);
			5429: out = 16'(-2015);
			5430: out = 16'(-7922);
			5431: out = 16'(1577);
			5432: out = 16'(17243);
			5433: out = 16'(18976);
			5434: out = 16'(5362);
			5435: out = 16'(-1924);
			5436: out = 16'(-12632);
			5437: out = 16'(-21702);
			5438: out = 16'(-16407);
			5439: out = 16'(1608);
			5440: out = 16'(11651);
			5441: out = 16'(11756);
			5442: out = 16'(8804);
			5443: out = 16'(2615);
			5444: out = 16'(-10454);
			5445: out = 16'(-13799);
			5446: out = 16'(2711);
			5447: out = 16'(6772);
			5448: out = 16'(10948);
			5449: out = 16'(8056);
			5450: out = 16'(222);
			5451: out = 16'(-3367);
			5452: out = 16'(-10894);
			5453: out = 16'(-4739);
			5454: out = 16'(6462);
			5455: out = 16'(4952);
			5456: out = 16'(-4845);
			5457: out = 16'(-4692);
			5458: out = 16'(5353);
			5459: out = 16'(8936);
			5460: out = 16'(11884);
			5461: out = 16'(8335);
			5462: out = 16'(2404);
			5463: out = 16'(-172);
			5464: out = 16'(-15946);
			5465: out = 16'(-9230);
			5466: out = 16'(3262);
			5467: out = 16'(9479);
			5468: out = 16'(4375);
			5469: out = 16'(12725);
			5470: out = 16'(11897);
			5471: out = 16'(525);
			5472: out = 16'(-22530);
			5473: out = 16'(-8596);
			5474: out = 16'(-3600);
			5475: out = 16'(-9418);
			5476: out = 16'(4744);
			5477: out = 16'(20341);
			5478: out = 16'(15748);
			5479: out = 16'(-9066);
			5480: out = 16'(-26284);
			5481: out = 16'(-13425);
			5482: out = 16'(6320);
			5483: out = 16'(8109);
			5484: out = 16'(-511);
			5485: out = 16'(-7195);
			5486: out = 16'(-8849);
			5487: out = 16'(-4725);
			5488: out = 16'(3870);
			5489: out = 16'(7190);
			5490: out = 16'(5110);
			5491: out = 16'(-3672);
			5492: out = 16'(-9158);
			5493: out = 16'(-1667);
			5494: out = 16'(-2108);
			5495: out = 16'(-3429);
			5496: out = 16'(-1060);
			5497: out = 16'(3801);
			5498: out = 16'(6745);
			5499: out = 16'(3505);
			5500: out = 16'(-1095);
			5501: out = 16'(-3351);
			5502: out = 16'(-8677);
			5503: out = 16'(-6179);
			5504: out = 16'(5951);
			5505: out = 16'(15683);
			5506: out = 16'(9143);
			5507: out = 16'(899);
			5508: out = 16'(390);
			5509: out = 16'(4805);
			5510: out = 16'(298);
			5511: out = 16'(-546);
			5512: out = 16'(2186);
			5513: out = 16'(4018);
			5514: out = 16'(-411);
			5515: out = 16'(-8545);
			5516: out = 16'(-8765);
			5517: out = 16'(-2647);
			5518: out = 16'(3860);
			5519: out = 16'(3865);
			5520: out = 16'(13889);
			5521: out = 16'(16489);
			5522: out = 16'(173);
			5523: out = 16'(-22589);
			5524: out = 16'(-28005);
			5525: out = 16'(-8104);
			5526: out = 16'(16095);
			5527: out = 16'(15912);
			5528: out = 16'(17224);
			5529: out = 16'(7175);
			5530: out = 16'(-7519);
			5531: out = 16'(-18762);
			5532: out = 16'(1075);
			5533: out = 16'(13409);
			5534: out = 16'(6699);
			5535: out = 16'(-4679);
			5536: out = 16'(-694);
			5537: out = 16'(1026);
			5538: out = 16'(-7144);
			5539: out = 16'(-13469);
			5540: out = 16'(13208);
			5541: out = 16'(13464);
			5542: out = 16'(-11585);
			5543: out = 16'(-28808);
			5544: out = 16'(-10216);
			5545: out = 16'(15207);
			5546: out = 16'(13102);
			5547: out = 16'(301);
			5548: out = 16'(1260);
			5549: out = 16'(6725);
			5550: out = 16'(172);
			5551: out = 16'(-6764);
			5552: out = 16'(12971);
			5553: out = 16'(20697);
			5554: out = 16'(11343);
			5555: out = 16'(-15493);
			5556: out = 16'(-26722);
			5557: out = 16'(-27988);
			5558: out = 16'(-2905);
			5559: out = 16'(11687);
			5560: out = 16'(7405);
			5561: out = 16'(-5199);
			5562: out = 16'(27);
			5563: out = 16'(6504);
			5564: out = 16'(3459);
			5565: out = 16'(2492);
			5566: out = 16'(3000);
			5567: out = 16'(6172);
			5568: out = 16'(3976);
			5569: out = 16'(-1493);
			5570: out = 16'(812);
			5571: out = 16'(7051);
			5572: out = 16'(5115);
			5573: out = 16'(-8816);
			5574: out = 16'(-26600);
			5575: out = 16'(-18226);
			5576: out = 16'(11064);
			5577: out = 16'(23961);
			5578: out = 16'(15429);
			5579: out = 16'(-8125);
			5580: out = 16'(-24905);
			5581: out = 16'(-22944);
			5582: out = 16'(-3469);
			5583: out = 16'(7972);
			5584: out = 16'(14107);
			5585: out = 16'(15055);
			5586: out = 16'(11529);
			5587: out = 16'(-7614);
			5588: out = 16'(-16641);
			5589: out = 16'(-10101);
			5590: out = 16'(243);
			5591: out = 16'(1690);
			5592: out = 16'(6358);
			5593: out = 16'(4676);
			5594: out = 16'(-14971);
			5595: out = 16'(836);
			5596: out = 16'(5594);
			5597: out = 16'(11547);
			5598: out = 16'(5015);
			5599: out = 16'(-6285);
			5600: out = 16'(-26254);
			5601: out = 16'(-14096);
			5602: out = 16'(13135);
			5603: out = 16'(15712);
			5604: out = 16'(4945);
			5605: out = 16'(3137);
			5606: out = 16'(2060);
			5607: out = 16'(-7968);
			5608: out = 16'(-23842);
			5609: out = 16'(-10372);
			5610: out = 16'(10008);
			5611: out = 16'(11749);
			5612: out = 16'(2284);
			5613: out = 16'(14011);
			5614: out = 16'(15393);
			5615: out = 16'(-5207);
			5616: out = 16'(-21386);
			5617: out = 16'(-4020);
			5618: out = 16'(7214);
			5619: out = 16'(-7193);
			5620: out = 16'(1588);
			5621: out = 16'(9040);
			5622: out = 16'(9328);
			5623: out = 16'(-5526);
			5624: out = 16'(-2430);
			5625: out = 16'(4027);
			5626: out = 16'(12690);
			5627: out = 16'(1441);
			5628: out = 16'(-14210);
			5629: out = 16'(-21156);
			5630: out = 16'(-7245);
			5631: out = 16'(124);
			5632: out = 16'(-1287);
			5633: out = 16'(9744);
			5634: out = 16'(17343);
			5635: out = 16'(4309);
			5636: out = 16'(-19366);
			5637: out = 16'(-22980);
			5638: out = 16'(-25);
			5639: out = 16'(16820);
			5640: out = 16'(13483);
			5641: out = 16'(5563);
			5642: out = 16'(1611);
			5643: out = 16'(-4366);
			5644: out = 16'(-5450);
			5645: out = 16'(9794);
			5646: out = 16'(11690);
			5647: out = 16'(3397);
			5648: out = 16'(-9343);
			5649: out = 16'(-12465);
			5650: out = 16'(-2152);
			5651: out = 16'(4214);
			5652: out = 16'(4244);
			5653: out = 16'(1187);
			5654: out = 16'(1155);
			5655: out = 16'(-9474);
			5656: out = 16'(-9947);
			5657: out = 16'(2866);
			5658: out = 16'(7157);
			5659: out = 16'(-2999);
			5660: out = 16'(-5294);
			5661: out = 16'(12219);
			5662: out = 16'(22121);
			5663: out = 16'(16918);
			5664: out = 16'(-10259);
			5665: out = 16'(-30016);
			5666: out = 16'(-27869);
			5667: out = 16'(-21420);
			5668: out = 16'(-8233);
			5669: out = 16'(11605);
			5670: out = 16'(28064);
			5671: out = 16'(14995);
			5672: out = 16'(-3810);
			5673: out = 16'(-23314);
			5674: out = 16'(-26743);
			5675: out = 16'(-13391);
			5676: out = 16'(10818);
			5677: out = 16'(22262);
			5678: out = 16'(18433);
			5679: out = 16'(2144);
			5680: out = 16'(-13287);
			5681: out = 16'(-17976);
			5682: out = 16'(922);
			5683: out = 16'(24094);
			5684: out = 16'(18952);
			5685: out = 16'(-7069);
			5686: out = 16'(-27256);
			5687: out = 16'(-16243);
			5688: out = 16'(-5855);
			5689: out = 16'(12935);
			5690: out = 16'(23809);
			5691: out = 16'(16979);
			5692: out = 16'(-21240);
			5693: out = 16'(-32118);
			5694: out = 16'(-17225);
			5695: out = 16'(13308);
			5696: out = 16'(15870);
			5697: out = 16'(22499);
			5698: out = 16'(18158);
			5699: out = 16'(1098);
			5700: out = 16'(-25462);
			5701: out = 16'(-23463);
			5702: out = 16'(-2515);
			5703: out = 16'(12422);
			5704: out = 16'(9258);
			5705: out = 16'(6472);
			5706: out = 16'(5555);
			5707: out = 16'(3062);
			5708: out = 16'(-3685);
			5709: out = 16'(-9258);
			5710: out = 16'(-197);
			5711: out = 16'(7365);
			5712: out = 16'(3015);
			5713: out = 16'(-8286);
			5714: out = 16'(1120);
			5715: out = 16'(9093);
			5716: out = 16'(40);
			5717: out = 16'(-16762);
			5718: out = 16'(-12903);
			5719: out = 16'(6316);
			5720: out = 16'(17841);
			5721: out = 16'(13831);
			5722: out = 16'(3385);
			5723: out = 16'(-8143);
			5724: out = 16'(-12937);
			5725: out = 16'(-3616);
			5726: out = 16'(8203);
			5727: out = 16'(16850);
			5728: out = 16'(7157);
			5729: out = 16'(-12184);
			5730: out = 16'(-16321);
			5731: out = 16'(-10662);
			5732: out = 16'(-199);
			5733: out = 16'(6513);
			5734: out = 16'(5120);
			5735: out = 16'(2987);
			5736: out = 16'(-3261);
			5737: out = 16'(-5475);
			5738: out = 16'(-4019);
			5739: out = 16'(19577);
			5740: out = 16'(13569);
			5741: out = 16'(-6356);
			5742: out = 16'(-18978);
			5743: out = 16'(6452);
			5744: out = 16'(10880);
			5745: out = 16'(1438);
			5746: out = 16'(-5727);
			5747: out = 16'(3231);
			5748: out = 16'(1569);
			5749: out = 16'(-211);
			5750: out = 16'(-3435);
			5751: out = 16'(-11623);
			5752: out = 16'(-9345);
			5753: out = 16'(9607);
			5754: out = 16'(19747);
			5755: out = 16'(8312);
			5756: out = 16'(-2169);
			5757: out = 16'(5313);
			5758: out = 16'(6237);
			5759: out = 16'(-19872);
			5760: out = 16'(-19024);
			5761: out = 16'(8332);
			5762: out = 16'(27527);
			5763: out = 16'(7175);
			5764: out = 16'(-9317);
			5765: out = 16'(-27362);
			5766: out = 16'(-21962);
			5767: out = 16'(-6049);
			5768: out = 16'(16130);
			5769: out = 16'(17554);
			5770: out = 16'(13440);
			5771: out = 16'(1617);
			5772: out = 16'(626);
			5773: out = 16'(-11977);
			5774: out = 16'(3596);
			5775: out = 16'(20867);
			5776: out = 16'(15859);
			5777: out = 16'(-13264);
			5778: out = 16'(-27326);
			5779: out = 16'(-19259);
			5780: out = 16'(-1176);
			5781: out = 16'(6456);
			5782: out = 16'(15126);
			5783: out = 16'(9913);
			5784: out = 16'(-4118);
			5785: out = 16'(-3367);
			5786: out = 16'(3397);
			5787: out = 16'(122);
			5788: out = 16'(-5148);
			5789: out = 16'(19379);
			5790: out = 16'(16664);
			5791: out = 16'(844);
			5792: out = 16'(-19397);
			5793: out = 16'(-16136);
			5794: out = 16'(-20295);
			5795: out = 16'(-9134);
			5796: out = 16'(8100);
			5797: out = 16'(18622);
			5798: out = 16'(-1600);
			5799: out = 16'(-15004);
			5800: out = 16'(-9859);
			5801: out = 16'(8213);
			5802: out = 16'(2620);
			5803: out = 16'(91);
			5804: out = 16'(953);
			5805: out = 16'(5810);
			5806: out = 16'(321);
			5807: out = 16'(-8061);
			5808: out = 16'(-18486);
			5809: out = 16'(-16397);
			5810: out = 16'(2468);
			5811: out = 16'(1077);
			5812: out = 16'(1342);
			5813: out = 16'(13322);
			5814: out = 16'(27058);
			5815: out = 16'(6373);
			5816: out = 16'(-18147);
			5817: out = 16'(-27593);
			5818: out = 16'(-8635);
			5819: out = 16'(16498);
			5820: out = 16'(24299);
			5821: out = 16'(13613);
			5822: out = 16'(-908);
			5823: out = 16'(-4146);
			5824: out = 16'(-500);
			5825: out = 16'(2892);
			5826: out = 16'(-791);
			5827: out = 16'(-12598);
			5828: out = 16'(-9956);
			5829: out = 16'(-5513);
			5830: out = 16'(-3343);
			5831: out = 16'(2658);
			5832: out = 16'(16331);
			5833: out = 16'(23054);
			5834: out = 16'(14302);
			5835: out = 16'(-1802);
			5836: out = 16'(-27113);
			5837: out = 16'(-15125);
			5838: out = 16'(10930);
			5839: out = 16'(18021);
			5840: out = 16'(3209);
			5841: out = 16'(26);
			5842: out = 16'(-2672);
			5843: out = 16'(-10988);
			5844: out = 16'(-19710);
			5845: out = 16'(-5975);
			5846: out = 16'(13578);
			5847: out = 16'(17568);
			5848: out = 16'(5017);
			5849: out = 16'(2308);
			5850: out = 16'(7439);
			5851: out = 16'(14387);
			5852: out = 16'(7237);
			5853: out = 16'(-11225);
			5854: out = 16'(-26750);
			5855: out = 16'(-13284);
			5856: out = 16'(11320);
			5857: out = 16'(9622);
			5858: out = 16'(-17694);
			5859: out = 16'(-23560);
			5860: out = 16'(7616);
			5861: out = 16'(22894);
			5862: out = 16'(19233);
			5863: out = 16'(8263);
			5864: out = 16'(501);
			5865: out = 16'(-14449);
			5866: out = 16'(-26969);
			5867: out = 16'(-23175);
			5868: out = 16'(1342);
			5869: out = 16'(15561);
			5870: out = 16'(18122);
			5871: out = 16'(6418);
			5872: out = 16'(-1529);
			5873: out = 16'(-2910);
			5874: out = 16'(2244);
			5875: out = 16'(-5086);
			5876: out = 16'(-10917);
			5877: out = 16'(-8923);
			5878: out = 16'(-7795);
			5879: out = 16'(-782);
			5880: out = 16'(9075);
			5881: out = 16'(15497);
			5882: out = 16'(12041);
			5883: out = 16'(103);
			5884: out = 16'(-8429);
			5885: out = 16'(-9153);
			5886: out = 16'(-7604);
			5887: out = 16'(-692);
			5888: out = 16'(6332);
			5889: out = 16'(9794);
			5890: out = 16'(4178);
			5891: out = 16'(638);
			5892: out = 16'(-7334);
			5893: out = 16'(-6633);
			5894: out = 16'(3055);
			5895: out = 16'(587);
			5896: out = 16'(6738);
			5897: out = 16'(12832);
			5898: out = 16'(15781);
			5899: out = 16'(11236);
			5900: out = 16'(5602);
			5901: out = 16'(-11345);
			5902: out = 16'(-29972);
			5903: out = 16'(-26744);
			5904: out = 16'(-9590);
			5905: out = 16'(15527);
			5906: out = 16'(23884);
			5907: out = 16'(19258);
			5908: out = 16'(10144);
			5909: out = 16'(6573);
			5910: out = 16'(-4038);
			5911: out = 16'(-19131);
			5912: out = 16'(-15787);
			5913: out = 16'(6790);
			5914: out = 16'(17468);
			5915: out = 16'(3734);
			5916: out = 16'(-23430);
			5917: out = 16'(-15720);
			5918: out = 16'(6790);
			5919: out = 16'(11118);
			5920: out = 16'(1416);
			5921: out = 16'(-9325);
			5922: out = 16'(-9056);
			5923: out = 16'(-899);
			5924: out = 16'(10024);
			5925: out = 16'(10502);
			5926: out = 16'(11948);
			5927: out = 16'(9302);
			5928: out = 16'(438);
			5929: out = 16'(-11084);
			5930: out = 16'(-10768);
			5931: out = 16'(2696);
			5932: out = 16'(12654);
			5933: out = 16'(8898);
			5934: out = 16'(-16101);
			5935: out = 16'(-30204);
			5936: out = 16'(-14676);
			5937: out = 16'(6895);
			5938: out = 16'(18217);
			5939: out = 16'(10043);
			5940: out = 16'(533);
			5941: out = 16'(-3561);
			5942: out = 16'(-1800);
			5943: out = 16'(-10614);
			5944: out = 16'(-13975);
			5945: out = 16'(2347);
			5946: out = 16'(17344);
			5947: out = 16'(16650);
			5948: out = 16'(8863);
			5949: out = 16'(4570);
			5950: out = 16'(2313);
			5951: out = 16'(-9362);
			5952: out = 16'(-24200);
			5953: out = 16'(-28509);
			5954: out = 16'(-8648);
			5955: out = 16'(7400);
			5956: out = 16'(19846);
			5957: out = 16'(23303);
			5958: out = 16'(13487);
			5959: out = 16'(-9729);
			5960: out = 16'(-16447);
			5961: out = 16'(-4529);
			5962: out = 16'(-1095);
			5963: out = 16'(-2760);
			5964: out = 16'(-3353);
			5965: out = 16'(3211);
			5966: out = 16'(4147);
			5967: out = 16'(-733);
			5968: out = 16'(-886);
			5969: out = 16'(10418);
			5970: out = 16'(14016);
			5971: out = 16'(-9577);
			5972: out = 16'(-29225);
			5973: out = 16'(-20257);
			5974: out = 16'(10561);
			5975: out = 16'(21090);
			5976: out = 16'(12651);
			5977: out = 16'(1135);
			5978: out = 16'(-9921);
			5979: out = 16'(-17303);
			5980: out = 16'(-2228);
			5981: out = 16'(22472);
			5982: out = 16'(21341);
			5983: out = 16'(-10127);
			5984: out = 16'(-26623);
			5985: out = 16'(-14863);
			5986: out = 16'(5562);
			5987: out = 16'(3272);
			5988: out = 16'(15552);
			5989: out = 16'(13724);
			5990: out = 16'(10163);
			5991: out = 16'(-739);
			5992: out = 16'(-3286);
			5993: out = 16'(-6779);
			5994: out = 16'(-966);
			5995: out = 16'(379);
			5996: out = 16'(-326);
			5997: out = 16'(-2256);
			5998: out = 16'(11181);
			5999: out = 16'(18665);
			6000: out = 16'(10419);
			6001: out = 16'(-9927);
			6002: out = 16'(-8604);
			6003: out = 16'(2438);
			6004: out = 16'(-203);
			6005: out = 16'(-11347);
			6006: out = 16'(-2726);
			6007: out = 16'(14481);
			6008: out = 16'(11841);
			6009: out = 16'(2871);
			6010: out = 16'(-18442);
			6011: out = 16'(-16092);
			6012: out = 16'(3219);
			6013: out = 16'(5309);
			6014: out = 16'(-1198);
			6015: out = 16'(-5533);
			6016: out = 16'(2204);
			6017: out = 16'(8190);
			6018: out = 16'(12924);
			6019: out = 16'(1929);
			6020: out = 16'(-4127);
			6021: out = 16'(5356);
			6022: out = 16'(4419);
			6023: out = 16'(-2061);
			6024: out = 16'(-7008);
			6025: out = 16'(1814);
			6026: out = 16'(4075);
			6027: out = 16'(3956);
			6028: out = 16'(-7319);
			6029: out = 16'(-12458);
			6030: out = 16'(-6983);
			6031: out = 16'(6293);
			6032: out = 16'(1683);
			6033: out = 16'(-2980);
			6034: out = 16'(8313);
			6035: out = 16'(3548);
			6036: out = 16'(-13906);
			6037: out = 16'(-17383);
			6038: out = 16'(10549);
			6039: out = 16'(9628);
			6040: out = 16'(2495);
			6041: out = 16'(260);
			6042: out = 16'(8064);
			6043: out = 16'(6769);
			6044: out = 16'(-11183);
			6045: out = 16'(-22293);
			6046: out = 16'(-10005);
			6047: out = 16'(447);
			6048: out = 16'(1994);
			6049: out = 16'(3424);
			6050: out = 16'(11761);
			6051: out = 16'(11702);
			6052: out = 16'(-3405);
			6053: out = 16'(-13650);
			6054: out = 16'(-2440);
			6055: out = 16'(14218);
			6056: out = 16'(1405);
			6057: out = 16'(-9998);
			6058: out = 16'(-1998);
			6059: out = 16'(15239);
			6060: out = 16'(1961);
			6061: out = 16'(-1956);
			6062: out = 16'(6132);
			6063: out = 16'(13636);
			6064: out = 16'(-3777);
			6065: out = 16'(-9998);
			6066: out = 16'(-6249);
			6067: out = 16'(136);
			6068: out = 16'(-4901);
			6069: out = 16'(-4236);
			6070: out = 16'(1565);
			6071: out = 16'(5603);
			6072: out = 16'(-2122);
			6073: out = 16'(-4224);
			6074: out = 16'(-468);
			6075: out = 16'(7559);
			6076: out = 16'(7352);
			6077: out = 16'(-1773);
			6078: out = 16'(-14698);
			6079: out = 16'(-14996);
			6080: out = 16'(1709);
			6081: out = 16'(11118);
			6082: out = 16'(21957);
			6083: out = 16'(20328);
			6084: out = 16'(7116);
			6085: out = 16'(-19106);
			6086: out = 16'(-21974);
			6087: out = 16'(-12797);
			6088: out = 16'(-3563);
			6089: out = 16'(-4805);
			6090: out = 16'(9897);
			6091: out = 16'(13159);
			6092: out = 16'(6531);
			6093: out = 16'(-5294);
			6094: out = 16'(-134);
			6095: out = 16'(-5382);
			6096: out = 16'(-9651);
			6097: out = 16'(-41);
			6098: out = 16'(21108);
			6099: out = 16'(18160);
			6100: out = 16'(232);
			6101: out = 16'(-16988);
			6102: out = 16'(-19133);
			6103: out = 16'(-9367);
			6104: out = 16'(4768);
			6105: out = 16'(12238);
			6106: out = 16'(11472);
			6107: out = 16'(2700);
			6108: out = 16'(-925);
			6109: out = 16'(-71);
			6110: out = 16'(-47);
			6111: out = 16'(-263);
			6112: out = 16'(2582);
			6113: out = 16'(3591);
			6114: out = 16'(-894);
			6115: out = 16'(-3527);
			6116: out = 16'(4974);
			6117: out = 16'(11440);
			6118: out = 16'(-718);
			6119: out = 16'(-22271);
			6120: out = 16'(-32118);
			6121: out = 16'(-17912);
			6122: out = 16'(3331);
			6123: out = 16'(9670);
			6124: out = 16'(8796);
			6125: out = 16'(14673);
			6126: out = 16'(16392);
			6127: out = 16'(741);
			6128: out = 16'(-13123);
			6129: out = 16'(-18026);
			6130: out = 16'(-12943);
			6131: out = 16'(-7482);
			6132: out = 16'(-781);
			6133: out = 16'(10170);
			6134: out = 16'(16714);
			6135: out = 16'(11037);
			6136: out = 16'(1957);
			6137: out = 16'(-9941);
			6138: out = 16'(-18714);
			6139: out = 16'(-17603);
			6140: out = 16'(3444);
			6141: out = 16'(8984);
			6142: out = 16'(3880);
			6143: out = 16'(-686);
			6144: out = 16'(3437);
			6145: out = 16'(3220);
			6146: out = 16'(45);
			6147: out = 16'(5004);
			6148: out = 16'(18077);
			6149: out = 16'(2307);
			6150: out = 16'(-18838);
			6151: out = 16'(-21920);
			6152: out = 16'(4546);
			6153: out = 16'(9505);
			6154: out = 16'(9771);
			6155: out = 16'(7432);
			6156: out = 16'(7049);
			6157: out = 16'(-902);
			6158: out = 16'(-6733);
			6159: out = 16'(-5812);
			6160: out = 16'(2064);
			6161: out = 16'(8537);
			6162: out = 16'(-6544);
			6163: out = 16'(-15082);
			6164: out = 16'(-2458);
			6165: out = 16'(18436);
			6166: out = 16'(6185);
			6167: out = 16'(138);
			6168: out = 16'(8840);
			6169: out = 16'(16665);
			6170: out = 16'(-5872);
			6171: out = 16'(-23550);
			6172: out = 16'(-18384);
			6173: out = 16'(6214);
			6174: out = 16'(12874);
			6175: out = 16'(19256);
			6176: out = 16'(19502);
			6177: out = 16'(13060);
			6178: out = 16'(-379);
			6179: out = 16'(-22938);
			6180: out = 16'(-30390);
			6181: out = 16'(-25500);
			6182: out = 16'(-2223);
			6183: out = 16'(15754);
			6184: out = 16'(21062);
			6185: out = 16'(13654);
			6186: out = 16'(-2299);
			6187: out = 16'(-7802);
			6188: out = 16'(-5357);
			6189: out = 16'(-523);
			6190: out = 16'(-440);
			6191: out = 16'(1912);
			6192: out = 16'(456);
			6193: out = 16'(308);
			6194: out = 16'(1989);
			6195: out = 16'(1477);
			6196: out = 16'(742);
			6197: out = 16'(1281);
			6198: out = 16'(6066);
			6199: out = 16'(6050);
			6200: out = 16'(-338);
			6201: out = 16'(-14156);
			6202: out = 16'(-15535);
			6203: out = 16'(-990);
			6204: out = 16'(2953);
			6205: out = 16'(-7365);
			6206: out = 16'(-10850);
			6207: out = 16'(-1104);
			6208: out = 16'(5759);
			6209: out = 16'(-3666);
			6210: out = 16'(-1769);
			6211: out = 16'(15217);
			6212: out = 16'(20935);
			6213: out = 16'(-3702);
			6214: out = 16'(-19109);
			6215: out = 16'(-4552);
			6216: out = 16'(9773);
			6217: out = 16'(15751);
			6218: out = 16'(12015);
			6219: out = 16'(3133);
			6220: out = 16'(-9862);
			6221: out = 16'(-26520);
			6222: out = 16'(-16822);
			6223: out = 16'(6802);
			6224: out = 16'(11843);
			6225: out = 16'(4141);
			6226: out = 16'(4152);
			6227: out = 16'(7746);
			6228: out = 16'(780);
			6229: out = 16'(-11003);
			6230: out = 16'(-14190);
			6231: out = 16'(-6999);
			6232: out = 16'(2336);
			6233: out = 16'(12481);
			6234: out = 16'(20138);
			6235: out = 16'(17378);
			6236: out = 16'(2699);
			6237: out = 16'(-16048);
			6238: out = 16'(-14142);
			6239: out = 16'(45);
			6240: out = 16'(9990);
			6241: out = 16'(4386);
			6242: out = 16'(-419);
			6243: out = 16'(-16742);
			6244: out = 16'(-27095);
			6245: out = 16'(-18359);
			6246: out = 16'(3011);
			6247: out = 16'(14268);
			6248: out = 16'(15490);
			6249: out = 16'(11765);
			6250: out = 16'(5785);
			6251: out = 16'(-3500);
			6252: out = 16'(-7414);
			6253: out = 16'(-6421);
			6254: out = 16'(-4675);
			6255: out = 16'(-10171);
			6256: out = 16'(-6560);
			6257: out = 16'(3780);
			6258: out = 16'(9223);
			6259: out = 16'(9290);
			6260: out = 16'(11469);
			6261: out = 16'(10552);
			6262: out = 16'(-712);
			6263: out = 16'(-22402);
			6264: out = 16'(-27906);
			6265: out = 16'(-15204);
			6266: out = 16'(1344);
			6267: out = 16'(14931);
			6268: out = 16'(17782);
			6269: out = 16'(12566);
			6270: out = 16'(3355);
			6271: out = 16'(2315);
			6272: out = 16'(-6462);
			6273: out = 16'(-15515);
			6274: out = 16'(-19178);
			6275: out = 16'(-3758);
			6276: out = 16'(361);
			6277: out = 16'(9092);
			6278: out = 16'(13828);
			6279: out = 16'(11083);
			6280: out = 16'(-1880);
			6281: out = 16'(-6958);
			6282: out = 16'(-3823);
			6283: out = 16'(2656);
			6284: out = 16'(1705);
			6285: out = 16'(2438);
			6286: out = 16'(-498);
			6287: out = 16'(-2493);
			6288: out = 16'(-107);
			6289: out = 16'(3420);
			6290: out = 16'(1615);
			6291: out = 16'(1845);
			6292: out = 16'(8128);
			6293: out = 16'(5135);
			6294: out = 16'(-8772);
			6295: out = 16'(-14251);
			6296: out = 16'(2507);
			6297: out = 16'(13156);
			6298: out = 16'(4547);
			6299: out = 16'(-7292);
			6300: out = 16'(-3200);
			6301: out = 16'(5770);
			6302: out = 16'(4945);
			6303: out = 16'(-323);
			6304: out = 16'(94);
			6305: out = 16'(-1913);
			6306: out = 16'(-6198);
			6307: out = 16'(-6208);
			6308: out = 16'(1455);
			6309: out = 16'(-250);
			6310: out = 16'(1851);
			6311: out = 16'(6995);
			6312: out = 16'(16142);
			6313: out = 16'(10355);
			6314: out = 16'(3301);
			6315: out = 16'(-18165);
			6316: out = 16'(-26721);
			6317: out = 16'(-12041);
			6318: out = 16'(8990);
			6319: out = 16'(13448);
			6320: out = 16'(12983);
			6321: out = 16'(9288);
			6322: out = 16'(-766);
			6323: out = 16'(-21107);
			6324: out = 16'(-19682);
			6325: out = 16'(5820);
			6326: out = 16'(4921);
			6327: out = 16'(3052);
			6328: out = 16'(706);
			6329: out = 16'(5949);
			6330: out = 16'(-1047);
			6331: out = 16'(1578);
			6332: out = 16'(-1282);
			6333: out = 16'(3254);
			6334: out = 16'(4611);
			6335: out = 16'(6030);
			6336: out = 16'(-13421);
			6337: out = 16'(-28597);
			6338: out = 16'(-26342);
			6339: out = 16'(-6626);
			6340: out = 16'(3173);
			6341: out = 16'(14977);
			6342: out = 16'(22846);
			6343: out = 16'(16057);
			6344: out = 16'(-3389);
			6345: out = 16'(-4744);
			6346: out = 16'(7372);
			6347: out = 16'(102);
			6348: out = 16'(-13899);
			6349: out = 16'(-10279);
			6350: out = 16'(11034);
			6351: out = 16'(12547);
			6352: out = 16'(13792);
			6353: out = 16'(7583);
			6354: out = 16'(4349);
			6355: out = 16'(-5839);
			6356: out = 16'(-20179);
			6357: out = 16'(-28780);
			6358: out = 16'(-16735);
			6359: out = 16'(3589);
			6360: out = 16'(19159);
			6361: out = 16'(14094);
			6362: out = 16'(9305);
			6363: out = 16'(7180);
			6364: out = 16'(5419);
			6365: out = 16'(-9369);
			6366: out = 16'(-14560);
			6367: out = 16'(-2171);
			6368: out = 16'(14816);
			6369: out = 16'(12723);
			6370: out = 16'(-893);
			6371: out = 16'(-19417);
			6372: out = 16'(-26704);
			6373: out = 16'(-9987);
			6374: out = 16'(14073);
			6375: out = 16'(14998);
			6376: out = 16'(2289);
			6377: out = 16'(1043);
			6378: out = 16'(13245);
			6379: out = 16'(9416);
			6380: out = 16'(-11176);
			6381: out = 16'(-21343);
			6382: out = 16'(-1844);
			6383: out = 16'(14410);
			6384: out = 16'(8253);
			6385: out = 16'(-1781);
			6386: out = 16'(-5965);
			6387: out = 16'(-9844);
			6388: out = 16'(-14964);
			6389: out = 16'(-8144);
			6390: out = 16'(4590);
			6391: out = 16'(12296);
			6392: out = 16'(10201);
			6393: out = 16'(4925);
			6394: out = 16'(2854);
			6395: out = 16'(-2127);
			6396: out = 16'(-3510);
			6397: out = 16'(1635);
			6398: out = 16'(7487);
			6399: out = 16'(-4923);
			6400: out = 16'(-14432);
			6401: out = 16'(-2928);
			6402: out = 16'(10863);
			6403: out = 16'(6730);
			6404: out = 16'(-8653);
			6405: out = 16'(-6741);
			6406: out = 16'(15304);
			6407: out = 16'(10372);
			6408: out = 16'(-16827);
			6409: out = 16'(-28705);
			6410: out = 16'(-6886);
			6411: out = 16'(19984);
			6412: out = 16'(11612);
			6413: out = 16'(-3342);
			6414: out = 16'(-2099);
			6415: out = 16'(13813);
			6416: out = 16'(1137);
			6417: out = 16'(-17440);
			6418: out = 16'(-11219);
			6419: out = 16'(12456);
			6420: out = 16'(18195);
			6421: out = 16'(3635);
			6422: out = 16'(-11968);
			6423: out = 16'(-16265);
			6424: out = 16'(-1237);
			6425: out = 16'(16829);
			6426: out = 16'(23987);
			6427: out = 16'(13497);
			6428: out = 16'(153);
			6429: out = 16'(-15984);
			6430: out = 16'(-17885);
			6431: out = 16'(-3892);
			6432: out = 16'(1412);
			6433: out = 16'(1279);
			6434: out = 16'(119);
			6435: out = 16'(1884);
			6436: out = 16'(13852);
			6437: out = 16'(8114);
			6438: out = 16'(4793);
			6439: out = 16'(8064);
			6440: out = 16'(6669);
			6441: out = 16'(-9818);
			6442: out = 16'(-21189);
			6443: out = 16'(-11577);
			6444: out = 16'(3486);
			6445: out = 16'(6749);
			6446: out = 16'(631);
			6447: out = 16'(4695);
			6448: out = 16'(14360);
			6449: out = 16'(8927);
			6450: out = 16'(-11898);
			6451: out = 16'(-20971);
			6452: out = 16'(-1722);
			6453: out = 16'(6944);
			6454: out = 16'(5116);
			6455: out = 16'(-6097);
			6456: out = 16'(-9970);
			6457: out = 16'(-934);
			6458: out = 16'(7422);
			6459: out = 16'(10679);
			6460: out = 16'(11885);
			6461: out = 16'(11000);
			6462: out = 16'(8657);
			6463: out = 16'(277);
			6464: out = 16'(-11234);
			6465: out = 16'(-19082);
			6466: out = 16'(-20321);
			6467: out = 16'(-9856);
			6468: out = 16'(4664);
			6469: out = 16'(13200);
			6470: out = 16'(8387);
			6471: out = 16'(6116);
			6472: out = 16'(-298);
			6473: out = 16'(-15929);
			6474: out = 16'(-28802);
			6475: out = 16'(-18967);
			6476: out = 16'(8178);
			6477: out = 16'(22570);
			6478: out = 16'(19279);
			6479: out = 16'(10623);
			6480: out = 16'(1064);
			6481: out = 16'(-11736);
			6482: out = 16'(-23901);
			6483: out = 16'(-24988);
			6484: out = 16'(-9513);
			6485: out = 16'(6210);
			6486: out = 16'(12454);
			6487: out = 16'(2084);
			6488: out = 16'(6475);
			6489: out = 16'(9249);
			6490: out = 16'(4098);
			6491: out = 16'(-3842);
			6492: out = 16'(-3922);
			6493: out = 16'(-9839);
			6494: out = 16'(-17329);
			6495: out = 16'(-4235);
			6496: out = 16'(14701);
			6497: out = 16'(19340);
			6498: out = 16'(9321);
			6499: out = 16'(-627);
			6500: out = 16'(-1582);
			6501: out = 16'(-3406);
			6502: out = 16'(-7873);
			6503: out = 16'(-10648);
			6504: out = 16'(-741);
			6505: out = 16'(-3447);
			6506: out = 16'(-7315);
			6507: out = 16'(700);
			6508: out = 16'(16795);
			6509: out = 16'(21802);
			6510: out = 16'(17592);
			6511: out = 16'(6749);
			6512: out = 16'(-8038);
			6513: out = 16'(-15678);
			6514: out = 16'(-8131);
			6515: out = 16'(-326);
			6516: out = 16'(-7418);
			6517: out = 16'(-17012);
			6518: out = 16'(-2382);
			6519: out = 16'(24094);
			6520: out = 16'(25407);
			6521: out = 16'(8095);
			6522: out = 16'(-9375);
			6523: out = 16'(-11737);
			6524: out = 16'(-7992);
			6525: out = 16'(674);
			6526: out = 16'(3);
			6527: out = 16'(3704);
			6528: out = 16'(4914);
			6529: out = 16'(-4291);
			6530: out = 16'(-9436);
			6531: out = 16'(3500);
			6532: out = 16'(17751);
			6533: out = 16'(8747);
			6534: out = 16'(2409);
			6535: out = 16'(-539);
			6536: out = 16'(-1949);
			6537: out = 16'(-11392);
			6538: out = 16'(-5051);
			6539: out = 16'(2433);
			6540: out = 16'(3165);
			6541: out = 16'(-4715);
			6542: out = 16'(-507);
			6543: out = 16'(3795);
			6544: out = 16'(3355);
			6545: out = 16'(-1431);
			6546: out = 16'(1716);
			6547: out = 16'(7218);
			6548: out = 16'(6698);
			6549: out = 16'(-2596);
			6550: out = 16'(-12027);
			6551: out = 16'(-8656);
			6552: out = 16'(5409);
			6553: out = 16'(18220);
			6554: out = 16'(17010);
			6555: out = 16'(5773);
			6556: out = 16'(-16156);
			6557: out = 16'(-25687);
			6558: out = 16'(-9146);
			6559: out = 16'(752);
			6560: out = 16'(-3046);
			6561: out = 16'(-6393);
			6562: out = 16'(5038);
			6563: out = 16'(16338);
			6564: out = 16'(3869);
			6565: out = 16'(-18111);
			6566: out = 16'(-21589);
			6567: out = 16'(-807);
			6568: out = 16'(12200);
			6569: out = 16'(6734);
			6570: out = 16'(189);
			6571: out = 16'(-1686);
			6572: out = 16'(10356);
			6573: out = 16'(4031);
			6574: out = 16'(-9168);
			6575: out = 16'(-9734);
			6576: out = 16'(9075);
			6577: out = 16'(8976);
			6578: out = 16'(-5417);
			6579: out = 16'(-11523);
			6580: out = 16'(-8167);
			6581: out = 16'(-447);
			6582: out = 16'(2460);
			6583: out = 16'(9285);
			6584: out = 16'(14138);
			6585: out = 16'(17836);
			6586: out = 16'(5422);
			6587: out = 16'(-9119);
			6588: out = 16'(-4871);
			6589: out = 16'(4802);
			6590: out = 16'(5556);
			6591: out = 16'(-3022);
			6592: out = 16'(-10864);
			6593: out = 16'(-5550);
			6594: out = 16'(1702);
			6595: out = 16'(6698);
			6596: out = 16'(9033);
			6597: out = 16'(12959);
			6598: out = 16'(1938);
			6599: out = 16'(-12477);
			6600: out = 16'(-17930);
			6601: out = 16'(-6701);
			6602: out = 16'(-1060);
			6603: out = 16'(3385);
			6604: out = 16'(12402);
			6605: out = 16'(24041);
			6606: out = 16'(8442);
			6607: out = 16'(-13053);
			6608: out = 16'(-24143);
			6609: out = 16'(-8401);
			6610: out = 16'(-12207);
			6611: out = 16'(-7587);
			6612: out = 16'(6379);
			6613: out = 16'(18148);
			6614: out = 16'(14134);
			6615: out = 16'(8456);
			6616: out = 16'(351);
			6617: out = 16'(-8657);
			6618: out = 16'(-7161);
			6619: out = 16'(-3217);
			6620: out = 16'(-2828);
			6621: out = 16'(-6207);
			6622: out = 16'(356);
			6623: out = 16'(1683);
			6624: out = 16'(1559);
			6625: out = 16'(-310);
			6626: out = 16'(-972);
			6627: out = 16'(9324);
			6628: out = 16'(12908);
			6629: out = 16'(-928);
			6630: out = 16'(-26746);
			6631: out = 16'(-15715);
			6632: out = 16'(1080);
			6633: out = 16'(1638);
			6634: out = 16'(-9889);
			6635: out = 16'(9074);
			6636: out = 16'(17916);
			6637: out = 16'(13376);
			6638: out = 16'(2577);
			6639: out = 16'(4968);
			6640: out = 16'(-5248);
			6641: out = 16'(-17779);
			6642: out = 16'(-21123);
			6643: out = 16'(-12261);
			6644: out = 16'(7068);
			6645: out = 16'(14994);
			6646: out = 16'(13556);
			6647: out = 16'(7712);
			6648: out = 16'(16904);
			6649: out = 16'(5861);
			6650: out = 16'(-17017);
			6651: out = 16'(-28469);
			6652: out = 16'(-13674);
			6653: out = 16'(1891);
			6654: out = 16'(7060);
			6655: out = 16'(10345);
			6656: out = 16'(12917);
			6657: out = 16'(1947);
			6658: out = 16'(-12785);
			6659: out = 16'(-13094);
			6660: out = 16'(7307);
			6661: out = 16'(12289);
			6662: out = 16'(5469);
			6663: out = 16'(179);
			6664: out = 16'(1703);
			6665: out = 16'(4797);
			6666: out = 16'(2312);
			6667: out = 16'(783);
			6668: out = 16'(4333);
			6669: out = 16'(-3861);
			6670: out = 16'(-13619);
			6671: out = 16'(-12671);
			6672: out = 16'(2835);
			6673: out = 16'(-6869);
			6674: out = 16'(-4805);
			6675: out = 16'(6797);
			6676: out = 16'(20021);
			6677: out = 16'(8930);
			6678: out = 16'(7697);
			6679: out = 16'(3644);
			6680: out = 16'(965);
			6681: out = 16'(-5604);
			6682: out = 16'(-4356);
			6683: out = 16'(-8142);
			6684: out = 16'(-7938);
			6685: out = 16'(707);
			6686: out = 16'(15479);
			6687: out = 16'(15168);
			6688: out = 16'(9511);
			6689: out = 16'(6382);
			6690: out = 16'(1296);
			6691: out = 16'(-17684);
			6692: out = 16'(-30714);
			6693: out = 16'(-23185);
			6694: out = 16'(-4523);
			6695: out = 16'(4844);
			6696: out = 16'(8209);
			6697: out = 16'(17994);
			6698: out = 16'(23424);
			6699: out = 16'(21515);
			6700: out = 16'(1628);
			6701: out = 16'(-24093);
			6702: out = 16'(-29792);
			6703: out = 16'(-22674);
			6704: out = 16'(-6320);
			6705: out = 16'(7729);
			6706: out = 16'(18616);
			6707: out = 16'(18377);
			6708: out = 16'(10859);
			6709: out = 16'(-884);
			6710: out = 16'(-10294);
			6711: out = 16'(-8876);
			6712: out = 16'(-5929);
			6713: out = 16'(-4587);
			6714: out = 16'(-3243);
			6715: out = 16'(7548);
			6716: out = 16'(10992);
			6717: out = 16'(9076);
			6718: out = 16'(1150);
			6719: out = 16'(1123);
			6720: out = 16'(-4236);
			6721: out = 16'(1548);
			6722: out = 16'(3636);
			6723: out = 16'(1930);
			6724: out = 16'(-22035);
			6725: out = 16'(-11272);
			6726: out = 16'(11756);
			6727: out = 16'(13270);
			6728: out = 16'(2332);
			6729: out = 16'(1640);
			6730: out = 16'(4864);
			6731: out = 16'(-400);
			6732: out = 16'(-3944);
			6733: out = 16'(-2418);
			6734: out = 16'(-820);
			6735: out = 16'(-6811);
			6736: out = 16'(-8569);
			6737: out = 16'(-3558);
			6738: out = 16'(7401);
			6739: out = 16'(9823);
			6740: out = 16'(1574);
			6741: out = 16'(-3520);
			6742: out = 16'(-7703);
			6743: out = 16'(-10080);
			6744: out = 16'(-6731);
			6745: out = 16'(2741);
			6746: out = 16'(8777);
			6747: out = 16'(8268);
			6748: out = 16'(7898);
			6749: out = 16'(4090);
			6750: out = 16'(2017);
			6751: out = 16'(-11063);
			6752: out = 16'(-24085);
			6753: out = 16'(-13840);
			6754: out = 16'(4856);
			6755: out = 16'(12205);
			6756: out = 16'(6352);
			6757: out = 16'(-3989);
			6758: out = 16'(3206);
			6759: out = 16'(1056);
			6760: out = 16'(-3906);
			6761: out = 16'(7093);
			6762: out = 16'(17698);
			6763: out = 16'(13951);
			6764: out = 16'(-4863);
			6765: out = 16'(-18168);
			6766: out = 16'(-23806);
			6767: out = 16'(-13678);
			6768: out = 16'(-7602);
			6769: out = 16'(-814);
			6770: out = 16'(10245);
			6771: out = 16'(23201);
			6772: out = 16'(14320);
			6773: out = 16'(-2988);
			6774: out = 16'(-7303);
			6775: out = 16'(8094);
			6776: out = 16'(7519);
			6777: out = 16'(-8700);
			6778: out = 16'(-14619);
			6779: out = 16'(-271);
			6780: out = 16'(9900);
			6781: out = 16'(7107);
			6782: out = 16'(7248);
			6783: out = 16'(3686);
			6784: out = 16'(7509);
			6785: out = 16'(3239);
			6786: out = 16'(-7807);
			6787: out = 16'(-27985);
			6788: out = 16'(-18828);
			6789: out = 16'(1262);
			6790: out = 16'(15943);
			6791: out = 16'(19497);
			6792: out = 16'(17187);
			6793: out = 16'(2287);
			6794: out = 16'(-12063);
			6795: out = 16'(-12788);
			6796: out = 16'(-1275);
			6797: out = 16'(1893);
			6798: out = 16'(24);
			6799: out = 16'(2456);
			6800: out = 16'(11659);
			6801: out = 16'(-533);
			6802: out = 16'(-19258);
			6803: out = 16'(-18789);
			6804: out = 16'(733);
			6805: out = 16'(15310);
			6806: out = 16'(12422);
			6807: out = 16'(3187);
			6808: out = 16'(-4002);
			6809: out = 16'(-8308);
			6810: out = 16'(-8625);
			6811: out = 16'(-164);
			6812: out = 16'(14265);
			6813: out = 16'(5579);
			6814: out = 16'(-10199);
			6815: out = 16'(-15222);
			6816: out = 16'(2620);
			6817: out = 16'(-320);
			6818: out = 16'(-5532);
			6819: out = 16'(-8793);
			6820: out = 16'(-409);
			6821: out = 16'(9185);
			6822: out = 16'(19192);
			6823: out = 16'(17257);
			6824: out = 16'(7802);
			6825: out = 16'(-8442);
			6826: out = 16'(-10319);
			6827: out = 16'(-12194);
			6828: out = 16'(-16775);
			6829: out = 16'(-12599);
			6830: out = 16'(-1938);
			6831: out = 16'(7866);
			6832: out = 16'(14816);
			6833: out = 16'(23676);
			6834: out = 16'(17081);
			6835: out = 16'(5445);
			6836: out = 16'(-7081);
			6837: out = 16'(-9824);
			6838: out = 16'(-22926);
			6839: out = 16'(-16700);
			6840: out = 16'(-991);
			6841: out = 16'(7919);
			6842: out = 16'(7120);
			6843: out = 16'(5107);
			6844: out = 16'(5367);
			6845: out = 16'(3571);
			6846: out = 16'(-1985);
			6847: out = 16'(-5277);
			6848: out = 16'(407);
			6849: out = 16'(5814);
			6850: out = 16'(-1398);
			6851: out = 16'(-4003);
			6852: out = 16'(-3722);
			6853: out = 16'(-4411);
			6854: out = 16'(-9879);
			6855: out = 16'(8001);
			6856: out = 16'(21708);
			6857: out = 16'(17466);
			6858: out = 16'(-2516);
			6859: out = 16'(-19015);
			6860: out = 16'(-18471);
			6861: out = 16'(-4841);
			6862: out = 16'(1981);
			6863: out = 16'(5622);
			6864: out = 16'(-3672);
			6865: out = 16'(-8685);
			6866: out = 16'(-2704);
			6867: out = 16'(13482);
			6868: out = 16'(13069);
			6869: out = 16'(6796);
			6870: out = 16'(485);
			6871: out = 16'(68);
			6872: out = 16'(-5715);
			6873: out = 16'(-2477);
			6874: out = 16'(8092);
			6875: out = 16'(16211);
			6876: out = 16'(146);
			6877: out = 16'(-13596);
			6878: out = 16'(-19336);
			6879: out = 16'(-13616);
			6880: out = 16'(-6328);
			6881: out = 16'(6541);
			6882: out = 16'(16153);
			6883: out = 16'(19421);
			6884: out = 16'(13417);
			6885: out = 16'(3289);
			6886: out = 16'(-9084);
			6887: out = 16'(-11155);
			6888: out = 16'(202);
			6889: out = 16'(3048);
			6890: out = 16'(-7208);
			6891: out = 16'(-13614);
			6892: out = 16'(-599);
			6893: out = 16'(7395);
			6894: out = 16'(4950);
			6895: out = 16'(-1030);
			6896: out = 16'(3359);
			6897: out = 16'(12809);
			6898: out = 16'(14868);
			6899: out = 16'(5457);
			6900: out = 16'(-8290);
			6901: out = 16'(-23439);
			6902: out = 16'(-24023);
			6903: out = 16'(-14247);
			6904: out = 16'(-274);
			6905: out = 16'(15341);
			6906: out = 16'(16580);
			6907: out = 16'(15488);
			6908: out = 16'(11819);
			6909: out = 16'(6412);
			6910: out = 16'(-15490);
			6911: out = 16'(-21803);
			6912: out = 16'(-12625);
			6913: out = 16'(-5217);
			6914: out = 16'(-5213);
			6915: out = 16'(-2536);
			6916: out = 16'(10712);
			6917: out = 16'(23698);
			6918: out = 16'(22182);
			6919: out = 16'(8991);
			6920: out = 16'(-11443);
			6921: out = 16'(-28539);
			6922: out = 16'(-22663);
			6923: out = 16'(-19208);
			6924: out = 16'(-10404);
			6925: out = 16'(-1550);
			6926: out = 16'(6294);
			6927: out = 16'(10487);
			6928: out = 16'(13679);
			6929: out = 16'(7435);
			6930: out = 16'(-2574);
			6931: out = 16'(-12653);
			6932: out = 16'(-411);
			6933: out = 16'(7985);
			6934: out = 16'(-719);
			6935: out = 16'(-3393);
			6936: out = 16'(-300);
			6937: out = 16'(1017);
			6938: out = 16'(-5131);
			6939: out = 16'(-2053);
			6940: out = 16'(4699);
			6941: out = 16'(8550);
			6942: out = 16'(2112);
			6943: out = 16'(-5095);
			6944: out = 16'(-10765);
			6945: out = 16'(-5890);
			6946: out = 16'(5334);
			6947: out = 16'(15500);
			6948: out = 16'(10744);
			6949: out = 16'(1077);
			6950: out = 16'(-4816);
			6951: out = 16'(1762);
			6952: out = 16'(796);
			6953: out = 16'(2035);
			6954: out = 16'(-3391);
			6955: out = 16'(-3946);
			6956: out = 16'(7187);
			6957: out = 16'(7443);
			6958: out = 16'(-6018);
			6959: out = 16'(-10231);
			6960: out = 16'(13917);
			6961: out = 16'(12944);
			6962: out = 16'(-8887);
			6963: out = 16'(-26163);
			6964: out = 16'(-6427);
			6965: out = 16'(8687);
			6966: out = 16'(7308);
			6967: out = 16'(1312);
			6968: out = 16'(13914);
			6969: out = 16'(11008);
			6970: out = 16'(8272);
			6971: out = 16'(-8095);
			6972: out = 16'(-22166);
			6973: out = 16'(-22057);
			6974: out = 16'(190);
			6975: out = 16'(11999);
			6976: out = 16'(7107);
			6977: out = 16'(1222);
			6978: out = 16'(2034);
			6979: out = 16'(4737);
			6980: out = 16'(5866);
			6981: out = 16'(12980);
			6982: out = 16'(1813);
			6983: out = 16'(1503);
			6984: out = 16'(5197);
			6985: out = 16'(2585);
			6986: out = 16'(-20109);
			6987: out = 16'(-24843);
			6988: out = 16'(-5943);
			6989: out = 16'(9659);
			6990: out = 16'(2626);
			6991: out = 16'(-3236);
			6992: out = 16'(9063);
			6993: out = 16'(20937);
			6994: out = 16'(1011);
			6995: out = 16'(-17724);
			6996: out = 16'(-21264);
			6997: out = 16'(-5426);
			6998: out = 16'(-387);
			6999: out = 16'(11333);
			7000: out = 16'(14646);
			7001: out = 16'(13672);
			7002: out = 16'(5237);
			7003: out = 16'(8852);
			7004: out = 16'(-837);
			7005: out = 16'(-17576);
			7006: out = 16'(-28392);
			7007: out = 16'(-21350);
			7008: out = 16'(-5184);
			7009: out = 16'(5112);
			7010: out = 16'(4772);
			7011: out = 16'(1436);
			7012: out = 16'(10233);
			7013: out = 16'(19198);
			7014: out = 16'(12191);
			7015: out = 16'(-10703);
			7016: out = 16'(-11950);
			7017: out = 16'(1477);
			7018: out = 16'(3644);
			7019: out = 16'(-16019);
			7020: out = 16'(-22255);
			7021: out = 16'(-10532);
			7022: out = 16'(5399);
			7023: out = 16'(8114);
			7024: out = 16'(9771);
			7025: out = 16'(11263);
			7026: out = 16'(9356);
			7027: out = 16'(928);
			7028: out = 16'(-2105);
			7029: out = 16'(-1370);
			7030: out = 16'(273);
			7031: out = 16'(-1799);
			7032: out = 16'(-871);
			7033: out = 16'(4847);
			7034: out = 16'(9727);
			7035: out = 16'(6667);
			7036: out = 16'(-1302);
			7037: out = 16'(-10618);
			7038: out = 16'(-13466);
			7039: out = 16'(-7064);
			7040: out = 16'(5964);
			7041: out = 16'(13975);
			7042: out = 16'(12924);
			7043: out = 16'(4748);
			7044: out = 16'(-1018);
			7045: out = 16'(3280);
			7046: out = 16'(4143);
			7047: out = 16'(-5291);
			7048: out = 16'(-16481);
			7049: out = 16'(-5684);
			7050: out = 16'(2377);
			7051: out = 16'(6929);
			7052: out = 16'(10843);
			7053: out = 16'(17785);
			7054: out = 16'(5590);
			7055: out = 16'(-11447);
			7056: out = 16'(-20284);
			7057: out = 16'(-9264);
			7058: out = 16'(1695);
			7059: out = 16'(12005);
			7060: out = 16'(17109);
			7061: out = 16'(12413);
			7062: out = 16'(-5776);
			7063: out = 16'(-13696);
			7064: out = 16'(-745);
			7065: out = 16'(12644);
			7066: out = 16'(4787);
			7067: out = 16'(-12911);
			7068: out = 16'(-16067);
			7069: out = 16'(-4662);
			7070: out = 16'(1320);
			7071: out = 16'(-13326);
			7072: out = 16'(-11281);
			7073: out = 16'(9785);
			7074: out = 16'(17460);
			7075: out = 16'(10524);
			7076: out = 16'(7951);
			7077: out = 16'(10422);
			7078: out = 16'(-1358);
			7079: out = 16'(-12459);
			7080: out = 16'(-26011);
			7081: out = 16'(-22662);
			7082: out = 16'(-4933);
			7083: out = 16'(17168);
			7084: out = 16'(14120);
			7085: out = 16'(3228);
			7086: out = 16'(-1470);
			7087: out = 16'(11725);
			7088: out = 16'(1833);
			7089: out = 16'(-16183);
			7090: out = 16'(-25207);
			7091: out = 16'(-2973);
			7092: out = 16'(49);
			7093: out = 16'(3188);
			7094: out = 16'(6890);
			7095: out = 16'(12310);
			7096: out = 16'(13175);
			7097: out = 16'(13265);
			7098: out = 16'(904);
			7099: out = 16'(-23452);
			7100: out = 16'(-18124);
			7101: out = 16'(-7230);
			7102: out = 16'(-374);
			7103: out = 16'(-5502);
			7104: out = 16'(-2984);
			7105: out = 16'(3714);
			7106: out = 16'(16148);
			7107: out = 16'(11800);
			7108: out = 16'(-15465);
			7109: out = 16'(-20453);
			7110: out = 16'(434);
			7111: out = 16'(16554);
			7112: out = 16'(8503);
			7113: out = 16'(-8562);
			7114: out = 16'(-7747);
			7115: out = 16'(3824);
			7116: out = 16'(4538);
			7117: out = 16'(2862);
			7118: out = 16'(9065);
			7119: out = 16'(14211);
			7120: out = 16'(3405);
			7121: out = 16'(-18052);
			7122: out = 16'(-30231);
			7123: out = 16'(-22336);
			7124: out = 16'(-2311);
			7125: out = 16'(17811);
			7126: out = 16'(16686);
			7127: out = 16'(10252);
			7128: out = 16'(3743);
			7129: out = 16'(482);
			7130: out = 16'(-5967);
			7131: out = 16'(-7100);
			7132: out = 16'(-215);
			7133: out = 16'(9561);
			7134: out = 16'(9629);
			7135: out = 16'(8094);
			7136: out = 16'(7946);
			7137: out = 16'(6172);
			7138: out = 16'(-1394);
			7139: out = 16'(-18463);
			7140: out = 16'(-29425);
			7141: out = 16'(-20889);
			7142: out = 16'(3206);
			7143: out = 16'(11963);
			7144: out = 16'(11897);
			7145: out = 16'(13643);
			7146: out = 16'(18323);
			7147: out = 16'(5556);
			7148: out = 16'(-6756);
			7149: out = 16'(-6662);
			7150: out = 16'(4272);
			7151: out = 16'(-563);
			7152: out = 16'(-14343);
			7153: out = 16'(-18798);
			7154: out = 16'(3775);
			7155: out = 16'(8992);
			7156: out = 16'(17584);
			7157: out = 16'(9190);
			7158: out = 16'(-3595);
			7159: out = 16'(-5496);
			7160: out = 16'(4114);
			7161: out = 16'(-1099);
			7162: out = 16'(-16536);
			7163: out = 16'(-12270);
			7164: out = 16'(-3265);
			7165: out = 16'(520);
			7166: out = 16'(-1628);
			7167: out = 16'(9817);
			7168: out = 16'(12294);
			7169: out = 16'(17709);
			7170: out = 16'(14923);
			7171: out = 16'(7141);
			7172: out = 16'(-17806);
			7173: out = 16'(-26701);
			7174: out = 16'(-21063);
			7175: out = 16'(-6870);
			7176: out = 16'(3770);
			7177: out = 16'(16749);
			7178: out = 16'(19360);
			7179: out = 16'(11045);
			7180: out = 16'(-414);
			7181: out = 16'(-5765);
			7182: out = 16'(-6877);
			7183: out = 16'(-10185);
			7184: out = 16'(-19479);
			7185: out = 16'(-8805);
			7186: out = 16'(4123);
			7187: out = 16'(6284);
			7188: out = 16'(-4461);
			7189: out = 16'(-3997);
			7190: out = 16'(3352);
			7191: out = 16'(12090);
			7192: out = 16'(7114);
			7193: out = 16'(3624);
			7194: out = 16'(-5139);
			7195: out = 16'(3882);
			7196: out = 16'(12066);
			7197: out = 16'(-3772);
			7198: out = 16'(-26103);
			7199: out = 16'(-17061);
			7200: out = 16'(12652);
			7201: out = 16'(10884);
			7202: out = 16'(-4681);
			7203: out = 16'(-5087);
			7204: out = 16'(10960);
			7205: out = 16'(5475);
			7206: out = 16'(2836);
			7207: out = 16'(-6353);
			7208: out = 16'(-1606);
			7209: out = 16'(5537);
			7210: out = 16'(20198);
			7211: out = 16'(10307);
			7212: out = 16'(2493);
			7213: out = 16'(167);
			7214: out = 16'(7948);
			7215: out = 16'(-14301);
			7216: out = 16'(-28410);
			7217: out = 16'(-15920);
			7218: out = 16'(10450);
			7219: out = 16'(11327);
			7220: out = 16'(6952);
			7221: out = 16'(4101);
			7222: out = 16'(295);
			7223: out = 16'(-4075);
			7224: out = 16'(399);
			7225: out = 16'(4659);
			7226: out = 16'(-1622);
			7227: out = 16'(6746);
			7228: out = 16'(7017);
			7229: out = 16'(-2034);
			7230: out = 16'(-15257);
			7231: out = 16'(11821);
			7232: out = 16'(14006);
			7233: out = 16'(2163);
			7234: out = 16'(-14811);
			7235: out = 16'(-7393);
			7236: out = 16'(-3112);
			7237: out = 16'(2228);
			7238: out = 16'(-2623);
			7239: out = 16'(-5638);
			7240: out = 16'(-2750);
			7241: out = 16'(14610);
			7242: out = 16'(16268);
			7243: out = 16'(2158);
			7244: out = 16'(-5553);
			7245: out = 16'(9340);
			7246: out = 16'(11976);
			7247: out = 16'(-11343);
			7248: out = 16'(-27117);
			7249: out = 16'(-14339);
			7250: out = 16'(3509);
			7251: out = 16'(2314);
			7252: out = 16'(14631);
			7253: out = 16'(18132);
			7254: out = 16'(15858);
			7255: out = 16'(2510);
			7256: out = 16'(-12777);
			7257: out = 16'(-27791);
			7258: out = 16'(-29138);
			7259: out = 16'(-17069);
			7260: out = 16'(16254);
			7261: out = 16'(24095);
			7262: out = 16'(24514);
			7263: out = 16'(16619);
			7264: out = 16'(9486);
			7265: out = 16'(-21160);
			7266: out = 16'(-30342);
			7267: out = 16'(-23433);
			7268: out = 16'(-4858);
			7269: out = 16'(759);
			7270: out = 16'(10586);
			7271: out = 16'(9977);
			7272: out = 16'(8039);
			7273: out = 16'(14364);
			7274: out = 16'(7792);
			7275: out = 16'(-13476);
			7276: out = 16'(-25994);
			7277: out = 16'(249);
			7278: out = 16'(3373);
			7279: out = 16'(-4480);
			7280: out = 16'(-8027);
			7281: out = 16'(6897);
			7282: out = 16'(16379);
			7283: out = 16'(10336);
			7284: out = 16'(-3161);
			7285: out = 16'(-6180);
			7286: out = 16'(1741);
			7287: out = 16'(1059);
			7288: out = 16'(-5042);
			7289: out = 16'(-2566);
			7290: out = 16'(-725);
			7291: out = 16'(2314);
			7292: out = 16'(-5788);
			7293: out = 16'(-10513);
			7294: out = 16'(1941);
			7295: out = 16'(15385);
			7296: out = 16'(11936);
			7297: out = 16'(-2019);
			7298: out = 16'(-6355);
			7299: out = 16'(-3760);
			7300: out = 16'(2844);
			7301: out = 16'(2698);
			7302: out = 16'(2821);
			7303: out = 16'(3500);
			7304: out = 16'(9749);
			7305: out = 16'(4196);
			7306: out = 16'(-10934);
			7307: out = 16'(-12654);
			7308: out = 16'(-4750);
			7309: out = 16'(3485);
			7310: out = 16'(5420);
			7311: out = 16'(7904);
			7312: out = 16'(14084);
			7313: out = 16'(14732);
			7314: out = 16'(5978);
			7315: out = 16'(-4629);
			7316: out = 16'(-17590);
			7317: out = 16'(-19662);
			7318: out = 16'(-10284);
			7319: out = 16'(797);
			7320: out = 16'(7272);
			7321: out = 16'(6914);
			7322: out = 16'(7080);
			7323: out = 16'(8509);
			7324: out = 16'(6593);
			7325: out = 16'(-336);
			7326: out = 16'(-4238);
			7327: out = 16'(-3131);
			7328: out = 16'(114);
			7329: out = 16'(-10326);
			7330: out = 16'(-13781);
			7331: out = 16'(-2429);
			7332: out = 16'(6499);
			7333: out = 16'(6718);
			7334: out = 16'(2283);
			7335: out = 16'(3511);
			7336: out = 16'(6741);
			7337: out = 16'(2213);
			7338: out = 16'(-1725);
			7339: out = 16'(4870);
			7340: out = 16'(13259);
			7341: out = 16'(-9091);
			7342: out = 16'(-29149);
			7343: out = 16'(-21825);
			7344: out = 16'(15818);
			7345: out = 16'(27754);
			7346: out = 16'(11008);
			7347: out = 16'(-2525);
			7348: out = 16'(2935);
			7349: out = 16'(9027);
			7350: out = 16'(-959);
			7351: out = 16'(-20938);
			7352: out = 16'(-25550);
			7353: out = 16'(-10588);
			7354: out = 16'(7232);
			7355: out = 16'(5014);
			7356: out = 16'(753);
			7357: out = 16'(4055);
			7358: out = 16'(14665);
			7359: out = 16'(2157);
			7360: out = 16'(-11634);
			7361: out = 16'(-6842);
			7362: out = 16'(10201);
			7363: out = 16'(7469);
			7364: out = 16'(-5481);
			7365: out = 16'(-13189);
			7366: out = 16'(-11572);
			7367: out = 16'(-819);
			7368: out = 16'(8300);
			7369: out = 16'(8883);
			7370: out = 16'(2168);
			7371: out = 16'(2065);
			7372: out = 16'(7299);
			7373: out = 16'(4619);
			7374: out = 16'(-10584);
			7375: out = 16'(-23763);
			7376: out = 16'(-13127);
			7377: out = 16'(6683);
			7378: out = 16'(7449);
			7379: out = 16'(1243);
			7380: out = 16'(4118);
			7381: out = 16'(17202);
			7382: out = 16'(15627);
			7383: out = 16'(-1685);
			7384: out = 16'(-21692);
			7385: out = 16'(-17502);
			7386: out = 16'(3668);
			7387: out = 16'(14662);
			7388: out = 16'(6738);
			7389: out = 16'(219);
			7390: out = 16'(-2504);
			7391: out = 16'(-4646);
			7392: out = 16'(-12053);
			7393: out = 16'(-3553);
			7394: out = 16'(7913);
			7395: out = 16'(6449);
			7396: out = 16'(150);
			7397: out = 16'(7528);
			7398: out = 16'(19038);
			7399: out = 16'(14001);
			7400: out = 16'(-1975);
			7401: out = 16'(-15456);
			7402: out = 16'(-11904);
			7403: out = 16'(-2309);
			7404: out = 16'(-5);
			7405: out = 16'(-869);
			7406: out = 16'(6504);
			7407: out = 16'(14783);
			7408: out = 16'(12255);
			7409: out = 16'(1248);
			7410: out = 16'(-3285);
			7411: out = 16'(3289);
			7412: out = 16'(9957);
			7413: out = 16'(7820);
			7414: out = 16'(-7108);
			7415: out = 16'(-22045);
			7416: out = 16'(-19458);
			7417: out = 16'(-2177);
			7418: out = 16'(8955);
			7419: out = 16'(3941);
			7420: out = 16'(3142);
			7421: out = 16'(17746);
			7422: out = 16'(17622);
			7423: out = 16'(-5185);
			7424: out = 16'(-26054);
			7425: out = 16'(-13624);
			7426: out = 16'(-1493);
			7427: out = 16'(-10128);
			7428: out = 16'(-20052);
			7429: out = 16'(4047);
			7430: out = 16'(25148);
			7431: out = 16'(23885);
			7432: out = 16'(4284);
			7433: out = 16'(-11080);
			7434: out = 16'(-6520);
			7435: out = 16'(-11677);
			7436: out = 16'(-26098);
			7437: out = 16'(-26583);
			7438: out = 16'(8000);
			7439: out = 16'(23740);
			7440: out = 16'(12636);
			7441: out = 16'(-804);
			7442: out = 16'(588);
			7443: out = 16'(1725);
			7444: out = 16'(-1048);
			7445: out = 16'(-4750);
			7446: out = 16'(-865);
			7447: out = 16'(-293);
			7448: out = 16'(1045);
			7449: out = 16'(-3429);
			7450: out = 16'(-12340);
			7451: out = 16'(-1456);
			7452: out = 16'(2346);
			7453: out = 16'(984);
			7454: out = 16'(-594);
			7455: out = 16'(4588);
			7456: out = 16'(9652);
			7457: out = 16'(9865);
			7458: out = 16'(1663);
			7459: out = 16'(-6398);
			7460: out = 16'(-15261);
			7461: out = 16'(-11010);
			7462: out = 16'(2124);
			7463: out = 16'(16303);
			7464: out = 16'(7191);
			7465: out = 16'(31);
			7466: out = 16'(-7047);
			7467: out = 16'(-8450);
			7468: out = 16'(-15154);
			7469: out = 16'(1224);
			7470: out = 16'(15032);
			7471: out = 16'(13735);
			7472: out = 16'(1454);
			7473: out = 16'(4076);
			7474: out = 16'(3323);
			7475: out = 16'(-4840);
			7476: out = 16'(-12619);
			7477: out = 16'(-8734);
			7478: out = 16'(-10867);
			7479: out = 16'(-9454);
			7480: out = 16'(13858);
			7481: out = 16'(25678);
			7482: out = 16'(12454);
			7483: out = 16'(-7536);
			7484: out = 16'(-8789);
			7485: out = 16'(-5377);
			7486: out = 16'(-14331);
			7487: out = 16'(-20798);
			7488: out = 16'(2431);
			7489: out = 16'(3020);
			7490: out = 16'(11053);
			7491: out = 16'(11599);
			7492: out = 16'(13109);
			7493: out = 16'(6830);
			7494: out = 16'(2661);
			7495: out = 16'(-7965);
			7496: out = 16'(-9637);
			7497: out = 16'(6139);
			7498: out = 16'(7286);
			7499: out = 16'(-4936);
			7500: out = 16'(-13831);
			7501: out = 16'(-4007);
			7502: out = 16'(2417);
			7503: out = 16'(2816);
			7504: out = 16'(5452);
			7505: out = 16'(17266);
			7506: out = 16'(19200);
			7507: out = 16'(10163);
			7508: out = 16'(-7922);
			7509: out = 16'(-22805);
			7510: out = 16'(-23000);
			7511: out = 16'(-15503);
			7512: out = 16'(-4204);
			7513: out = 16'(7386);
			7514: out = 16'(10998);
			7515: out = 16'(12048);
			7516: out = 16'(11016);
			7517: out = 16'(9771);
			7518: out = 16'(-622);
			7519: out = 16'(3126);
			7520: out = 16'(-2610);
			7521: out = 16'(-10142);
			7522: out = 16'(-12667);
			7523: out = 16'(-3425);
			7524: out = 16'(787);
			7525: out = 16'(4210);
			7526: out = 16'(8567);
			7527: out = 16'(3949);
			7528: out = 16'(-327);
			7529: out = 16'(-1357);
			7530: out = 16'(872);
			7531: out = 16'(11042);
			7532: out = 16'(-2345);
			7533: out = 16'(-8144);
			7534: out = 16'(-988);
			7535: out = 16'(3812);
			7536: out = 16'(-12037);
			7537: out = 16'(-13296);
			7538: out = 16'(8865);
			7539: out = 16'(16417);
			7540: out = 16'(10397);
			7541: out = 16'(-14041);
			7542: out = 16'(-22715);
			7543: out = 16'(-8316);
			7544: out = 16'(10273);
			7545: out = 16'(241);
			7546: out = 16'(-6630);
			7547: out = 16'(4756);
			7548: out = 16'(12596);
			7549: out = 16'(5663);
			7550: out = 16'(-5827);
			7551: out = 16'(-10674);
			7552: out = 16'(-4396);
			7553: out = 16'(-4998);
			7554: out = 16'(871);
			7555: out = 16'(7231);
			7556: out = 16'(8207);
			7557: out = 16'(10588);
			7558: out = 16'(14411);
			7559: out = 16'(-2254);
			7560: out = 16'(-29392);
			7561: out = 16'(-26649);
			7562: out = 16'(-2096);
			7563: out = 16'(11937);
			7564: out = 16'(-298);
			7565: out = 16'(11813);
			7566: out = 16'(17331);
			7567: out = 16'(16592);
			7568: out = 16'(1988);
			7569: out = 16'(-2850);
			7570: out = 16'(-9118);
			7571: out = 16'(-4593);
			7572: out = 16'(-2414);
			7573: out = 16'(-4202);
			7574: out = 16'(-9020);
			7575: out = 16'(-7071);
			7576: out = 16'(-3128);
			7577: out = 16'(1137);
			7578: out = 16'(9332);
			7579: out = 16'(11891);
			7580: out = 16'(1877);
			7581: out = 16'(-11713);
			7582: out = 16'(1962);
			7583: out = 16'(7377);
			7584: out = 16'(-6656);
			7585: out = 16'(-27177);
			7586: out = 16'(-6019);
			7587: out = 16'(3367);
			7588: out = 16'(7857);
			7589: out = 16'(15476);
			7590: out = 16'(25801);
			7591: out = 16'(15969);
			7592: out = 16'(-9850);
			7593: out = 16'(-29454);
			7594: out = 16'(-21581);
			7595: out = 16'(-8039);
			7596: out = 16'(-888);
			7597: out = 16'(4621);
			7598: out = 16'(16765);
			7599: out = 16'(20795);
			7600: out = 16'(9705);
			7601: out = 16'(-7001);
			7602: out = 16'(-13525);
			7603: out = 16'(-4661);
			7604: out = 16'(-6980);
			7605: out = 16'(-11896);
			7606: out = 16'(-1980);
			7607: out = 16'(18032);
			7608: out = 16'(18387);
			7609: out = 16'(5420);
			7610: out = 16'(-2570);
			7611: out = 16'(4092);
			7612: out = 16'(-3005);
			7613: out = 16'(-16474);
			7614: out = 16'(-20212);
			7615: out = 16'(2092);
			7616: out = 16'(1099);
			7617: out = 16'(8367);
			7618: out = 16'(12816);
			7619: out = 16'(12965);
			7620: out = 16'(2605);
			7621: out = 16'(-4218);
			7622: out = 16'(-11729);
			7623: out = 16'(-12932);
			7624: out = 16'(-4134);
			7625: out = 16'(11049);
			7626: out = 16'(15791);
			7627: out = 16'(11342);
			7628: out = 16'(940);
			7629: out = 16'(-4100);
			7630: out = 16'(-10008);
			7631: out = 16'(-3869);
			7632: out = 16'(13101);
			7633: out = 16'(13176);
			7634: out = 16'(-9079);
			7635: out = 16'(-25126);
			7636: out = 16'(-4749);
			7637: out = 16'(-2206);
			7638: out = 16'(2416);
			7639: out = 16'(-2126);
			7640: out = 16'(1663);
			7641: out = 16'(8949);
			7642: out = 16'(20208);
			7643: out = 16'(7777);
			7644: out = 16'(-16638);
			7645: out = 16'(-28625);
			7646: out = 16'(-12172);
			7647: out = 16'(5644);
			7648: out = 16'(5808);
			7649: out = 16'(-72);
			7650: out = 16'(6535);
			7651: out = 16'(12285);
			7652: out = 16'(4520);
			7653: out = 16'(-16557);
			7654: out = 16'(-4621);
			7655: out = 16'(-1208);
			7656: out = 16'(-1885);
			7657: out = 16'(-4218);
			7658: out = 16'(745);
			7659: out = 16'(48);
			7660: out = 16'(5695);
			7661: out = 16'(9809);
			7662: out = 16'(-6534);
			7663: out = 16'(-3337);
			7664: out = 16'(9140);
			7665: out = 16'(14919);
			7666: out = 16'(4401);
			7667: out = 16'(-6913);
			7668: out = 16'(-5813);
			7669: out = 16'(-70);
			7670: out = 16'(-8693);
			7671: out = 16'(-420);
			7672: out = 16'(1236);
			7673: out = 16'(2307);
			7674: out = 16'(2521);
			7675: out = 16'(15234);
			7676: out = 16'(9645);
			7677: out = 16'(-2777);
			7678: out = 16'(-12804);
			7679: out = 16'(-1996);
			7680: out = 16'(-5928);
			7681: out = 16'(-4671);
			7682: out = 16'(9648);
			7683: out = 16'(25734);
			7684: out = 16'(24397);
			7685: out = 16'(6692);
			7686: out = 16'(-14085);
			7687: out = 16'(-21163);
			7688: out = 16'(-13554);
			7689: out = 16'(-2950);
			7690: out = 16'(74);
			7691: out = 16'(1138);
			7692: out = 16'(9571);
			7693: out = 16'(8686);
			7694: out = 16'(-2602);
			7695: out = 16'(-11209);
			7696: out = 16'(5228);
			7697: out = 16'(9954);
			7698: out = 16'(-141);
			7699: out = 16'(-14237);
			7700: out = 16'(-9093);
			7701: out = 16'(7059);
			7702: out = 16'(17457);
			7703: out = 16'(11255);
			7704: out = 16'(750);
			7705: out = 16'(-1743);
			7706: out = 16'(749);
			7707: out = 16'(-5331);
			7708: out = 16'(-16109);
			7709: out = 16'(-15169);
			7710: out = 16'(-1573);
			7711: out = 16'(4408);
			7712: out = 16'(-375);
			7713: out = 16'(-3275);
			7714: out = 16'(11927);
			7715: out = 16'(18678);
			7716: out = 16'(6290);
			7717: out = 16'(-7744);
			7718: out = 16'(-8286);
			7719: out = 16'(-3231);
			7720: out = 16'(-7225);
			7721: out = 16'(-9605);
			7722: out = 16'(-10466);
			7723: out = 16'(4332);
			7724: out = 16'(18378);
			7725: out = 16'(20475);
			7726: out = 16'(235);
			7727: out = 16'(-13448);
			7728: out = 16'(-13248);
			7729: out = 16'(331);
			7730: out = 16'(-15303);
			7731: out = 16'(-2761);
			7732: out = 16'(13746);
			7733: out = 16'(14893);
			7734: out = 16'(1644);
			7735: out = 16'(1913);
			7736: out = 16'(5047);
			7737: out = 16'(99);
			7738: out = 16'(-8697);
			7739: out = 16'(-9935);
			7740: out = 16'(-3844);
			7741: out = 16'(1080);
			7742: out = 16'(6309);
			7743: out = 16'(1972);
			7744: out = 16'(1242);
			7745: out = 16'(-2891);
			7746: out = 16'(-7719);
			7747: out = 16'(-13246);
			7748: out = 16'(-4001);
			7749: out = 16'(2657);
			7750: out = 16'(-904);
			7751: out = 16'(-9878);
			7752: out = 16'(-1378);
			7753: out = 16'(9107);
			7754: out = 16'(11178);
			7755: out = 16'(11087);
			7756: out = 16'(2813);
			7757: out = 16'(-7593);
			7758: out = 16'(-7900);
			7759: out = 16'(6258);
			7760: out = 16'(9165);
			7761: out = 16'(-6052);
			7762: out = 16'(-22016);
			7763: out = 16'(-16538);
			7764: out = 16'(3096);
			7765: out = 16'(12091);
			7766: out = 16'(14723);
			7767: out = 16'(18672);
			7768: out = 16'(9016);
			7769: out = 16'(-9806);
			7770: out = 16'(-21962);
			7771: out = 16'(-12186);
			7772: out = 16'(-6497);
			7773: out = 16'(-1226);
			7774: out = 16'(332);
			7775: out = 16'(8283);
			7776: out = 16'(16215);
			7777: out = 16'(20024);
			7778: out = 16'(12005);
			7779: out = 16'(352);
			7780: out = 16'(-8018);
			7781: out = 16'(1038);
			7782: out = 16'(3457);
			7783: out = 16'(-6554);
			7784: out = 16'(-17111);
			7785: out = 16'(2138);
			7786: out = 16'(12037);
			7787: out = 16'(-1063);
			7788: out = 16'(-21521);
			7789: out = 16'(-3123);
			7790: out = 16'(14741);
			7791: out = 16'(15044);
			7792: out = 16'(82);
			7793: out = 16'(-13381);
			7794: out = 16'(-8234);
			7795: out = 16'(-1314);
			7796: out = 16'(-5997);
			7797: out = 16'(-9716);
			7798: out = 16'(-3847);
			7799: out = 16'(9865);
			7800: out = 16'(13783);
			7801: out = 16'(7949);
			7802: out = 16'(-3217);
			7803: out = 16'(-3175);
			7804: out = 16'(640);
			7805: out = 16'(-2623);
			7806: out = 16'(-25952);
			7807: out = 16'(-22103);
			7808: out = 16'(-2546);
			7809: out = 16'(10726);
			7810: out = 16'(13886);
			7811: out = 16'(8283);
			7812: out = 16'(-1766);
			7813: out = 16'(-10256);
			7814: out = 16'(-6995);
			7815: out = 16'(5682);
			7816: out = 16'(14898);
			7817: out = 16'(11877);
			7818: out = 16'(3192);
			7819: out = 16'(197);
			7820: out = 16'(-2117);
			7821: out = 16'(-7313);
			7822: out = 16'(-9316);
			7823: out = 16'(-13534);
			7824: out = 16'(-3740);
			7825: out = 16'(4792);
			7826: out = 16'(7798);
			7827: out = 16'(1702);
			7828: out = 16'(14980);
			7829: out = 16'(16155);
			7830: out = 16'(2455);
			7831: out = 16'(-11823);
			7832: out = 16'(-4838);
			7833: out = 16'(1534);
			7834: out = 16'(-1447);
			7835: out = 16'(348);
			7836: out = 16'(-9747);
			7837: out = 16'(-9523);
			7838: out = 16'(-2232);
			7839: out = 16'(8472);
			7840: out = 16'(10448);
			7841: out = 16'(11097);
			7842: out = 16'(6784);
			7843: out = 16'(74);
			7844: out = 16'(-9162);
			7845: out = 16'(-8416);
			7846: out = 16'(-6533);
			7847: out = 16'(-8718);
			7848: out = 16'(-7229);
			7849: out = 16'(2318);
			7850: out = 16'(15571);
			7851: out = 16'(18783);
			7852: out = 16'(13290);
			7853: out = 16'(1544);
			7854: out = 16'(-1010);
			7855: out = 16'(-3320);
			7856: out = 16'(-12686);
			7857: out = 16'(-26492);
			7858: out = 16'(-16868);
			7859: out = 16'(6622);
			7860: out = 16'(14971);
			7861: out = 16'(6704);
			7862: out = 16'(5769);
			7863: out = 16'(12158);
			7864: out = 16'(10045);
			7865: out = 16'(-6371);
			7866: out = 16'(-10279);
			7867: out = 16'(-4263);
			7868: out = 16'(-3564);
			7869: out = 16'(-6658);
			7870: out = 16'(-9953);
			7871: out = 16'(4221);
			7872: out = 16'(13621);
			7873: out = 16'(6979);
			7874: out = 16'(214);
			7875: out = 16'(7766);
			7876: out = 16'(11228);
			7877: out = 16'(-1529);
			7878: out = 16'(-17698);
			7879: out = 16'(-15841);
			7880: out = 16'(-6489);
			7881: out = 16'(-4331);
			7882: out = 16'(314);
			7883: out = 16'(12456);
			7884: out = 16'(15314);
			7885: out = 16'(2564);
			7886: out = 16'(-9718);
			7887: out = 16'(-10236);
			7888: out = 16'(-7527);
			7889: out = 16'(-10111);
			7890: out = 16'(-4485);
			7891: out = 16'(-675);
			7892: out = 16'(10113);
			7893: out = 16'(13508);
			7894: out = 16'(10896);
			7895: out = 16'(970);
			7896: out = 16'(2279);
			7897: out = 16'(-2415);
			7898: out = 16'(-17757);
			7899: out = 16'(-12770);
			7900: out = 16'(-2947);
			7901: out = 16'(10187);
			7902: out = 16'(14933);
			7903: out = 16'(15215);
			7904: out = 16'(8837);
			7905: out = 16'(3227);
			7906: out = 16'(-4541);
			7907: out = 16'(-7477);
			7908: out = 16'(-17407);
			7909: out = 16'(-11640);
			7910: out = 16'(1492);
			7911: out = 16'(10354);
			7912: out = 16'(7445);
			7913: out = 16'(8519);
			7914: out = 16'(5789);
			7915: out = 16'(-1112);
			7916: out = 16'(-15568);
			7917: out = 16'(-4053);
			7918: out = 16'(5781);
			7919: out = 16'(-3582);
			7920: out = 16'(-19243);
			7921: out = 16'(-2359);
			7922: out = 16'(20045);
			7923: out = 16'(12327);
			7924: out = 16'(-13088);
			7925: out = 16'(-15518);
			7926: out = 16'(7847);
			7927: out = 16'(16033);
			7928: out = 16'(-2095);
			7929: out = 16'(-17592);
			7930: out = 16'(-13595);
			7931: out = 16'(-5171);
			7932: out = 16'(-6002);
			7933: out = 16'(14259);
			7934: out = 16'(22101);
			7935: out = 16'(9198);
			7936: out = 16'(-11564);
			7937: out = 16'(-4587);
			7938: out = 16'(6671);
			7939: out = 16'(-140);
			7940: out = 16'(-17605);
			7941: out = 16'(-10759);
			7942: out = 16'(10857);
			7943: out = 16'(12544);
			7944: out = 16'(-2746);
			7945: out = 16'(2560);
			7946: out = 16'(7842);
			7947: out = 16'(8072);
			7948: out = 16'(-5457);
			7949: out = 16'(-9391);
			7950: out = 16'(-18100);
			7951: out = 16'(2283);
			7952: out = 16'(15523);
			7953: out = 16'(7707);
			7954: out = 16'(519);
			7955: out = 16'(-6079);
			7956: out = 16'(-3588);
			7957: out = 16'(2321);
			7958: out = 16'(5799);
			7959: out = 16'(2972);
			7960: out = 16'(1631);
			7961: out = 16'(4336);
			7962: out = 16'(7762);
			7963: out = 16'(170);
			7964: out = 16'(-12195);
			7965: out = 16'(-15088);
			7966: out = 16'(6110);
			7967: out = 16'(4746);
			7968: out = 16'(8382);
			7969: out = 16'(7756);
			7970: out = 16'(7892);
			7971: out = 16'(-13628);
			7972: out = 16'(-10013);
			7973: out = 16'(-8392);
			7974: out = 16'(-12167);
			7975: out = 16'(-5917);
			7976: out = 16'(9891);
			7977: out = 16'(7871);
			7978: out = 16'(-8020);
			7979: out = 16'(-15017);
			7980: out = 16'(5150);
			7981: out = 16'(12515);
			7982: out = 16'(-1156);
			7983: out = 16'(-12298);
			7984: out = 16'(2026);
			7985: out = 16'(11531);
			7986: out = 16'(3172);
			7987: out = 16'(-6477);
			7988: out = 16'(761);
			7989: out = 16'(11435);
			7990: out = 16'(9778);
			7991: out = 16'(-2079);
			7992: out = 16'(-8479);
			7993: out = 16'(-9454);
			7994: out = 16'(-6079);
			7995: out = 16'(-3730);
			7996: out = 16'(3980);
			7997: out = 16'(3728);
			7998: out = 16'(8873);
			7999: out = 16'(7922);
			8000: out = 16'(-7611);
			8001: out = 16'(-11459);
			8002: out = 16'(-1203);
			8003: out = 16'(13237);
			8004: out = 16'(15103);
			8005: out = 16'(-10248);
			8006: out = 16'(-18168);
			8007: out = 16'(-4528);
			8008: out = 16'(9520);
			8009: out = 16'(13943);
			8010: out = 16'(13182);
			8011: out = 16'(12485);
			8012: out = 16'(4484);
			8013: out = 16'(-11425);
			8014: out = 16'(-28691);
			8015: out = 16'(-23583);
			8016: out = 16'(-3710);
			8017: out = 16'(8172);
			8018: out = 16'(9091);
			8019: out = 16'(17412);
			8020: out = 16'(20879);
			8021: out = 16'(12951);
			8022: out = 16'(-18158);
			8023: out = 16'(-24372);
			8024: out = 16'(-11631);
			8025: out = 16'(-5383);
			8026: out = 16'(-11266);
			8027: out = 16'(-655);
			8028: out = 16'(17779);
			8029: out = 16'(22694);
			8030: out = 16'(12044);
			8031: out = 16'(6105);
			8032: out = 16'(-532);
			8033: out = 16'(-11847);
			8034: out = 16'(-24139);
			8035: out = 16'(-11862);
			8036: out = 16'(1549);
			8037: out = 16'(-1330);
			8038: out = 16'(-8583);
			8039: out = 16'(10581);
			8040: out = 16'(26780);
			8041: out = 16'(14482);
			8042: out = 16'(-17641);
			8043: out = 16'(-25337);
			8044: out = 16'(-11026);
			8045: out = 16'(3358);
			8046: out = 16'(-452);
			8047: out = 16'(2908);
			8048: out = 16'(3165);
			8049: out = 16'(7189);
			8050: out = 16'(6369);
			8051: out = 16'(2842);
			8052: out = 16'(2976);
			8053: out = 16'(7275);
			8054: out = 16'(3268);
			8055: out = 16'(-12280);
			8056: out = 16'(-22742);
			8057: out = 16'(-13169);
			8058: out = 16'(8108);
			8059: out = 16'(16328);
			8060: out = 16'(7784);
			8061: out = 16'(3019);
			8062: out = 16'(7003);
			8063: out = 16'(4800);
			8064: out = 16'(-4480);
			8065: out = 16'(-20535);
			8066: out = 16'(-18768);
			8067: out = 16'(-62);
			8068: out = 16'(16585);
			8069: out = 16'(8864);
			8070: out = 16'(3838);
			8071: out = 16'(4323);
			8072: out = 16'(238);
			8073: out = 16'(-10867);
			8074: out = 16'(-12594);
			8075: out = 16'(-5002);
			8076: out = 16'(-918);
			8077: out = 16'(6130);
			8078: out = 16'(15148);
			8079: out = 16'(17538);
			8080: out = 16'(5938);
			8081: out = 16'(-9442);
			8082: out = 16'(-7313);
			8083: out = 16'(6963);
			8084: out = 16'(7100);
			8085: out = 16'(-14177);
			8086: out = 16'(-18980);
			8087: out = 16'(-2959);
			8088: out = 16'(9269);
			8089: out = 16'(8247);
			8090: out = 16'(-1212);
			8091: out = 16'(-693);
			8092: out = 16'(749);
			8093: out = 16'(-445);
			8094: out = 16'(-4329);
			8095: out = 16'(9190);
			8096: out = 16'(14993);
			8097: out = 16'(3108);
			8098: out = 16'(-10972);
			8099: out = 16'(-3815);
			8100: out = 16'(2049);
			8101: out = 16'(-6721);
			8102: out = 16'(-549);
			8103: out = 16'(13502);
			8104: out = 16'(14643);
			8105: out = 16'(-3748);
			8106: out = 16'(-17618);
			8107: out = 16'(-15621);
			8108: out = 16'(-7145);
			8109: out = 16'(-4703);
			8110: out = 16'(5855);
			8111: out = 16'(2235);
			8112: out = 16'(1570);
			8113: out = 16'(695);
			8114: out = 16'(5690);
			8115: out = 16'(2782);
			8116: out = 16'(8173);
			8117: out = 16'(11552);
			8118: out = 16'(9233);
			8119: out = 16'(-6137);
			8120: out = 16'(-7272);
			8121: out = 16'(-2362);
			8122: out = 16'(-844);
			8123: out = 16'(-4093);
			8124: out = 16'(2992);
			8125: out = 16'(9704);
			8126: out = 16'(5627);
			8127: out = 16'(962);
			8128: out = 16'(-12876);
			8129: out = 16'(-7269);
			8130: out = 16'(2962);
			8131: out = 16'(-132);
			8132: out = 16'(-174);
			8133: out = 16'(4784);
			8134: out = 16'(8371);
			8135: out = 16'(3463);
			8136: out = 16'(-830);
			8137: out = 16'(777);
			8138: out = 16'(2816);
			8139: out = 16'(-894);
			8140: out = 16'(-2685);
			8141: out = 16'(1308);
			8142: out = 16'(6372);
			8143: out = 16'(6485);
			8144: out = 16'(7052);
			8145: out = 16'(10971);
			8146: out = 16'(8258);
			8147: out = 16'(-7315);
			8148: out = 16'(-23475);
			8149: out = 16'(-25473);
			8150: out = 16'(-8691);
			8151: out = 16'(3813);
			8152: out = 16'(5280);
			8153: out = 16'(9297);
			8154: out = 16'(17188);
			8155: out = 16'(11120);
			8156: out = 16'(-10778);
			8157: out = 16'(-15035);
			8158: out = 16'(-14435);
			8159: out = 16'(-5775);
			8160: out = 16'(3668);
			8161: out = 16'(8964);
			8162: out = 16'(5093);
			8163: out = 16'(-5461);
			8164: out = 16'(-8648);
			8165: out = 16'(2403);
			8166: out = 16'(10802);
			8167: out = 16'(-228);
			8168: out = 16'(-14079);
			8169: out = 16'(-5882);
			8170: out = 16'(10591);
			8171: out = 16'(9454);
			8172: out = 16'(-8171);
			8173: out = 16'(-19784);
			8174: out = 16'(-11081);
			8175: out = 16'(7554);
			8176: out = 16'(12437);
			8177: out = 16'(2508);
			8178: out = 16'(-2556);
			8179: out = 16'(-17);
			8180: out = 16'(12070);
			8181: out = 16'(13456);
			8182: out = 16'(-1641);
			8183: out = 16'(-16901);
			8184: out = 16'(-13680);
			8185: out = 16'(-3521);
			8186: out = 16'(-7191);
			8187: out = 16'(-1654);
			8188: out = 16'(13087);
			8189: out = 16'(22577);
			8190: out = 16'(14569);
			8191: out = 16'(1452);
			8192: out = 16'(-8333);
			8193: out = 16'(-11997);
			8194: out = 16'(-10614);
			8195: out = 16'(-16490);
			8196: out = 16'(4194);
			8197: out = 16'(17750);
			8198: out = 16'(8372);
			8199: out = 16'(-16622);
			8200: out = 16'(-13414);
			8201: out = 16'(-1421);
			8202: out = 16'(1357);
			8203: out = 16'(1106);
			8204: out = 16'(6576);
			8205: out = 16'(9077);
			8206: out = 16'(1929);
			8207: out = 16'(-8269);
			8208: out = 16'(399);
			8209: out = 16'(7318);
			8210: out = 16'(3196);
			8211: out = 16'(-7774);
			8212: out = 16'(-2207);
			8213: out = 16'(21);
			8214: out = 16'(-1268);
			8215: out = 16'(-3901);
			8216: out = 16'(4624);
			8217: out = 16'(7124);
			8218: out = 16'(10474);
			8219: out = 16'(8368);
			8220: out = 16'(-2492);
			8221: out = 16'(-17590);
			8222: out = 16'(-18400);
			8223: out = 16'(-5444);
			8224: out = 16'(-117);
			8225: out = 16'(3720);
			8226: out = 16'(6844);
			8227: out = 16'(14898);
			8228: out = 16'(17791);
			8229: out = 16'(12692);
			8230: out = 16'(690);
			8231: out = 16'(-9752);
			8232: out = 16'(-18517);
			8233: out = 16'(-3737);
			8234: out = 16'(-9734);
			8235: out = 16'(-8987);
			8236: out = 16'(5109);
			8237: out = 16'(23965);
			8238: out = 16'(9507);
			8239: out = 16'(-1865);
			8240: out = 16'(-1896);
			8241: out = 16'(3932);
			8242: out = 16'(-5280);
			8243: out = 16'(-10457);
			8244: out = 16'(-10877);
			8245: out = 16'(-6542);
			8246: out = 16'(-1040);
			8247: out = 16'(15563);
			8248: out = 16'(16889);
			8249: out = 16'(-2966);
			8250: out = 16'(-17336);
			8251: out = 16'(-8448);
			8252: out = 16'(6384);
			8253: out = 16'(1781);
			8254: out = 16'(-2248);
			8255: out = 16'(-3219);
			8256: out = 16'(6504);
			8257: out = 16'(7659);
			8258: out = 16'(982);
			8259: out = 16'(-11218);
			8260: out = 16'(-6175);
			8261: out = 16'(2932);
			8262: out = 16'(-229);
			8263: out = 16'(-3512);
			8264: out = 16'(-2247);
			8265: out = 16'(1265);
			8266: out = 16'(207);
			8267: out = 16'(1884);
			8268: out = 16'(5201);
			8269: out = 16'(6826);
			8270: out = 16'(1825);
			8271: out = 16'(804);
			8272: out = 16'(-1263);
			8273: out = 16'(3395);
			8274: out = 16'(6042);
			8275: out = 16'(-1597);
			8276: out = 16'(-7967);
			8277: out = 16'(-8305);
			8278: out = 16'(-2918);
			8279: out = 16'(-371);
			8280: out = 16'(4219);
			8281: out = 16'(4503);
			8282: out = 16'(4764);
			8283: out = 16'(3137);
			8284: out = 16'(-10980);
			8285: out = 16'(-15280);
			8286: out = 16'(-547);
			8287: out = 16'(17856);
			8288: out = 16'(13731);
			8289: out = 16'(1574);
			8290: out = 16'(-8441);
			8291: out = 16'(-8932);
			8292: out = 16'(-6680);
			8293: out = 16'(-7270);
			8294: out = 16'(-3468);
			8295: out = 16'(5516);
			8296: out = 16'(3475);
			8297: out = 16'(4053);
			8298: out = 16'(-4922);
			8299: out = 16'(-7399);
			8300: out = 16'(1076);
			8301: out = 16'(10298);
			8302: out = 16'(4308);
			8303: out = 16'(-1429);
			8304: out = 16'(5708);
			8305: out = 16'(-341);
			8306: out = 16'(-85);
			8307: out = 16'(-4275);
			8308: out = 16'(-4521);
			8309: out = 16'(3366);
			8310: out = 16'(8673);
			8311: out = 16'(2322);
			8312: out = 16'(-8335);
			8313: out = 16'(-10598);
			8314: out = 16'(-11376);
			8315: out = 16'(-5528);
			8316: out = 16'(7586);
			8317: out = 16'(18245);
			8318: out = 16'(10590);
			8319: out = 16'(-5858);
			8320: out = 16'(-13170);
			8321: out = 16'(-1064);
			8322: out = 16'(7149);
			8323: out = 16'(6148);
			8324: out = 16'(2524);
			8325: out = 16'(4523);
			8326: out = 16'(-4731);
			8327: out = 16'(-2404);
			8328: out = 16'(-1586);
			8329: out = 16'(-1414);
			8330: out = 16'(-1441);
			8331: out = 16'(9606);
			8332: out = 16'(14947);
			8333: out = 16'(9297);
			8334: out = 16'(-1925);
			8335: out = 16'(-11437);
			8336: out = 16'(-10669);
			8337: out = 16'(-3615);
			8338: out = 16'(1580);
			8339: out = 16'(1722);
			8340: out = 16'(766);
			8341: out = 16'(1);
			8342: out = 16'(-1128);
			8343: out = 16'(-19564);
			8344: out = 16'(-11628);
			8345: out = 16'(8031);
			8346: out = 16'(19609);
			8347: out = 16'(14084);
			8348: out = 16'(4926);
			8349: out = 16'(-8222);
			8350: out = 16'(-18140);
			8351: out = 16'(-23176);
			8352: out = 16'(-5388);
			8353: out = 16'(9144);
			8354: out = 16'(13394);
			8355: out = 16'(6117);
			8356: out = 16'(3741);
			8357: out = 16'(-5218);
			8358: out = 16'(-4926);
			8359: out = 16'(1060);
			8360: out = 16'(1968);
			8361: out = 16'(-7394);
			8362: out = 16'(-1139);
			8363: out = 16'(14296);
			8364: out = 16'(10558);
			8365: out = 16'(-9709);
			8366: out = 16'(-12990);
			8367: out = 16'(6891);
			8368: out = 16'(12968);
			8369: out = 16'(1216);
			8370: out = 16'(-5124);
			8371: out = 16'(3734);
			8372: out = 16'(5599);
			8373: out = 16'(4833);
			8374: out = 16'(142);
			8375: out = 16'(-1929);
			8376: out = 16'(-10688);
			8377: out = 16'(-1557);
			8378: out = 16'(-5880);
			8379: out = 16'(-5602);
			8380: out = 16'(1482);
			8381: out = 16'(9421);
			8382: out = 16'(14269);
			8383: out = 16'(18975);
			8384: out = 16'(15141);
			8385: out = 16'(-4387);
			8386: out = 16'(-26050);
			8387: out = 16'(-25136);
			8388: out = 16'(-6927);
			8389: out = 16'(1081);
			8390: out = 16'(4289);
			8391: out = 16'(7048);
			8392: out = 16'(7264);
			8393: out = 16'(1391);
			8394: out = 16'(1374);
			8395: out = 16'(3656);
			8396: out = 16'(1085);
			8397: out = 16'(-8832);
			8398: out = 16'(-10787);
			8399: out = 16'(-1390);
			8400: out = 16'(5362);
			8401: out = 16'(-3147);
			8402: out = 16'(-11858);
			8403: out = 16'(-5459);
			8404: out = 16'(12768);
			8405: out = 16'(16346);
			8406: out = 16'(5375);
			8407: out = 16'(-6441);
			8408: out = 16'(-4014);
			8409: out = 16'(-553);
			8410: out = 16'(-4363);
			8411: out = 16'(-10968);
			8412: out = 16'(1485);
			8413: out = 16'(11716);
			8414: out = 16'(2759);
			8415: out = 16'(-1469);
			8416: out = 16'(-1127);
			8417: out = 16'(3654);
			8418: out = 16'(3839);
			8419: out = 16'(1645);
			8420: out = 16'(-601);
			8421: out = 16'(-5174);
			8422: out = 16'(-7641);
			8423: out = 16'(6749);
			8424: out = 16'(3098);
			8425: out = 16'(-10744);
			8426: out = 16'(-22958);
			8427: out = 16'(-4138);
			8428: out = 16'(-683);
			8429: out = 16'(10007);
			8430: out = 16'(13908);
			8431: out = 16'(13270);
			8432: out = 16'(946);
			8433: out = 16'(-600);
			8434: out = 16'(-6978);
			8435: out = 16'(-17323);
			8436: out = 16'(-4884);
			8437: out = 16'(7561);
			8438: out = 16'(10588);
			8439: out = 16'(6520);
			8440: out = 16'(4324);
			8441: out = 16'(3060);
			8442: out = 16'(-6816);
			8443: out = 16'(-15267);
			8444: out = 16'(-1207);
			8445: out = 16'(1579);
			8446: out = 16'(-2565);
			8447: out = 16'(-6092);
			8448: out = 16'(6389);
			8449: out = 16'(8551);
			8450: out = 16'(8335);
			8451: out = 16'(970);
			8452: out = 16'(-2293);
			8453: out = 16'(-2791);
			8454: out = 16'(2477);
			8455: out = 16'(1546);
			8456: out = 16'(898);
			8457: out = 16'(3382);
			8458: out = 16'(11118);
			8459: out = 16'(5733);
			8460: out = 16'(-4513);
			8461: out = 16'(-1710);
			8462: out = 16'(-602);
			8463: out = 16'(-2664);
			8464: out = 16'(-4371);
			8465: out = 16'(103);
			8466: out = 16'(8984);
			8467: out = 16'(10320);
			8468: out = 16'(8924);
			8469: out = 16'(6245);
			8470: out = 16'(-4005);
			8471: out = 16'(-20622);
			8472: out = 16'(-23413);
			8473: out = 16'(-5521);
			8474: out = 16'(-948);
			8475: out = 16'(5155);
			8476: out = 16'(11687);
			8477: out = 16'(14981);
			8478: out = 16'(14);
			8479: out = 16'(-4187);
			8480: out = 16'(-1610);
			8481: out = 16'(6316);
			8482: out = 16'(8431);
			8483: out = 16'(1784);
			8484: out = 16'(-4790);
			8485: out = 16'(-8500);
			8486: out = 16'(-13160);
			8487: out = 16'(-5022);
			8488: out = 16'(1416);
			8489: out = 16'(5799);
			8490: out = 16'(6950);
			8491: out = 16'(10517);
			8492: out = 16'(-3761);
			8493: out = 16'(-20557);
			8494: out = 16'(-21469);
			8495: out = 16'(-2458);
			8496: out = 16'(8494);
			8497: out = 16'(4395);
			8498: out = 16'(2290);
			8499: out = 16'(10443);
			8500: out = 16'(15757);
			8501: out = 16'(7305);
			8502: out = 16'(-3299);
			8503: out = 16'(-8327);
			8504: out = 16'(3086);
			8505: out = 16'(-5878);
			8506: out = 16'(-16447);
			8507: out = 16'(-11045);
			8508: out = 16'(1548);
			8509: out = 16'(-947);
			8510: out = 16'(-2590);
			8511: out = 16'(7288);
			8512: out = 16'(14805);
			8513: out = 16'(2276);
			8514: out = 16'(-7391);
			8515: out = 16'(-3152);
			8516: out = 16'(-4336);
			8517: out = 16'(-7175);
			8518: out = 16'(-6686);
			8519: out = 16'(4175);
			8520: out = 16'(4008);
			8521: out = 16'(6001);
			8522: out = 16'(-6318);
			8523: out = 16'(-8199);
			8524: out = 16'(708);
			8525: out = 16'(16525);
			8526: out = 16'(617);
			8527: out = 16'(-16488);
			8528: out = 16'(-17867);
			8529: out = 16'(-1216);
			8530: out = 16'(3328);
			8531: out = 16'(11355);
			8532: out = 16'(15685);
			8533: out = 16'(-3561);
			8534: out = 16'(-10720);
			8535: out = 16'(-1752);
			8536: out = 16'(8565);
			8537: out = 16'(-1892);
			8538: out = 16'(-9447);
			8539: out = 16'(3302);
			8540: out = 16'(23212);
			8541: out = 16'(17844);
			8542: out = 16'(-1834);
			8543: out = 16'(-16478);
			8544: out = 16'(-11680);
			8545: out = 16'(-3199);
			8546: out = 16'(1942);
			8547: out = 16'(2463);
			8548: out = 16'(9023);
			8549: out = 16'(13026);
			8550: out = 16'(14824);
			8551: out = 16'(-4557);
			8552: out = 16'(-12593);
			8553: out = 16'(-5094);
			8554: out = 16'(3530);
			8555: out = 16'(-4778);
			8556: out = 16'(-8928);
			8557: out = 16'(-3360);
			8558: out = 16'(3105);
			8559: out = 16'(6684);
			8560: out = 16'(9232);
			8561: out = 16'(10160);
			8562: out = 16'(5279);
			8563: out = 16'(-1997);
			8564: out = 16'(-7551);
			8565: out = 16'(-7334);
			8566: out = 16'(-4321);
			8567: out = 16'(-233);
			8568: out = 16'(2976);
			8569: out = 16'(4282);
			8570: out = 16'(2297);
			8571: out = 16'(4686);
			8572: out = 16'(-1285);
			8573: out = 16'(835);
			8574: out = 16'(3570);
			8575: out = 16'(-1382);
			8576: out = 16'(-13601);
			8577: out = 16'(-14925);
			8578: out = 16'(-6143);
			8579: out = 16'(-1216);
			8580: out = 16'(13637);
			8581: out = 16'(7383);
			8582: out = 16'(-2970);
			8583: out = 16'(-6033);
			8584: out = 16'(9315);
			8585: out = 16'(9424);
			8586: out = 16'(188);
			8587: out = 16'(-11533);
			8588: out = 16'(-11946);
			8589: out = 16'(-9356);
			8590: out = 16'(2580);
			8591: out = 16'(12640);
			8592: out = 16'(12637);
			8593: out = 16'(2962);
			8594: out = 16'(-2069);
			8595: out = 16'(-778);
			8596: out = 16'(1635);
			8597: out = 16'(6054);
			8598: out = 16'(3777);
			8599: out = 16'(-7968);
			8600: out = 16'(-23576);
			8601: out = 16'(-11438);
			8602: out = 16'(-1521);
			8603: out = 16'(2924);
			8604: out = 16'(970);
			8605: out = 16'(-3540);
			8606: out = 16'(-705);
			8607: out = 16'(7780);
			8608: out = 16'(13569);
			8609: out = 16'(7844);
			8610: out = 16'(2715);
			8611: out = 16'(-3417);
			8612: out = 16'(-3126);
			8613: out = 16'(701);
			8614: out = 16'(-10409);
			8615: out = 16'(-14890);
			8616: out = 16'(885);
			8617: out = 16'(17776);
			8618: out = 16'(6963);
			8619: out = 16'(-15448);
			8620: out = 16'(-18468);
			8621: out = 16'(4548);
			8622: out = 16'(6622);
			8623: out = 16'(-1659);
			8624: out = 16'(-7878);
			8625: out = 16'(853);
			8626: out = 16'(10023);
			8627: out = 16'(7473);
			8628: out = 16'(1720);
			8629: out = 16'(-1031);
			8630: out = 16'(-7702);
			8631: out = 16'(-128);
			8632: out = 16'(5470);
			8633: out = 16'(6020);
			8634: out = 16'(-349);
			8635: out = 16'(1602);
			8636: out = 16'(2598);
			8637: out = 16'(1662);
			8638: out = 16'(-4074);
			8639: out = 16'(-5396);
			8640: out = 16'(-9600);
			8641: out = 16'(-9128);
			8642: out = 16'(-2360);
			8643: out = 16'(4104);
			8644: out = 16'(12516);
			8645: out = 16'(14035);
			8646: out = 16'(7729);
			8647: out = 16'(-4280);
			8648: out = 16'(-5271);
			8649: out = 16'(-2534);
			8650: out = 16'(2230);
			8651: out = 16'(6749);
			8652: out = 16'(5446);
			8653: out = 16'(-4063);
			8654: out = 16'(-12220);
			8655: out = 16'(-5363);
			8656: out = 16'(7655);
			8657: out = 16'(17169);
			8658: out = 16'(14387);
			8659: out = 16'(8521);
			8660: out = 16'(2229);
			8661: out = 16'(-3413);
			8662: out = 16'(-18980);
			8663: out = 16'(-28907);
			8664: out = 16'(-22660);
			8665: out = 16'(6888);
			8666: out = 16'(20667);
			8667: out = 16'(17715);
			8668: out = 16'(12874);
			8669: out = 16'(8308);
			8670: out = 16'(-2114);
			8671: out = 16'(-13222);
			8672: out = 16'(-16282);
			8673: out = 16'(-9603);
			8674: out = 16'(-6207);
			8675: out = 16'(61);
			8676: out = 16'(10433);
			8677: out = 16'(7326);
			8678: out = 16'(2975);
			8679: out = 16'(4351);
			8680: out = 16'(10968);
			8681: out = 16'(6291);
			8682: out = 16'(-5900);
			8683: out = 16'(-12812);
			8684: out = 16'(-5392);
			8685: out = 16'(-1783);
			8686: out = 16'(1862);
			8687: out = 16'(1536);
			8688: out = 16'(6082);
			8689: out = 16'(3754);
			8690: out = 16'(6188);
			8691: out = 16'(-6954);
			8692: out = 16'(-13732);
			8693: out = 16'(-13181);
			8694: out = 16'(-27);
			8695: out = 16'(-8228);
			8696: out = 16'(-3069);
			8697: out = 16'(14721);
			8698: out = 16'(20692);
			8699: out = 16'(-3824);
			8700: out = 16'(-15460);
			8701: out = 16'(-5613);
			8702: out = 16'(-5283);
			8703: out = 16'(-962);
			8704: out = 16'(7580);
			8705: out = 16'(10547);
			8706: out = 16'(-6746);
			8707: out = 16'(-5596);
			8708: out = 16'(8106);
			8709: out = 16'(18609);
			8710: out = 16'(6979);
			8711: out = 16'(-14767);
			8712: out = 16'(-23443);
			8713: out = 16'(-14867);
			8714: out = 16'(-7079);
			8715: out = 16'(416);
			8716: out = 16'(1461);
			8717: out = 16'(3700);
			8718: out = 16'(5786);
			8719: out = 16'(10164);
			8720: out = 16'(10110);
			8721: out = 16'(6586);
			8722: out = 16'(-1813);
			8723: out = 16'(-10589);
			8724: out = 16'(-13212);
			8725: out = 16'(-6170);
			8726: out = 16'(4728);
			8727: out = 16'(11133);
			8728: out = 16'(13718);
			8729: out = 16'(5601);
			8730: out = 16'(-4152);
			8731: out = 16'(-7550);
			8732: out = 16'(-5369);
			8733: out = 16'(-286);
			8734: out = 16'(4253);
			8735: out = 16'(6526);
			8736: out = 16'(-1675);
			8737: out = 16'(-381);
			8738: out = 16'(-981);
			8739: out = 16'(-741);
			8740: out = 16'(3184);
			8741: out = 16'(8294);
			8742: out = 16'(11346);
			8743: out = 16'(13747);
			8744: out = 16'(13038);
			8745: out = 16'(-6487);
			8746: out = 16'(-19335);
			8747: out = 16'(-12969);
			8748: out = 16'(4756);
			8749: out = 16'(515);
			8750: out = 16'(-3735);
			8751: out = 16'(-924);
			8752: out = 16'(7568);
			8753: out = 16'(3757);
			8754: out = 16'(-5923);
			8755: out = 16'(-13344);
			8756: out = 16'(-7863);
			8757: out = 16'(255);
			8758: out = 16'(7972);
			8759: out = 16'(4158);
			8760: out = 16'(-331);
			8761: out = 16'(1774);
			8762: out = 16'(3656);
			8763: out = 16'(2169);
			8764: out = 16'(-3113);
			8765: out = 16'(-8201);
			8766: out = 16'(-10774);
			8767: out = 16'(-4574);
			8768: out = 16'(5064);
			8769: out = 16'(8762);
			8770: out = 16'(2519);
			8771: out = 16'(-2422);
			8772: out = 16'(420);
			8773: out = 16'(4708);
			8774: out = 16'(-7889);
			8775: out = 16'(-5478);
			8776: out = 16'(-978);
			8777: out = 16'(3545);
			8778: out = 16'(-1955);
			8779: out = 16'(12545);
			8780: out = 16'(7488);
			8781: out = 16'(-5747);
			8782: out = 16'(-14617);
			8783: out = 16'(7144);
			8784: out = 16'(9368);
			8785: out = 16'(2492);
			8786: out = 16'(305);
			8787: out = 16'(-2130);
			8788: out = 16'(-1403);
			8789: out = 16'(-3554);
			8790: out = 16'(-6459);
			8791: out = 16'(-5732);
			8792: out = 16'(4679);
			8793: out = 16'(15758);
			8794: out = 16'(14958);
			8795: out = 16'(1282);
			8796: out = 16'(-10428);
			8797: out = 16'(-7707);
			8798: out = 16'(2221);
			8799: out = 16'(-235);
			8800: out = 16'(875);
			8801: out = 16'(-3217);
			8802: out = 16'(-792);
			8803: out = 16'(4247);
			8804: out = 16'(6871);
			8805: out = 16'(-665);
			8806: out = 16'(-6749);
			8807: out = 16'(-5106);
			8808: out = 16'(2110);
			8809: out = 16'(1198);
			8810: out = 16'(-520);
			8811: out = 16'(-164);
			8812: out = 16'(-3602);
			8813: out = 16'(-3006);
			8814: out = 16'(-4278);
			8815: out = 16'(-3607);
			8816: out = 16'(453);
			8817: out = 16'(5929);
			8818: out = 16'(4615);
			8819: out = 16'(-1085);
			8820: out = 16'(-2345);
			8821: out = 16'(-251);
			8822: out = 16'(5292);
			8823: out = 16'(-660);
			8824: out = 16'(-14628);
			8825: out = 16'(-3547);
			8826: out = 16'(4660);
			8827: out = 16'(9505);
			8828: out = 16'(3758);
			8829: out = 16'(-6163);
			8830: out = 16'(-11840);
			8831: out = 16'(-633);
			8832: out = 16'(12261);
			8833: out = 16'(7312);
			8834: out = 16'(8505);
			8835: out = 16'(8263);
			8836: out = 16'(7459);
			8837: out = 16'(-1876);
			8838: out = 16'(-3371);
			8839: out = 16'(-8596);
			8840: out = 16'(-3873);
			8841: out = 16'(3467);
			8842: out = 16'(899);
			8843: out = 16'(-11742);
			8844: out = 16'(-10472);
			8845: out = 16'(7866);
			8846: out = 16'(12359);
			8847: out = 16'(5189);
			8848: out = 16'(-7780);
			8849: out = 16'(-12425);
			8850: out = 16'(-11523);
			8851: out = 16'(-2061);
			8852: out = 16'(414);
			8853: out = 16'(1228);
			8854: out = 16'(4979);
			8855: out = 16'(14803);
			8856: out = 16'(9326);
			8857: out = 16'(-5980);
			8858: out = 16'(-17155);
			8859: out = 16'(-11524);
			8860: out = 16'(-2482);
			8861: out = 16'(-229);
			8862: out = 16'(-945);
			8863: out = 16'(-442);
			8864: out = 16'(8363);
			8865: out = 16'(7416);
			8866: out = 16'(-1855);
			8867: out = 16'(-684);
			8868: out = 16'(2138);
			8869: out = 16'(6716);
			8870: out = 16'(5270);
			8871: out = 16'(1339);
			8872: out = 16'(-10113);
			8873: out = 16'(-13755);
			8874: out = 16'(-9385);
			8875: out = 16'(1946);
			8876: out = 16'(14042);
			8877: out = 16'(21139);
			8878: out = 16'(15316);
			8879: out = 16'(866);
			8880: out = 16'(-17705);
			8881: out = 16'(-14061);
			8882: out = 16'(-4266);
			8883: out = 16'(-4325);
			8884: out = 16'(-3444);
			8885: out = 16'(-2363);
			8886: out = 16'(7259);
			8887: out = 16'(13422);
			8888: out = 16'(12533);
			8889: out = 16'(-3822);
			8890: out = 16'(-8960);
			8891: out = 16'(-4348);
			8892: out = 16'(-1136);
			8893: out = 16'(-13298);
			8894: out = 16'(-9149);
			8895: out = 16'(10043);
			8896: out = 16'(20407);
			8897: out = 16'(3700);
			8898: out = 16'(-2030);
			8899: out = 16'(5455);
			8900: out = 16'(10078);
			8901: out = 16'(-11150);
			8902: out = 16'(-19285);
			8903: out = 16'(-12286);
			8904: out = 16'(3907);
			8905: out = 16'(6994);
			8906: out = 16'(4543);
			8907: out = 16'(-6764);
			8908: out = 16'(-9818);
			8909: out = 16'(3591);
			8910: out = 16'(813);
			8911: out = 16'(73);
			8912: out = 16'(1656);
			8913: out = 16'(4416);
			8914: out = 16'(2083);
			8915: out = 16'(-2100);
			8916: out = 16'(-5723);
			8917: out = 16'(-5610);
			8918: out = 16'(-4699);
			8919: out = 16'(-1284);
			8920: out = 16'(3193);
			8921: out = 16'(8374);
			8922: out = 16'(7765);
			8923: out = 16'(11915);
			8924: out = 16'(4500);
			8925: out = 16'(-8792);
			8926: out = 16'(-14754);
			8927: out = 16'(-883);
			8928: out = 16'(11504);
			8929: out = 16'(9589);
			8930: out = 16'(759);
			8931: out = 16'(-3388);
			8932: out = 16'(-1178);
			8933: out = 16'(-3545);
			8934: out = 16'(-10734);
			8935: out = 16'(-1125);
			8936: out = 16'(6066);
			8937: out = 16'(5533);
			8938: out = 16'(-3245);
			8939: out = 16'(807);
			8940: out = 16'(-2616);
			8941: out = 16'(2817);
			8942: out = 16'(6494);
			8943: out = 16'(4289);
			8944: out = 16'(-4743);
			8945: out = 16'(-2337);
			8946: out = 16'(4207);
			8947: out = 16'(3366);
			8948: out = 16'(-3285);
			8949: out = 16'(-3968);
			8950: out = 16'(-578);
			8951: out = 16'(120);
			8952: out = 16'(5127);
			8953: out = 16'(2188);
			8954: out = 16'(-3847);
			8955: out = 16'(-8206);
			8956: out = 16'(-8131);
			8957: out = 16'(-5381);
			8958: out = 16'(-3109);
			8959: out = 16'(3322);
			8960: out = 16'(13626);
			8961: out = 16'(18738);
			8962: out = 16'(9138);
			8963: out = 16'(-3785);
			8964: out = 16'(-6144);
			8965: out = 16'(-4312);
			8966: out = 16'(-6973);
			8967: out = 16'(-13126);
			8968: out = 16'(-12957);
			8969: out = 16'(-2157);
			8970: out = 16'(5970);
			8971: out = 16'(11714);
			8972: out = 16'(16457);
			8973: out = 16'(12656);
			8974: out = 16'(1053);
			8975: out = 16'(-8077);
			8976: out = 16'(-4495);
			8977: out = 16'(-2022);
			8978: out = 16'(-1134);
			8979: out = 16'(-7475);
			8980: out = 16'(-3192);
			8981: out = 16'(10734);
			8982: out = 16'(12194);
			8983: out = 16'(-1334);
			8984: out = 16'(-9580);
			8985: out = 16'(-3244);
			8986: out = 16'(254);
			8987: out = 16'(-8077);
			8988: out = 16'(-8707);
			8989: out = 16'(6641);
			8990: out = 16'(11957);
			8991: out = 16'(3726);
			8992: out = 16'(-2319);
			8993: out = 16'(5186);
			8994: out = 16'(8823);
			8995: out = 16'(432);
			8996: out = 16'(-10215);
			8997: out = 16'(-9905);
			8998: out = 16'(-8889);
			8999: out = 16'(2579);
			9000: out = 16'(2402);
			9001: out = 16'(-2246);
			9002: out = 16'(-7609);
			9003: out = 16'(5134);
			9004: out = 16'(4534);
			9005: out = 16'(55);
			9006: out = 16'(1149);
			9007: out = 16'(13493);
			9008: out = 16'(8386);
			9009: out = 16'(-4740);
			9010: out = 16'(-11014);
			9011: out = 16'(6588);
			9012: out = 16'(6022);
			9013: out = 16'(-545);
			9014: out = 16'(-5057);
			9015: out = 16'(-477);
			9016: out = 16'(1536);
			9017: out = 16'(1504);
			9018: out = 16'(-8228);
			9019: out = 16'(-26415);
			9020: out = 16'(-7371);
			9021: out = 16'(17297);
			9022: out = 16'(22179);
			9023: out = 16'(7318);
			9024: out = 16'(-12518);
			9025: out = 16'(-13968);
			9026: out = 16'(-3379);
			9027: out = 16'(-702);
			9028: out = 16'(1010);
			9029: out = 16'(5344);
			9030: out = 16'(11791);
			9031: out = 16'(4502);
			9032: out = 16'(-8548);
			9033: out = 16'(-22829);
			9034: out = 16'(-10743);
			9035: out = 16'(8148);
			9036: out = 16'(11517);
			9037: out = 16'(-1767);
			9038: out = 16'(1361);
			9039: out = 16'(8990);
			9040: out = 16'(2307);
			9041: out = 16'(-15552);
			9042: out = 16'(-10796);
			9043: out = 16'(7895);
			9044: out = 16'(10420);
			9045: out = 16'(-1675);
			9046: out = 16'(-8537);
			9047: out = 16'(-4564);
			9048: out = 16'(-1093);
			9049: out = 16'(4980);
			9050: out = 16'(-6033);
			9051: out = 16'(-14024);
			9052: out = 16'(-10525);
			9053: out = 16'(16628);
			9054: out = 16'(14712);
			9055: out = 16'(17203);
			9056: out = 16'(11600);
			9057: out = 16'(82);
			9058: out = 16'(-10607);
			9059: out = 16'(-5242);
			9060: out = 16'(-7082);
			9061: out = 16'(-24158);
			9062: out = 16'(-14699);
			9063: out = 16'(7241);
			9064: out = 16'(17129);
			9065: out = 16'(6293);
			9066: out = 16'(-8419);
			9067: out = 16'(1117);
			9068: out = 16'(10075);
			9069: out = 16'(-471);
			9070: out = 16'(-13165);
			9071: out = 16'(-6335);
			9072: out = 16'(10838);
			9073: out = 16'(12322);
			9074: out = 16'(2044);
			9075: out = 16'(-9294);
			9076: out = 16'(-5588);
			9077: out = 16'(1210);
			9078: out = 16'(583);
			9079: out = 16'(6146);
			9080: out = 16'(8071);
			9081: out = 16'(1218);
			9082: out = 16'(-13466);
			9083: out = 16'(-10287);
			9084: out = 16'(-6387);
			9085: out = 16'(4280);
			9086: out = 16'(15151);
			9087: out = 16'(17882);
			9088: out = 16'(13192);
			9089: out = 16'(5408);
			9090: out = 16'(-137);
			9091: out = 16'(-5336);
			9092: out = 16'(-4604);
			9093: out = 16'(-8273);
			9094: out = 16'(-10734);
			9095: out = 16'(-7444);
			9096: out = 16'(441);
			9097: out = 16'(896);
			9098: out = 16'(2615);
			9099: out = 16'(11357);
			9100: out = 16'(9156);
			9101: out = 16'(4415);
			9102: out = 16'(-708);
			9103: out = 16'(328);
			9104: out = 16'(-1194);
			9105: out = 16'(53);
			9106: out = 16'(706);
			9107: out = 16'(5326);
			9108: out = 16'(5111);
			9109: out = 16'(587);
			9110: out = 16'(-13481);
			9111: out = 16'(-21227);
			9112: out = 16'(-16067);
			9113: out = 16'(1423);
			9114: out = 16'(4385);
			9115: out = 16'(5373);
			9116: out = 16'(12036);
			9117: out = 16'(14623);
			9118: out = 16'(-761);
			9119: out = 16'(-13045);
			9120: out = 16'(-5770);
			9121: out = 16'(-71);
			9122: out = 16'(2282);
			9123: out = 16'(2062);
			9124: out = 16'(4229);
			9125: out = 16'(-469);
			9126: out = 16'(-10151);
			9127: out = 16'(-12507);
			9128: out = 16'(359);
			9129: out = 16'(7994);
			9130: out = 16'(8398);
			9131: out = 16'(-3872);
			9132: out = 16'(-11362);
			9133: out = 16'(-9197);
			9134: out = 16'(-864);
			9135: out = 16'(-1774);
			9136: out = 16'(252);
			9137: out = 16'(9910);
			9138: out = 16'(14769);
			9139: out = 16'(7998);
			9140: out = 16'(-1325);
			9141: out = 16'(-4618);
			9142: out = 16'(-3643);
			9143: out = 16'(-4070);
			9144: out = 16'(-5480);
			9145: out = 16'(-6482);
			9146: out = 16'(-7145);
			9147: out = 16'(127);
			9148: out = 16'(10023);
			9149: out = 16'(14056);
			9150: out = 16'(10048);
			9151: out = 16'(2759);
			9152: out = 16'(197);
			9153: out = 16'(-2656);
			9154: out = 16'(-8471);
			9155: out = 16'(-12450);
			9156: out = 16'(-4995);
			9157: out = 16'(1837);
			9158: out = 16'(-787);
			9159: out = 16'(-3599);
			9160: out = 16'(62);
			9161: out = 16'(6086);
			9162: out = 16'(5922);
			9163: out = 16'(2224);
			9164: out = 16'(2863);
			9165: out = 16'(7967);
			9166: out = 16'(8569);
			9167: out = 16'(-1224);
			9168: out = 16'(-10295);
			9169: out = 16'(-10506);
			9170: out = 16'(-461);
			9171: out = 16'(3378);
			9172: out = 16'(8147);
			9173: out = 16'(-574);
			9174: out = 16'(-123);
			9175: out = 16'(6333);
			9176: out = 16'(3936);
			9177: out = 16'(-13950);
			9178: out = 16'(-18661);
			9179: out = 16'(-1475);
			9180: out = 16'(11830);
			9181: out = 16'(-2055);
			9182: out = 16'(-8720);
			9183: out = 16'(7824);
			9184: out = 16'(20777);
			9185: out = 16'(10252);
			9186: out = 16'(-12510);
			9187: out = 16'(-25778);
			9188: out = 16'(-20242);
			9189: out = 16'(705);
			9190: out = 16'(5964);
			9191: out = 16'(-533);
			9192: out = 16'(-6158);
			9193: out = 16'(7242);
			9194: out = 16'(4627);
			9195: out = 16'(-5202);
			9196: out = 16'(-7530);
			9197: out = 16'(12286);
			9198: out = 16'(15986);
			9199: out = 16'(10240);
			9200: out = 16'(277);
			9201: out = 16'(-3966);
			9202: out = 16'(-4605);
			9203: out = 16'(-1361);
			9204: out = 16'(-5870);
			9205: out = 16'(-18383);
			9206: out = 16'(-2977);
			9207: out = 16'(11175);
			9208: out = 16'(8006);
			9209: out = 16'(-5765);
			9210: out = 16'(2990);
			9211: out = 16'(9203);
			9212: out = 16'(4188);
			9213: out = 16'(-6452);
			9214: out = 16'(-605);
			9215: out = 16'(11924);
			9216: out = 16'(12538);
			9217: out = 16'(-6567);
			9218: out = 16'(-28068);
			9219: out = 16'(-13976);
			9220: out = 16'(11913);
			9221: out = 16'(15155);
			9222: out = 16'(286);
			9223: out = 16'(-1895);
			9224: out = 16'(2089);
			9225: out = 16'(2352);
			9226: out = 16'(-7314);
			9227: out = 16'(-12602);
			9228: out = 16'(-6356);
			9229: out = 16'(10149);
			9230: out = 16'(15372);
			9231: out = 16'(4382);
			9232: out = 16'(-12910);
			9233: out = 16'(-10720);
			9234: out = 16'(9065);
			9235: out = 16'(18934);
			9236: out = 16'(1111);
			9237: out = 16'(-14254);
			9238: out = 16'(-9361);
			9239: out = 16'(5760);
			9240: out = 16'(-7909);
			9241: out = 16'(-16902);
			9242: out = 16'(-2335);
			9243: out = 16'(17743);
			9244: out = 16'(4941);
			9245: out = 16'(-12821);
			9246: out = 16'(-14175);
			9247: out = 16'(4766);
			9248: out = 16'(14313);
			9249: out = 16'(11441);
			9250: out = 16'(1153);
			9251: out = 16'(-8725);
			9252: out = 16'(-8416);
			9253: out = 16'(-6901);
			9254: out = 16'(3014);
			9255: out = 16'(9670);
			9256: out = 16'(4946);
			9257: out = 16'(-761);
			9258: out = 16'(4118);
			9259: out = 16'(9280);
			9260: out = 16'(2120);
			9261: out = 16'(-7010);
			9262: out = 16'(-9101);
			9263: out = 16'(-8668);
			9264: out = 16'(-13799);
			9265: out = 16'(-8176);
			9266: out = 16'(4381);
			9267: out = 16'(14938);
			9268: out = 16'(13688);
			9269: out = 16'(1449);
			9270: out = 16'(-4313);
			9271: out = 16'(-8177);
			9272: out = 16'(-8867);
			9273: out = 16'(1687);
			9274: out = 16'(5808);
			9275: out = 16'(2842);
			9276: out = 16'(-259);
			9277: out = 16'(7711);
			9278: out = 16'(8379);
			9279: out = 16'(1507);
			9280: out = 16'(-8599);
			9281: out = 16'(-6193);
			9282: out = 16'(-6037);
			9283: out = 16'(-396);
			9284: out = 16'(-1274);
			9285: out = 16'(-1207);
			9286: out = 16'(4404);
			9287: out = 16'(12548);
			9288: out = 16'(7779);
			9289: out = 16'(-3127);
			9290: out = 16'(-7392);
			9291: out = 16'(5607);
			9292: out = 16'(11094);
			9293: out = 16'(2812);
			9294: out = 16'(-10133);
			9295: out = 16'(-6800);
			9296: out = 16'(-342);
			9297: out = 16'(5514);
			9298: out = 16'(10262);
			9299: out = 16'(8106);
			9300: out = 16'(-1834);
			9301: out = 16'(-8968);
			9302: out = 16'(-6016);
			9303: out = 16'(-7822);
			9304: out = 16'(-5595);
			9305: out = 16'(3600);
			9306: out = 16'(15965);
			9307: out = 16'(17835);
			9308: out = 16'(7793);
			9309: out = 16'(-1089);
			9310: out = 16'(-2330);
			9311: out = 16'(-7270);
			9312: out = 16'(-10795);
			9313: out = 16'(-12847);
			9314: out = 16'(-6130);
			9315: out = 16'(933);
			9316: out = 16'(9111);
			9317: out = 16'(8492);
			9318: out = 16'(8875);
			9319: out = 16'(7233);
			9320: out = 16'(-8752);
			9321: out = 16'(-18238);
			9322: out = 16'(-4948);
			9323: out = 16'(16218);
			9324: out = 16'(10866);
			9325: out = 16'(-438);
			9326: out = 16'(-1909);
			9327: out = 16'(7608);
			9328: out = 16'(16);
			9329: out = 16'(-1999);
			9330: out = 16'(-3097);
			9331: out = 16'(-1414);
			9332: out = 16'(-12058);
			9333: out = 16'(-9346);
			9334: out = 16'(-5894);
			9335: out = 16'(3780);
			9336: out = 16'(5875);
			9337: out = 16'(14313);
			9338: out = 16'(-4202);
			9339: out = 16'(-18441);
			9340: out = 16'(-11005);
			9341: out = 16'(12826);
			9342: out = 16'(8783);
			9343: out = 16'(-121);
			9344: out = 16'(1487);
			9345: out = 16'(3281);
			9346: out = 16'(-1055);
			9347: out = 16'(-9464);
			9348: out = 16'(-11005);
			9349: out = 16'(-2907);
			9350: out = 16'(7810);
			9351: out = 16'(12097);
			9352: out = 16'(2069);
			9353: out = 16'(-22179);
			9354: out = 16'(-1407);
			9355: out = 16'(13845);
			9356: out = 16'(7922);
			9357: out = 16'(-13727);
			9358: out = 16'(-10901);
			9359: out = 16'(-4349);
			9360: out = 16'(1784);
			9361: out = 16'(-128);
			9362: out = 16'(2701);
			9363: out = 16'(148);
			9364: out = 16'(3528);
			9365: out = 16'(8113);
			9366: out = 16'(10643);
			9367: out = 16'(5885);
			9368: out = 16'(85);
			9369: out = 16'(-7273);
			9370: out = 16'(-9657);
			9371: out = 16'(-3511);
			9372: out = 16'(11787);
			9373: out = 16'(13817);
			9374: out = 16'(-1647);
			9375: out = 16'(-10921);
			9376: out = 16'(-7137);
			9377: out = 16'(-235);
			9378: out = 16'(-3836);
			9379: out = 16'(1021);
			9380: out = 16'(-3970);
			9381: out = 16'(-7935);
			9382: out = 16'(-8625);
			9383: out = 16'(7557);
			9384: out = 16'(5255);
			9385: out = 16'(6891);
			9386: out = 16'(11394);
			9387: out = 16'(15718);
			9388: out = 16'(-3855);
			9389: out = 16'(-14502);
			9390: out = 16'(-10753);
			9391: out = 16'(672);
			9392: out = 16'(8288);
			9393: out = 16'(10518);
			9394: out = 16'(4706);
			9395: out = 16'(-7150);
			9396: out = 16'(-1733);
			9397: out = 16'(-5693);
			9398: out = 16'(-9123);
			9399: out = 16'(-6868);
			9400: out = 16'(10167);
			9401: out = 16'(11024);
			9402: out = 16'(9095);
			9403: out = 16'(5382);
			9404: out = 16'(3022);
			9405: out = 16'(-1637);
			9406: out = 16'(-373);
			9407: out = 16'(-486);
			9408: out = 16'(-4942);
			9409: out = 16'(-10496);
			9410: out = 16'(-2798);
			9411: out = 16'(6018);
			9412: out = 16'(2173);
			9413: out = 16'(-11329);
			9414: out = 16'(-4948);
			9415: out = 16'(12326);
			9416: out = 16'(14302);
			9417: out = 16'(4795);
			9418: out = 16'(-2476);
			9419: out = 16'(623);
			9420: out = 16'(-1392);
			9421: out = 16'(-6080);
			9422: out = 16'(-13939);
			9423: out = 16'(-897);
			9424: out = 16'(9018);
			9425: out = 16'(4195);
			9426: out = 16'(-13514);
			9427: out = 16'(-4091);
			9428: out = 16'(7322);
			9429: out = 16'(-1775);
			9430: out = 16'(-13907);
			9431: out = 16'(-507);
			9432: out = 16'(12740);
			9433: out = 16'(4551);
			9434: out = 16'(1494);
			9435: out = 16'(9376);
			9436: out = 16'(14132);
			9437: out = 16'(474);
			9438: out = 16'(-20463);
			9439: out = 16'(-17978);
			9440: out = 16'(-4743);
			9441: out = 16'(1528);
			9442: out = 16'(7670);
			9443: out = 16'(6465);
			9444: out = 16'(3755);
			9445: out = 16'(-7942);
			9446: out = 16'(-21270);
			9447: out = 16'(-4488);
			9448: out = 16'(8363);
			9449: out = 16'(6636);
			9450: out = 16'(553);
			9451: out = 16'(1183);
			9452: out = 16'(5931);
			9453: out = 16'(4674);
			9454: out = 16'(-428);
			9455: out = 16'(-1537);
			9456: out = 16'(-311);
			9457: out = 16'(-1508);
			9458: out = 16'(-2273);
			9459: out = 16'(1441);
			9460: out = 16'(2079);
			9461: out = 16'(135);
			9462: out = 16'(2041);
			9463: out = 16'(7427);
			9464: out = 16'(2211);
			9465: out = 16'(-5113);
			9466: out = 16'(-1395);
			9467: out = 16'(8597);
			9468: out = 16'(1810);
			9469: out = 16'(-15614);
			9470: out = 16'(-16460);
			9471: out = 16'(7042);
			9472: out = 16'(8776);
			9473: out = 16'(5846);
			9474: out = 16'(-2028);
			9475: out = 16'(-2829);
			9476: out = 16'(-8287);
			9477: out = 16'(-1184);
			9478: out = 16'(2820);
			9479: out = 16'(10968);
			9480: out = 16'(16590);
			9481: out = 16'(8229);
			9482: out = 16'(-12376);
			9483: out = 16'(-21747);
			9484: out = 16'(-1274);
			9485: out = 16'(11798);
			9486: out = 16'(11883);
			9487: out = 16'(-4499);
			9488: out = 16'(-17631);
			9489: out = 16'(-3937);
			9490: out = 16'(6830);
			9491: out = 16'(5141);
			9492: out = 16'(-1490);
			9493: out = 16'(-11984);
			9494: out = 16'(2180);
			9495: out = 16'(5714);
			9496: out = 16'(-4052);
			9497: out = 16'(-14216);
			9498: out = 16'(1833);
			9499: out = 16'(10778);
			9500: out = 16'(6717);
			9501: out = 16'(2146);
			9502: out = 16'(3409);
			9503: out = 16'(4971);
			9504: out = 16'(1382);
			9505: out = 16'(-5247);
			9506: out = 16'(-5702);
			9507: out = 16'(-8389);
			9508: out = 16'(-7312);
			9509: out = 16'(-1079);
			9510: out = 16'(6578);
			9511: out = 16'(1481);
			9512: out = 16'(-769);
			9513: out = 16'(5098);
			9514: out = 16'(5776);
			9515: out = 16'(1645);
			9516: out = 16'(-6164);
			9517: out = 16'(-5521);
			9518: out = 16'(-1854);
			9519: out = 16'(10063);
			9520: out = 16'(2942);
			9521: out = 16'(-2879);
			9522: out = 16'(1672);
			9523: out = 16'(3208);
			9524: out = 16'(-3800);
			9525: out = 16'(-5093);
			9526: out = 16'(5079);
			9527: out = 16'(10707);
			9528: out = 16'(5935);
			9529: out = 16'(2139);
			9530: out = 16'(4166);
			9531: out = 16'(428);
			9532: out = 16'(-7606);
			9533: out = 16'(-9949);
			9534: out = 16'(-1606);
			9535: out = 16'(1898);
			9536: out = 16'(7002);
			9537: out = 16'(2140);
			9538: out = 16'(-4425);
			9539: out = 16'(-10537);
			9540: out = 16'(1237);
			9541: out = 16'(1812);
			9542: out = 16'(-537);
			9543: out = 16'(817);
			9544: out = 16'(8387);
			9545: out = 16'(4630);
			9546: out = 16'(-2903);
			9547: out = 16'(-5117);
			9548: out = 16'(2157);
			9549: out = 16'(5944);
			9550: out = 16'(5095);
			9551: out = 16'(1554);
			9552: out = 16'(39);
			9553: out = 16'(-671);
			9554: out = 16'(-1547);
			9555: out = 16'(-5097);
			9556: out = 16'(-6876);
			9557: out = 16'(156);
			9558: out = 16'(7480);
			9559: out = 16'(2042);
			9560: out = 16'(-12512);
			9561: out = 16'(-6068);
			9562: out = 16'(10311);
			9563: out = 16'(18132);
			9564: out = 16'(7131);
			9565: out = 16'(-4140);
			9566: out = 16'(-6764);
			9567: out = 16'(-477);
			9568: out = 16'(-3005);
			9569: out = 16'(-3028);
			9570: out = 16'(-15746);
			9571: out = 16'(-2755);
			9572: out = 16'(13883);
			9573: out = 16'(11512);
			9574: out = 16'(-917);
			9575: out = 16'(-507);
			9576: out = 16'(3981);
			9577: out = 16'(268);
			9578: out = 16'(-4672);
			9579: out = 16'(347);
			9580: out = 16'(1418);
			9581: out = 16'(-8062);
			9582: out = 16'(-12265);
			9583: out = 16'(-108);
			9584: out = 16'(6875);
			9585: out = 16'(-695);
			9586: out = 16'(572);
			9587: out = 16'(1233);
			9588: out = 16'(-798);
			9589: out = 16'(-9693);
			9590: out = 16'(-2867);
			9591: out = 16'(-2776);
			9592: out = 16'(7881);
			9593: out = 16'(9999);
			9594: out = 16'(6804);
			9595: out = 16'(-656);
			9596: out = 16'(3494);
			9597: out = 16'(-3733);
			9598: out = 16'(-21253);
			9599: out = 16'(-10031);
			9600: out = 16'(5740);
			9601: out = 16'(5839);
			9602: out = 16'(-8154);
			9603: out = 16'(-6848);
			9604: out = 16'(-2527);
			9605: out = 16'(-848);
			9606: out = 16'(-4306);
			9607: out = 16'(2503);
			9608: out = 16'(423);
			9609: out = 16'(335);
			9610: out = 16'(2845);
			9611: out = 16'(11997);
			9612: out = 16'(2978);
			9613: out = 16'(-1483);
			9614: out = 16'(-2284);
			9615: out = 16'(2014);
			9616: out = 16'(-471);
			9617: out = 16'(60);
			9618: out = 16'(-1476);
			9619: out = 16'(-2844);
			9620: out = 16'(4);
			9621: out = 16'(1007);
			9622: out = 16'(3765);
			9623: out = 16'(6600);
			9624: out = 16'(852);
			9625: out = 16'(-501);
			9626: out = 16'(-2231);
			9627: out = 16'(4194);
			9628: out = 16'(13496);
			9629: out = 16'(2374);
			9630: out = 16'(-13699);
			9631: out = 16'(-13675);
			9632: out = 16'(8089);
			9633: out = 16'(3913);
			9634: out = 16'(1503);
			9635: out = 16'(-536);
			9636: out = 16'(1213);
			9637: out = 16'(-4706);
			9638: out = 16'(-1090);
			9639: out = 16'(5823);
			9640: out = 16'(11658);
			9641: out = 16'(8237);
			9642: out = 16'(2225);
			9643: out = 16'(-5905);
			9644: out = 16'(-11304);
			9645: out = 16'(-15743);
			9646: out = 16'(-121);
			9647: out = 16'(8434);
			9648: out = 16'(6770);
			9649: out = 16'(-630);
			9650: out = 16'(-140);
			9651: out = 16'(-4958);
			9652: out = 16'(-8014);
			9653: out = 16'(-3094);
			9654: out = 16'(2837);
			9655: out = 16'(8416);
			9656: out = 16'(7252);
			9657: out = 16'(2623);
			9658: out = 16'(-3255);
			9659: out = 16'(-3700);
			9660: out = 16'(-2545);
			9661: out = 16'(863);
			9662: out = 16'(3403);
			9663: out = 16'(5579);
			9664: out = 16'(-26);
			9665: out = 16'(-7051);
			9666: out = 16'(-11133);
			9667: out = 16'(-10507);
			9668: out = 16'(-9884);
			9669: out = 16'(-1428);
			9670: out = 16'(11805);
			9671: out = 16'(16800);
			9672: out = 16'(3865);
			9673: out = 16'(-10461);
			9674: out = 16'(-11153);
			9675: out = 16'(7995);
			9676: out = 16'(-1524);
			9677: out = 16'(-7402);
			9678: out = 16'(5132);
			9679: out = 16'(13763);
			9680: out = 16'(9194);
			9681: out = 16'(-9211);
			9682: out = 16'(-18253);
			9683: out = 16'(-9175);
			9684: out = 16'(-776);
			9685: out = 16'(-2005);
			9686: out = 16'(1961);
			9687: out = 16'(14720);
			9688: out = 16'(13189);
			9689: out = 16'(2033);
			9690: out = 16'(-5119);
			9691: out = 16'(1452);
			9692: out = 16'(-1321);
			9693: out = 16'(-216);
			9694: out = 16'(-5661);
			9695: out = 16'(-11543);
			9696: out = 16'(-15072);
			9697: out = 16'(-1320);
			9698: out = 16'(11923);
			9699: out = 16'(12428);
			9700: out = 16'(358);
			9701: out = 16'(-590);
			9702: out = 16'(5492);
			9703: out = 16'(10649);
			9704: out = 16'(5206);
			9705: out = 16'(-1259);
			9706: out = 16'(-2316);
			9707: out = 16'(5571);
			9708: out = 16'(8376);
			9709: out = 16'(1623);
			9710: out = 16'(-7974);
			9711: out = 16'(-6415);
			9712: out = 16'(-491);
			9713: out = 16'(10);
			9714: out = 16'(-5882);
			9715: out = 16'(-100);
			9716: out = 16'(7006);
			9717: out = 16'(-3565);
			9718: out = 16'(-7507);
			9719: out = 16'(-1060);
			9720: out = 16'(8248);
			9721: out = 16'(5611);
			9722: out = 16'(2217);
			9723: out = 16'(3510);
			9724: out = 16'(5805);
			9725: out = 16'(46);
			9726: out = 16'(2702);
			9727: out = 16'(1026);
			9728: out = 16'(501);
			9729: out = 16'(-1592);
			9730: out = 16'(-3378);
			9731: out = 16'(-14027);
			9732: out = 16'(-23318);
			9733: out = 16'(-18393);
			9734: out = 16'(1745);
			9735: out = 16'(10552);
			9736: out = 16'(5360);
			9737: out = 16'(305);
			9738: out = 16'(4590);
			9739: out = 16'(13674);
			9740: out = 16'(6023);
			9741: out = 16'(-7476);
			9742: out = 16'(-9617);
			9743: out = 16'(-2356);
			9744: out = 16'(-2310);
			9745: out = 16'(-9010);
			9746: out = 16'(-7871);
			9747: out = 16'(7259);
			9748: out = 16'(13400);
			9749: out = 16'(7703);
			9750: out = 16'(-2173);
			9751: out = 16'(-10043);
			9752: out = 16'(-7182);
			9753: out = 16'(-878);
			9754: out = 16'(967);
			9755: out = 16'(-2704);
			9756: out = 16'(-777);
			9757: out = 16'(4160);
			9758: out = 16'(6805);
			9759: out = 16'(3804);
			9760: out = 16'(697);
			9761: out = 16'(650);
			9762: out = 16'(68);
			9763: out = 16'(-5181);
			9764: out = 16'(-1636);
			9765: out = 16'(846);
			9766: out = 16'(4152);
			9767: out = 16'(3791);
			9768: out = 16'(8469);
			9769: out = 16'(-1740);
			9770: out = 16'(-3844);
			9771: out = 16'(19);
			9772: out = 16'(-438);
			9773: out = 16'(-624);
			9774: out = 16'(6109);
			9775: out = 16'(13186);
			9776: out = 16'(8210);
			9777: out = 16'(-7965);
			9778: out = 16'(-14862);
			9779: out = 16'(-5091);
			9780: out = 16'(4273);
			9781: out = 16'(-1223);
			9782: out = 16'(-10469);
			9783: out = 16'(-7422);
			9784: out = 16'(5985);
			9785: out = 16'(7296);
			9786: out = 16'(7456);
			9787: out = 16'(6088);
			9788: out = 16'(6805);
			9789: out = 16'(6981);
			9790: out = 16'(-6626);
			9791: out = 16'(-17431);
			9792: out = 16'(-9354);
			9793: out = 16'(11354);
			9794: out = 16'(-949);
			9795: out = 16'(-15998);
			9796: out = 16'(-11391);
			9797: out = 16'(13554);
			9798: out = 16'(5374);
			9799: out = 16'(1687);
			9800: out = 16'(4012);
			9801: out = 16'(8409);
			9802: out = 16'(575);
			9803: out = 16'(-8980);
			9804: out = 16'(-11631);
			9805: out = 16'(-3312);
			9806: out = 16'(8387);
			9807: out = 16'(4113);
			9808: out = 16'(-339);
			9809: out = 16'(0);
			9810: out = 16'(-304);
			9811: out = 16'(-1373);
			9812: out = 16'(-62);
			9813: out = 16'(5084);
			9814: out = 16'(9503);
			9815: out = 16'(1219);
			9816: out = 16'(-4779);
			9817: out = 16'(-5531);
			9818: out = 16'(667);
			9819: out = 16'(2524);
			9820: out = 16'(8456);
			9821: out = 16'(2934);
			9822: out = 16'(-8795);
			9823: out = 16'(-3660);
			9824: out = 16'(-765);
			9825: out = 16'(-3075);
			9826: out = 16'(-7999);
			9827: out = 16'(-3027);
			9828: out = 16'(-3088);
			9829: out = 16'(-5109);
			9830: out = 16'(-8064);
			9831: out = 16'(-6673);
			9832: out = 16'(4575);
			9833: out = 16'(8231);
			9834: out = 16'(5950);
			9835: out = 16'(6367);
			9836: out = 16'(11505);
			9837: out = 16'(9748);
			9838: out = 16'(1281);
			9839: out = 16'(-8037);
			9840: out = 16'(-16959);
			9841: out = 16'(-9218);
			9842: out = 16'(3301);
			9843: out = 16'(7543);
			9844: out = 16'(5848);
			9845: out = 16'(-11475);
			9846: out = 16'(-16380);
			9847: out = 16'(-3195);
			9848: out = 16'(9820);
			9849: out = 16'(7658);
			9850: out = 16'(3065);
			9851: out = 16'(4817);
			9852: out = 16'(6586);
			9853: out = 16'(-8685);
			9854: out = 16'(-8537);
			9855: out = 16'(10843);
			9856: out = 16'(21067);
			9857: out = 16'(9387);
			9858: out = 16'(-10760);
			9859: out = 16'(-8823);
			9860: out = 16'(7324);
			9861: out = 16'(-257);
			9862: out = 16'(-15437);
			9863: out = 16'(-15077);
			9864: out = 16'(6794);
			9865: out = 16'(14636);
			9866: out = 16'(-16);
			9867: out = 16'(-19239);
			9868: out = 16'(-18659);
			9869: out = 16'(1128);
			9870: out = 16'(10734);
			9871: out = 16'(10215);
			9872: out = 16'(7945);
			9873: out = 16'(8977);
			9874: out = 16'(191);
			9875: out = 16'(-2325);
			9876: out = 16'(-3154);
			9877: out = 16'(1082);
			9878: out = 16'(2657);
			9879: out = 16'(5707);
			9880: out = 16'(-5316);
			9881: out = 16'(-20173);
			9882: out = 16'(-27028);
			9883: out = 16'(3045);
			9884: out = 16'(17163);
			9885: out = 16'(6555);
			9886: out = 16'(-9159);
			9887: out = 16'(5377);
			9888: out = 16'(7881);
			9889: out = 16'(-6802);
			9890: out = 16'(-21938);
			9891: out = 16'(-1122);
			9892: out = 16'(9839);
			9893: out = 16'(4668);
			9894: out = 16'(-3405);
			9895: out = 16'(8782);
			9896: out = 16'(8553);
			9897: out = 16'(1262);
			9898: out = 16'(-9115);
			9899: out = 16'(-6382);
			9900: out = 16'(-6623);
			9901: out = 16'(3985);
			9902: out = 16'(9881);
			9903: out = 16'(3044);
			9904: out = 16'(-8565);
			9905: out = 16'(867);
			9906: out = 16'(15719);
			9907: out = 16'(6986);
			9908: out = 16'(-6997);
			9909: out = 16'(-17888);
			9910: out = 16'(-7742);
			9911: out = 16'(3973);
			9912: out = 16'(1886);
			9913: out = 16'(-6585);
			9914: out = 16'(-78);
			9915: out = 16'(11230);
			9916: out = 16'(7246);
			9917: out = 16'(-9168);
			9918: out = 16'(-15574);
			9919: out = 16'(-7063);
			9920: out = 16'(243);
			9921: out = 16'(-319);
			9922: out = 16'(1632);
			9923: out = 16'(6513);
			9924: out = 16'(8519);
			9925: out = 16'(6997);
			9926: out = 16'(10904);
			9927: out = 16'(8603);
			9928: out = 16'(-7170);
			9929: out = 16'(-16813);
			9930: out = 16'(-15840);
			9931: out = 16'(-4238);
			9932: out = 16'(2565);
			9933: out = 16'(7767);
			9934: out = 16'(9092);
			9935: out = 16'(12737);
			9936: out = 16'(10513);
			9937: out = 16'(3330);
			9938: out = 16'(-8159);
			9939: out = 16'(-9468);
			9940: out = 16'(-3855);
			9941: out = 16'(1859);
			9942: out = 16'(192);
			9943: out = 16'(2810);
			9944: out = 16'(3353);
			9945: out = 16'(-97);
			9946: out = 16'(-224);
			9947: out = 16'(7548);
			9948: out = 16'(11039);
			9949: out = 16'(5022);
			9950: out = 16'(1714);
			9951: out = 16'(-3402);
			9952: out = 16'(-5154);
			9953: out = 16'(-823);
			9954: out = 16'(9127);
			9955: out = 16'(7685);
			9956: out = 16'(-3859);
			9957: out = 16'(-12240);
			9958: out = 16'(-3052);
			9959: out = 16'(-451);
			9960: out = 16'(-3082);
			9961: out = 16'(-5608);
			9962: out = 16'(371);
			9963: out = 16'(-242);
			9964: out = 16'(3020);
			9965: out = 16'(7986);
			9966: out = 16'(10264);
			9967: out = 16'(1007);
			9968: out = 16'(-571);
			9969: out = 16'(4042);
			9970: out = 16'(4835);
			9971: out = 16'(743);
			9972: out = 16'(-14971);
			9973: out = 16'(-15749);
			9974: out = 16'(-2918);
			9975: out = 16'(3691);
			9976: out = 16'(2012);
			9977: out = 16'(3028);
			9978: out = 16'(492);
			9979: out = 16'(-15000);
			9980: out = 16'(-27479);
			9981: out = 16'(-15990);
			9982: out = 16'(10339);
			9983: out = 16'(17558);
			9984: out = 16'(11913);
			9985: out = 16'(2309);
			9986: out = 16'(43);
			9987: out = 16'(748);
			9988: out = 16'(8132);
			9989: out = 16'(4393);
			9990: out = 16'(-65);
			9991: out = 16'(-5340);
			9992: out = 16'(546);
			9993: out = 16'(-21692);
			9994: out = 16'(-22029);
			9995: out = 16'(1280);
			9996: out = 16'(16387);
			9997: out = 16'(10286);
			9998: out = 16'(1289);
			9999: out = 16'(-1040);
			10000: out = 16'(-405);
			10001: out = 16'(-2118);
			10002: out = 16'(-3557);
			10003: out = 16'(-130);
			10004: out = 16'(4547);
			10005: out = 16'(2086);
			10006: out = 16'(403);
			10007: out = 16'(622);
			10008: out = 16'(1912);
			10009: out = 16'(2995);
			10010: out = 16'(-6505);
			10011: out = 16'(-8277);
			10012: out = 16'(6668);
			10013: out = 16'(19960);
			10014: out = 16'(15842);
			10015: out = 16'(-6881);
			10016: out = 16'(-24024);
			10017: out = 16'(-12171);
			10018: out = 16'(-2681);
			10019: out = 16'(7565);
			10020: out = 16'(11627);
			10021: out = 16'(10405);
			10022: out = 16'(-5);
			10023: out = 16'(-6632);
			10024: out = 16'(-4337);
			10025: out = 16'(3730);
			10026: out = 16'(1139);
			10027: out = 16'(510);
			10028: out = 16'(-445);
			10029: out = 16'(-546);
			10030: out = 16'(-6214);
			10031: out = 16'(1720);
			10032: out = 16'(6772);
			10033: out = 16'(7007);
			10034: out = 16'(2154);
			10035: out = 16'(1923);
			10036: out = 16'(-5427);
			10037: out = 16'(-11729);
			10038: out = 16'(-6548);
			10039: out = 16'(-7346);
			10040: out = 16'(2684);
			10041: out = 16'(8217);
			10042: out = 16'(7293);
			10043: out = 16'(-37);
			10044: out = 16'(2903);
			10045: out = 16'(1180);
			10046: out = 16'(-6489);
			10047: out = 16'(-8771);
			10048: out = 16'(-8607);
			10049: out = 16'(-4097);
			10050: out = 16'(4655);
			10051: out = 16'(17106);
			10052: out = 16'(11937);
			10053: out = 16'(2847);
			10054: out = 16'(-6958);
			10055: out = 16'(-12248);
			10056: out = 16'(-7361);
			10057: out = 16'(-4097);
			10058: out = 16'(-618);
			10059: out = 16'(5382);
			10060: out = 16'(6403);
			10061: out = 16'(7233);
			10062: out = 16'(6357);
			10063: out = 16'(7053);
			10064: out = 16'(7098);
			10065: out = 16'(-1412);
			10066: out = 16'(-16523);
			10067: out = 16'(-24898);
			10068: out = 16'(-10192);
			10069: out = 16'(-3545);
			10070: out = 16'(4457);
			10071: out = 16'(10712);
			10072: out = 16'(13407);
			10073: out = 16'(3774);
			10074: out = 16'(-5214);
			10075: out = 16'(-9160);
			10076: out = 16'(-4462);
			10077: out = 16'(529);
			10078: out = 16'(2055);
			10079: out = 16'(-2666);
			10080: out = 16'(-3787);
			10081: out = 16'(5904);
			10082: out = 16'(10817);
			10083: out = 16'(2847);
			10084: out = 16'(-9506);
			10085: out = 16'(-9639);
			10086: out = 16'(-4929);
			10087: out = 16'(-1773);
			10088: out = 16'(-2496);
			10089: out = 16'(1797);
			10090: out = 16'(8495);
			10091: out = 16'(10251);
			10092: out = 16'(1679);
			10093: out = 16'(-6684);
			10094: out = 16'(-2886);
			10095: out = 16'(2871);
			10096: out = 16'(-699);
			10097: out = 16'(-6645);
			10098: out = 16'(-688);
			10099: out = 16'(7687);
			10100: out = 16'(5572);
			10101: out = 16'(-2355);
			10102: out = 16'(717);
			10103: out = 16'(12686);
			10104: out = 16'(16827);
			10105: out = 16'(6013);
			10106: out = 16'(-10338);
			10107: out = 16'(-13104);
			10108: out = 16'(-5816);
			10109: out = 16'(1523);
			10110: out = 16'(1296);
			10111: out = 16'(7777);
			10112: out = 16'(3011);
			10113: out = 16'(-1203);
			10114: out = 16'(-1953);
			10115: out = 16'(-2986);
			10116: out = 16'(-1759);
			10117: out = 16'(2156);
			10118: out = 16'(3622);
			10119: out = 16'(3275);
			10120: out = 16'(-5642);
			10121: out = 16'(-4103);
			10122: out = 16'(3367);
			10123: out = 16'(6358);
			10124: out = 16'(-5022);
			10125: out = 16'(-106);
			10126: out = 16'(11986);
			10127: out = 16'(7696);
			10128: out = 16'(2443);
			10129: out = 16'(-10542);
			10130: out = 16'(-17377);
			10131: out = 16'(-18033);
			10132: out = 16'(-5320);
			10133: out = 16'(-1171);
			10134: out = 16'(2924);
			10135: out = 16'(6350);
			10136: out = 16'(8339);
			10137: out = 16'(4259);
			10138: out = 16'(3390);
			10139: out = 16'(3197);
			10140: out = 16'(-3032);
			10141: out = 16'(-7732);
			10142: out = 16'(-6639);
			10143: out = 16'(-677);
			10144: out = 16'(1357);
			10145: out = 16'(940);
			10146: out = 16'(-683);
			10147: out = 16'(3095);
			10148: out = 16'(9508);
			10149: out = 16'(8110);
			10150: out = 16'(-233);
			10151: out = 16'(-9919);
			10152: out = 16'(-9743);
			10153: out = 16'(1329);
			10154: out = 16'(8798);
			10155: out = 16'(6322);
			10156: out = 16'(3319);
			10157: out = 16'(5888);
			10158: out = 16'(-339);
			10159: out = 16'(-14607);
			10160: out = 16'(-17490);
			10161: out = 16'(7582);
			10162: out = 16'(8226);
			10163: out = 16'(3801);
			10164: out = 16'(1090);
			10165: out = 16'(6920);
			10166: out = 16'(-809);
			10167: out = 16'(-3803);
			10168: out = 16'(-2500);
			10169: out = 16'(3949);
			10170: out = 16'(5924);
			10171: out = 16'(4610);
			10172: out = 16'(-643);
			10173: out = 16'(-5175);
			10174: out = 16'(-5785);
			10175: out = 16'(2776);
			10176: out = 16'(10185);
			10177: out = 16'(9560);
			10178: out = 16'(6471);
			10179: out = 16'(-5736);
			10180: out = 16'(-5172);
			10181: out = 16'(2141);
			10182: out = 16'(6472);
			10183: out = 16'(-16404);
			10184: out = 16'(-16305);
			10185: out = 16'(825);
			10186: out = 16'(12129);
			10187: out = 16'(7215);
			10188: out = 16'(5120);
			10189: out = 16'(5475);
			10190: out = 16'(5914);
			10191: out = 16'(1988);
			10192: out = 16'(912);
			10193: out = 16'(-8455);
			10194: out = 16'(-21296);
			10195: out = 16'(-21556);
			10196: out = 16'(-8690);
			10197: out = 16'(6786);
			10198: out = 16'(14684);
			10199: out = 16'(17366);
			10200: out = 16'(12398);
			10201: out = 16'(270);
			10202: out = 16'(-15458);
			10203: out = 16'(-22017);
			10204: out = 16'(-10708);
			10205: out = 16'(1012);
			10206: out = 16'(2157);
			10207: out = 16'(510);
			10208: out = 16'(-577);
			10209: out = 16'(7408);
			10210: out = 16'(6492);
			10211: out = 16'(448);
			10212: out = 16'(128);
			10213: out = 16'(650);
			10214: out = 16'(-4360);
			10215: out = 16'(-7390);
			10216: out = 16'(3446);
			10217: out = 16'(4147);
			10218: out = 16'(2070);
			10219: out = 16'(1077);
			10220: out = 16'(5477);
			10221: out = 16'(512);
			10222: out = 16'(-3136);
			10223: out = 16'(-4223);
			10224: out = 16'(-2865);
			10225: out = 16'(118);
			10226: out = 16'(-7174);
			10227: out = 16'(-6127);
			10228: out = 16'(7667);
			10229: out = 16'(10967);
			10230: out = 16'(6007);
			10231: out = 16'(-7909);
			10232: out = 16'(-14076);
			10233: out = 16'(-4122);
			10234: out = 16'(5872);
			10235: out = 16'(8425);
			10236: out = 16'(5000);
			10237: out = 16'(1547);
			10238: out = 16'(87);
			10239: out = 16'(168);
			10240: out = 16'(-69);
			10241: out = 16'(205);
			10242: out = 16'(-107);
			10243: out = 16'(-2372);
			10244: out = 16'(-6517);
			10245: out = 16'(-6119);
			10246: out = 16'(-616);
			10247: out = 16'(5803);
			10248: out = 16'(5178);
			10249: out = 16'(2687);
			10250: out = 16'(1132);
			10251: out = 16'(8333);
			10252: out = 16'(127);
			10253: out = 16'(-11859);
			10254: out = 16'(-2619);
			10255: out = 16'(1456);
			10256: out = 16'(8635);
			10257: out = 16'(6057);
			10258: out = 16'(-211);
			10259: out = 16'(-3308);
			10260: out = 16'(-1267);
			10261: out = 16'(-321);
			10262: out = 16'(703);
			10263: out = 16'(3209);
			10264: out = 16'(2085);
			10265: out = 16'(-5572);
			10266: out = 16'(-9172);
			10267: out = 16'(-974);
			10268: out = 16'(7963);
			10269: out = 16'(3209);
			10270: out = 16'(-6593);
			10271: out = 16'(-6433);
			10272: out = 16'(10309);
			10273: out = 16'(13536);
			10274: out = 16'(4710);
			10275: out = 16'(182);
			10276: out = 16'(2398);
			10277: out = 16'(2257);
			10278: out = 16'(-4693);
			10279: out = 16'(-8410);
			10280: out = 16'(-729);
			10281: out = 16'(3124);
			10282: out = 16'(-322);
			10283: out = 16'(-2396);
			10284: out = 16'(3139);
			10285: out = 16'(1637);
			10286: out = 16'(-5042);
			10287: out = 16'(-4746);
			10288: out = 16'(8346);
			10289: out = 16'(7809);
			10290: out = 16'(-2984);
			10291: out = 16'(-9577);
			10292: out = 16'(3621);
			10293: out = 16'(-575);
			10294: out = 16'(43);
			10295: out = 16'(-1043);
			10296: out = 16'(-615);
			10297: out = 16'(-7526);
			10298: out = 16'(-3180);
			10299: out = 16'(1092);
			10300: out = 16'(1050);
			10301: out = 16'(9);
			10302: out = 16'(-5436);
			10303: out = 16'(-5831);
			10304: out = 16'(4706);
			10305: out = 16'(17941);
			10306: out = 16'(9889);
			10307: out = 16'(-7309);
			10308: out = 16'(-16897);
			10309: out = 16'(-6982);
			10310: out = 16'(-519);
			10311: out = 16'(3308);
			10312: out = 16'(5046);
			10313: out = 16'(5723);
			10314: out = 16'(-2899);
			10315: out = 16'(-9270);
			10316: out = 16'(-8650);
			10317: out = 16'(-4717);
			10318: out = 16'(-9499);
			10319: out = 16'(-8144);
			10320: out = 16'(603);
			10321: out = 16'(6683);
			10322: out = 16'(681);
			10323: out = 16'(-2820);
			10324: out = 16'(4612);
			10325: out = 16'(14864);
			10326: out = 16'(14779);
			10327: out = 16'(4173);
			10328: out = 16'(-591);
			10329: out = 16'(-1205);
			10330: out = 16'(-5720);
			10331: out = 16'(-15206);
			10332: out = 16'(-13014);
			10333: out = 16'(-1603);
			10334: out = 16'(6260);
			10335: out = 16'(9271);
			10336: out = 16'(6196);
			10337: out = 16'(2064);
			10338: out = 16'(346);
			10339: out = 16'(1057);
			10340: out = 16'(1940);
			10341: out = 16'(-1437);
			10342: out = 16'(-5245);
			10343: out = 16'(-7679);
			10344: out = 16'(-2294);
			10345: out = 16'(-1296);
			10346: out = 16'(4870);
			10347: out = 16'(17931);
			10348: out = 16'(18268);
			10349: out = 16'(1757);
			10350: out = 16'(-16426);
			10351: out = 16'(-16818);
			10352: out = 16'(-4535);
			10353: out = 16'(1143);
			10354: out = 16'(-2076);
			10355: out = 16'(-1315);
			10356: out = 16'(3292);
			10357: out = 16'(9618);
			10358: out = 16'(6125);
			10359: out = 16'(-1070);
			10360: out = 16'(135);
			10361: out = 16'(-6246);
			10362: out = 16'(-5896);
			10363: out = 16'(-2179);
			10364: out = 16'(-2795);
			10365: out = 16'(8449);
			10366: out = 16'(10418);
			10367: out = 16'(6159);
			10368: out = 16'(-946);
			10369: out = 16'(167);
			10370: out = 16'(-729);
			10371: out = 16'(433);
			10372: out = 16'(719);
			10373: out = 16'(446);
			10374: out = 16'(-3251);
			10375: out = 16'(2326);
			10376: out = 16'(12580);
			10377: out = 16'(11968);
			10378: out = 16'(-1651);
			10379: out = 16'(-17194);
			10380: out = 16'(-20874);
			10381: out = 16'(-7814);
			10382: out = 16'(-12460);
			10383: out = 16'(-9384);
			10384: out = 16'(4151);
			10385: out = 16'(17274);
			10386: out = 16'(15064);
			10387: out = 16'(9238);
			10388: out = 16'(659);
			10389: out = 16'(-5786);
			10390: out = 16'(1759);
			10391: out = 16'(-2889);
			10392: out = 16'(-14505);
			10393: out = 16'(-20087);
			10394: out = 16'(-2410);
			10395: out = 16'(5902);
			10396: out = 16'(5434);
			10397: out = 16'(4949);
			10398: out = 16'(14725);
			10399: out = 16'(7603);
			10400: out = 16'(-1609);
			10401: out = 16'(-7869);
			10402: out = 16'(-2515);
			10403: out = 16'(-9731);
			10404: out = 16'(-7185);
			10405: out = 16'(-1871);
			10406: out = 16'(2395);
			10407: out = 16'(3865);
			10408: out = 16'(8123);
			10409: out = 16'(5719);
			10410: out = 16'(-5569);
			10411: out = 16'(-13395);
			10412: out = 16'(-6495);
			10413: out = 16'(7098);
			10414: out = 16'(5764);
			10415: out = 16'(-5265);
			10416: out = 16'(-14183);
			10417: out = 16'(-1045);
			10418: out = 16'(11992);
			10419: out = 16'(8465);
			10420: out = 16'(-15987);
			10421: out = 16'(-15616);
			10422: out = 16'(5024);
			10423: out = 16'(16946);
			10424: out = 16'(15489);
			10425: out = 16'(10041);
			10426: out = 16'(2230);
			10427: out = 16'(-5387);
			10428: out = 16'(-13498);
			10429: out = 16'(-7979);
			10430: out = 16'(-7643);
			10431: out = 16'(-10087);
			10432: out = 16'(150);
			10433: out = 16'(11822);
			10434: out = 16'(10064);
			10435: out = 16'(5181);
			10436: out = 16'(12661);
			10437: out = 16'(18064);
			10438: out = 16'(3307);
			10439: out = 16'(-17108);
			10440: out = 16'(-14779);
			10441: out = 16'(-1301);
			10442: out = 16'(3552);
			10443: out = 16'(-1931);
			10444: out = 16'(2539);
			10445: out = 16'(5763);
			10446: out = 16'(10449);
			10447: out = 16'(5476);
			10448: out = 16'(1227);
			10449: out = 16'(-18858);
			10450: out = 16'(-5194);
			10451: out = 16'(1264);
			10452: out = 16'(-407);
			10453: out = 16'(-6058);
			10454: out = 16'(8725);
			10455: out = 16'(6533);
			10456: out = 16'(-904);
			10457: out = 16'(-174);
			10458: out = 16'(4272);
			10459: out = 16'(-2290);
			10460: out = 16'(-1684);
			10461: out = 16'(11262);
			10462: out = 16'(5530);
			10463: out = 16'(-10083);
			10464: out = 16'(-12120);
			10465: out = 16'(5635);
			10466: out = 16'(-3238);
			10467: out = 16'(-10091);
			10468: out = 16'(-10889);
			10469: out = 16'(-1198);
			10470: out = 16'(-4787);
			10471: out = 16'(2434);
			10472: out = 16'(9044);
			10473: out = 16'(10936);
			10474: out = 16'(-225);
			10475: out = 16'(993);
			10476: out = 16'(4696);
			10477: out = 16'(2456);
			10478: out = 16'(-15093);
			10479: out = 16'(-13225);
			10480: out = 16'(-11564);
			10481: out = 16'(-5051);
			10482: out = 16'(2480);
			10483: out = 16'(15142);
			10484: out = 16'(17465);
			10485: out = 16'(11881);
			10486: out = 16'(-1218);
			10487: out = 16'(-15249);
			10488: out = 16'(-14284);
			10489: out = 16'(-3800);
			10490: out = 16'(-1311);
			10491: out = 16'(-8931);
			10492: out = 16'(-3243);
			10493: out = 16'(10913);
			10494: out = 16'(16689);
			10495: out = 16'(10741);
			10496: out = 16'(1292);
			10497: out = 16'(-1741);
			10498: out = 16'(-7790);
			10499: out = 16'(-18824);
			10500: out = 16'(-14530);
			10501: out = 16'(1120);
			10502: out = 16'(10253);
			10503: out = 16'(5786);
			10504: out = 16'(5457);
			10505: out = 16'(5641);
			10506: out = 16'(7772);
			10507: out = 16'(4680);
			10508: out = 16'(-2792);
			10509: out = 16'(-12514);
			10510: out = 16'(-14006);
			10511: out = 16'(-3680);
			10512: out = 16'(6528);
			10513: out = 16'(10435);
			10514: out = 16'(1221);
			10515: out = 16'(-3740);
			10516: out = 16'(512);
			10517: out = 16'(1014);
			10518: out = 16'(-8434);
			10519: out = 16'(-10912);
			10520: out = 16'(1854);
			10521: out = 16'(10606);
			10522: out = 16'(9201);
			10523: out = 16'(6047);
			10524: out = 16'(7363);
			10525: out = 16'(7425);
			10526: out = 16'(-3311);
			10527: out = 16'(-9352);
			10528: out = 16'(-5939);
			10529: out = 16'(-4956);
			10530: out = 16'(-74);
			10531: out = 16'(-1777);
			10532: out = 16'(-834);
			10533: out = 16'(6566);
			10534: out = 16'(8376);
			10535: out = 16'(9891);
			10536: out = 16'(6023);
			10537: out = 16'(265);
			10538: out = 16'(-3355);
			10539: out = 16'(-2911);
			10540: out = 16'(-6476);
			10541: out = 16'(-8718);
			10542: out = 16'(6305);
			10543: out = 16'(13045);
			10544: out = 16'(11012);
			10545: out = 16'(1989);
			10546: out = 16'(-2900);
			10547: out = 16'(-7623);
			10548: out = 16'(-7745);
			10549: out = 16'(-7632);
			10550: out = 16'(-5477);
			10551: out = 16'(-5148);
			10552: out = 16'(2938);
			10553: out = 16'(11999);
			10554: out = 16'(16159);
			10555: out = 16'(9233);
			10556: out = 16'(3130);
			10557: out = 16'(-5532);
			10558: out = 16'(-13392);
			10559: out = 16'(-15573);
			10560: out = 16'(-4910);
			10561: out = 16'(3670);
			10562: out = 16'(2539);
			10563: out = 16'(-2312);
			10564: out = 16'(927);
			10565: out = 16'(5853);
			10566: out = 16'(4901);
			10567: out = 16'(-203);
			10568: out = 16'(-360);
			10569: out = 16'(355);
			10570: out = 16'(-2313);
			10571: out = 16'(-5446);
			10572: out = 16'(-987);
			10573: out = 16'(6475);
			10574: out = 16'(8028);
			10575: out = 16'(1690);
			10576: out = 16'(-10895);
			10577: out = 16'(-9934);
			10578: out = 16'(-3993);
			10579: out = 16'(1812);
			10580: out = 16'(8870);
			10581: out = 16'(1630);
			10582: out = 16'(-4455);
			10583: out = 16'(-957);
			10584: out = 16'(8630);
			10585: out = 16'(5930);
			10586: out = 16'(-2260);
			10587: out = 16'(-4438);
			10588: out = 16'(1889);
			10589: out = 16'(6507);
			10590: out = 16'(-1862);
			10591: out = 16'(-6976);
			10592: out = 16'(2221);
			10593: out = 16'(10906);
			10594: out = 16'(-340);
			10595: out = 16'(-14978);
			10596: out = 16'(-10906);
			10597: out = 16'(4500);
			10598: out = 16'(9034);
			10599: out = 16'(18);
			10600: out = 16'(-1387);
			10601: out = 16'(9111);
			10602: out = 16'(9085);
			10603: out = 16'(-7467);
			10604: out = 16'(-16629);
			10605: out = 16'(1702);
			10606: out = 16'(5527);
			10607: out = 16'(395);
			10608: out = 16'(-7698);
			10609: out = 16'(-2711);
			10610: out = 16'(-2959);
			10611: out = 16'(3312);
			10612: out = 16'(4362);
			10613: out = 16'(5564);
			10614: out = 16'(-547);
			10615: out = 16'(2909);
			10616: out = 16'(-242);
			10617: out = 16'(-2503);
			10618: out = 16'(-620);
			10619: out = 16'(13901);
			10620: out = 16'(11172);
			10621: out = 16'(359);
			10622: out = 16'(-4372);
			10623: out = 16'(2380);
			10624: out = 16'(-3187);
			10625: out = 16'(-13775);
			10626: out = 16'(-12195);
			10627: out = 16'(-5179);
			10628: out = 16'(1007);
			10629: out = 16'(2934);
			10630: out = 16'(7776);
			10631: out = 16'(5725);
			10632: out = 16'(7533);
			10633: out = 16'(2074);
			10634: out = 16'(-4436);
			10635: out = 16'(-9106);
			10636: out = 16'(4441);
			10637: out = 16'(9088);
			10638: out = 16'(739);
			10639: out = 16'(-11387);
			10640: out = 16'(-3218);
			10641: out = 16'(2324);
			10642: out = 16'(-890);
			10643: out = 16'(-3922);
			10644: out = 16'(-4100);
			10645: out = 16'(1093);
			10646: out = 16'(3156);
			10647: out = 16'(3844);
			10648: out = 16'(-5911);
			10649: out = 16'(2332);
			10650: out = 16'(7959);
			10651: out = 16'(6568);
			10652: out = 16'(-231);
			10653: out = 16'(-1967);
			10654: out = 16'(-5687);
			10655: out = 16'(-4512);
			10656: out = 16'(-1719);
			10657: out = 16'(1614);
			10658: out = 16'(-10229);
			10659: out = 16'(-12873);
			10660: out = 16'(5232);
			10661: out = 16'(20184);
			10662: out = 16'(9059);
			10663: out = 16'(-1964);
			10664: out = 16'(-872);
			10665: out = 16'(-8609);
			10666: out = 16'(-19341);
			10667: out = 16'(-7869);
			10668: out = 16'(16981);
			10669: out = 16'(1658);
			10670: out = 16'(-5472);
			10671: out = 16'(-676);
			10672: out = 16'(10474);
			10673: out = 16'(-776);
			10674: out = 16'(-4031);
			10675: out = 16'(1571);
			10676: out = 16'(4388);
			10677: out = 16'(-17764);
			10678: out = 16'(-12215);
			10679: out = 16'(5064);
			10680: out = 16'(18291);
			10681: out = 16'(6074);
			10682: out = 16'(5407);
			10683: out = 16'(-2812);
			10684: out = 16'(-1354);
			10685: out = 16'(-842);
			10686: out = 16'(2109);
			10687: out = 16'(-5967);
			10688: out = 16'(-5228);
			10689: out = 16'(-3035);
			10690: out = 16'(-12505);
			10691: out = 16'(2610);
			10692: out = 16'(18643);
			10693: out = 16'(11295);
			10694: out = 16'(-13842);
			10695: out = 16'(-19929);
			10696: out = 16'(1600);
			10697: out = 16'(12024);
			10698: out = 16'(-6770);
			10699: out = 16'(-996);
			10700: out = 16'(8929);
			10701: out = 16'(5286);
			10702: out = 16'(-17192);
			10703: out = 16'(-11998);
			10704: out = 16'(354);
			10705: out = 16'(6931);
			10706: out = 16'(-1451);
			10707: out = 16'(1616);
			10708: out = 16'(1462);
			10709: out = 16'(3893);
			10710: out = 16'(3568);
			10711: out = 16'(10827);
			10712: out = 16'(6949);
			10713: out = 16'(2170);
			10714: out = 16'(-5373);
			10715: out = 16'(-3707);
			10716: out = 16'(-12222);
			10717: out = 16'(-5998);
			10718: out = 16'(696);
			10719: out = 16'(4837);
			10720: out = 16'(-546);
			10721: out = 16'(8099);
			10722: out = 16'(8502);
			10723: out = 16'(-52);
			10724: out = 16'(-312);
			10725: out = 16'(488);
			10726: out = 16'(-5264);
			10727: out = 16'(-10179);
			10728: out = 16'(6719);
			10729: out = 16'(9123);
			10730: out = 16'(1555);
			10731: out = 16'(-9180);
			10732: out = 16'(-3172);
			10733: out = 16'(-1939);
			10734: out = 16'(1971);
			10735: out = 16'(851);
			10736: out = 16'(2036);
			10737: out = 16'(-4484);
			10738: out = 16'(-1394);
			10739: out = 16'(-246);
			10740: out = 16'(434);
			10741: out = 16'(-911);
			10742: out = 16'(8654);
			10743: out = 16'(8072);
			10744: out = 16'(-1286);
			10745: out = 16'(-6964);
			10746: out = 16'(1669);
			10747: out = 16'(5043);
			10748: out = 16'(-1057);
			10749: out = 16'(-3572);
			10750: out = 16'(1503);
			10751: out = 16'(4303);
			10752: out = 16'(-3559);
			10753: out = 16'(-12902);
			10754: out = 16'(-5573);
			10755: out = 16'(2023);
			10756: out = 16'(1536);
			10757: out = 16'(750);
			10758: out = 16'(3093);
			10759: out = 16'(5292);
			10760: out = 16'(1364);
			10761: out = 16'(1158);
			10762: out = 16'(2409);
			10763: out = 16'(8043);
			10764: out = 16'(-4243);
			10765: out = 16'(-13329);
			10766: out = 16'(2249);
			10767: out = 16'(9462);
			10768: out = 16'(-2976);
			10769: out = 16'(-11011);
			10770: out = 16'(7973);
			10771: out = 16'(13762);
			10772: out = 16'(1382);
			10773: out = 16'(-9406);
			10774: out = 16'(4020);
			10775: out = 16'(7813);
			10776: out = 16'(2255);
			10777: out = 16'(-8808);
			10778: out = 16'(-5068);
			10779: out = 16'(-830);
			10780: out = 16'(5014);
			10781: out = 16'(-1104);
			10782: out = 16'(-6524);
			10783: out = 16'(-9472);
			10784: out = 16'(3617);
			10785: out = 16'(5591);
			10786: out = 16'(1557);
			10787: out = 16'(40);
			10788: out = 16'(7566);
			10789: out = 16'(4597);
			10790: out = 16'(-2756);
			10791: out = 16'(-3891);
			10792: out = 16'(1251);
			10793: out = 16'(-773);
			10794: out = 16'(-9104);
			10795: out = 16'(-12831);
			10796: out = 16'(-6982);
			10797: out = 16'(8485);
			10798: out = 16'(19373);
			10799: out = 16'(17329);
			10800: out = 16'(-201);
			10801: out = 16'(-14537);
			10802: out = 16'(-17802);
			10803: out = 16'(-6361);
			10804: out = 16'(-1036);
			10805: out = 16'(10101);
			10806: out = 16'(4133);
			10807: out = 16'(-549);
			10808: out = 16'(-406);
			10809: out = 16'(11105);
			10810: out = 16'(-3546);
			10811: out = 16'(-14668);
			10812: out = 16'(-5217);
			10813: out = 16'(2800);
			10814: out = 16'(-1574);
			10815: out = 16'(-5495);
			10816: out = 16'(1872);
			10817: out = 16'(1946);
			10818: out = 16'(4554);
			10819: out = 16'(5113);
			10820: out = 16'(9547);
			10821: out = 16'(11163);
			10822: out = 16'(4122);
			10823: out = 16'(-6125);
			10824: out = 16'(-12569);
			10825: out = 16'(-16891);
			10826: out = 16'(-2437);
			10827: out = 16'(2071);
			10828: out = 16'(-492);
			10829: out = 16'(-5349);
			10830: out = 16'(6183);
			10831: out = 16'(1275);
			10832: out = 16'(-6560);
			10833: out = 16'(-8427);
			10834: out = 16'(6437);
			10835: out = 16'(8811);
			10836: out = 16'(8639);
			10837: out = 16'(6240);
			10838: out = 16'(10946);
			10839: out = 16'(3720);
			10840: out = 16'(6443);
			10841: out = 16'(-1512);
			10842: out = 16'(-26349);
			10843: out = 16'(-30840);
			10844: out = 16'(-6035);
			10845: out = 16'(17064);
			10846: out = 16'(7808);
			10847: out = 16'(-12861);
			10848: out = 16'(-10809);
			10849: out = 16'(10518);
			10850: out = 16'(12310);
			10851: out = 16'(3836);
			10852: out = 16'(-19226);
			10853: out = 16'(-15346);
			10854: out = 16'(6472);
			10855: out = 16'(3786);
			10856: out = 16'(5226);
			10857: out = 16'(6391);
			10858: out = 16'(10387);
			10859: out = 16'(8177);
			10860: out = 16'(3006);
			10861: out = 16'(-6457);
			10862: out = 16'(-8371);
			10863: out = 16'(682);
			10864: out = 16'(2593);
			10865: out = 16'(1808);
			10866: out = 16'(-330);
			10867: out = 16'(1091);
			10868: out = 16'(6932);
			10869: out = 16'(4076);
			10870: out = 16'(-5029);
			10871: out = 16'(-8893);
			10872: out = 16'(-1080);
			10873: out = 16'(7762);
			10874: out = 16'(6122);
			10875: out = 16'(-327);
			10876: out = 16'(-4385);
			10877: out = 16'(-722);
			10878: out = 16'(-3540);
			10879: out = 16'(-6484);
			10880: out = 16'(1078);
			10881: out = 16'(8455);
			10882: out = 16'(11006);
			10883: out = 16'(8095);
			10884: out = 16'(3140);
			10885: out = 16'(498);
			10886: out = 16'(-5770);
			10887: out = 16'(-5066);
			10888: out = 16'(1589);
			10889: out = 16'(-2940);
			10890: out = 16'(-9311);
			10891: out = 16'(-9783);
			10892: out = 16'(678);
			10893: out = 16'(9185);
			10894: out = 16'(6656);
			10895: out = 16'(969);
			10896: out = 16'(489);
			10897: out = 16'(1089);
			10898: out = 16'(6089);
			10899: out = 16'(3764);
			10900: out = 16'(-1556);
			10901: out = 16'(-7604);
			10902: out = 16'(167);
			10903: out = 16'(408);
			10904: out = 16'(-385);
			10905: out = 16'(15);
			10906: out = 16'(5161);
			10907: out = 16'(3204);
			10908: out = 16'(3295);
			10909: out = 16'(1927);
			10910: out = 16'(-8135);
			10911: out = 16'(-8417);
			10912: out = 16'(1734);
			10913: out = 16'(8111);
			10914: out = 16'(-394);
			10915: out = 16'(-3144);
			10916: out = 16'(1806);
			10917: out = 16'(6702);
			10918: out = 16'(2936);
			10919: out = 16'(-5948);
			10920: out = 16'(-7535);
			10921: out = 16'(-6672);
			10922: out = 16'(-9343);
			10923: out = 16'(-10471);
			10924: out = 16'(455);
			10925: out = 16'(9674);
			10926: out = 16'(7430);
			10927: out = 16'(942);
			10928: out = 16'(2305);
			10929: out = 16'(4253);
			10930: out = 16'(1537);
			10931: out = 16'(3);
			10932: out = 16'(-801);
			10933: out = 16'(539);
			10934: out = 16'(1888);
			10935: out = 16'(3414);
			10936: out = 16'(-5424);
			10937: out = 16'(-10485);
			10938: out = 16'(-8304);
			10939: out = 16'(-2709);
			10940: out = 16'(3002);
			10941: out = 16'(-5142);
			10942: out = 16'(-8113);
			10943: out = 16'(5244);
			10944: out = 16'(12801);
			10945: out = 16'(11014);
			10946: out = 16'(65);
			10947: out = 16'(-2921);
			10948: out = 16'(1483);
			10949: out = 16'(7240);
			10950: out = 16'(-1469);
			10951: out = 16'(-8651);
			10952: out = 16'(-1525);
			10953: out = 16'(4672);
			10954: out = 16'(2215);
			10955: out = 16'(2036);
			10956: out = 16'(8960);
			10957: out = 16'(9268);
			10958: out = 16'(-1499);
			10959: out = 16'(-8513);
			10960: out = 16'(-4524);
			10961: out = 16'(-7544);
			10962: out = 16'(-10423);
			10963: out = 16'(-2986);
			10964: out = 16'(12179);
			10965: out = 16'(7863);
			10966: out = 16'(7547);
			10967: out = 16'(5243);
			10968: out = 16'(1741);
			10969: out = 16'(-16302);
			10970: out = 16'(-11905);
			10971: out = 16'(-5778);
			10972: out = 16'(4372);
			10973: out = 16'(10412);
			10974: out = 16'(7760);
			10975: out = 16'(3627);
			10976: out = 16'(5114);
			10977: out = 16'(4137);
			10978: out = 16'(-5619);
			10979: out = 16'(-15098);
			10980: out = 16'(-9958);
			10981: out = 16'(459);
			10982: out = 16'(301);
			10983: out = 16'(-7746);
			10984: out = 16'(-104);
			10985: out = 16'(13754);
			10986: out = 16'(5246);
			10987: out = 16'(1946);
			10988: out = 16'(-2290);
			10989: out = 16'(-5697);
			10990: out = 16'(-15117);
			10991: out = 16'(818);
			10992: out = 16'(7319);
			10993: out = 16'(2205);
			10994: out = 16'(-6526);
			10995: out = 16'(6973);
			10996: out = 16'(9296);
			10997: out = 16'(-2350);
			10998: out = 16'(-17510);
			10999: out = 16'(-10997);
			11000: out = 16'(356);
			11001: out = 16'(4090);
			11002: out = 16'(-1545);
			11003: out = 16'(-6436);
			11004: out = 16'(3176);
			11005: out = 16'(9114);
			11006: out = 16'(5224);
			11007: out = 16'(-2640);
			11008: out = 16'(1667);
			11009: out = 16'(3556);
			11010: out = 16'(-509);
			11011: out = 16'(-10637);
			11012: out = 16'(2278);
			11013: out = 16'(-3270);
			11014: out = 16'(-6083);
			11015: out = 16'(2328);
			11016: out = 16'(12772);
			11017: out = 16'(5090);
			11018: out = 16'(-3089);
			11019: out = 16'(-4217);
			11020: out = 16'(-4300);
			11021: out = 16'(-1361);
			11022: out = 16'(6659);
			11023: out = 16'(11369);
			11024: out = 16'(402);
			11025: out = 16'(-982);
			11026: out = 16'(332);
			11027: out = 16'(1883);
			11028: out = 16'(-5613);
			11029: out = 16'(-7804);
			11030: out = 16'(-4659);
			11031: out = 16'(2692);
			11032: out = 16'(-645);
			11033: out = 16'(-2136);
			11034: out = 16'(-3834);
			11035: out = 16'(7826);
			11036: out = 16'(13955);
			11037: out = 16'(18040);
			11038: out = 16'(-8193);
			11039: out = 16'(-10976);
			11040: out = 16'(1571);
			11041: out = 16'(2644);
			11042: out = 16'(-5249);
			11043: out = 16'(2925);
			11044: out = 16'(8395);
			11045: out = 16'(-8153);
			11046: out = 16'(-7368);
			11047: out = 16'(8428);
			11048: out = 16'(14268);
			11049: out = 16'(-4768);
			11050: out = 16'(-11883);
			11051: out = 16'(-7499);
			11052: out = 16'(-700);
			11053: out = 16'(-5176);
			11054: out = 16'(648);
			11055: out = 16'(875);
			11056: out = 16'(783);
			11057: out = 16'(2408);
			11058: out = 16'(12801);
			11059: out = 16'(12888);
			11060: out = 16'(-1157);
			11061: out = 16'(-14122);
			11062: out = 16'(-2177);
			11063: out = 16'(489);
			11064: out = 16'(-4871);
			11065: out = 16'(-13036);
			11066: out = 16'(-4843);
			11067: out = 16'(3917);
			11068: out = 16'(8825);
			11069: out = 16'(3202);
			11070: out = 16'(1441);
			11071: out = 16'(7273);
			11072: out = 16'(9072);
			11073: out = 16'(-1333);
			11074: out = 16'(-9718);
			11075: out = 16'(-1159);
			11076: out = 16'(10042);
			11077: out = 16'(5711);
			11078: out = 16'(-8999);
			11079: out = 16'(-15778);
			11080: out = 16'(-8609);
			11081: out = 16'(5125);
			11082: out = 16'(12599);
			11083: out = 16'(11478);
			11084: out = 16'(9755);
			11085: out = 16'(1178);
			11086: out = 16'(-3892);
			11087: out = 16'(-414);
			11088: out = 16'(-4930);
			11089: out = 16'(-6655);
			11090: out = 16'(-7833);
			11091: out = 16'(-5279);
			11092: out = 16'(-3471);
			11093: out = 16'(4643);
			11094: out = 16'(12568);
			11095: out = 16'(14160);
			11096: out = 16'(-910);
			11097: out = 16'(-6899);
			11098: out = 16'(-7704);
			11099: out = 16'(1398);
			11100: out = 16'(691);
			11101: out = 16'(10364);
			11102: out = 16'(-5957);
			11103: out = 16'(-12623);
			11104: out = 16'(2563);
			11105: out = 16'(9596);
			11106: out = 16'(-2884);
			11107: out = 16'(-9151);
			11108: out = 16'(2912);
			11109: out = 16'(3087);
			11110: out = 16'(-2690);
			11111: out = 16'(-4171);
			11112: out = 16'(3878);
			11113: out = 16'(-1368);
			11114: out = 16'(-1987);
			11115: out = 16'(-1968);
			11116: out = 16'(2246);
			11117: out = 16'(-1339);
			11118: out = 16'(-741);
			11119: out = 16'(-1755);
			11120: out = 16'(1995);
			11121: out = 16'(3357);
			11122: out = 16'(6992);
			11123: out = 16'(157);
			11124: out = 16'(-4714);
			11125: out = 16'(-6457);
			11126: out = 16'(-2856);
			11127: out = 16'(-10565);
			11128: out = 16'(-10851);
			11129: out = 16'(-151);
			11130: out = 16'(5973);
			11131: out = 16'(7348);
			11132: out = 16'(6183);
			11133: out = 16'(8130);
			11134: out = 16'(13947);
			11135: out = 16'(2848);
			11136: out = 16'(-6068);
			11137: out = 16'(-14431);
			11138: out = 16'(-22916);
			11139: out = 16'(-16119);
			11140: out = 16'(-303);
			11141: out = 16'(13032);
			11142: out = 16'(15462);
			11143: out = 16'(1620);
			11144: out = 16'(-937);
			11145: out = 16'(815);
			11146: out = 16'(789);
			11147: out = 16'(-5680);
			11148: out = 16'(-5740);
			11149: out = 16'(-6177);
			11150: out = 16'(-4219);
			11151: out = 16'(82);
			11152: out = 16'(11673);
			11153: out = 16'(9848);
			11154: out = 16'(758);
			11155: out = 16'(-7410);
			11156: out = 16'(-624);
			11157: out = 16'(-4598);
			11158: out = 16'(-7537);
			11159: out = 16'(1637);
			11160: out = 16'(8264);
			11161: out = 16'(4262);
			11162: out = 16'(-1588);
			11163: out = 16'(2108);
			11164: out = 16'(12337);
			11165: out = 16'(5238);
			11166: out = 16'(-6326);
			11167: out = 16'(-8038);
			11168: out = 16'(6123);
			11169: out = 16'(1912);
			11170: out = 16'(1936);
			11171: out = 16'(8933);
			11172: out = 16'(10762);
			11173: out = 16'(1565);
			11174: out = 16'(-7051);
			11175: out = 16'(-5516);
			11176: out = 16'(-386);
			11177: out = 16'(2711);
			11178: out = 16'(249);
			11179: out = 16'(-289);
			11180: out = 16'(-519);
			11181: out = 16'(1550);
			11182: out = 16'(5743);
			11183: out = 16'(13462);
			11184: out = 16'(9470);
			11185: out = 16'(-5686);
			11186: out = 16'(-23534);
			11187: out = 16'(-14157);
			11188: out = 16'(5122);
			11189: out = 16'(3160);
			11190: out = 16'(-12791);
			11191: out = 16'(-8675);
			11192: out = 16'(8937);
			11193: out = 16'(8111);
			11194: out = 16'(3762);
			11195: out = 16'(-874);
			11196: out = 16'(-93);
			11197: out = 16'(-4794);
			11198: out = 16'(-8943);
			11199: out = 16'(-11853);
			11200: out = 16'(-5544);
			11201: out = 16'(1683);
			11202: out = 16'(-5434);
			11203: out = 16'(1296);
			11204: out = 16'(6587);
			11205: out = 16'(5628);
			11206: out = 16'(320);
			11207: out = 16'(227);
			11208: out = 16'(-3438);
			11209: out = 16'(-7824);
			11210: out = 16'(-4796);
			11211: out = 16'(35);
			11212: out = 16'(6972);
			11213: out = 16'(7560);
			11214: out = 16'(-911);
			11215: out = 16'(-1574);
			11216: out = 16'(-6516);
			11217: out = 16'(-4481);
			11218: out = 16'(960);
			11219: out = 16'(3384);
			11220: out = 16'(-2042);
			11221: out = 16'(-2973);
			11222: out = 16'(1563);
			11223: out = 16'(7069);
			11224: out = 16'(4535);
			11225: out = 16'(6887);
			11226: out = 16'(7448);
			11227: out = 16'(-79);
			11228: out = 16'(-4147);
			11229: out = 16'(-2063);
			11230: out = 16'(-1948);
			11231: out = 16'(-7250);
			11232: out = 16'(-5586);
			11233: out = 16'(6053);
			11234: out = 16'(9643);
			11235: out = 16'(-828);
			11236: out = 16'(-11939);
			11237: out = 16'(-1362);
			11238: out = 16'(10678);
			11239: out = 16'(6350);
			11240: out = 16'(1488);
			11241: out = 16'(-8393);
			11242: out = 16'(-10341);
			11243: out = 16'(-6192);
			11244: out = 16'(6146);
			11245: out = 16'(10020);
			11246: out = 16'(10132);
			11247: out = 16'(2732);
			11248: out = 16'(-4410);
			11249: out = 16'(-14499);
			11250: out = 16'(-10283);
			11251: out = 16'(-3672);
			11252: out = 16'(-173);
			11253: out = 16'(8186);
			11254: out = 16'(8991);
			11255: out = 16'(1545);
			11256: out = 16'(-6065);
			11257: out = 16'(-6164);
			11258: out = 16'(3844);
			11259: out = 16'(5282);
			11260: out = 16'(2214);
			11261: out = 16'(8956);
			11262: out = 16'(5941);
			11263: out = 16'(-5805);
			11264: out = 16'(-14355);
			11265: out = 16'(1440);
			11266: out = 16'(2623);
			11267: out = 16'(4633);
			11268: out = 16'(962);
			11269: out = 16'(1523);
			11270: out = 16'(6945);
			11271: out = 16'(10630);
			11272: out = 16'(1880);
			11273: out = 16'(-10035);
			11274: out = 16'(-11003);
			11275: out = 16'(435);
			11276: out = 16'(6238);
			11277: out = 16'(2223);
			11278: out = 16'(-2711);
			11279: out = 16'(-1143);
			11280: out = 16'(152);
			11281: out = 16'(-73);
			11282: out = 16'(2876);
			11283: out = 16'(1524);
			11284: out = 16'(408);
			11285: out = 16'(1403);
			11286: out = 16'(6698);
			11287: out = 16'(3889);
			11288: out = 16'(2098);
			11289: out = 16'(48);
			11290: out = 16'(-848);
			11291: out = 16'(-10027);
			11292: out = 16'(-4336);
			11293: out = 16'(3352);
			11294: out = 16'(3453);
			11295: out = 16'(-5138);
			11296: out = 16'(-7210);
			11297: out = 16'(927);
			11298: out = 16'(9964);
			11299: out = 16'(5405);
			11300: out = 16'(1993);
			11301: out = 16'(-4070);
			11302: out = 16'(-7333);
			11303: out = 16'(-12522);
			11304: out = 16'(-3766);
			11305: out = 16'(-4020);
			11306: out = 16'(-1516);
			11307: out = 16'(4566);
			11308: out = 16'(7195);
			11309: out = 16'(-2630);
			11310: out = 16'(-3852);
			11311: out = 16'(8119);
			11312: out = 16'(643);
			11313: out = 16'(1024);
			11314: out = 16'(-997);
			11315: out = 16'(-1105);
			11316: out = 16'(-12454);
			11317: out = 16'(-4431);
			11318: out = 16'(-2815);
			11319: out = 16'(-790);
			11320: out = 16'(4425);
			11321: out = 16'(11021);
			11322: out = 16'(5589);
			11323: out = 16'(-2331);
			11324: out = 16'(-5582);
			11325: out = 16'(-118);
			11326: out = 16'(-7257);
			11327: out = 16'(-15609);
			11328: out = 16'(-11715);
			11329: out = 16'(7619);
			11330: out = 16'(12151);
			11331: out = 16'(11682);
			11332: out = 16'(12890);
			11333: out = 16'(11701);
			11334: out = 16'(1857);
			11335: out = 16'(-11696);
			11336: out = 16'(-16428);
			11337: out = 16'(637);
			11338: out = 16'(5064);
			11339: out = 16'(6909);
			11340: out = 16'(480);
			11341: out = 16'(-5503);
			11342: out = 16'(-24909);
			11343: out = 16'(-7402);
			11344: out = 16'(17857);
			11345: out = 16'(17484);
			11346: out = 16'(-8817);
			11347: out = 16'(-8185);
			11348: out = 16'(9667);
			11349: out = 16'(12776);
			11350: out = 16'(-10727);
			11351: out = 16'(-5906);
			11352: out = 16'(12123);
			11353: out = 16'(14164);
			11354: out = 16'(-2236);
			11355: out = 16'(-20981);
			11356: out = 16'(-17933);
			11357: out = 16'(745);
			11358: out = 16'(11117);
			11359: out = 16'(10074);
			11360: out = 16'(7537);
			11361: out = 16'(5421);
			11362: out = 16'(1349);
			11363: out = 16'(-17552);
			11364: out = 16'(-11810);
			11365: out = 16'(3610);
			11366: out = 16'(4138);
			11367: out = 16'(-9094);
			11368: out = 16'(-12987);
			11369: out = 16'(-800);
			11370: out = 16'(9481);
			11371: out = 16'(2157);
			11372: out = 16'(7099);
			11373: out = 16'(11668);
			11374: out = 16'(7428);
			11375: out = 16'(-5823);
			11376: out = 16'(-7860);
			11377: out = 16'(-6689);
			11378: out = 16'(-10235);
			11379: out = 16'(-14606);
			11380: out = 16'(7160);
			11381: out = 16'(18194);
			11382: out = 16'(8133);
			11383: out = 16'(-6082);
			11384: out = 16'(9150);
			11385: out = 16'(15970);
			11386: out = 16'(585);
			11387: out = 16'(-25903);
			11388: out = 16'(-27978);
			11389: out = 16'(-11145);
			11390: out = 16'(4253);
			11391: out = 16'(5892);
			11392: out = 16'(7579);
			11393: out = 16'(3197);
			11394: out = 16'(-1590);
			11395: out = 16'(-644);
			11396: out = 16'(12744);
			11397: out = 16'(11293);
			11398: out = 16'(3995);
			11399: out = 16'(-7292);
			11400: out = 16'(-8403);
			11401: out = 16'(758);
			11402: out = 16'(4912);
			11403: out = 16'(-2694);
			11404: out = 16'(-8651);
			11405: out = 16'(3438);
			11406: out = 16'(6555);
			11407: out = 16'(-250);
			11408: out = 16'(-5498);
			11409: out = 16'(9835);
			11410: out = 16'(7084);
			11411: out = 16'(3695);
			11412: out = 16'(-869);
			11413: out = 16'(1504);
			11414: out = 16'(-10701);
			11415: out = 16'(-9901);
			11416: out = 16'(-4901);
			11417: out = 16'(1407);
			11418: out = 16'(-599);
			11419: out = 16'(8464);
			11420: out = 16'(8385);
			11421: out = 16'(-216);
			11422: out = 16'(-9559);
			11423: out = 16'(4630);
			11424: out = 16'(11671);
			11425: out = 16'(2003);
			11426: out = 16'(-12200);
			11427: out = 16'(-10761);
			11428: out = 16'(-7221);
			11429: out = 16'(-5759);
			11430: out = 16'(1726);
			11431: out = 16'(13878);
			11432: out = 16'(12972);
			11433: out = 16'(922);
			11434: out = 16'(-6905);
			11435: out = 16'(-13429);
			11436: out = 16'(-5434);
			11437: out = 16'(5103);
			11438: out = 16'(10791);
			11439: out = 16'(727);
			11440: out = 16'(-7249);
			11441: out = 16'(-13609);
			11442: out = 16'(-7775);
			11443: out = 16'(2997);
			11444: out = 16'(11747);
			11445: out = 16'(6139);
			11446: out = 16'(3291);
			11447: out = 16'(8270);
			11448: out = 16'(13476);
			11449: out = 16'(-3993);
			11450: out = 16'(-19668);
			11451: out = 16'(-10104);
			11452: out = 16'(-966);
			11453: out = 16'(-10808);
			11454: out = 16'(-21102);
			11455: out = 16'(-2667);
			11456: out = 16'(11447);
			11457: out = 16'(19425);
			11458: out = 16'(10512);
			11459: out = 16'(4135);
			11460: out = 16'(-3572);
			11461: out = 16'(8930);
			11462: out = 16'(5791);
			11463: out = 16'(-7060);
			11464: out = 16'(-21030);
			11465: out = 16'(-8173);
			11466: out = 16'(1193);
			11467: out = 16'(9086);
			11468: out = 16'(18904);
			11469: out = 16'(14077);
			11470: out = 16'(-1652);
			11471: out = 16'(-14346);
			11472: out = 16'(-11685);
			11473: out = 16'(-5323);
			11474: out = 16'(-1);
			11475: out = 16'(3384);
			11476: out = 16'(4001);
			11477: out = 16'(4088);
			11478: out = 16'(-6911);
			11479: out = 16'(-2667);
			11480: out = 16'(11855);
			11481: out = 16'(10101);
			11482: out = 16'(-4114);
			11483: out = 16'(-10479);
			11484: out = 16'(-3337);
			11485: out = 16'(-6786);
			11486: out = 16'(-312);
			11487: out = 16'(-1238);
			11488: out = 16'(3903);
			11489: out = 16'(5867);
			11490: out = 16'(8667);
			11491: out = 16'(-7084);
			11492: out = 16'(-13626);
			11493: out = 16'(-5150);
			11494: out = 16'(493);
			11495: out = 16'(2107);
			11496: out = 16'(10023);
			11497: out = 16'(18864);
			11498: out = 16'(14932);
			11499: out = 16'(1909);
			11500: out = 16'(-7025);
			11501: out = 16'(-9500);
			11502: out = 16'(-11417);
			11503: out = 16'(-13424);
			11504: out = 16'(-5008);
			11505: out = 16'(3524);
			11506: out = 16'(1925);
			11507: out = 16'(4081);
			11508: out = 16'(12782);
			11509: out = 16'(16086);
			11510: out = 16'(4516);
			11511: out = 16'(-8931);
			11512: out = 16'(-13298);
			11513: out = 16'(-10516);
			11514: out = 16'(-11412);
			11515: out = 16'(-2986);
			11516: out = 16'(371);
			11517: out = 16'(9984);
			11518: out = 16'(14269);
			11519: out = 16'(11370);
			11520: out = 16'(-157);
			11521: out = 16'(-3405);
			11522: out = 16'(-3688);
			11523: out = 16'(-6933);
			11524: out = 16'(-6249);
			11525: out = 16'(542);
			11526: out = 16'(4581);
			11527: out = 16'(747);
			11528: out = 16'(-3228);
			11529: out = 16'(-658);
			11530: out = 16'(3517);
			11531: out = 16'(4388);
			11532: out = 16'(4261);
			11533: out = 16'(3905);
			11534: out = 16'(-1841);
			11535: out = 16'(-7636);
			11536: out = 16'(4660);
			11537: out = 16'(1281);
			11538: out = 16'(-611);
			11539: out = 16'(170);
			11540: out = 16'(6854);
			11541: out = 16'(-2380);
			11542: out = 16'(-2205);
			11543: out = 16'(4497);
			11544: out = 16'(7719);
			11545: out = 16'(-7003);
			11546: out = 16'(-6511);
			11547: out = 16'(8097);
			11548: out = 16'(13077);
			11549: out = 16'(-9387);
			11550: out = 16'(-18883);
			11551: out = 16'(-3484);
			11552: out = 16'(13197);
			11553: out = 16'(747);
			11554: out = 16'(-5198);
			11555: out = 16'(1929);
			11556: out = 16'(12500);
			11557: out = 16'(9880);
			11558: out = 16'(-14452);
			11559: out = 16'(-19983);
			11560: out = 16'(-1165);
			11561: out = 16'(14043);
			11562: out = 16'(14205);
			11563: out = 16'(5428);
			11564: out = 16'(-5080);
			11565: out = 16'(-11441);
			11566: out = 16'(-9830);
			11567: out = 16'(5532);
			11568: out = 16'(13183);
			11569: out = 16'(4970);
			11570: out = 16'(-13033);
			11571: out = 16'(-12017);
			11572: out = 16'(-3858);
			11573: out = 16'(564);
			11574: out = 16'(524);
			11575: out = 16'(16035);
			11576: out = 16'(16678);
			11577: out = 16'(-147);
			11578: out = 16'(-23854);
			11579: out = 16'(-17929);
			11580: out = 16'(-6423);
			11581: out = 16'(2781);
			11582: out = 16'(10469);
			11583: out = 16'(15759);
			11584: out = 16'(9765);
			11585: out = 16'(-1968);
			11586: out = 16'(-8117);
			11587: out = 16'(-3803);
			11588: out = 16'(-4671);
			11589: out = 16'(-10717);
			11590: out = 16'(-10588);
			11591: out = 16'(10);
			11592: out = 16'(9969);
			11593: out = 16'(9163);
			11594: out = 16'(4312);
			11595: out = 16'(1370);
			11596: out = 16'(4104);
			11597: out = 16'(1773);
			11598: out = 16'(-478);
			11599: out = 16'(-2262);
			11600: out = 16'(-2759);
			11601: out = 16'(-12737);
			11602: out = 16'(-9884);
			11603: out = 16'(9614);
			11604: out = 16'(11398);
			11605: out = 16'(6890);
			11606: out = 16'(5);
			11607: out = 16'(-2279);
			11608: out = 16'(-11539);
			11609: out = 16'(-3215);
			11610: out = 16'(2612);
			11611: out = 16'(3334);
			11612: out = 16'(7578);
			11613: out = 16'(5552);
			11614: out = 16'(11194);
			11615: out = 16'(9444);
			11616: out = 16'(-2656);
			11617: out = 16'(-17993);
			11618: out = 16'(-9853);
			11619: out = 16'(2734);
			11620: out = 16'(-1712);
			11621: out = 16'(-2660);
			11622: out = 16'(-727);
			11623: out = 16'(6951);
			11624: out = 16'(7383);
			11625: out = 16'(988);
			11626: out = 16'(778);
			11627: out = 16'(6987);
			11628: out = 16'(7797);
			11629: out = 16'(-1559);
			11630: out = 16'(-6729);
			11631: out = 16'(-4186);
			11632: out = 16'(1579);
			11633: out = 16'(2562);
			11634: out = 16'(8127);
			11635: out = 16'(5083);
			11636: out = 16'(-2898);
			11637: out = 16'(-10160);
			11638: out = 16'(-4139);
			11639: out = 16'(-2402);
			11640: out = 16'(-4827);
			11641: out = 16'(-6333);
			11642: out = 16'(1043);
			11643: out = 16'(1012);
			11644: out = 16'(-1243);
			11645: out = 16'(182);
			11646: out = 16'(6222);
			11647: out = 16'(7017);
			11648: out = 16'(3859);
			11649: out = 16'(-441);
			11650: out = 16'(-7905);
			11651: out = 16'(-6673);
			11652: out = 16'(-10247);
			11653: out = 16'(-9296);
			11654: out = 16'(-1200);
			11655: out = 16'(15127);
			11656: out = 16'(8463);
			11657: out = 16'(-3334);
			11658: out = 16'(-7466);
			11659: out = 16'(3435);
			11660: out = 16'(5946);
			11661: out = 16'(7416);
			11662: out = 16'(3220);
			11663: out = 16'(-11574);
			11664: out = 16'(-14307);
			11665: out = 16'(-647);
			11666: out = 16'(8542);
			11667: out = 16'(596);
			11668: out = 16'(-8877);
			11669: out = 16'(1159);
			11670: out = 16'(11917);
			11671: out = 16'(2073);
			11672: out = 16'(-15492);
			11673: out = 16'(-13369);
			11674: out = 16'(3146);
			11675: out = 16'(8877);
			11676: out = 16'(9845);
			11677: out = 16'(9536);
			11678: out = 16'(7097);
			11679: out = 16'(-3295);
			11680: out = 16'(-13361);
			11681: out = 16'(-7691);
			11682: out = 16'(827);
			11683: out = 16'(-702);
			11684: out = 16'(1817);
			11685: out = 16'(-993);
			11686: out = 16'(5067);
			11687: out = 16'(3985);
			11688: out = 16'(-3302);
			11689: out = 16'(-2002);
			11690: out = 16'(9411);
			11691: out = 16'(8651);
			11692: out = 16'(-7715);
			11693: out = 16'(-19687);
			11694: out = 16'(-9455);
			11695: out = 16'(8176);
			11696: out = 16'(13405);
			11697: out = 16'(14658);
			11698: out = 16'(7287);
			11699: out = 16'(-2960);
			11700: out = 16'(-13844);
			11701: out = 16'(-15920);
			11702: out = 16'(-13390);
			11703: out = 16'(-5648);
			11704: out = 16'(6315);
			11705: out = 16'(19690);
			11706: out = 16'(7847);
			11707: out = 16'(-6187);
			11708: out = 16'(-11585);
			11709: out = 16'(581);
			11710: out = 16'(3011);
			11711: out = 16'(6942);
			11712: out = 16'(4794);
			11713: out = 16'(1447);
			11714: out = 16'(170);
			11715: out = 16'(-3222);
			11716: out = 16'(-7408);
			11717: out = 16'(-4439);
			11718: out = 16'(4702);
			11719: out = 16'(15012);
			11720: out = 16'(10293);
			11721: out = 16'(-2468);
			11722: out = 16'(-9476);
			11723: out = 16'(-9801);
			11724: out = 16'(-4286);
			11725: out = 16'(4257);
			11726: out = 16'(13062);
			11727: out = 16'(1851);
			11728: out = 16'(-5825);
			11729: out = 16'(-8647);
			11730: out = 16'(-4209);
			11731: out = 16'(1994);
			11732: out = 16'(6205);
			11733: out = 16'(5845);
			11734: out = 16'(3660);
			11735: out = 16'(1514);
			11736: out = 16'(-6258);
			11737: out = 16'(-12992);
			11738: out = 16'(-9756);
			11739: out = 16'(2724);
			11740: out = 16'(2895);
			11741: out = 16'(1621);
			11742: out = 16'(5551);
			11743: out = 16'(7771);
			11744: out = 16'(-508);
			11745: out = 16'(-13017);
			11746: out = 16'(-10796);
			11747: out = 16'(3617);
			11748: out = 16'(1528);
			11749: out = 16'(-9624);
			11750: out = 16'(-9000);
			11751: out = 16'(6971);
			11752: out = 16'(3987);
			11753: out = 16'(4190);
			11754: out = 16'(5882);
			11755: out = 16'(10091);
			11756: out = 16'(-231);
			11757: out = 16'(-215);
			11758: out = 16'(-1367);
			11759: out = 16'(950);
			11760: out = 16'(-493);
			11761: out = 16'(4339);
			11762: out = 16'(2498);
			11763: out = 16'(192);
			11764: out = 16'(-4784);
			11765: out = 16'(860);
			11766: out = 16'(-4610);
			11767: out = 16'(-4998);
			11768: out = 16'(1315);
			11769: out = 16'(9036);
			11770: out = 16'(2938);
			11771: out = 16'(210);
			11772: out = 16'(1350);
			11773: out = 16'(-714);
			11774: out = 16'(-1652);
			11775: out = 16'(7896);
			11776: out = 16'(9809);
			11777: out = 16'(-16357);
			11778: out = 16'(-18896);
			11779: out = 16'(-5292);
			11780: out = 16'(8466);
			11781: out = 16'(-1040);
			11782: out = 16'(7235);
			11783: out = 16'(7136);
			11784: out = 16'(6671);
			11785: out = 16'(-1709);
			11786: out = 16'(248);
			11787: out = 16'(-10911);
			11788: out = 16'(-11473);
			11789: out = 16'(812);
			11790: out = 16'(13569);
			11791: out = 16'(3639);
			11792: out = 16'(-9089);
			11793: out = 16'(-10157);
			11794: out = 16'(3043);
			11795: out = 16'(11771);
			11796: out = 16'(11212);
			11797: out = 16'(2815);
			11798: out = 16'(-5524);
			11799: out = 16'(-17788);
			11800: out = 16'(-13199);
			11801: out = 16'(-923);
			11802: out = 16'(3722);
			11803: out = 16'(13041);
			11804: out = 16'(18204);
			11805: out = 16'(18767);
			11806: out = 16'(6965);
			11807: out = 16'(-422);
			11808: out = 16'(-20590);
			11809: out = 16'(-23992);
			11810: out = 16'(-10947);
			11811: out = 16'(5512);
			11812: out = 16'(6141);
			11813: out = 16'(11405);
			11814: out = 16'(11662);
			11815: out = 16'(206);
			11816: out = 16'(-13067);
			11817: out = 16'(-1661);
			11818: out = 16'(16311);
			11819: out = 16'(10821);
			11820: out = 16'(-10668);
			11821: out = 16'(-20370);
			11822: out = 16'(-8634);
			11823: out = 16'(5613);
			11824: out = 16'(14147);
			11825: out = 16'(11660);
			11826: out = 16'(5152);
			11827: out = 16'(-5862);
			11828: out = 16'(-12070);
			11829: out = 16'(-19256);
			11830: out = 16'(-15594);
			11831: out = 16'(-4070);
			11832: out = 16'(9738);
			11833: out = 16'(15445);
			11834: out = 16'(11594);
			11835: out = 16'(-6965);
			11836: out = 16'(-27670);
			11837: out = 16'(-10773);
			11838: out = 16'(9290);
			11839: out = 16'(4512);
			11840: out = 16'(-12428);
			11841: out = 16'(-8259);
			11842: out = 16'(5859);
			11843: out = 16'(3977);
			11844: out = 16'(-9831);
			11845: out = 16'(-2246);
			11846: out = 16'(10449);
			11847: out = 16'(8439);
			11848: out = 16'(-6902);
			11849: out = 16'(-7836);
			11850: out = 16'(-2364);
			11851: out = 16'(4961);
			11852: out = 16'(7264);
			11853: out = 16'(11633);
			11854: out = 16'(-2156);
			11855: out = 16'(-8934);
			11856: out = 16'(-5404);
			11857: out = 16'(4544);
			11858: out = 16'(-10184);
			11859: out = 16'(-9816);
			11860: out = 16'(5272);
			11861: out = 16'(18009);
			11862: out = 16'(2129);
			11863: out = 16'(-582);
			11864: out = 16'(7538);
			11865: out = 16'(14490);
			11866: out = 16'(-1373);
			11867: out = 16'(-6768);
			11868: out = 16'(-3126);
			11869: out = 16'(10450);
			11870: out = 16'(14665);
			11871: out = 16'(4772);
			11872: out = 16'(-11132);
			11873: out = 16'(-12089);
			11874: out = 16'(3765);
			11875: out = 16'(802);
			11876: out = 16'(1);
			11877: out = 16'(2796);
			11878: out = 16'(5695);
			11879: out = 16'(-7136);
			11880: out = 16'(-4466);
			11881: out = 16'(9439);
			11882: out = 16'(20043);
			11883: out = 16'(12389);
			11884: out = 16'(-1258);
			11885: out = 16'(-14782);
			11886: out = 16'(-15654);
			11887: out = 16'(-1156);
			11888: out = 16'(12332);
			11889: out = 16'(14949);
			11890: out = 16'(2712);
			11891: out = 16'(-20579);
			11892: out = 16'(-16281);
			11893: out = 16'(-11859);
			11894: out = 16'(-7172);
			11895: out = 16'(1463);
			11896: out = 16'(13981);
			11897: out = 16'(15943);
			11898: out = 16'(6573);
			11899: out = 16'(-3445);
			11900: out = 16'(-1726);
			11901: out = 16'(-1849);
			11902: out = 16'(-6101);
			11903: out = 16'(-5426);
			11904: out = 16'(9931);
			11905: out = 16'(6315);
			11906: out = 16'(-4073);
			11907: out = 16'(-12291);
			11908: out = 16'(-7420);
			11909: out = 16'(-421);
			11910: out = 16'(4125);
			11911: out = 16'(4352);
			11912: out = 16'(4270);
			11913: out = 16'(2026);
			11914: out = 16'(-1048);
			11915: out = 16'(-3312);
			11916: out = 16'(-1337);
			11917: out = 16'(6263);
			11918: out = 16'(5359);
			11919: out = 16'(2464);
			11920: out = 16'(-1338);
			11921: out = 16'(-8227);
			11922: out = 16'(-9040);
			11923: out = 16'(-5589);
			11924: out = 16'(-1372);
			11925: out = 16'(959);
			11926: out = 16'(4608);
			11927: out = 16'(8311);
			11928: out = 16'(8203);
			11929: out = 16'(4383);
			11930: out = 16'(-12239);
			11931: out = 16'(-7581);
			11932: out = 16'(7252);
			11933: out = 16'(13699);
			11934: out = 16'(7287);
			11935: out = 16'(1010);
			11936: out = 16'(-4777);
			11937: out = 16'(-9459);
			11938: out = 16'(-11150);
			11939: out = 16'(-2043);
			11940: out = 16'(4595);
			11941: out = 16'(2878);
			11942: out = 16'(-599);
			11943: out = 16'(-340);
			11944: out = 16'(1798);
			11945: out = 16'(982);
			11946: out = 16'(1080);
			11947: out = 16'(7139);
			11948: out = 16'(10607);
			11949: out = 16'(2359);
			11950: out = 16'(-10063);
			11951: out = 16'(-4124);
			11952: out = 16'(6989);
			11953: out = 16'(9626);
			11954: out = 16'(1152);
			11955: out = 16'(-9020);
			11956: out = 16'(-8102);
			11957: out = 16'(-2690);
			11958: out = 16'(402);
			11959: out = 16'(1520);
			11960: out = 16'(1702);
			11961: out = 16'(557);
			11962: out = 16'(540);
			11963: out = 16'(2860);
			11964: out = 16'(6086);
			11965: out = 16'(2992);
			11966: out = 16'(-1492);
			11967: out = 16'(-3346);
			11968: out = 16'(-6786);
			11969: out = 16'(-4677);
			11970: out = 16'(3228);
			11971: out = 16'(7951);
			11972: out = 16'(1152);
			11973: out = 16'(-2458);
			11974: out = 16'(5016);
			11975: out = 16'(12566);
			11976: out = 16'(4647);
			11977: out = 16'(-11206);
			11978: out = 16'(-16400);
			11979: out = 16'(-6237);
			11980: out = 16'(892);
			11981: out = 16'(12668);
			11982: out = 16'(13055);
			11983: out = 16'(6778);
			11984: out = 16'(-4502);
			11985: out = 16'(-11676);
			11986: out = 16'(-17241);
			11987: out = 16'(-15422);
			11988: out = 16'(-3968);
			11989: out = 16'(9339);
			11990: out = 16'(17550);
			11991: out = 16'(11669);
			11992: out = 16'(-1823);
			11993: out = 16'(-9190);
			11994: out = 16'(-797);
			11995: out = 16'(7141);
			11996: out = 16'(3560);
			11997: out = 16'(-3429);
			11998: out = 16'(1001);
			11999: out = 16'(7158);
			12000: out = 16'(-253);
			12001: out = 16'(-19500);
			12002: out = 16'(-6964);
			12003: out = 16'(4624);
			12004: out = 16'(2917);
			12005: out = 16'(-6565);
			12006: out = 16'(-12978);
			12007: out = 16'(-3178);
			12008: out = 16'(5779);
			12009: out = 16'(4166);
			12010: out = 16'(-1830);
			12011: out = 16'(1665);
			12012: out = 16'(7961);
			12013: out = 16'(11646);
			12014: out = 16'(11180);
			12015: out = 16'(323);
			12016: out = 16'(-13400);
			12017: out = 16'(-14089);
			12018: out = 16'(4188);
			12019: out = 16'(1315);
			12020: out = 16'(-5755);
			12021: out = 16'(-4900);
			12022: out = 16'(7229);
			12023: out = 16'(2029);
			12024: out = 16'(-5970);
			12025: out = 16'(-6827);
			12026: out = 16'(7767);
			12027: out = 16'(14308);
			12028: out = 16'(9224);
			12029: out = 16'(-9082);
			12030: out = 16'(-20228);
			12031: out = 16'(-4916);
			12032: out = 16'(2972);
			12033: out = 16'(5263);
			12034: out = 16'(10146);
			12035: out = 16'(19608);
			12036: out = 16'(108);
			12037: out = 16'(-22127);
			12038: out = 16'(-26024);
			12039: out = 16'(972);
			12040: out = 16'(10358);
			12041: out = 16'(13272);
			12042: out = 16'(6928);
			12043: out = 16'(-1587);
			12044: out = 16'(-19837);
			12045: out = 16'(-8933);
			12046: out = 16'(10386);
			12047: out = 16'(16009);
			12048: out = 16'(529);
			12049: out = 16'(-3616);
			12050: out = 16'(-2204);
			12051: out = 16'(1962);
			12052: out = 16'(-695);
			12053: out = 16'(968);
			12054: out = 16'(476);
			12055: out = 16'(6674);
			12056: out = 16'(11333);
			12057: out = 16'(-1127);
			12058: out = 16'(-18409);
			12059: out = 16'(-13717);
			12060: out = 16'(11522);
			12061: out = 16'(5921);
			12062: out = 16'(-1390);
			12063: out = 16'(914);
			12064: out = 16'(13208);
			12065: out = 16'(5703);
			12066: out = 16'(-6635);
			12067: out = 16'(-16332);
			12068: out = 16'(-10044);
			12069: out = 16'(-3975);
			12070: out = 16'(4166);
			12071: out = 16'(2652);
			12072: out = 16'(2405);
			12073: out = 16'(2320);
			12074: out = 16'(1694);
			12075: out = 16'(-3938);
			12076: out = 16'(-2481);
			12077: out = 16'(5737);
			12078: out = 16'(3487);
			12079: out = 16'(-946);
			12080: out = 16'(-2150);
			12081: out = 16'(-354);
			12082: out = 16'(-4908);
			12083: out = 16'(-1677);
			12084: out = 16'(8904);
			12085: out = 16'(12458);
			12086: out = 16'(-7902);
			12087: out = 16'(-12853);
			12088: out = 16'(-4614);
			12089: out = 16'(7204);
			12090: out = 16'(1783);
			12091: out = 16'(5906);
			12092: out = 16'(1622);
			12093: out = 16'(-4405);
			12094: out = 16'(-12813);
			12095: out = 16'(-1067);
			12096: out = 16'(256);
			12097: out = 16'(3033);
			12098: out = 16'(9855);
			12099: out = 16'(10568);
			12100: out = 16'(3906);
			12101: out = 16'(-1884);
			12102: out = 16'(901);
			12103: out = 16'(-1525);
			12104: out = 16'(-1565);
			12105: out = 16'(-11144);
			12106: out = 16'(-12526);
			12107: out = 16'(4171);
			12108: out = 16'(18518);
			12109: out = 16'(10868);
			12110: out = 16'(-5366);
			12111: out = 16'(-11917);
			12112: out = 16'(-2475);
			12113: out = 16'(1477);
			12114: out = 16'(-1251);
			12115: out = 16'(-2009);
			12116: out = 16'(3448);
			12117: out = 16'(1978);
			12118: out = 16'(-26);
			12119: out = 16'(2291);
			12120: out = 16'(5884);
			12121: out = 16'(2420);
			12122: out = 16'(-3570);
			12123: out = 16'(-7198);
			12124: out = 16'(-3545);
			12125: out = 16'(3326);
			12126: out = 16'(12626);
			12127: out = 16'(14152);
			12128: out = 16'(7228);
			12129: out = 16'(-14945);
			12130: out = 16'(-19031);
			12131: out = 16'(-6359);
			12132: out = 16'(6281);
			12133: out = 16'(-4485);
			12134: out = 16'(1173);
			12135: out = 16'(9665);
			12136: out = 16'(7687);
			12137: out = 16'(-14108);
			12138: out = 16'(-9867);
			12139: out = 16'(2117);
			12140: out = 16'(5615);
			12141: out = 16'(0);
			12142: out = 16'(-5010);
			12143: out = 16'(-11133);
			12144: out = 16'(-12005);
			12145: out = 16'(1511);
			12146: out = 16'(7431);
			12147: out = 16'(9751);
			12148: out = 16'(9939);
			12149: out = 16'(15082);
			12150: out = 16'(3411);
			12151: out = 16'(-4376);
			12152: out = 16'(-14284);
			12153: out = 16'(-13826);
			12154: out = 16'(-5530);
			12155: out = 16'(11756);
			12156: out = 16'(10760);
			12157: out = 16'(738);
			12158: out = 16'(-8586);
			12159: out = 16'(3175);
			12160: out = 16'(2900);
			12161: out = 16'(-2632);
			12162: out = 16'(2547);
			12163: out = 16'(6875);
			12164: out = 16'(-5456);
			12165: out = 16'(-13831);
			12166: out = 16'(5885);
			12167: out = 16'(6661);
			12168: out = 16'(1527);
			12169: out = 16'(-5681);
			12170: out = 16'(-1069);
			12171: out = 16'(5009);
			12172: out = 16'(3200);
			12173: out = 16'(-1230);
			12174: out = 16'(7);
			12175: out = 16'(-4652);
			12176: out = 16'(-2239);
			12177: out = 16'(538);
			12178: out = 16'(1159);
			12179: out = 16'(-11375);
			12180: out = 16'(-2978);
			12181: out = 16'(6392);
			12182: out = 16'(10476);
			12183: out = 16'(2819);
			12184: out = 16'(2590);
			12185: out = 16'(-2598);
			12186: out = 16'(-3969);
			12187: out = 16'(-3705);
			12188: out = 16'(-8366);
			12189: out = 16'(-9640);
			12190: out = 16'(1361);
			12191: out = 16'(12789);
			12192: out = 16'(892);
			12193: out = 16'(-2782);
			12194: out = 16'(2692);
			12195: out = 16'(9287);
			12196: out = 16'(-1728);
			12197: out = 16'(-2556);
			12198: out = 16'(288);
			12199: out = 16'(3322);
			12200: out = 16'(-6243);
			12201: out = 16'(1934);
			12202: out = 16'(2755);
			12203: out = 16'(2750);
			12204: out = 16'(232);
			12205: out = 16'(-1378);
			12206: out = 16'(-10670);
			12207: out = 16'(-10490);
			12208: out = 16'(4012);
			12209: out = 16'(6556);
			12210: out = 16'(3780);
			12211: out = 16'(-2429);
			12212: out = 16'(1444);
			12213: out = 16'(8060);
			12214: out = 16'(7521);
			12215: out = 16'(-4286);
			12216: out = 16'(-6698);
			12217: out = 16'(5180);
			12218: out = 16'(6601);
			12219: out = 16'(-9540);
			12220: out = 16'(-13971);
			12221: out = 16'(12269);
			12222: out = 16'(11885);
			12223: out = 16'(1087);
			12224: out = 16'(-7587);
			12225: out = 16'(1539);
			12226: out = 16'(1369);
			12227: out = 16'(232);
			12228: out = 16'(-7139);
			12229: out = 16'(-10290);
			12230: out = 16'(-696);
			12231: out = 16'(2085);
			12232: out = 16'(6313);
			12233: out = 16'(11302);
			12234: out = 16'(8827);
			12235: out = 16'(-717);
			12236: out = 16'(-8053);
			12237: out = 16'(-7320);
			12238: out = 16'(-3221);
			12239: out = 16'(-5998);
			12240: out = 16'(-6890);
			12241: out = 16'(-2494);
			12242: out = 16'(5047);
			12243: out = 16'(8063);
			12244: out = 16'(8739);
			12245: out = 16'(4550);
			12246: out = 16'(-491);
			12247: out = 16'(-4285);
			12248: out = 16'(-597);
			12249: out = 16'(854);
			12250: out = 16'(-265);
			12251: out = 16'(-98);
			12252: out = 16'(2386);
			12253: out = 16'(-551);
			12254: out = 16'(-4190);
			12255: out = 16'(-131);
			12256: out = 16'(398);
			12257: out = 16'(-4480);
			12258: out = 16'(-7469);
			12259: out = 16'(1507);
			12260: out = 16'(5140);
			12261: out = 16'(5009);
			12262: out = 16'(2628);
			12263: out = 16'(6931);
			12264: out = 16'(-634);
			12265: out = 16'(689);
			12266: out = 16'(-2441);
			12267: out = 16'(-2242);
			12268: out = 16'(-5686);
			12269: out = 16'(6810);
			12270: out = 16'(408);
			12271: out = 16'(-13176);
			12272: out = 16'(-10944);
			12273: out = 16'(-192);
			12274: out = 16'(2418);
			12275: out = 16'(126);
			12276: out = 16'(2931);
			12277: out = 16'(2246);
			12278: out = 16'(-2471);
			12279: out = 16'(-464);
			12280: out = 16'(8252);
			12281: out = 16'(-2098);
			12282: out = 16'(-11604);
			12283: out = 16'(-3444);
			12284: out = 16'(16986);
			12285: out = 16'(11151);
			12286: out = 16'(-1869);
			12287: out = 16'(-10302);
			12288: out = 16'(-3564);
			12289: out = 16'(-4118);
			12290: out = 16'(531);
			12291: out = 16'(-311);
			12292: out = 16'(-823);
			12293: out = 16'(-7147);
			12294: out = 16'(6666);
			12295: out = 16'(10558);
			12296: out = 16'(9289);
			12297: out = 16'(2608);
			12298: out = 16'(3671);
			12299: out = 16'(-7644);
			12300: out = 16'(-12957);
			12301: out = 16'(-4531);
			12302: out = 16'(9341);
			12303: out = 16'(-1418);
			12304: out = 16'(-17365);
			12305: out = 16'(-16616);
			12306: out = 16'(5425);
			12307: out = 16'(15228);
			12308: out = 16'(14389);
			12309: out = 16'(9649);
			12310: out = 16'(731);
			12311: out = 16'(632);
			12312: out = 16'(-5233);
			12313: out = 16'(-8542);
			12314: out = 16'(-5003);
			12315: out = 16'(2890);
			12316: out = 16'(2964);
			12317: out = 16'(562);
			12318: out = 16'(516);
			12319: out = 16'(8146);
			12320: out = 16'(3108);
			12321: out = 16'(-3692);
			12322: out = 16'(-8069);
			12323: out = 16'(-9392);
			12324: out = 16'(-9939);
			12325: out = 16'(-348);
			12326: out = 16'(10684);
			12327: out = 16'(8849);
			12328: out = 16'(-690);
			12329: out = 16'(-6678);
			12330: out = 16'(-2483);
			12331: out = 16'(5085);
			12332: out = 16'(1061);
			12333: out = 16'(-407);
			12334: out = 16'(394);
			12335: out = 16'(455);
			12336: out = 16'(-8899);
			12337: out = 16'(-4488);
			12338: out = 16'(3756);
			12339: out = 16'(6356);
			12340: out = 16'(6562);
			12341: out = 16'(-785);
			12342: out = 16'(-8950);
			12343: out = 16'(-11381);
			12344: out = 16'(476);
			12345: out = 16'(8411);
			12346: out = 16'(13786);
			12347: out = 16'(11105);
			12348: out = 16'(1588);
			12349: out = 16'(-12804);
			12350: out = 16'(-16822);
			12351: out = 16'(-5757);
			12352: out = 16'(9429);
			12353: out = 16'(6926);
			12354: out = 16'(-709);
			12355: out = 16'(-7238);
			12356: out = 16'(-2987);
			12357: out = 16'(6086);
			12358: out = 16'(11461);
			12359: out = 16'(5806);
			12360: out = 16'(-792);
			12361: out = 16'(-582);
			12362: out = 16'(-800);
			12363: out = 16'(-4360);
			12364: out = 16'(-3836);
			12365: out = 16'(1851);
			12366: out = 16'(-8831);
			12367: out = 16'(-16177);
			12368: out = 16'(-1986);
			12369: out = 16'(20077);
			12370: out = 16'(11469);
			12371: out = 16'(-7810);
			12372: out = 16'(-12361);
			12373: out = 16'(2840);
			12374: out = 16'(-3750);
			12375: out = 16'(-6716);
			12376: out = 16'(1861);
			12377: out = 16'(16213);
			12378: out = 16'(5563);
			12379: out = 16'(2260);
			12380: out = 16'(-621);
			12381: out = 16'(-2419);
			12382: out = 16'(-15917);
			12383: out = 16'(-1275);
			12384: out = 16'(9130);
			12385: out = 16'(6600);
			12386: out = 16'(-9249);
			12387: out = 16'(-11950);
			12388: out = 16'(-7668);
			12389: out = 16'(3233);
			12390: out = 16'(10996);
			12391: out = 16'(2464);
			12392: out = 16'(4602);
			12393: out = 16'(8116);
			12394: out = 16'(6270);
			12395: out = 16'(-13519);
			12396: out = 16'(-2855);
			12397: out = 16'(6428);
			12398: out = 16'(4478);
			12399: out = 16'(-2474);
			12400: out = 16'(-2886);
			12401: out = 16'(-2843);
			12402: out = 16'(-1527);
			12403: out = 16'(1793);
			12404: out = 16'(6110);
			12405: out = 16'(3691);
			12406: out = 16'(95);
			12407: out = 16'(-1310);
			12408: out = 16'(5139);
			12409: out = 16'(-2533);
			12410: out = 16'(-6128);
			12411: out = 16'(2271);
			12412: out = 16'(10797);
			12413: out = 16'(1663);
			12414: out = 16'(-8719);
			12415: out = 16'(-7753);
			12416: out = 16'(471);
			12417: out = 16'(-6315);
			12418: out = 16'(-7258);
			12419: out = 16'(6545);
			12420: out = 16'(15125);
			12421: out = 16'(10235);
			12422: out = 16'(-6092);
			12423: out = 16'(-10554);
			12424: out = 16'(464);
			12425: out = 16'(6242);
			12426: out = 16'(-3035);
			12427: out = 16'(-12418);
			12428: out = 16'(-11197);
			12429: out = 16'(441);
			12430: out = 16'(1189);
			12431: out = 16'(1812);
			12432: out = 16'(5341);
			12433: out = 16'(11019);
			12434: out = 16'(554);
			12435: out = 16'(-2966);
			12436: out = 16'(-2462);
			12437: out = 16'(-8171);
			12438: out = 16'(-10345);
			12439: out = 16'(1141);
			12440: out = 16'(13827);
			12441: out = 16'(11720);
			12442: out = 16'(5769);
			12443: out = 16'(142);
			12444: out = 16'(-1796);
			12445: out = 16'(225);
			12446: out = 16'(-3724);
			12447: out = 16'(4130);
			12448: out = 16'(1534);
			12449: out = 16'(-10999);
			12450: out = 16'(-22988);
			12451: out = 16'(-1322);
			12452: out = 16'(12546);
			12453: out = 16'(6825);
			12454: out = 16'(7553);
			12455: out = 16'(5964);
			12456: out = 16'(-148);
			12457: out = 16'(-14478);
			12458: out = 16'(-17141);
			12459: out = 16'(-6419);
			12460: out = 16'(7754);
			12461: out = 16'(4751);
			12462: out = 16'(-2381);
			12463: out = 16'(6277);
			12464: out = 16'(14768);
			12465: out = 16'(4437);
			12466: out = 16'(-13649);
			12467: out = 16'(-9120);
			12468: out = 16'(5585);
			12469: out = 16'(10697);
			12470: out = 16'(4776);
			12471: out = 16'(1574);
			12472: out = 16'(1723);
			12473: out = 16'(-5056);
			12474: out = 16'(-14801);
			12475: out = 16'(-13535);
			12476: out = 16'(-2702);
			12477: out = 16'(4345);
			12478: out = 16'(6402);
			12479: out = 16'(7122);
			12480: out = 16'(-1883);
			12481: out = 16'(-5054);
			12482: out = 16'(4650);
			12483: out = 16'(15873);
			12484: out = 16'(11694);
			12485: out = 16'(-3017);
			12486: out = 16'(-6947);
			12487: out = 16'(1083);
			12488: out = 16'(-181);
			12489: out = 16'(-6526);
			12490: out = 16'(-3812);
			12491: out = 16'(5039);
			12492: out = 16'(-711);
			12493: out = 16'(-1863);
			12494: out = 16'(-1711);
			12495: out = 16'(-2261);
			12496: out = 16'(-12525);
			12497: out = 16'(7747);
			12498: out = 16'(11560);
			12499: out = 16'(2497);
			12500: out = 16'(-9879);
			12501: out = 16'(-3728);
			12502: out = 16'(1473);
			12503: out = 16'(3207);
			12504: out = 16'(5116);
			12505: out = 16'(7612);
			12506: out = 16'(11494);
			12507: out = 16'(1094);
			12508: out = 16'(-13985);
			12509: out = 16'(-14143);
			12510: out = 16'(-3416);
			12511: out = 16'(-248);
			12512: out = 16'(-5469);
			12513: out = 16'(-4284);
			12514: out = 16'(77);
			12515: out = 16'(5834);
			12516: out = 16'(8582);
			12517: out = 16'(7960);
			12518: out = 16'(2858);
			12519: out = 16'(-7886);
			12520: out = 16'(-12491);
			12521: out = 16'(-4894);
			12522: out = 16'(792);
			12523: out = 16'(-1145);
			12524: out = 16'(-5084);
			12525: out = 16'(-1452);
			12526: out = 16'(4883);
			12527: out = 16'(10715);
			12528: out = 16'(6260);
			12529: out = 16'(-2365);
			12530: out = 16'(-4911);
			12531: out = 16'(-8465);
			12532: out = 16'(-3955);
			12533: out = 16'(2737);
			12534: out = 16'(6583);
			12535: out = 16'(1110);
			12536: out = 16'(442);
			12537: out = 16'(-1628);
			12538: out = 16'(-7176);
			12539: out = 16'(-5160);
			12540: out = 16'(-1345);
			12541: out = 16'(971);
			12542: out = 16'(-1394);
			12543: out = 16'(1416);
			12544: out = 16'(1707);
			12545: out = 16'(7594);
			12546: out = 16'(11308);
			12547: out = 16'(10824);
			12548: out = 16'(1990);
			12549: out = 16'(-909);
			12550: out = 16'(-3925);
			12551: out = 16'(-11400);
			12552: out = 16'(-9346);
			12553: out = 16'(1687);
			12554: out = 16'(12604);
			12555: out = 16'(12121);
			12556: out = 16'(2124);
			12557: out = 16'(-8347);
			12558: out = 16'(-8762);
			12559: out = 16'(3302);
			12560: out = 16'(11152);
			12561: out = 16'(10210);
			12562: out = 16'(-4285);
			12563: out = 16'(-12559);
			12564: out = 16'(3679);
			12565: out = 16'(8442);
			12566: out = 16'(3351);
			12567: out = 16'(-1364);
			12568: out = 16'(3861);
			12569: out = 16'(1777);
			12570: out = 16'(-2504);
			12571: out = 16'(-3524);
			12572: out = 16'(-537);
			12573: out = 16'(-4590);
			12574: out = 16'(-8259);
			12575: out = 16'(395);
			12576: out = 16'(12578);
			12577: out = 16'(2075);
			12578: out = 16'(-6630);
			12579: out = 16'(-2520);
			12580: out = 16'(10080);
			12581: out = 16'(5050);
			12582: out = 16'(-363);
			12583: out = 16'(-4415);
			12584: out = 16'(-3513);
			12585: out = 16'(-9311);
			12586: out = 16'(-1503);
			12587: out = 16'(80);
			12588: out = 16'(-393);
			12589: out = 16'(15);
			12590: out = 16'(-227);
			12591: out = 16'(3939);
			12592: out = 16'(7176);
			12593: out = 16'(5868);
			12594: out = 16'(-8906);
			12595: out = 16'(-1796);
			12596: out = 16'(7664);
			12597: out = 16'(4854);
			12598: out = 16'(-14966);
			12599: out = 16'(-11087);
			12600: out = 16'(-2329);
			12601: out = 16'(-732);
			12602: out = 16'(-4984);
			12603: out = 16'(-236);
			12604: out = 16'(5552);
			12605: out = 16'(6923);
			12606: out = 16'(2350);
			12607: out = 16'(6354);
			12608: out = 16'(-1944);
			12609: out = 16'(-11406);
			12610: out = 16'(-8946);
			12611: out = 16'(6332);
			12612: out = 16'(5955);
			12613: out = 16'(-4376);
			12614: out = 16'(-5976);
			12615: out = 16'(3494);
			12616: out = 16'(8360);
			12617: out = 16'(-2817);
			12618: out = 16'(-11596);
			12619: out = 16'(101);
			12620: out = 16'(7320);
			12621: out = 16'(-607);
			12622: out = 16'(-9512);
			12623: out = 16'(1263);
			12624: out = 16'(-24);
			12625: out = 16'(582);
			12626: out = 16'(720);
			12627: out = 16'(4052);
			12628: out = 16'(13047);
			12629: out = 16'(6201);
			12630: out = 16'(-5626);
			12631: out = 16'(-10228);
			12632: out = 16'(577);
			12633: out = 16'(5290);
			12634: out = 16'(5570);
			12635: out = 16'(207);
			12636: out = 16'(-5974);
			12637: out = 16'(-8648);
			12638: out = 16'(2560);
			12639: out = 16'(10378);
			12640: out = 16'(2261);
			12641: out = 16'(-1130);
			12642: out = 16'(4020);
			12643: out = 16'(7418);
			12644: out = 16'(-1330);
			12645: out = 16'(-4786);
			12646: out = 16'(-2136);
			12647: out = 16'(2074);
			12648: out = 16'(-1379);
			12649: out = 16'(-6086);
			12650: out = 16'(-723);
			12651: out = 16'(7509);
			12652: out = 16'(7599);
			12653: out = 16'(7960);
			12654: out = 16'(2876);
			12655: out = 16'(2561);
			12656: out = 16'(1252);
			12657: out = 16'(-19);
			12658: out = 16'(-10055);
			12659: out = 16'(-6871);
			12660: out = 16'(1905);
			12661: out = 16'(1943);
			12662: out = 16'(5110);
			12663: out = 16'(1287);
			12664: out = 16'(-6000);
			12665: out = 16'(-13878);
			12666: out = 16'(4651);
			12667: out = 16'(4674);
			12668: out = 16'(-294);
			12669: out = 16'(-4972);
			12670: out = 16'(-5263);
			12671: out = 16'(-1444);
			12672: out = 16'(6556);
			12673: out = 16'(9460);
			12674: out = 16'(2423);
			12675: out = 16'(-4068);
			12676: out = 16'(-7679);
			12677: out = 16'(-8553);
			12678: out = 16'(-5066);
			12679: out = 16'(-7522);
			12680: out = 16'(-383);
			12681: out = 16'(4989);
			12682: out = 16'(3418);
			12683: out = 16'(-5813);
			12684: out = 16'(-5978);
			12685: out = 16'(-7259);
			12686: out = 16'(-9786);
			12687: out = 16'(356);
			12688: out = 16'(13845);
			12689: out = 16'(12299);
			12690: out = 16'(-1655);
			12691: out = 16'(-6974);
			12692: out = 16'(-1781);
			12693: out = 16'(3920);
			12694: out = 16'(1462);
			12695: out = 16'(-456);
			12696: out = 16'(4604);
			12697: out = 16'(4748);
			12698: out = 16'(-4407);
			12699: out = 16'(-11309);
			12700: out = 16'(-365);
			12701: out = 16'(8734);
			12702: out = 16'(4000);
			12703: out = 16'(-5036);
			12704: out = 16'(456);
			12705: out = 16'(8846);
			12706: out = 16'(6394);
			12707: out = 16'(-3965);
			12708: out = 16'(338);
			12709: out = 16'(1658);
			12710: out = 16'(1059);
			12711: out = 16'(-3948);
			12712: out = 16'(-473);
			12713: out = 16'(-3851);
			12714: out = 16'(5599);
			12715: out = 16'(14095);
			12716: out = 16'(11427);
			12717: out = 16'(1830);
			12718: out = 16'(1955);
			12719: out = 16'(6076);
			12720: out = 16'(-1734);
			12721: out = 16'(-6409);
			12722: out = 16'(-13621);
			12723: out = 16'(-3828);
			12724: out = 16'(9090);
			12725: out = 16'(12968);
			12726: out = 16'(372);
			12727: out = 16'(-3001);
			12728: out = 16'(-1757);
			12729: out = 16'(-4119);
			12730: out = 16'(-17659);
			12731: out = 16'(-11167);
			12732: out = 16'(5931);
			12733: out = 16'(13385);
			12734: out = 16'(1430);
			12735: out = 16'(6468);
			12736: out = 16'(11735);
			12737: out = 16'(4473);
			12738: out = 16'(-5699);
			12739: out = 16'(4031);
			12740: out = 16'(4112);
			12741: out = 16'(-19771);
			12742: out = 16'(-28175);
			12743: out = 16'(-13435);
			12744: out = 16'(10434);
			12745: out = 16'(12166);
			12746: out = 16'(2365);
			12747: out = 16'(-405);
			12748: out = 16'(-2948);
			12749: out = 16'(-12593);
			12750: out = 16'(-20382);
			12751: out = 16'(3176);
			12752: out = 16'(19041);
			12753: out = 16'(12530);
			12754: out = 16'(-19);
			12755: out = 16'(-7129);
			12756: out = 16'(-3605);
			12757: out = 16'(-2118);
			12758: out = 16'(-4174);
			12759: out = 16'(-5607);
			12760: out = 16'(-3274);
			12761: out = 16'(-1854);
			12762: out = 16'(1337);
			12763: out = 16'(1926);
			12764: out = 16'(4297);
			12765: out = 16'(-2528);
			12766: out = 16'(-4385);
			12767: out = 16'(4191);
			12768: out = 16'(4318);
			12769: out = 16'(-14476);
			12770: out = 16'(-24546);
			12771: out = 16'(188);
			12772: out = 16'(15111);
			12773: out = 16'(12116);
			12774: out = 16'(1323);
			12775: out = 16'(-1326);
			12776: out = 16'(7886);
			12777: out = 16'(-421);
			12778: out = 16'(-8313);
			12779: out = 16'(-2979);
			12780: out = 16'(3365);
			12781: out = 16'(4426);
			12782: out = 16'(8779);
			12783: out = 16'(16381);
			12784: out = 16'(8805);
			12785: out = 16'(298);
			12786: out = 16'(-11497);
			12787: out = 16'(-11396);
			12788: out = 16'(-4);
			12789: out = 16'(4714);
			12790: out = 16'(2420);
			12791: out = 16'(-1593);
			12792: out = 16'(-2311);
			12793: out = 16'(670);
			12794: out = 16'(4881);
			12795: out = 16'(4488);
			12796: out = 16'(-355);
			12797: out = 16'(5158);
			12798: out = 16'(1886);
			12799: out = 16'(1990);
			12800: out = 16'(3975);
			12801: out = 16'(5866);
			12802: out = 16'(5434);
			12803: out = 16'(4696);
			12804: out = 16'(-2902);
			12805: out = 16'(-19328);
			12806: out = 16'(-19411);
			12807: out = 16'(-8212);
			12808: out = 16'(2633);
			12809: out = 16'(4319);
			12810: out = 16'(13698);
			12811: out = 16'(10325);
			12812: out = 16'(-684);
			12813: out = 16'(-11374);
			12814: out = 16'(-5042);
			12815: out = 16'(-596);
			12816: out = 16'(-2355);
			12817: out = 16'(-6941);
			12818: out = 16'(-2510);
			12819: out = 16'(-275);
			12820: out = 16'(-93);
			12821: out = 16'(-879);
			12822: out = 16'(2156);
			12823: out = 16'(8962);
			12824: out = 16'(7816);
			12825: out = 16'(-2651);
			12826: out = 16'(-13815);
			12827: out = 16'(-13507);
			12828: out = 16'(-4075);
			12829: out = 16'(3847);
			12830: out = 16'(4228);
			12831: out = 16'(8910);
			12832: out = 16'(8456);
			12833: out = 16'(6362);
			12834: out = 16'(-3505);
			12835: out = 16'(-14825);
			12836: out = 16'(-25160);
			12837: out = 16'(-13117);
			12838: out = 16'(7970);
			12839: out = 16'(14539);
			12840: out = 16'(6024);
			12841: out = 16'(2251);
			12842: out = 16'(3077);
			12843: out = 16'(1864);
			12844: out = 16'(2344);
			12845: out = 16'(7877);
			12846: out = 16'(9282);
			12847: out = 16'(2483);
			12848: out = 16'(-9575);
			12849: out = 16'(-5081);
			12850: out = 16'(2034);
			12851: out = 16'(971);
			12852: out = 16'(289);
			12853: out = 16'(2170);
			12854: out = 16'(-976);
			12855: out = 16'(-10047);
			12856: out = 16'(-11408);
			12857: out = 16'(-1479);
			12858: out = 16'(7790);
			12859: out = 16'(7040);
			12860: out = 16'(1935);
			12861: out = 16'(2293);
			12862: out = 16'(3798);
			12863: out = 16'(3001);
			12864: out = 16'(-117);
			12865: out = 16'(149);
			12866: out = 16'(-3355);
			12867: out = 16'(-6773);
			12868: out = 16'(-7523);
			12869: out = 16'(-16);
			12870: out = 16'(3434);
			12871: out = 16'(8184);
			12872: out = 16'(9663);
			12873: out = 16'(5428);
			12874: out = 16'(-8220);
			12875: out = 16'(-12485);
			12876: out = 16'(-5694);
			12877: out = 16'(-251);
			12878: out = 16'(554);
			12879: out = 16'(3264);
			12880: out = 16'(7334);
			12881: out = 16'(5426);
			12882: out = 16'(1565);
			12883: out = 16'(-2889);
			12884: out = 16'(-3797);
			12885: out = 16'(-2943);
			12886: out = 16'(-6381);
			12887: out = 16'(-2803);
			12888: out = 16'(2865);
			12889: out = 16'(5701);
			12890: out = 16'(8491);
			12891: out = 16'(6204);
			12892: out = 16'(1178);
			12893: out = 16'(-5918);
			12894: out = 16'(-7421);
			12895: out = 16'(82);
			12896: out = 16'(7903);
			12897: out = 16'(1750);
			12898: out = 16'(-14777);
			12899: out = 16'(-7619);
			12900: out = 16'(7357);
			12901: out = 16'(10932);
			12902: out = 16'(3369);
			12903: out = 16'(896);
			12904: out = 16'(4957);
			12905: out = 16'(1165);
			12906: out = 16'(-11256);
			12907: out = 16'(-13959);
			12908: out = 16'(2958);
			12909: out = 16'(15924);
			12910: out = 16'(11254);
			12911: out = 16'(3226);
			12912: out = 16'(-10533);
			12913: out = 16'(-17545);
			12914: out = 16'(-13977);
			12915: out = 16'(537);
			12916: out = 16'(630);
			12917: out = 16'(2639);
			12918: out = 16'(7291);
			12919: out = 16'(7162);
			12920: out = 16'(19);
			12921: out = 16'(-10487);
			12922: out = 16'(-7784);
			12923: out = 16'(3825);
			12924: out = 16'(6600);
			12925: out = 16'(1600);
			12926: out = 16'(1306);
			12927: out = 16'(1080);
			12928: out = 16'(-5369);
			12929: out = 16'(-18456);
			12930: out = 16'(-10174);
			12931: out = 16'(7078);
			12932: out = 16'(4950);
			12933: out = 16'(73);
			12934: out = 16'(6099);
			12935: out = 16'(11732);
			12936: out = 16'(-1595);
			12937: out = 16'(-12569);
			12938: out = 16'(-8421);
			12939: out = 16'(5411);
			12940: out = 16'(5362);
			12941: out = 16'(8850);
			12942: out = 16'(5195);
			12943: out = 16'(4227);
			12944: out = 16'(-1675);
			12945: out = 16'(43);
			12946: out = 16'(-266);
			12947: out = 16'(9829);
			12948: out = 16'(10798);
			12949: out = 16'(-6269);
			12950: out = 16'(-16470);
			12951: out = 16'(-9403);
			12952: out = 16'(2954);
			12953: out = 16'(3835);
			12954: out = 16'(6017);
			12955: out = 16'(7415);
			12956: out = 16'(4690);
			12957: out = 16'(-1715);
			12958: out = 16'(-2127);
			12959: out = 16'(3064);
			12960: out = 16'(3372);
			12961: out = 16'(-1290);
			12962: out = 16'(-8546);
			12963: out = 16'(-2213);
			12964: out = 16'(-1346);
			12965: out = 16'(-3432);
			12966: out = 16'(-527);
			12967: out = 16'(8041);
			12968: out = 16'(-708);
			12969: out = 16'(-10638);
			12970: out = 16'(957);
			12971: out = 16'(11059);
			12972: out = 16'(2426);
			12973: out = 16'(-11497);
			12974: out = 16'(-7379);
			12975: out = 16'(7653);
			12976: out = 16'(6072);
			12977: out = 16'(-2880);
			12978: out = 16'(-1003);
			12979: out = 16'(3701);
			12980: out = 16'(2514);
			12981: out = 16'(-1617);
			12982: out = 16'(756);
			12983: out = 16'(-743);
			12984: out = 16'(4383);
			12985: out = 16'(2950);
			12986: out = 16'(-2789);
			12987: out = 16'(-14139);
			12988: out = 16'(-8792);
			12989: out = 16'(-2708);
			12990: out = 16'(2175);
			12991: out = 16'(5224);
			12992: out = 16'(4354);
			12993: out = 16'(3166);
			12994: out = 16'(1971);
			12995: out = 16'(-414);
			12996: out = 16'(365);
			12997: out = 16'(2011);
			12998: out = 16'(5864);
			12999: out = 16'(6489);
			13000: out = 16'(5442);
			13001: out = 16'(-4369);
			13002: out = 16'(-5097);
			13003: out = 16'(555);
			13004: out = 16'(-3475);
			13005: out = 16'(-3734);
			13006: out = 16'(-2564);
			13007: out = 16'(736);
			13008: out = 16'(-1978);
			13009: out = 16'(3754);
			13010: out = 16'(1506);
			13011: out = 16'(-265);
			13012: out = 16'(691);
			13013: out = 16'(9713);
			13014: out = 16'(1267);
			13015: out = 16'(-10337);
			13016: out = 16'(-9783);
			13017: out = 16'(7362);
			13018: out = 16'(9051);
			13019: out = 16'(-2440);
			13020: out = 16'(-12387);
			13021: out = 16'(-1359);
			13022: out = 16'(-121);
			13023: out = 16'(-218);
			13024: out = 16'(-1950);
			13025: out = 16'(-2554);
			13026: out = 16'(-4972);
			13027: out = 16'(-5410);
			13028: out = 16'(-4054);
			13029: out = 16'(1546);
			13030: out = 16'(9034);
			13031: out = 16'(14547);
			13032: out = 16'(9803);
			13033: out = 16'(-2847);
			13034: out = 16'(-17288);
			13035: out = 16'(-7579);
			13036: out = 16'(9435);
			13037: out = 16'(11105);
			13038: out = 16'(1136);
			13039: out = 16'(-4673);
			13040: out = 16'(1155);
			13041: out = 16'(5244);
			13042: out = 16'(-1711);
			13043: out = 16'(-8422);
			13044: out = 16'(-5588);
			13045: out = 16'(4563);
			13046: out = 16'(12503);
			13047: out = 16'(8756);
			13048: out = 16'(5088);
			13049: out = 16'(-2088);
			13050: out = 16'(-9894);
			13051: out = 16'(-5305);
			13052: out = 16'(-728);
			13053: out = 16'(-1627);
			13054: out = 16'(-3192);
			13055: out = 16'(3065);
			13056: out = 16'(2333);
			13057: out = 16'(-5360);
			13058: out = 16'(-6802);
			13059: out = 16'(6912);
			13060: out = 16'(13460);
			13061: out = 16'(5151);
			13062: out = 16'(-4711);
			13063: out = 16'(-4071);
			13064: out = 16'(1875);
			13065: out = 16'(-4858);
			13066: out = 16'(-12855);
			13067: out = 16'(-9658);
			13068: out = 16'(3711);
			13069: out = 16'(2407);
			13070: out = 16'(2982);
			13071: out = 16'(9418);
			13072: out = 16'(475);
			13073: out = 16'(-9032);
			13074: out = 16'(-9197);
			13075: out = 16'(2722);
			13076: out = 16'(2889);
			13077: out = 16'(1893);
			13078: out = 16'(-1072);
			13079: out = 16'(1018);
			13080: out = 16'(601);
			13081: out = 16'(1060);
			13082: out = 16'(-370);
			13083: out = 16'(814);
			13084: out = 16'(-621);
			13085: out = 16'(-3917);
			13086: out = 16'(-4794);
			13087: out = 16'(210);
			13088: out = 16'(506);
			13089: out = 16'(-805);
			13090: out = 16'(-6098);
			13091: out = 16'(2851);
			13092: out = 16'(13107);
			13093: out = 16'(8837);
			13094: out = 16'(-467);
			13095: out = 16'(-1156);
			13096: out = 16'(90);
			13097: out = 16'(-6391);
			13098: out = 16'(-5911);
			13099: out = 16'(6524);
			13100: out = 16'(12018);
			13101: out = 16'(884);
			13102: out = 16'(-22386);
			13103: out = 16'(-15540);
			13104: out = 16'(2838);
			13105: out = 16'(-166);
			13106: out = 16'(-455);
			13107: out = 16'(5257);
			13108: out = 16'(17045);
			13109: out = 16'(13921);
			13110: out = 16'(9243);
			13111: out = 16'(-7797);
			13112: out = 16'(-8755);
			13113: out = 16'(-4635);
			13114: out = 16'(-7726);
			13115: out = 16'(-11615);
			13116: out = 16'(1070);
			13117: out = 16'(14963);
			13118: out = 16'(8484);
			13119: out = 16'(-3892);
			13120: out = 16'(-12811);
			13121: out = 16'(-9162);
			13122: out = 16'(-1601);
			13123: out = 16'(8069);
			13124: out = 16'(9063);
			13125: out = 16'(6829);
			13126: out = 16'(2088);
			13127: out = 16'(5574);
			13128: out = 16'(-3577);
			13129: out = 16'(-5595);
			13130: out = 16'(3306);
			13131: out = 16'(13485);
			13132: out = 16'(7228);
			13133: out = 16'(-4189);
			13134: out = 16'(-14070);
			13135: out = 16'(-20011);
			13136: out = 16'(-4373);
			13137: out = 16'(6871);
			13138: out = 16'(6656);
			13139: out = 16'(-67);
			13140: out = 16'(-2116);
			13141: out = 16'(-3424);
			13142: out = 16'(-3730);
			13143: out = 16'(-830);
			13144: out = 16'(9534);
			13145: out = 16'(11714);
			13146: out = 16'(5386);
			13147: out = 16'(-4973);
			13148: out = 16'(-10302);
			13149: out = 16'(-14915);
			13150: out = 16'(-12291);
			13151: out = 16'(-3119);
			13152: out = 16'(3849);
			13153: out = 16'(4406);
			13154: out = 16'(266);
			13155: out = 16'(1404);
			13156: out = 16'(7386);
			13157: out = 16'(3224);
			13158: out = 16'(-5027);
			13159: out = 16'(-4235);
			13160: out = 16'(7240);
			13161: out = 16'(2063);
			13162: out = 16'(-3460);
			13163: out = 16'(-6197);
			13164: out = 16'(-1018);
			13165: out = 16'(-90);
			13166: out = 16'(2020);
			13167: out = 16'(1925);
			13168: out = 16'(4466);
			13169: out = 16'(7979);
			13170: out = 16'(-1063);
			13171: out = 16'(-11351);
			13172: out = 16'(-10765);
			13173: out = 16'(2377);
			13174: out = 16'(9605);
			13175: out = 16'(10327);
			13176: out = 16'(6033);
			13177: out = 16'(-880);
			13178: out = 16'(-3231);
			13179: out = 16'(-6524);
			13180: out = 16'(-4112);
			13181: out = 16'(2847);
			13182: out = 16'(7024);
			13183: out = 16'(6870);
			13184: out = 16'(4774);
			13185: out = 16'(1117);
			13186: out = 16'(-3630);
			13187: out = 16'(-1909);
			13188: out = 16'(4065);
			13189: out = 16'(3002);
			13190: out = 16'(-9515);
			13191: out = 16'(-10861);
			13192: out = 16'(2055);
			13193: out = 16'(12718);
			13194: out = 16'(4272);
			13195: out = 16'(4182);
			13196: out = 16'(-1794);
			13197: out = 16'(-3470);
			13198: out = 16'(-6725);
			13199: out = 16'(-5834);
			13200: out = 16'(-12834);
			13201: out = 16'(-8262);
			13202: out = 16'(6696);
			13203: out = 16'(16310);
			13204: out = 16'(5691);
			13205: out = 16'(-5141);
			13206: out = 16'(-4120);
			13207: out = 16'(5905);
			13208: out = 16'(4810);
			13209: out = 16'(1877);
			13210: out = 16'(1095);
			13211: out = 16'(146);
			13212: out = 16'(-6421);
			13213: out = 16'(-13772);
			13214: out = 16'(-12543);
			13215: out = 16'(-662);
			13216: out = 16'(4246);
			13217: out = 16'(7108);
			13218: out = 16'(4006);
			13219: out = 16'(-586);
			13220: out = 16'(-6362);
			13221: out = 16'(2455);
			13222: out = 16'(8942);
			13223: out = 16'(6241);
			13224: out = 16'(-2409);
			13225: out = 16'(-3164);
			13226: out = 16'(-1928);
			13227: out = 16'(-562);
			13228: out = 16'(3430);
			13229: out = 16'(7244);
			13230: out = 16'(9336);
			13231: out = 16'(5341);
			13232: out = 16'(-1170);
			13233: out = 16'(-9173);
			13234: out = 16'(-7575);
			13235: out = 16'(-4723);
			13236: out = 16'(-3854);
			13237: out = 16'(-2841);
			13238: out = 16'(5379);
			13239: out = 16'(8905);
			13240: out = 16'(3341);
			13241: out = 16'(-6154);
			13242: out = 16'(-2492);
			13243: out = 16'(5082);
			13244: out = 16'(8507);
			13245: out = 16'(6600);
			13246: out = 16'(1519);
			13247: out = 16'(-8634);
			13248: out = 16'(-18951);
			13249: out = 16'(-16378);
			13250: out = 16'(4314);
			13251: out = 16'(13089);
			13252: out = 16'(3799);
			13253: out = 16'(-3046);
			13254: out = 16'(12258);
			13255: out = 16'(11697);
			13256: out = 16'(-10416);
			13257: out = 16'(-27556);
			13258: out = 16'(-4368);
			13259: out = 16'(11136);
			13260: out = 16'(6577);
			13261: out = 16'(-2286);
			13262: out = 16'(-1546);
			13263: out = 16'(1344);
			13264: out = 16'(-10230);
			13265: out = 16'(-15486);
			13266: out = 16'(4592);
			13267: out = 16'(20266);
			13268: out = 16'(10684);
			13269: out = 16'(-5763);
			13270: out = 16'(-8671);
			13271: out = 16'(-10031);
			13272: out = 16'(-6706);
			13273: out = 16'(1351);
			13274: out = 16'(11250);
			13275: out = 16'(55);
			13276: out = 16'(-5000);
			13277: out = 16'(-8260);
			13278: out = 16'(-1621);
			13279: out = 16'(5956);
			13280: out = 16'(3813);
			13281: out = 16'(-43);
			13282: out = 16'(3688);
			13283: out = 16'(9666);
			13284: out = 16'(-9093);
			13285: out = 16'(-16026);
			13286: out = 16'(-3724);
			13287: out = 16'(11323);
			13288: out = 16'(9773);
			13289: out = 16'(4930);
			13290: out = 16'(6324);
			13291: out = 16'(5797);
			13292: out = 16'(-13244);
			13293: out = 16'(-17071);
			13294: out = 16'(-64);
			13295: out = 16'(17077);
			13296: out = 16'(7762);
			13297: out = 16'(2559);
			13298: out = 16'(-3210);
			13299: out = 16'(-6516);
			13300: out = 16'(-8683);
			13301: out = 16'(-2400);
			13302: out = 16'(9690);
			13303: out = 16'(13953);
			13304: out = 16'(6716);
			13305: out = 16'(-12792);
			13306: out = 16'(-7937);
			13307: out = 16'(3844);
			13308: out = 16'(3017);
			13309: out = 16'(4751);
			13310: out = 16'(1060);
			13311: out = 16'(-1887);
			13312: out = 16'(-4945);
			13313: out = 16'(4317);
			13314: out = 16'(-4137);
			13315: out = 16'(-5061);
			13316: out = 16'(4522);
			13317: out = 16'(14562);
			13318: out = 16'(3990);
			13319: out = 16'(-8608);
			13320: out = 16'(-9884);
			13321: out = 16'(524);
			13322: out = 16'(680);
			13323: out = 16'(-2640);
			13324: out = 16'(-1963);
			13325: out = 16'(3086);
			13326: out = 16'(3168);
			13327: out = 16'(-5284);
			13328: out = 16'(-8803);
			13329: out = 16'(-1844);
			13330: out = 16'(2277);
			13331: out = 16'(1656);
			13332: out = 16'(893);
			13333: out = 16'(4408);
			13334: out = 16'(6986);
			13335: out = 16'(114);
			13336: out = 16'(-4000);
			13337: out = 16'(177);
			13338: out = 16'(5797);
			13339: out = 16'(-673);
			13340: out = 16'(-3876);
			13341: out = 16'(9);
			13342: out = 16'(3504);
			13343: out = 16'(1194);
			13344: out = 16'(-2387);
			13345: out = 16'(-403);
			13346: out = 16'(1417);
			13347: out = 16'(-9672);
			13348: out = 16'(-13271);
			13349: out = 16'(-5440);
			13350: out = 16'(6383);
			13351: out = 16'(7420);
			13352: out = 16'(11684);
			13353: out = 16'(15090);
			13354: out = 16'(13718);
			13355: out = 16'(974);
			13356: out = 16'(-10518);
			13357: out = 16'(-20167);
			13358: out = 16'(-14998);
			13359: out = 16'(4913);
			13360: out = 16'(12909);
			13361: out = 16'(12501);
			13362: out = 16'(1613);
			13363: out = 16'(-8646);
			13364: out = 16'(-9181);
			13365: out = 16'(-200);
			13366: out = 16'(1250);
			13367: out = 16'(-2417);
			13368: out = 16'(2608);
			13369: out = 16'(6037);
			13370: out = 16'(574);
			13371: out = 16'(-6822);
			13372: out = 16'(2752);
			13373: out = 16'(9966);
			13374: out = 16'(9891);
			13375: out = 16'(-1972);
			13376: out = 16'(-10446);
			13377: out = 16'(-18074);
			13378: out = 16'(-4770);
			13379: out = 16'(8157);
			13380: out = 16'(9971);
			13381: out = 16'(4448);
			13382: out = 16'(5320);
			13383: out = 16'(3092);
			13384: out = 16'(-7673);
			13385: out = 16'(-21598);
			13386: out = 16'(-18840);
			13387: out = 16'(-4995);
			13388: out = 16'(4906);
			13389: out = 16'(7986);
			13390: out = 16'(5100);
			13391: out = 16'(3109);
			13392: out = 16'(1300);
			13393: out = 16'(1612);
			13394: out = 16'(-6989);
			13395: out = 16'(-2443);
			13396: out = 16'(6785);
			13397: out = 16'(9602);
			13398: out = 16'(-3241);
			13399: out = 16'(-5089);
			13400: out = 16'(3538);
			13401: out = 16'(13513);
			13402: out = 16'(8851);
			13403: out = 16'(6224);
			13404: out = 16'(-1062);
			13405: out = 16'(-6514);
			13406: out = 16'(-11688);
			13407: out = 16'(-4168);
			13408: out = 16'(-4106);
			13409: out = 16'(-2922);
			13410: out = 16'(5369);
			13411: out = 16'(16405);
			13412: out = 16'(3860);
			13413: out = 16'(-10895);
			13414: out = 16'(-3027);
			13415: out = 16'(5764);
			13416: out = 16'(5299);
			13417: out = 16'(-4139);
			13418: out = 16'(-2683);
			13419: out = 16'(7830);
			13420: out = 16'(11475);
			13421: out = 16'(-2451);
			13422: out = 16'(-15626);
			13423: out = 16'(-4893);
			13424: out = 16'(40);
			13425: out = 16'(-4159);
			13426: out = 16'(-10084);
			13427: out = 16'(-7345);
			13428: out = 16'(4518);
			13429: out = 16'(8786);
			13430: out = 16'(4987);
			13431: out = 16'(-2087);
			13432: out = 16'(-8798);
			13433: out = 16'(-13064);
			13434: out = 16'(-5587);
			13435: out = 16'(9083);
			13436: out = 16'(11443);
			13437: out = 16'(4359);
			13438: out = 16'(-1108);
			13439: out = 16'(1685);
			13440: out = 16'(5606);
			13441: out = 16'(-2336);
			13442: out = 16'(-9487);
			13443: out = 16'(-7286);
			13444: out = 16'(-1359);
			13445: out = 16'(6924);
			13446: out = 16'(9237);
			13447: out = 16'(6599);
			13448: out = 16'(1111);
			13449: out = 16'(-2036);
			13450: out = 16'(-2941);
			13451: out = 16'(-1932);
			13452: out = 16'(249);
			13453: out = 16'(-334);
			13454: out = 16'(688);
			13455: out = 16'(-1519);
			13456: out = 16'(-3303);
			13457: out = 16'(-201);
			13458: out = 16'(9347);
			13459: out = 16'(11299);
			13460: out = 16'(3251);
			13461: out = 16'(-11817);
			13462: out = 16'(-3900);
			13463: out = 16'(2450);
			13464: out = 16'(2123);
			13465: out = 16'(3142);
			13466: out = 16'(8509);
			13467: out = 16'(9908);
			13468: out = 16'(4315);
			13469: out = 16'(-4033);
			13470: out = 16'(-11602);
			13471: out = 16'(-8228);
			13472: out = 16'(3865);
			13473: out = 16'(11090);
			13474: out = 16'(927);
			13475: out = 16'(-5633);
			13476: out = 16'(-4921);
			13477: out = 16'(1275);
			13478: out = 16'(6711);
			13479: out = 16'(3323);
			13480: out = 16'(2930);
			13481: out = 16'(4698);
			13482: out = 16'(3880);
			13483: out = 16'(-9369);
			13484: out = 16'(-11299);
			13485: out = 16'(-664);
			13486: out = 16'(7634);
			13487: out = 16'(7393);
			13488: out = 16'(3601);
			13489: out = 16'(1090);
			13490: out = 16'(-898);
			13491: out = 16'(-1670);
			13492: out = 16'(-6388);
			13493: out = 16'(-10013);
			13494: out = 16'(-7835);
			13495: out = 16'(2841);
			13496: out = 16'(7509);
			13497: out = 16'(4217);
			13498: out = 16'(-3826);
			13499: out = 16'(-5027);
			13500: out = 16'(-14126);
			13501: out = 16'(-11562);
			13502: out = 16'(-785);
			13503: out = 16'(8612);
			13504: out = 16'(10215);
			13505: out = 16'(6931);
			13506: out = 16'(137);
			13507: out = 16'(-5781);
			13508: out = 16'(-8345);
			13509: out = 16'(-3006);
			13510: out = 16'(2312);
			13511: out = 16'(2865);
			13512: out = 16'(-4908);
			13513: out = 16'(-8144);
			13514: out = 16'(-9054);
			13515: out = 16'(-3716);
			13516: out = 16'(3259);
			13517: out = 16'(5685);
			13518: out = 16'(-3555);
			13519: out = 16'(-9637);
			13520: out = 16'(-1716);
			13521: out = 16'(6816);
			13522: out = 16'(522);
			13523: out = 16'(-5550);
			13524: out = 16'(5163);
			13525: out = 16'(8154);
			13526: out = 16'(6728);
			13527: out = 16'(403);
			13528: out = 16'(1476);
			13529: out = 16'(-1025);
			13530: out = 16'(2445);
			13531: out = 16'(-2881);
			13532: out = 16'(-7015);
			13533: out = 16'(-428);
			13534: out = 16'(2109);
			13535: out = 16'(-402);
			13536: out = 16'(1905);
			13537: out = 16'(12032);
			13538: out = 16'(8198);
			13539: out = 16'(-2448);
			13540: out = 16'(-7159);
			13541: out = 16'(1050);
			13542: out = 16'(6459);
			13543: out = 16'(-307);
			13544: out = 16'(-9430);
			13545: out = 16'(-7347);
			13546: out = 16'(1270);
			13547: out = 16'(3838);
			13548: out = 16'(2150);
			13549: out = 16'(3339);
			13550: out = 16'(2227);
			13551: out = 16'(3139);
			13552: out = 16'(1672);
			13553: out = 16'(1460);
			13554: out = 16'(-284);
			13555: out = 16'(2442);
			13556: out = 16'(925);
			13557: out = 16'(-323);
			13558: out = 16'(-818);
			13559: out = 16'(-5370);
			13560: out = 16'(-7147);
			13561: out = 16'(-2086);
			13562: out = 16'(2799);
			13563: out = 16'(8592);
			13564: out = 16'(3988);
			13565: out = 16'(2798);
			13566: out = 16'(1021);
			13567: out = 16'(-1310);
			13568: out = 16'(-12362);
			13569: out = 16'(-5835);
			13570: out = 16'(7729);
			13571: out = 16'(7146);
			13572: out = 16'(529);
			13573: out = 16'(7752);
			13574: out = 16'(14372);
			13575: out = 16'(436);
			13576: out = 16'(-19284);
			13577: out = 16'(-22994);
			13578: out = 16'(-10039);
			13579: out = 16'(-1698);
			13580: out = 16'(11262);
			13581: out = 16'(15823);
			13582: out = 16'(10295);
			13583: out = 16'(-5223);
			13584: out = 16'(-9638);
			13585: out = 16'(-4725);
			13586: out = 16'(3978);
			13587: out = 16'(2946);
			13588: out = 16'(-4330);
			13589: out = 16'(-2461);
			13590: out = 16'(2926);
			13591: out = 16'(2749);
			13592: out = 16'(587);
			13593: out = 16'(-512);
			13594: out = 16'(-1228);
			13595: out = 16'(-7807);
			13596: out = 16'(-16106);
			13597: out = 16'(-11177);
			13598: out = 16'(1519);
			13599: out = 16'(11115);
			13600: out = 16'(14051);
			13601: out = 16'(6587);
			13602: out = 16'(2476);
			13603: out = 16'(-3113);
			13604: out = 16'(-4584);
			13605: out = 16'(-3719);
			13606: out = 16'(2621);
			13607: out = 16'(-2341);
			13608: out = 16'(-6909);
			13609: out = 16'(-464);
			13610: out = 16'(11499);
			13611: out = 16'(352);
			13612: out = 16'(-16035);
			13613: out = 16'(-8754);
			13614: out = 16'(3202);
			13615: out = 16'(4819);
			13616: out = 16'(-486);
			13617: out = 16'(4776);
			13618: out = 16'(8840);
			13619: out = 16'(7748);
			13620: out = 16'(-423);
			13621: out = 16'(-2865);
			13622: out = 16'(289);
			13623: out = 16'(4160);
			13624: out = 16'(-544);
			13625: out = 16'(-7983);
			13626: out = 16'(-10400);
			13627: out = 16'(-5167);
			13628: out = 16'(3347);
			13629: out = 16'(10303);
			13630: out = 16'(11651);
			13631: out = 16'(5856);
			13632: out = 16'(-3216);
			13633: out = 16'(-10928);
			13634: out = 16'(-15621);
			13635: out = 16'(-15369);
			13636: out = 16'(-6532);
			13637: out = 16'(11443);
			13638: out = 16'(23074);
			13639: out = 16'(16820);
			13640: out = 16'(-1739);
			13641: out = 16'(-17673);
			13642: out = 16'(-18616);
			13643: out = 16'(-987);
			13644: out = 16'(-2870);
			13645: out = 16'(-5002);
			13646: out = 16'(1144);
			13647: out = 16'(10440);
			13648: out = 16'(10275);
			13649: out = 16'(5361);
			13650: out = 16'(-626);
			13651: out = 16'(-3585);
			13652: out = 16'(-3382);
			13653: out = 16'(-346);
			13654: out = 16'(-2506);
			13655: out = 16'(-7242);
			13656: out = 16'(1620);
			13657: out = 16'(10198);
			13658: out = 16'(9835);
			13659: out = 16'(-735);
			13660: out = 16'(-15285);
			13661: out = 16'(-9199);
			13662: out = 16'(2268);
			13663: out = 16'(4274);
			13664: out = 16'(1268);
			13665: out = 16'(7648);
			13666: out = 16'(13152);
			13667: out = 16'(8843);
			13668: out = 16'(972);
			13669: out = 16'(-7804);
			13670: out = 16'(-2382);
			13671: out = 16'(2904);
			13672: out = 16'(-1892);
			13673: out = 16'(-14981);
			13674: out = 16'(-8088);
			13675: out = 16'(6870);
			13676: out = 16'(9075);
			13677: out = 16'(8620);
			13678: out = 16'(-1057);
			13679: out = 16'(-613);
			13680: out = 16'(2796);
			13681: out = 16'(5030);
			13682: out = 16'(-14547);
			13683: out = 16'(-17582);
			13684: out = 16'(-1675);
			13685: out = 16'(9820);
			13686: out = 16'(8746);
			13687: out = 16'(3941);
			13688: out = 16'(3239);
			13689: out = 16'(3971);
			13690: out = 16'(-6384);
			13691: out = 16'(-13583);
			13692: out = 16'(-13079);
			13693: out = 16'(-2980);
			13694: out = 16'(408);
			13695: out = 16'(7858);
			13696: out = 16'(5653);
			13697: out = 16'(2018);
			13698: out = 16'(4588);
			13699: out = 16'(7782);
			13700: out = 16'(-18);
			13701: out = 16'(-9150);
			13702: out = 16'(-6437);
			13703: out = 16'(-1917);
			13704: out = 16'(-5245);
			13705: out = 16'(-7848);
			13706: out = 16'(1888);
			13707: out = 16'(11050);
			13708: out = 16'(9143);
			13709: out = 16'(2322);
			13710: out = 16'(-217);
			13711: out = 16'(-3700);
			13712: out = 16'(-9393);
			13713: out = 16'(-10147);
			13714: out = 16'(1835);
			13715: out = 16'(13204);
			13716: out = 16'(18932);
			13717: out = 16'(11300);
			13718: out = 16'(-2267);
			13719: out = 16'(-15005);
			13720: out = 16'(-14179);
			13721: out = 16'(-7117);
			13722: out = 16'(-439);
			13723: out = 16'(3443);
			13724: out = 16'(9438);
			13725: out = 16'(8984);
			13726: out = 16'(1072);
			13727: out = 16'(-8491);
			13728: out = 16'(-7104);
			13729: out = 16'(-3491);
			13730: out = 16'(-4269);
			13731: out = 16'(-6166);
			13732: out = 16'(9285);
			13733: out = 16'(14123);
			13734: out = 16'(12257);
			13735: out = 16'(2467);
			13736: out = 16'(-4245);
			13737: out = 16'(-6922);
			13738: out = 16'(102);
			13739: out = 16'(3077);
			13740: out = 16'(-97);
			13741: out = 16'(-8535);
			13742: out = 16'(-2925);
			13743: out = 16'(4353);
			13744: out = 16'(3308);
			13745: out = 16'(465);
			13746: out = 16'(154);
			13747: out = 16'(-1147);
			13748: out = 16'(-3671);
			13749: out = 16'(-1760);
			13750: out = 16'(3782);
			13751: out = 16'(2314);
			13752: out = 16'(-2837);
			13753: out = 16'(315);
			13754: out = 16'(3410);
			13755: out = 16'(310);
			13756: out = 16'(-2775);
			13757: out = 16'(6637);
			13758: out = 16'(6068);
			13759: out = 16'(405);
			13760: out = 16'(-7775);
			13761: out = 16'(-7065);
			13762: out = 16'(-3000);
			13763: out = 16'(3232);
			13764: out = 16'(6239);
			13765: out = 16'(7835);
			13766: out = 16'(342);
			13767: out = 16'(-4243);
			13768: out = 16'(-9332);
			13769: out = 16'(-10640);
			13770: out = 16'(-12424);
			13771: out = 16'(2410);
			13772: out = 16'(10717);
			13773: out = 16'(8807);
			13774: out = 16'(2964);
			13775: out = 16'(4373);
			13776: out = 16'(3136);
			13777: out = 16'(-4223);
			13778: out = 16'(-15037);
			13779: out = 16'(-7036);
			13780: out = 16'(5);
			13781: out = 16'(5845);
			13782: out = 16'(10536);
			13783: out = 16'(5403);
			13784: out = 16'(4867);
			13785: out = 16'(3472);
			13786: out = 16'(-2450);
			13787: out = 16'(-12587);
			13788: out = 16'(-12192);
			13789: out = 16'(-3639);
			13790: out = 16'(2795);
			13791: out = 16'(7925);
			13792: out = 16'(1164);
			13793: out = 16'(4415);
			13794: out = 16'(7484);
			13795: out = 16'(522);
			13796: out = 16'(-6671);
			13797: out = 16'(-6400);
			13798: out = 16'(-3053);
			13799: out = 16'(-1801);
			13800: out = 16'(4983);
			13801: out = 16'(11083);
			13802: out = 16'(9901);
			13803: out = 16'(3956);
			13804: out = 16'(-516);
			13805: out = 16'(1317);
			13806: out = 16'(-6280);
			13807: out = 16'(-16439);
			13808: out = 16'(-1281);
			13809: out = 16'(11477);
			13810: out = 16'(12590);
			13811: out = 16'(1825);
			13812: out = 16'(-4561);
			13813: out = 16'(-2417);
			13814: out = 16'(2181);
			13815: out = 16'(1275);
			13816: out = 16'(-42);
			13817: out = 16'(536);
			13818: out = 16'(941);
			13819: out = 16'(-3718);
			13820: out = 16'(-9033);
			13821: out = 16'(384);
			13822: out = 16'(8752);
			13823: out = 16'(12774);
			13824: out = 16'(5889);
			13825: out = 16'(-10843);
			13826: out = 16'(-15965);
			13827: out = 16'(-5293);
			13828: out = 16'(6948);
			13829: out = 16'(8752);
			13830: out = 16'(1711);
			13831: out = 16'(-73);
			13832: out = 16'(52);
			13833: out = 16'(-3417);
			13834: out = 16'(-10245);
			13835: out = 16'(-5336);
			13836: out = 16'(1620);
			13837: out = 16'(-1017);
			13838: out = 16'(-4256);
			13839: out = 16'(-4403);
			13840: out = 16'(-894);
			13841: out = 16'(-500);
			13842: out = 16'(-2038);
			13843: out = 16'(-1871);
			13844: out = 16'(-154);
			13845: out = 16'(1189);
			13846: out = 16'(5270);
			13847: out = 16'(5200);
			13848: out = 16'(1892);
			13849: out = 16'(-4913);
			13850: out = 16'(-6960);
			13851: out = 16'(-2020);
			13852: out = 16'(5205);
			13853: out = 16'(3425);
			13854: out = 16'(-4357);
			13855: out = 16'(-11568);
			13856: out = 16'(-6451);
			13857: out = 16'(407);
			13858: out = 16'(3960);
			13859: out = 16'(6949);
			13860: out = 16'(13171);
			13861: out = 16'(9446);
			13862: out = 16'(-3877);
			13863: out = 16'(-17106);
			13864: out = 16'(-12255);
			13865: out = 16'(1788);
			13866: out = 16'(14654);
			13867: out = 16'(20571);
			13868: out = 16'(8004);
			13869: out = 16'(-6745);
			13870: out = 16'(-10331);
			13871: out = 16'(261);
			13872: out = 16'(450);
			13873: out = 16'(-4231);
			13874: out = 16'(-4430);
			13875: out = 16'(4531);
			13876: out = 16'(11399);
			13877: out = 16'(5552);
			13878: out = 16'(-997);
			13879: out = 16'(1657);
			13880: out = 16'(9028);
			13881: out = 16'(-3084);
			13882: out = 16'(-16443);
			13883: out = 16'(-14868);
			13884: out = 16'(1188);
			13885: out = 16'(9227);
			13886: out = 16'(9612);
			13887: out = 16'(6570);
			13888: out = 16'(1903);
			13889: out = 16'(155);
			13890: out = 16'(-773);
			13891: out = 16'(960);
			13892: out = 16'(1815);
			13893: out = 16'(457);
			13894: out = 16'(-1881);
			13895: out = 16'(858);
			13896: out = 16'(3958);
			13897: out = 16'(-2615);
			13898: out = 16'(-5549);
			13899: out = 16'(-3508);
			13900: out = 16'(-142);
			13901: out = 16'(-441);
			13902: out = 16'(-6786);
			13903: out = 16'(-5113);
			13904: out = 16'(2427);
			13905: out = 16'(4108);
			13906: out = 16'(1140);
			13907: out = 16'(-1877);
			13908: out = 16'(-47);
			13909: out = 16'(2245);
			13910: out = 16'(1717);
			13911: out = 16'(-4657);
			13912: out = 16'(-8728);
			13913: out = 16'(-2845);
			13914: out = 16'(6680);
			13915: out = 16'(12490);
			13916: out = 16'(6900);
			13917: out = 16'(-1682);
			13918: out = 16'(-5819);
			13919: out = 16'(-10081);
			13920: out = 16'(-18541);
			13921: out = 16'(-19037);
			13922: out = 16'(1184);
			13923: out = 16'(14132);
			13924: out = 16'(12277);
			13925: out = 16'(2888);
			13926: out = 16'(927);
			13927: out = 16'(-1926);
			13928: out = 16'(-42);
			13929: out = 16'(-1614);
			13930: out = 16'(-3534);
			13931: out = 16'(-232);
			13932: out = 16'(3065);
			13933: out = 16'(3197);
			13934: out = 16'(1265);
			13935: out = 16'(2774);
			13936: out = 16'(4172);
			13937: out = 16'(3438);
			13938: out = 16'(-3715);
			13939: out = 16'(-13012);
			13940: out = 16'(-10781);
			13941: out = 16'(1809);
			13942: out = 16'(8063);
			13943: out = 16'(1013);
			13944: out = 16'(2731);
			13945: out = 16'(3004);
			13946: out = 16'(22);
			13947: out = 16'(-7266);
			13948: out = 16'(-6431);
			13949: out = 16'(-2487);
			13950: out = 16'(1964);
			13951: out = 16'(3722);
			13952: out = 16'(10465);
			13953: out = 16'(11793);
			13954: out = 16'(8862);
			13955: out = 16'(-2516);
			13956: out = 16'(-17196);
			13957: out = 16'(-10649);
			13958: out = 16'(5997);
			13959: out = 16'(10172);
			13960: out = 16'(-20);
			13961: out = 16'(-733);
			13962: out = 16'(3406);
			13963: out = 16'(1113);
			13964: out = 16'(-9695);
			13965: out = 16'(-1348);
			13966: out = 16'(1151);
			13967: out = 16'(-4800);
			13968: out = 16'(-13811);
			13969: out = 16'(-6950);
			13970: out = 16'(2006);
			13971: out = 16'(7414);
			13972: out = 16'(9705);
			13973: out = 16'(13845);
			13974: out = 16'(11958);
			13975: out = 16'(406);
			13976: out = 16'(-11386);
			13977: out = 16'(-7313);
			13978: out = 16'(-2243);
			13979: out = 16'(2746);
			13980: out = 16'(5179);
			13981: out = 16'(8972);
			13982: out = 16'(816);
			13983: out = 16'(-2936);
			13984: out = 16'(-3961);
			13985: out = 16'(-837);
			13986: out = 16'(1891);
			13987: out = 16'(-1413);
			13988: out = 16'(-6500);
			13989: out = 16'(-4881);
			13990: out = 16'(3185);
			13991: out = 16'(10790);
			13992: out = 16'(10257);
			13993: out = 16'(4968);
			13994: out = 16'(830);
			13995: out = 16'(-195);
			13996: out = 16'(-3405);
			13997: out = 16'(-9802);
			13998: out = 16'(-13202);
			13999: out = 16'(-5132);
			14000: out = 16'(4706);
			14001: out = 16'(9775);
			14002: out = 16'(9951);
			14003: out = 16'(-4390);
			14004: out = 16'(-5975);
			14005: out = 16'(-5627);
			14006: out = 16'(-4854);
			14007: out = 16'(-3134);
			14008: out = 16'(6488);
			14009: out = 16'(7372);
			14010: out = 16'(88);
			14011: out = 16'(-4644);
			14012: out = 16'(2833);
			14013: out = 16'(6760);
			14014: out = 16'(-3135);
			14015: out = 16'(-23851);
			14016: out = 16'(-8594);
			14017: out = 16'(5243);
			14018: out = 16'(6658);
			14019: out = 16'(126);
			14020: out = 16'(8687);
			14021: out = 16'(8280);
			14022: out = 16'(4487);
			14023: out = 16'(-1151);
			14024: out = 16'(303);
			14025: out = 16'(-6430);
			14026: out = 16'(-5453);
			14027: out = 16'(1492);
			14028: out = 16'(2229);
			14029: out = 16'(2594);
			14030: out = 16'(4672);
			14031: out = 16'(5987);
			14032: out = 16'(-2555);
			14033: out = 16'(-9863);
			14034: out = 16'(-10709);
			14035: out = 16'(193);
			14036: out = 16'(7247);
			14037: out = 16'(3542);
			14038: out = 16'(-4213);
			14039: out = 16'(-1699);
			14040: out = 16'(5198);
			14041: out = 16'(8686);
			14042: out = 16'(1626);
			14043: out = 16'(1608);
			14044: out = 16'(3721);
			14045: out = 16'(736);
			14046: out = 16'(-14836);
			14047: out = 16'(-11100);
			14048: out = 16'(6213);
			14049: out = 16'(7071);
			14050: out = 16'(4907);
			14051: out = 16'(4841);
			14052: out = 16'(4715);
			14053: out = 16'(-6409);
			14054: out = 16'(-1175);
			14055: out = 16'(3352);
			14056: out = 16'(4563);
			14057: out = 16'(-1309);
			14058: out = 16'(-436);
			14059: out = 16'(4679);
			14060: out = 16'(6262);
			14061: out = 16'(-3216);
			14062: out = 16'(-8201);
			14063: out = 16'(-12499);
			14064: out = 16'(-5960);
			14065: out = 16'(1191);
			14066: out = 16'(4998);
			14067: out = 16'(705);
			14068: out = 16'(2640);
			14069: out = 16'(6893);
			14070: out = 16'(7588);
			14071: out = 16'(3106);
			14072: out = 16'(635);
			14073: out = 16'(-3241);
			14074: out = 16'(-9925);
			14075: out = 16'(-6341);
			14076: out = 16'(-2321);
			14077: out = 16'(883);
			14078: out = 16'(3550);
			14079: out = 16'(11167);
			14080: out = 16'(4672);
			14081: out = 16'(-9303);
			14082: out = 16'(-18246);
			14083: out = 16'(-7489);
			14084: out = 16'(-3348);
			14085: out = 16'(-1344);
			14086: out = 16'(5360);
			14087: out = 16'(15153);
			14088: out = 16'(11602);
			14089: out = 16'(-4869);
			14090: out = 16'(-16181);
			14091: out = 16'(-5104);
			14092: out = 16'(3649);
			14093: out = 16'(3912);
			14094: out = 16'(-3598);
			14095: out = 16'(-6258);
			14096: out = 16'(-6222);
			14097: out = 16'(-2156);
			14098: out = 16'(-1015);
			14099: out = 16'(1683);
			14100: out = 16'(8498);
			14101: out = 16'(7490);
			14102: out = 16'(1481);
			14103: out = 16'(-3141);
			14104: out = 16'(-1468);
			14105: out = 16'(-4561);
			14106: out = 16'(-2309);
			14107: out = 16'(7822);
			14108: out = 16'(16693);
			14109: out = 16'(5345);
			14110: out = 16'(-9947);
			14111: out = 16'(-15493);
			14112: out = 16'(-3118);
			14113: out = 16'(1982);
			14114: out = 16'(4940);
			14115: out = 16'(1324);
			14116: out = 16'(1247);
			14117: out = 16'(6894);
			14118: out = 16'(10334);
			14119: out = 16'(4912);
			14120: out = 16'(-921);
			14121: out = 16'(-529);
			14122: out = 16'(848);
			14123: out = 16'(-3373);
			14124: out = 16'(-7670);
			14125: out = 16'(-6569);
			14126: out = 16'(2020);
			14127: out = 16'(1801);
			14128: out = 16'(-936);
			14129: out = 16'(861);
			14130: out = 16'(10688);
			14131: out = 16'(1854);
			14132: out = 16'(-11771);
			14133: out = 16'(-15142);
			14134: out = 16'(-1685);
			14135: out = 16'(3240);
			14136: out = 16'(4440);
			14137: out = 16'(6295);
			14138: out = 16'(6378);
			14139: out = 16'(1682);
			14140: out = 16'(-4773);
			14141: out = 16'(-8683);
			14142: out = 16'(-5869);
			14143: out = 16'(2961);
			14144: out = 16'(9309);
			14145: out = 16'(3542);
			14146: out = 16'(-10040);
			14147: out = 16'(-13865);
			14148: out = 16'(-5655);
			14149: out = 16'(1736);
			14150: out = 16'(52);
			14151: out = 16'(-7064);
			14152: out = 16'(3828);
			14153: out = 16'(12826);
			14154: out = 16'(5586);
			14155: out = 16'(-10267);
			14156: out = 16'(-10110);
			14157: out = 16'(1978);
			14158: out = 16'(6803);
			14159: out = 16'(-2665);
			14160: out = 16'(-3903);
			14161: out = 16'(-274);
			14162: out = 16'(2269);
			14163: out = 16'(-2766);
			14164: out = 16'(4510);
			14165: out = 16'(4378);
			14166: out = 16'(2718);
			14167: out = 16'(-721);
			14168: out = 16'(801);
			14169: out = 16'(-5632);
			14170: out = 16'(-5644);
			14171: out = 16'(2886);
			14172: out = 16'(11269);
			14173: out = 16'(2472);
			14174: out = 16'(-9104);
			14175: out = 16'(-12143);
			14176: out = 16'(-3638);
			14177: out = 16'(-543);
			14178: out = 16'(2414);
			14179: out = 16'(4432);
			14180: out = 16'(4131);
			14181: out = 16'(9267);
			14182: out = 16'(8078);
			14183: out = 16'(-2156);
			14184: out = 16'(-18294);
			14185: out = 16'(-5111);
			14186: out = 16'(4034);
			14187: out = 16'(11170);
			14188: out = 16'(10730);
			14189: out = 16'(8838);
			14190: out = 16'(-4733);
			14191: out = 16'(-11251);
			14192: out = 16'(-9158);
			14193: out = 16'(119);
			14194: out = 16'(-298);
			14195: out = 16'(2713);
			14196: out = 16'(1898);
			14197: out = 16'(-3156);
			14198: out = 16'(-5204);
			14199: out = 16'(7186);
			14200: out = 16'(12078);
			14201: out = 16'(1460);
			14202: out = 16'(23);
			14203: out = 16'(6364);
			14204: out = 16'(6637);
			14205: out = 16'(-5141);
			14206: out = 16'(-11279);
			14207: out = 16'(391);
			14208: out = 16'(11416);
			14209: out = 16'(6579);
			14210: out = 16'(-1804);
			14211: out = 16'(-4009);
			14212: out = 16'(-2756);
			14213: out = 16'(-5735);
			14214: out = 16'(-7153);
			14215: out = 16'(3206);
			14216: out = 16'(8470);
			14217: out = 16'(660);
			14218: out = 16'(-8317);
			14219: out = 16'(-2636);
			14220: out = 16'(8182);
			14221: out = 16'(7569);
			14222: out = 16'(-1419);
			14223: out = 16'(-6593);
			14224: out = 16'(-2581);
			14225: out = 16'(-853);
			14226: out = 16'(-2369);
			14227: out = 16'(2114);
			14228: out = 16'(6818);
			14229: out = 16'(5640);
			14230: out = 16'(1238);
			14231: out = 16'(-828);
			14232: out = 16'(-6744);
			14233: out = 16'(-14799);
			14234: out = 16'(-11044);
			14235: out = 16'(9425);
			14236: out = 16'(5999);
			14237: out = 16'(-889);
			14238: out = 16'(-1864);
			14239: out = 16'(4071);
			14240: out = 16'(-8346);
			14241: out = 16'(-18350);
			14242: out = 16'(-14097);
			14243: out = 16'(4537);
			14244: out = 16'(9392);
			14245: out = 16'(7486);
			14246: out = 16'(2903);
			14247: out = 16'(458);
			14248: out = 16'(-3408);
			14249: out = 16'(-4389);
			14250: out = 16'(3634);
			14251: out = 16'(12193);
			14252: out = 16'(6664);
			14253: out = 16'(-5238);
			14254: out = 16'(-9951);
			14255: out = 16'(-3139);
			14256: out = 16'(122);
			14257: out = 16'(10109);
			14258: out = 16'(5314);
			14259: out = 16'(1214);
			14260: out = 16'(-3156);
			14261: out = 16'(-13007);
			14262: out = 16'(-16904);
			14263: out = 16'(-5325);
			14264: out = 16'(11775);
			14265: out = 16'(18344);
			14266: out = 16'(9595);
			14267: out = 16'(2592);
			14268: out = 16'(510);
			14269: out = 16'(-475);
			14270: out = 16'(-12395);
			14271: out = 16'(-9194);
			14272: out = 16'(4167);
			14273: out = 16'(4804);
			14274: out = 16'(9229);
			14275: out = 16'(1832);
			14276: out = 16'(-2904);
			14277: out = 16'(-4688);
			14278: out = 16'(9462);
			14279: out = 16'(3360);
			14280: out = 16'(-2790);
			14281: out = 16'(-6162);
			14282: out = 16'(-5840);
			14283: out = 16'(-12688);
			14284: out = 16'(-4692);
			14285: out = 16'(12107);
			14286: out = 16'(14486);
			14287: out = 16'(9496);
			14288: out = 16'(2208);
			14289: out = 16'(-1289);
			14290: out = 16'(-3667);
			14291: out = 16'(-17713);
			14292: out = 16'(-16287);
			14293: out = 16'(1066);
			14294: out = 16'(13701);
			14295: out = 16'(8139);
			14296: out = 16'(5525);
			14297: out = 16'(5322);
			14298: out = 16'(99);
			14299: out = 16'(-6477);
			14300: out = 16'(-12673);
			14301: out = 16'(-4920);
			14302: out = 16'(6782);
			14303: out = 16'(8642);
			14304: out = 16'(2039);
			14305: out = 16'(-1888);
			14306: out = 16'(-4699);
			14307: out = 16'(-12007);
			14308: out = 16'(-9236);
			14309: out = 16'(-1475);
			14310: out = 16'(3110);
			14311: out = 16'(-334);
			14312: out = 16'(-1940);
			14313: out = 16'(1269);
			14314: out = 16'(6150);
			14315: out = 16'(8810);
			14316: out = 16'(11538);
			14317: out = 16'(8762);
			14318: out = 16'(-3271);
			14319: out = 16'(-18716);
			14320: out = 16'(-17319);
			14321: out = 16'(-5513);
			14322: out = 16'(7863);
			14323: out = 16'(10119);
			14324: out = 16'(5139);
			14325: out = 16'(2797);
			14326: out = 16'(504);
			14327: out = 16'(-6635);
			14328: out = 16'(-15628);
			14329: out = 16'(-2841);
			14330: out = 16'(4911);
			14331: out = 16'(1890);
			14332: out = 16'(-4547);
			14333: out = 16'(663);
			14334: out = 16'(6638);
			14335: out = 16'(7215);
			14336: out = 16'(3099);
			14337: out = 16'(2872);
			14338: out = 16'(2384);
			14339: out = 16'(1524);
			14340: out = 16'(-700);
			14341: out = 16'(-19);
			14342: out = 16'(-2473);
			14343: out = 16'(-1656);
			14344: out = 16'(770);
			14345: out = 16'(2270);
			14346: out = 16'(-624);
			14347: out = 16'(-2672);
			14348: out = 16'(-1142);
			14349: out = 16'(2999);
			14350: out = 16'(4477);
			14351: out = 16'(2798);
			14352: out = 16'(164);
			14353: out = 16'(44);
			14354: out = 16'(576);
			14355: out = 16'(3666);
			14356: out = 16'(4838);
			14357: out = 16'(3323);
			14358: out = 16'(-3048);
			14359: out = 16'(-1185);
			14360: out = 16'(280);
			14361: out = 16'(1451);
			14362: out = 16'(2102);
			14363: out = 16'(6107);
			14364: out = 16'(3168);
			14365: out = 16'(-4836);
			14366: out = 16'(-13772);
			14367: out = 16'(-1947);
			14368: out = 16'(-2665);
			14369: out = 16'(-7600);
			14370: out = 16'(-7975);
			14371: out = 16'(1657);
			14372: out = 16'(4711);
			14373: out = 16'(3198);
			14374: out = 16'(-513);
			14375: out = 16'(1652);
			14376: out = 16'(-5432);
			14377: out = 16'(-2791);
			14378: out = 16'(4133);
			14379: out = 16'(5557);
			14380: out = 16'(-197);
			14381: out = 16'(1212);
			14382: out = 16'(4761);
			14383: out = 16'(41);
			14384: out = 16'(1513);
			14385: out = 16'(151);
			14386: out = 16'(-1954);
			14387: out = 16'(-7332);
			14388: out = 16'(-2711);
			14389: out = 16'(-1469);
			14390: out = 16'(610);
			14391: out = 16'(-216);
			14392: out = 16'(3106);
			14393: out = 16'(-3707);
			14394: out = 16'(-3456);
			14395: out = 16'(1569);
			14396: out = 16'(7018);
			14397: out = 16'(-3902);
			14398: out = 16'(-3797);
			14399: out = 16'(4785);
			14400: out = 16'(9255);
			14401: out = 16'(1560);
			14402: out = 16'(-1299);
			14403: out = 16'(915);
			14404: out = 16'(1823);
			14405: out = 16'(-2263);
			14406: out = 16'(-1456);
			14407: out = 16'(456);
			14408: out = 16'(-408);
			14409: out = 16'(-25);
			14410: out = 16'(1307);
			14411: out = 16'(1962);
			14412: out = 16'(-1429);
			14413: out = 16'(-3386);
			14414: out = 16'(-1858);
			14415: out = 16'(3838);
			14416: out = 16'(3888);
			14417: out = 16'(-2983);
			14418: out = 16'(-6603);
			14419: out = 16'(-3109);
			14420: out = 16'(644);
			14421: out = 16'(-405);
			14422: out = 16'(-59);
			14423: out = 16'(4884);
			14424: out = 16'(7931);
			14425: out = 16'(1965);
			14426: out = 16'(-10513);
			14427: out = 16'(-9485);
			14428: out = 16'(1575);
			14429: out = 16'(7988);
			14430: out = 16'(5951);
			14431: out = 16'(2728);
			14432: out = 16'(1818);
			14433: out = 16'(-585);
			14434: out = 16'(-2488);
			14435: out = 16'(-5036);
			14436: out = 16'(3100);
			14437: out = 16'(8973);
			14438: out = 16'(4113);
			14439: out = 16'(-7546);
			14440: out = 16'(-5725);
			14441: out = 16'(2847);
			14442: out = 16'(3260);
			14443: out = 16'(611);
			14444: out = 16'(-1639);
			14445: out = 16'(2460);
			14446: out = 16'(5281);
			14447: out = 16'(4638);
			14448: out = 16'(253);
			14449: out = 16'(2033);
			14450: out = 16'(5242);
			14451: out = 16'(1408);
			14452: out = 16'(-2101);
			14453: out = 16'(-2865);
			14454: out = 16'(845);
			14455: out = 16'(2232);
			14456: out = 16'(-2662);
			14457: out = 16'(-10231);
			14458: out = 16'(-9685);
			14459: out = 16'(860);
			14460: out = 16'(-737);
			14461: out = 16'(227);
			14462: out = 16'(-1391);
			14463: out = 16'(-1033);
			14464: out = 16'(161);
			14465: out = 16'(2534);
			14466: out = 16'(647);
			14467: out = 16'(463);
			14468: out = 16'(2677);
			14469: out = 16'(1606);
			14470: out = 16'(-4768);
			14471: out = 16'(-3774);
			14472: out = 16'(6503);
			14473: out = 16'(10179);
			14474: out = 16'(70);
			14475: out = 16'(-8093);
			14476: out = 16'(-5339);
			14477: out = 16'(-2794);
			14478: out = 16'(-11555);
			14479: out = 16'(-14367);
			14480: out = 16'(-919);
			14481: out = 16'(6828);
			14482: out = 16'(3690);
			14483: out = 16'(-1204);
			14484: out = 16'(1276);
			14485: out = 16'(692);
			14486: out = 16'(1932);
			14487: out = 16'(492);
			14488: out = 16'(-170);
			14489: out = 16'(-2824);
			14490: out = 16'(-4596);
			14491: out = 16'(-2166);
			14492: out = 16'(3239);
			14493: out = 16'(3108);
			14494: out = 16'(3370);
			14495: out = 16'(1928);
			14496: out = 16'(2506);
			14497: out = 16'(-1218);
			14498: out = 16'(2087);
			14499: out = 16'(-6005);
			14500: out = 16'(-4307);
			14501: out = 16'(3586);
			14502: out = 16'(6020);
			14503: out = 16'(-1670);
			14504: out = 16'(-797);
			14505: out = 16'(4964);
			14506: out = 16'(-704);
			14507: out = 16'(-4363);
			14508: out = 16'(-775);
			14509: out = 16'(5179);
			14510: out = 16'(-958);
			14511: out = 16'(7346);
			14512: out = 16'(6707);
			14513: out = 16'(3112);
			14514: out = 16'(-3606);
			14515: out = 16'(-91);
			14516: out = 16'(-158);
			14517: out = 16'(2428);
			14518: out = 16'(3512);
			14519: out = 16'(-2523);
			14520: out = 16'(-7152);
			14521: out = 16'(-6868);
			14522: out = 16'(-120);
			14523: out = 16'(9190);
			14524: out = 16'(8746);
			14525: out = 16'(2407);
			14526: out = 16'(-5332);
			14527: out = 16'(-7847);
			14528: out = 16'(-6777);
			14529: out = 16'(-867);
			14530: out = 16'(3382);
			14531: out = 16'(4742);
			14532: out = 16'(6118);
			14533: out = 16'(7616);
			14534: out = 16'(4716);
			14535: out = 16'(-1224);
			14536: out = 16'(1738);
			14537: out = 16'(478);
			14538: out = 16'(-3893);
			14539: out = 16'(-8900);
			14540: out = 16'(-5520);
			14541: out = 16'(3976);
			14542: out = 16'(6999);
			14543: out = 16'(-2271);
			14544: out = 16'(-9557);
			14545: out = 16'(-7825);
			14546: out = 16'(6100);
			14547: out = 16'(10371);
			14548: out = 16'(4707);
			14549: out = 16'(-14818);
			14550: out = 16'(-5133);
			14551: out = 16'(8960);
			14552: out = 16'(3089);
			14553: out = 16'(-17462);
			14554: out = 16'(-15906);
			14555: out = 16'(112);
			14556: out = 16'(4314);
			14557: out = 16'(-1134);
			14558: out = 16'(-3468);
			14559: out = 16'(5870);
			14560: out = 16'(10802);
			14561: out = 16'(2283);
			14562: out = 16'(-4106);
			14563: out = 16'(-3238);
			14564: out = 16'(816);
			14565: out = 16'(-429);
			14566: out = 16'(160);
			14567: out = 16'(-3234);
			14568: out = 16'(-6017);
			14569: out = 16'(-3883);
			14570: out = 16'(5535);
			14571: out = 16'(6841);
			14572: out = 16'(1101);
			14573: out = 16'(-1643);
			14574: out = 16'(3548);
			14575: out = 16'(495);
			14576: out = 16'(-15245);
			14577: out = 16'(-24122);
			14578: out = 16'(1564);
			14579: out = 16'(15003);
			14580: out = 16'(12920);
			14581: out = 16'(2799);
			14582: out = 16'(-603);
			14583: out = 16'(3408);
			14584: out = 16'(2330);
			14585: out = 16'(-4528);
			14586: out = 16'(-7148);
			14587: out = 16'(-422);
			14588: out = 16'(2874);
			14589: out = 16'(1451);
			14590: out = 16'(-575);
			14591: out = 16'(-7502);
			14592: out = 16'(-2892);
			14593: out = 16'(3852);
			14594: out = 16'(3703);
			14595: out = 16'(-9874);
			14596: out = 16'(-6412);
			14597: out = 16'(2957);
			14598: out = 16'(8758);
			14599: out = 16'(5763);
			14600: out = 16'(7022);
			14601: out = 16'(3858);
			14602: out = 16'(-4948);
			14603: out = 16'(-16683);
			14604: out = 16'(-11871);
			14605: out = 16'(-3794);
			14606: out = 16'(2688);
			14607: out = 16'(6549);
			14608: out = 16'(15209);
			14609: out = 16'(15211);
			14610: out = 16'(8202);
			14611: out = 16'(-3480);
			14612: out = 16'(-12841);
			14613: out = 16'(-14777);
			14614: out = 16'(-9741);
			14615: out = 16'(-2842);
			14616: out = 16'(3054);
			14617: out = 16'(8202);
			14618: out = 16'(8338);
			14619: out = 16'(3834);
			14620: out = 16'(319);
			14621: out = 16'(-2754);
			14622: out = 16'(718);
			14623: out = 16'(1601);
			14624: out = 16'(-4164);
			14625: out = 16'(-14863);
			14626: out = 16'(-6658);
			14627: out = 16'(9903);
			14628: out = 16'(14299);
			14629: out = 16'(7032);
			14630: out = 16'(533);
			14631: out = 16'(2538);
			14632: out = 16'(3234);
			14633: out = 16'(-2465);
			14634: out = 16'(-15574);
			14635: out = 16'(-9546);
			14636: out = 16'(9216);
			14637: out = 16'(15268);
			14638: out = 16'(462);
			14639: out = 16'(-11446);
			14640: out = 16'(-11628);
			14641: out = 16'(-5875);
			14642: out = 16'(-273);
			14643: out = 16'(3095);
			14644: out = 16'(8003);
			14645: out = 16'(10690);
			14646: out = 16'(7234);
			14647: out = 16'(-2433);
			14648: out = 16'(-10060);
			14649: out = 16'(-12547);
			14650: out = 16'(-16161);
			14651: out = 16'(-224);
			14652: out = 16'(10644);
			14653: out = 16'(7559);
			14654: out = 16'(-6042);
			14655: out = 16'(-254);
			14656: out = 16'(4192);
			14657: out = 16'(5015);
			14658: out = 16'(5441);
			14659: out = 16'(8344);
			14660: out = 16'(3885);
			14661: out = 16'(-8315);
			14662: out = 16'(-17353);
			14663: out = 16'(-10409);
			14664: out = 16'(2402);
			14665: out = 16'(7150);
			14666: out = 16'(6539);
			14667: out = 16'(7935);
			14668: out = 16'(7371);
			14669: out = 16'(-626);
			14670: out = 16'(-9369);
			14671: out = 16'(-10156);
			14672: out = 16'(-1942);
			14673: out = 16'(1350);
			14674: out = 16'(3698);
			14675: out = 16'(9094);
			14676: out = 16'(7018);
			14677: out = 16'(-1864);
			14678: out = 16'(-5551);
			14679: out = 16'(937);
			14680: out = 16'(227);
			14681: out = 16'(-6615);
			14682: out = 16'(-8782);
			14683: out = 16'(2399);
			14684: out = 16'(11659);
			14685: out = 16'(5188);
			14686: out = 16'(-7135);
			14687: out = 16'(-10416);
			14688: out = 16'(-2835);
			14689: out = 16'(-777);
			14690: out = 16'(-805);
			14691: out = 16'(3149);
			14692: out = 16'(9274);
			14693: out = 16'(12150);
			14694: out = 16'(6747);
			14695: out = 16'(31);
			14696: out = 16'(-2823);
			14697: out = 16'(-5187);
			14698: out = 16'(-5330);
			14699: out = 16'(-4419);
			14700: out = 16'(-1833);
			14701: out = 16'(-329);
			14702: out = 16'(6589);
			14703: out = 16'(9239);
			14704: out = 16'(5028);
			14705: out = 16'(479);
			14706: out = 16'(-388);
			14707: out = 16'(4548);
			14708: out = 16'(4901);
			14709: out = 16'(-3224);
			14710: out = 16'(-12072);
			14711: out = 16'(-9089);
			14712: out = 16'(1556);
			14713: out = 16'(7200);
			14714: out = 16'(13284);
			14715: out = 16'(10467);
			14716: out = 16'(2549);
			14717: out = 16'(-8436);
			14718: out = 16'(-10288);
			14719: out = 16'(-6072);
			14720: out = 16'(4409);
			14721: out = 16'(9352);
			14722: out = 16'(7006);
			14723: out = 16'(-1153);
			14724: out = 16'(-1894);
			14725: out = 16'(1534);
			14726: out = 16'(1619);
			14727: out = 16'(-10633);
			14728: out = 16'(-10467);
			14729: out = 16'(2058);
			14730: out = 16'(6461);
			14731: out = 16'(2324);
			14732: out = 16'(-5028);
			14733: out = 16'(-1245);
			14734: out = 16'(6787);
			14735: out = 16'(7281);
			14736: out = 16'(-4943);
			14737: out = 16'(-12298);
			14738: out = 16'(-7288);
			14739: out = 16'(1628);
			14740: out = 16'(3642);
			14741: out = 16'(4078);
			14742: out = 16'(3534);
			14743: out = 16'(-2781);
			14744: out = 16'(956);
			14745: out = 16'(2158);
			14746: out = 16'(-3876);
			14747: out = 16'(-13177);
			14748: out = 16'(-12477);
			14749: out = 16'(736);
			14750: out = 16'(9479);
			14751: out = 16'(5998);
			14752: out = 16'(885);
			14753: out = 16'(3365);
			14754: out = 16'(5486);
			14755: out = 16'(889);
			14756: out = 16'(-3423);
			14757: out = 16'(-1054);
			14758: out = 16'(2968);
			14759: out = 16'(2354);
			14760: out = 16'(-2705);
			14761: out = 16'(-3822);
			14762: out = 16'(-4944);
			14763: out = 16'(-4156);
			14764: out = 16'(661);
			14765: out = 16'(11799);
			14766: out = 16'(9387);
			14767: out = 16'(-1173);
			14768: out = 16'(-7338);
			14769: out = 16'(-1711);
			14770: out = 16'(-879);
			14771: out = 16'(-3737);
			14772: out = 16'(-1221);
			14773: out = 16'(2272);
			14774: out = 16'(4225);
			14775: out = 16'(-3882);
			14776: out = 16'(-10860);
			14777: out = 16'(-95);
			14778: out = 16'(5676);
			14779: out = 16'(5140);
			14780: out = 16'(2585);
			14781: out = 16'(6743);
			14782: out = 16'(-934);
			14783: out = 16'(-6192);
			14784: out = 16'(-7143);
			14785: out = 16'(-1879);
			14786: out = 16'(3311);
			14787: out = 16'(7122);
			14788: out = 16'(6120);
			14789: out = 16'(1410);
			14790: out = 16'(62);
			14791: out = 16'(-2559);
			14792: out = 16'(-1901);
			14793: out = 16'(116);
			14794: out = 16'(1031);
			14795: out = 16'(15);
			14796: out = 16'(-32);
			14797: out = 16'(-1025);
			14798: out = 16'(-3795);
			14799: out = 16'(-5626);
			14800: out = 16'(-378);
			14801: out = 16'(6915);
			14802: out = 16'(9958);
			14803: out = 16'(1397);
			14804: out = 16'(-2202);
			14805: out = 16'(-4588);
			14806: out = 16'(-8109);
			14807: out = 16'(-5896);
			14808: out = 16'(2541);
			14809: out = 16'(7298);
			14810: out = 16'(2989);
			14811: out = 16'(493);
			14812: out = 16'(-1171);
			14813: out = 16'(270);
			14814: out = 16'(-2089);
			14815: out = 16'(-7178);
			14816: out = 16'(-2232);
			14817: out = 16'(6740);
			14818: out = 16'(7839);
			14819: out = 16'(919);
			14820: out = 16'(-4622);
			14821: out = 16'(-4075);
			14822: out = 16'(-3300);
			14823: out = 16'(-5196);
			14824: out = 16'(-5447);
			14825: out = 16'(1022);
			14826: out = 16'(6676);
			14827: out = 16'(7144);
			14828: out = 16'(1321);
			14829: out = 16'(674);
			14830: out = 16'(-3906);
			14831: out = 16'(-8930);
			14832: out = 16'(-2767);
			14833: out = 16'(1580);
			14834: out = 16'(441);
			14835: out = 16'(-2670);
			14836: out = 16'(427);
			14837: out = 16'(145);
			14838: out = 16'(-159);
			14839: out = 16'(1259);
			14840: out = 16'(4319);
			14841: out = 16'(-77);
			14842: out = 16'(-6759);
			14843: out = 16'(-6001);
			14844: out = 16'(3833);
			14845: out = 16'(5390);
			14846: out = 16'(1323);
			14847: out = 16'(-209);
			14848: out = 16'(6384);
			14849: out = 16'(6654);
			14850: out = 16'(3078);
			14851: out = 16'(-3084);
			14852: out = 16'(-279);
			14853: out = 16'(4337);
			14854: out = 16'(10460);
			14855: out = 16'(-3742);
			14856: out = 16'(-18086);
			14857: out = 16'(-8313);
			14858: out = 16'(4101);
			14859: out = 16'(11110);
			14860: out = 16'(5646);
			14861: out = 16'(-782);
			14862: out = 16'(-9126);
			14863: out = 16'(-3305);
			14864: out = 16'(968);
			14865: out = 16'(1434);
			14866: out = 16'(5190);
			14867: out = 16'(7595);
			14868: out = 16'(2365);
			14869: out = 16'(-7477);
			14870: out = 16'(-7154);
			14871: out = 16'(-2893);
			14872: out = 16'(4582);
			14873: out = 16'(4796);
			14874: out = 16'(-1601);
			14875: out = 16'(-3066);
			14876: out = 16'(170);
			14877: out = 16'(2036);
			14878: out = 16'(-617);
			14879: out = 16'(-3552);
			14880: out = 16'(-535);
			14881: out = 16'(3376);
			14882: out = 16'(550);
			14883: out = 16'(-6587);
			14884: out = 16'(-5048);
			14885: out = 16'(4291);
			14886: out = 16'(7147);
			14887: out = 16'(328);
			14888: out = 16'(-8965);
			14889: out = 16'(-5776);
			14890: out = 16'(3926);
			14891: out = 16'(7143);
			14892: out = 16'(-1455);
			14893: out = 16'(-4550);
			14894: out = 16'(-218);
			14895: out = 16'(4325);
			14896: out = 16'(-1824);
			14897: out = 16'(-716);
			14898: out = 16'(1586);
			14899: out = 16'(-1043);
			14900: out = 16'(-6906);
			14901: out = 16'(-3439);
			14902: out = 16'(2258);
			14903: out = 16'(1646);
			14904: out = 16'(868);
			14905: out = 16'(-528);
			14906: out = 16'(1401);
			14907: out = 16'(-259);
			14908: out = 16'(-4511);
			14909: out = 16'(-5882);
			14910: out = 16'(-59);
			14911: out = 16'(4499);
			14912: out = 16'(4411);
			14913: out = 16'(-4850);
			14914: out = 16'(-3600);
			14915: out = 16'(4048);
			14916: out = 16'(10405);
			14917: out = 16'(-1879);
			14918: out = 16'(-3232);
			14919: out = 16'(-5792);
			14920: out = 16'(-6376);
			14921: out = 16'(-1141);
			14922: out = 16'(11202);
			14923: out = 16'(8429);
			14924: out = 16'(-1584);
			14925: out = 16'(-2434);
			14926: out = 16'(2680);
			14927: out = 16'(-2118);
			14928: out = 16'(-9140);
			14929: out = 16'(-1510);
			14930: out = 16'(6240);
			14931: out = 16'(3713);
			14932: out = 16'(-2615);
			14933: out = 16'(741);
			14934: out = 16'(351);
			14935: out = 16'(1398);
			14936: out = 16'(2827);
			14937: out = 16'(6538);
			14938: out = 16'(-149);
			14939: out = 16'(-3875);
			14940: out = 16'(-3522);
			14941: out = 16'(2768);
			14942: out = 16'(3740);
			14943: out = 16'(6636);
			14944: out = 16'(5229);
			14945: out = 16'(3871);
			14946: out = 16'(1549);
			14947: out = 16'(320);
			14948: out = 16'(-4397);
			14949: out = 16'(-6473);
			14950: out = 16'(-2450);
			14951: out = 16'(-1030);
			14952: out = 16'(722);
			14953: out = 16'(942);
			14954: out = 16'(951);
			14955: out = 16'(-442);
			14956: out = 16'(-195);
			14957: out = 16'(-268);
			14958: out = 16'(37);
			14959: out = 16'(800);
			14960: out = 16'(353);
			14961: out = 16'(-691);
			14962: out = 16'(1431);
			14963: out = 16'(7116);
			14964: out = 16'(7015);
			14965: out = 16'(1462);
			14966: out = 16'(-5194);
			14967: out = 16'(-8353);
			14968: out = 16'(-9158);
			14969: out = 16'(-11182);
			14970: out = 16'(-9156);
			14971: out = 16'(2097);
			14972: out = 16'(8094);
			14973: out = 16'(11020);
			14974: out = 16'(4821);
			14975: out = 16'(-4705);
			14976: out = 16'(-16937);
			14977: out = 16'(-8256);
			14978: out = 16'(1632);
			14979: out = 16'(1033);
			14980: out = 16'(-4005);
			14981: out = 16'(-1939);
			14982: out = 16'(6489);
			14983: out = 16'(9976);
			14984: out = 16'(2867);
			14985: out = 16'(-2192);
			14986: out = 16'(-5600);
			14987: out = 16'(-2324);
			14988: out = 16'(4464);
			14989: out = 16'(-5034);
			14990: out = 16'(-5212);
			14991: out = 16'(2375);
			14992: out = 16'(9338);
			14993: out = 16'(-1928);
			14994: out = 16'(-3089);
			14995: out = 16'(-589);
			14996: out = 16'(2790);
			14997: out = 16'(-647);
			14998: out = 16'(-1260);
			14999: out = 16'(-5837);
			15000: out = 16'(-5089);
			15001: out = 16'(6247);
			15002: out = 16'(16575);
			15003: out = 16'(11449);
			15004: out = 16'(-1593);
			15005: out = 16'(-7403);
			15006: out = 16'(-7801);
			15007: out = 16'(-3822);
			15008: out = 16'(-1471);
			15009: out = 16'(4148);
			15010: out = 16'(9041);
			15011: out = 16'(10942);
			15012: out = 16'(-339);
			15013: out = 16'(-14749);
			15014: out = 16'(-12042);
			15015: out = 16'(-7078);
			15016: out = 16'(-3683);
			15017: out = 16'(-415);
			15018: out = 16'(7073);
			15019: out = 16'(12705);
			15020: out = 16'(9400);
			15021: out = 16'(2224);
			15022: out = 16'(-464);
			15023: out = 16'(-5832);
			15024: out = 16'(-8009);
			15025: out = 16'(-5618);
			15026: out = 16'(456);
			15027: out = 16'(-2288);
			15028: out = 16'(97);
			15029: out = 16'(6686);
			15030: out = 16'(10503);
			15031: out = 16'(271);
			15032: out = 16'(-8782);
			15033: out = 16'(-11662);
			15034: out = 16'(-4785);
			15035: out = 16'(4231);
			15036: out = 16'(2799);
			15037: out = 16'(-10);
			15038: out = 16'(2539);
			15039: out = 16'(9532);
			15040: out = 16'(1713);
			15041: out = 16'(-3451);
			15042: out = 16'(-5665);
			15043: out = 16'(-5349);
			15044: out = 16'(-11248);
			15045: out = 16'(-8107);
			15046: out = 16'(-1435);
			15047: out = 16'(2811);
			15048: out = 16'(-2050);
			15049: out = 16'(3391);
			15050: out = 16'(8335);
			15051: out = 16'(6570);
			15052: out = 16'(-8598);
			15053: out = 16'(-2232);
			15054: out = 16'(-207);
			15055: out = 16'(-2921);
			15056: out = 16'(-1336);
			15057: out = 16'(10872);
			15058: out = 16'(11895);
			15059: out = 16'(1518);
			15060: out = 16'(-6922);
			15061: out = 16'(-1546);
			15062: out = 16'(2092);
			15063: out = 16'(-1306);
			15064: out = 16'(-2871);
			15065: out = 16'(-1157);
			15066: out = 16'(7123);
			15067: out = 16'(6101);
			15068: out = 16'(353);
			15069: out = 16'(-2647);
			15070: out = 16'(7576);
			15071: out = 16'(7974);
			15072: out = 16'(-1040);
			15073: out = 16'(-7433);
			15074: out = 16'(-2114);
			15075: out = 16'(649);
			15076: out = 16'(515);
			15077: out = 16'(5105);
			15078: out = 16'(5907);
			15079: out = 16'(3137);
			15080: out = 16'(-4721);
			15081: out = 16'(-10687);
			15082: out = 16'(-8483);
			15083: out = 16'(-3068);
			15084: out = 16'(3614);
			15085: out = 16'(7505);
			15086: out = 16'(2375);
			15087: out = 16'(435);
			15088: out = 16'(679);
			15089: out = 16'(1863);
			15090: out = 16'(-3254);
			15091: out = 16'(-2377);
			15092: out = 16'(-5610);
			15093: out = 16'(-6744);
			15094: out = 16'(791);
			15095: out = 16'(5353);
			15096: out = 16'(7192);
			15097: out = 16'(2607);
			15098: out = 16'(-3304);
			15099: out = 16'(-12608);
			15100: out = 16'(-5809);
			15101: out = 16'(5153);
			15102: out = 16'(11487);
			15103: out = 16'(12794);
			15104: out = 16'(5620);
			15105: out = 16'(-8821);
			15106: out = 16'(-19017);
			15107: out = 16'(-7734);
			15108: out = 16'(4373);
			15109: out = 16'(8112);
			15110: out = 16'(475);
			15111: out = 16'(-11200);
			15112: out = 16'(-5829);
			15113: out = 16'(412);
			15114: out = 16'(4527);
			15115: out = 16'(9496);
			15116: out = 16'(11895);
			15117: out = 16'(5828);
			15118: out = 16'(-6567);
			15119: out = 16'(-14235);
			15120: out = 16'(-9058);
			15121: out = 16'(2047);
			15122: out = 16'(7517);
			15123: out = 16'(7379);
			15124: out = 16'(4264);
			15125: out = 16'(-1878);
			15126: out = 16'(-11502);
			15127: out = 16'(-13857);
			15128: out = 16'(180);
			15129: out = 16'(3437);
			15130: out = 16'(3096);
			15131: out = 16'(3660);
			15132: out = 16'(6624);
			15133: out = 16'(3406);
			15134: out = 16'(-2417);
			15135: out = 16'(-5216);
			15136: out = 16'(-4264);
			15137: out = 16'(-10622);
			15138: out = 16'(-7142);
			15139: out = 16'(6028);
			15140: out = 16'(12569);
			15141: out = 16'(-4661);
			15142: out = 16'(-10701);
			15143: out = 16'(-547);
			15144: out = 16'(10993);
			15145: out = 16'(-1725);
			15146: out = 16'(746);
			15147: out = 16'(5137);
			15148: out = 16'(8837);
			15149: out = 16'(3643);
			15150: out = 16'(-3189);
			15151: out = 16'(-2455);
			15152: out = 16'(7022);
			15153: out = 16'(10829);
			15154: out = 16'(-389);
			15155: out = 16'(-9961);
			15156: out = 16'(-9339);
			15157: out = 16'(-1978);
			15158: out = 16'(-3921);
			15159: out = 16'(-1122);
			15160: out = 16'(3651);
			15161: out = 16'(7465);
			15162: out = 16'(-1802);
			15163: out = 16'(5257);
			15164: out = 16'(5517);
			15165: out = 16'(1735);
			15166: out = 16'(-4145);
			15167: out = 16'(5179);
			15168: out = 16'(938);
			15169: out = 16'(-7811);
			15170: out = 16'(-6532);
			15171: out = 16'(4265);
			15172: out = 16'(5592);
			15173: out = 16'(-2237);
			15174: out = 16'(-7389);
			15175: out = 16'(-3674);
			15176: out = 16'(-271);
			15177: out = 16'(-1471);
			15178: out = 16'(-1443);
			15179: out = 16'(4264);
			15180: out = 16'(9645);
			15181: out = 16'(7375);
			15182: out = 16'(-542);
			15183: out = 16'(-6085);
			15184: out = 16'(-3466);
			15185: out = 16'(2416);
			15186: out = 16'(3597);
			15187: out = 16'(-186);
			15188: out = 16'(1679);
			15189: out = 16'(4319);
			15190: out = 16'(4066);
			15191: out = 16'(-1830);
			15192: out = 16'(-5778);
			15193: out = 16'(-5537);
			15194: out = 16'(1564);
			15195: out = 16'(6686);
			15196: out = 16'(7759);
			15197: out = 16'(-436);
			15198: out = 16'(-2869);
			15199: out = 16'(386);
			15200: out = 16'(3015);
			15201: out = 16'(-900);
			15202: out = 16'(-1373);
			15203: out = 16'(-298);
			15204: out = 16'(-907);
			15205: out = 16'(-10532);
			15206: out = 16'(-8230);
			15207: out = 16'(1428);
			15208: out = 16'(7928);
			15209: out = 16'(9185);
			15210: out = 16'(5451);
			15211: out = 16'(-3407);
			15212: out = 16'(-10481);
			15213: out = 16'(-5083);
			15214: out = 16'(1896);
			15215: out = 16'(1044);
			15216: out = 16'(-2851);
			15217: out = 16'(-328);
			15218: out = 16'(465);
			15219: out = 16'(-5605);
			15220: out = 16'(-9428);
			15221: out = 16'(-866);
			15222: out = 16'(8410);
			15223: out = 16'(2740);
			15224: out = 16'(-8535);
			15225: out = 16'(-8867);
			15226: out = 16'(417);
			15227: out = 16'(3750);
			15228: out = 16'(2614);
			15229: out = 16'(5294);
			15230: out = 16'(2076);
			15231: out = 16'(365);
			15232: out = 16'(-2318);
			15233: out = 16'(-535);
			15234: out = 16'(-866);
			15235: out = 16'(815);
			15236: out = 16'(-807);
			15237: out = 16'(2810);
			15238: out = 16'(9673);
			15239: out = 16'(3295);
			15240: out = 16'(-8524);
			15241: out = 16'(-11422);
			15242: out = 16'(-2405);
			15243: out = 16'(117);
			15244: out = 16'(-860);
			15245: out = 16'(5738);
			15246: out = 16'(15252);
			15247: out = 16'(7904);
			15248: out = 16'(-8922);
			15249: out = 16'(-14622);
			15250: out = 16'(-1170);
			15251: out = 16'(-1268);
			15252: out = 16'(3609);
			15253: out = 16'(2829);
			15254: out = 16'(1268);
			15255: out = 16'(-6859);
			15256: out = 16'(-5163);
			15257: out = 16'(-3299);
			15258: out = 16'(4108);
			15259: out = 16'(13621);
			15260: out = 16'(14476);
			15261: out = 16'(6239);
			15262: out = 16'(-5911);
			15263: out = 16'(-13451);
			15264: out = 16'(-12919);
			15265: out = 16'(-4276);
			15266: out = 16'(2907);
			15267: out = 16'(3787);
			15268: out = 16'(-4420);
			15269: out = 16'(1980);
			15270: out = 16'(8717);
			15271: out = 16'(5212);
			15272: out = 16'(-10957);
			15273: out = 16'(-6062);
			15274: out = 16'(3925);
			15275: out = 16'(6688);
			15276: out = 16'(-83);
			15277: out = 16'(707);
			15278: out = 16'(3588);
			15279: out = 16'(5362);
			15280: out = 16'(1698);
			15281: out = 16'(5687);
			15282: out = 16'(272);
			15283: out = 16'(-4988);
			15284: out = 16'(-6290);
			15285: out = 16'(-482);
			15286: out = 16'(-66);
			15287: out = 16'(-24);
			15288: out = 16'(-906);
			15289: out = 16'(-2340);
			15290: out = 16'(442);
			15291: out = 16'(5363);
			15292: out = 16'(4955);
			15293: out = 16'(100);
			15294: out = 16'(-583);
			15295: out = 16'(6846);
			15296: out = 16'(8333);
			15297: out = 16'(46);
			15298: out = 16'(-8589);
			15299: out = 16'(-1776);
			15300: out = 16'(4552);
			15301: out = 16'(-2419);
			15302: out = 16'(-6928);
			15303: out = 16'(-2485);
			15304: out = 16'(4925);
			15305: out = 16'(2606);
			15306: out = 16'(678);
			15307: out = 16'(-7182);
			15308: out = 16'(-4487);
			15309: out = 16'(1844);
			15310: out = 16'(1802);
			15311: out = 16'(-4389);
			15312: out = 16'(-7281);
			15313: out = 16'(-1705);
			15314: out = 16'(6540);
			15315: out = 16'(3401);
			15316: out = 16'(-1200);
			15317: out = 16'(-1515);
			15318: out = 16'(2301);
			15319: out = 16'(-1075);
			15320: out = 16'(-6593);
			15321: out = 16'(-7072);
			15322: out = 16'(2428);
			15323: out = 16'(4272);
			15324: out = 16'(6542);
			15325: out = 16'(-1624);
			15326: out = 16'(-7524);
			15327: out = 16'(-4304);
			15328: out = 16'(2865);
			15329: out = 16'(-40);
			15330: out = 16'(-2891);
			15331: out = 16'(2616);
			15332: out = 16'(6868);
			15333: out = 16'(-2446);
			15334: out = 16'(-11442);
			15335: out = 16'(-4940);
			15336: out = 16'(-2343);
			15337: out = 16'(1576);
			15338: out = 16'(6165);
			15339: out = 16'(12793);
			15340: out = 16'(3409);
			15341: out = 16'(2094);
			15342: out = 16'(220);
			15343: out = 16'(-959);
			15344: out = 16'(-7945);
			15345: out = 16'(-414);
			15346: out = 16'(6228);
			15347: out = 16'(7708);
			15348: out = 16'(1367);
			15349: out = 16'(-8610);
			15350: out = 16'(-13977);
			15351: out = 16'(-6575);
			15352: out = 16'(4774);
			15353: out = 16'(3531);
			15354: out = 16'(296);
			15355: out = 16'(3365);
			15356: out = 16'(8839);
			15357: out = 16'(9075);
			15358: out = 16'(560);
			15359: out = 16'(-1694);
			15360: out = 16'(2297);
			15361: out = 16'(-2810);
			15362: out = 16'(-7682);
			15363: out = 16'(-4093);
			15364: out = 16'(7463);
			15365: out = 16'(7129);
			15366: out = 16'(6511);
			15367: out = 16'(-1671);
			15368: out = 16'(-6234);
			15369: out = 16'(-8372);
			15370: out = 16'(-2987);
			15371: out = 16'(-3983);
			15372: out = 16'(-535);
			15373: out = 16'(7084);
			15374: out = 16'(6897);
			15375: out = 16'(308);
			15376: out = 16'(-1963);
			15377: out = 16'(2615);
			15378: out = 16'(-1891);
			15379: out = 16'(-916);
			15380: out = 16'(2353);
			15381: out = 16'(7000);
			15382: out = 16'(3396);
			15383: out = 16'(-1500);
			15384: out = 16'(-8018);
			15385: out = 16'(-8484);
			15386: out = 16'(-6452);
			15387: out = 16'(8331);
			15388: out = 16'(8636);
			15389: out = 16'(2501);
			15390: out = 16'(-2812);
			15391: out = 16'(3766);
			15392: out = 16'(186);
			15393: out = 16'(-4679);
			15394: out = 16'(-4350);
			15395: out = 16'(3795);
			15396: out = 16'(3056);
			15397: out = 16'(1466);
			15398: out = 16'(-406);
			15399: out = 16'(-5005);
			15400: out = 16'(-6241);
			15401: out = 16'(20);
			15402: out = 16'(5531);
			15403: out = 16'(624);
			15404: out = 16'(-2245);
			15405: out = 16'(1493);
			15406: out = 16'(8355);
			15407: out = 16'(6628);
			15408: out = 16'(-5167);
			15409: out = 16'(-10367);
			15410: out = 16'(-3002);
			15411: out = 16'(5103);
			15412: out = 16'(439);
			15413: out = 16'(-6063);
			15414: out = 16'(-5979);
			15415: out = 16'(1004);
			15416: out = 16'(1621);
			15417: out = 16'(1143);
			15418: out = 16'(-2312);
			15419: out = 16'(-1087);
			15420: out = 16'(3795);
			15421: out = 16'(-49);
			15422: out = 16'(-9976);
			15423: out = 16'(-12150);
			15424: out = 16'(951);
			15425: out = 16'(4157);
			15426: out = 16'(4613);
			15427: out = 16'(7250);
			15428: out = 16'(12757);
			15429: out = 16'(1256);
			15430: out = 16'(-8098);
			15431: out = 16'(-11290);
			15432: out = 16'(-3565);
			15433: out = 16'(-3793);
			15434: out = 16'(4989);
			15435: out = 16'(4935);
			15436: out = 16'(201);
			15437: out = 16'(-1105);
			15438: out = 16'(4404);
			15439: out = 16'(6636);
			15440: out = 16'(560);
			15441: out = 16'(-9996);
			15442: out = 16'(-5807);
			15443: out = 16'(490);
			15444: out = 16'(946);
			15445: out = 16'(-3428);
			15446: out = 16'(5451);
			15447: out = 16'(4834);
			15448: out = 16'(-1425);
			15449: out = 16'(-6345);
			15450: out = 16'(-5550);
			15451: out = 16'(3169);
			15452: out = 16'(7769);
			15453: out = 16'(4168);
			15454: out = 16'(-7141);
			15455: out = 16'(-3638);
			15456: out = 16'(1099);
			15457: out = 16'(2135);
			15458: out = 16'(1157);
			15459: out = 16'(2133);
			15460: out = 16'(518);
			15461: out = 16'(-2609);
			15462: out = 16'(-3914);
			15463: out = 16'(-6130);
			15464: out = 16'(-2984);
			15465: out = 16'(3782);
			15466: out = 16'(8232);
			15467: out = 16'(5017);
			15468: out = 16'(-2837);
			15469: out = 16'(-7958);
			15470: out = 16'(-6987);
			15471: out = 16'(-5075);
			15472: out = 16'(331);
			15473: out = 16'(8032);
			15474: out = 16'(13166);
			15475: out = 16'(6616);
			15476: out = 16'(3741);
			15477: out = 16'(-1111);
			15478: out = 16'(-4726);
			15479: out = 16'(-12705);
			15480: out = 16'(-10941);
			15481: out = 16'(-8706);
			15482: out = 16'(4567);
			15483: out = 16'(15540);
			15484: out = 16'(9517);
			15485: out = 16'(-6895);
			15486: out = 16'(-9935);
			15487: out = 16'(2010);
			15488: out = 16'(1878);
			15489: out = 16'(-2582);
			15490: out = 16'(-3303);
			15491: out = 16'(3281);
			15492: out = 16'(5078);
			15493: out = 16'(3387);
			15494: out = 16'(2519);
			15495: out = 16'(2726);
			15496: out = 16'(-1901);
			15497: out = 16'(-2516);
			15498: out = 16'(111);
			15499: out = 16'(1066);
			15500: out = 16'(-5675);
			15501: out = 16'(118);
			15502: out = 16'(444);
			15503: out = 16'(1096);
			15504: out = 16'(-417);
			15505: out = 16'(533);
			15506: out = 16'(-2248);
			15507: out = 16'(-1127);
			15508: out = 16'(1061);
			15509: out = 16'(84);
			15510: out = 16'(-3871);
			15511: out = 16'(-3452);
			15512: out = 16'(2153);
			15513: out = 16'(6258);
			15514: out = 16'(4362);
			15515: out = 16'(1094);
			15516: out = 16'(-697);
			15517: out = 16'(-3341);
			15518: out = 16'(-6750);
			15519: out = 16'(-7024);
			15520: out = 16'(-1341);
			15521: out = 16'(4013);
			15522: out = 16'(6939);
			15523: out = 16'(4794);
			15524: out = 16'(4915);
			15525: out = 16'(3004);
			15526: out = 16'(496);
			15527: out = 16'(-18831);
			15528: out = 16'(-20447);
			15529: out = 16'(-2035);
			15530: out = 16'(9811);
			15531: out = 16'(6966);
			15532: out = 16'(3573);
			15533: out = 16'(6206);
			15534: out = 16'(5446);
			15535: out = 16'(-199);
			15536: out = 16'(-9020);
			15537: out = 16'(-8756);
			15538: out = 16'(722);
			15539: out = 16'(9577);
			15540: out = 16'(9356);
			15541: out = 16'(4661);
			15542: out = 16'(206);
			15543: out = 16'(-1247);
			15544: out = 16'(1003);
			15545: out = 16'(2890);
			15546: out = 16'(721);
			15547: out = 16'(-3556);
			15548: out = 16'(-5487);
			15549: out = 16'(-2271);
			15550: out = 16'(273);
			15551: out = 16'(301);
			15552: out = 16'(-640);
			15553: out = 16'(6154);
			15554: out = 16'(9761);
			15555: out = 16'(2220);
			15556: out = 16'(-8188);
			15557: out = 16'(-8081);
			15558: out = 16'(766);
			15559: out = 16'(3153);
			15560: out = 16'(-1374);
			15561: out = 16'(-5786);
			15562: out = 16'(798);
			15563: out = 16'(7340);
			15564: out = 16'(1100);
			15565: out = 16'(-2107);
			15566: out = 16'(53);
			15567: out = 16'(3333);
			15568: out = 16'(-919);
			15569: out = 16'(-11357);
			15570: out = 16'(-11566);
			15571: out = 16'(2490);
			15572: out = 16'(13525);
			15573: out = 16'(9027);
			15574: out = 16'(605);
			15575: out = 16'(-3913);
			15576: out = 16'(-5486);
			15577: out = 16'(-4502);
			15578: out = 16'(-7476);
			15579: out = 16'(-2044);
			15580: out = 16'(8954);
			15581: out = 16'(11484);
			15582: out = 16'(5351);
			15583: out = 16'(-1156);
			15584: out = 16'(-3028);
			15585: out = 16'(-5495);
			15586: out = 16'(-2892);
			15587: out = 16'(-1565);
			15588: out = 16'(938);
			15589: out = 16'(2612);
			15590: out = 16'(12100);
			15591: out = 16'(7112);
			15592: out = 16'(-1595);
			15593: out = 16'(-4263);
			15594: out = 16'(5046);
			15595: out = 16'(2837);
			15596: out = 16'(-4551);
			15597: out = 16'(-7243);
			15598: out = 16'(-3524);
			15599: out = 16'(-474);
			15600: out = 16'(-797);
			15601: out = 16'(2353);
			15602: out = 16'(10504);
			15603: out = 16'(12609);
			15604: out = 16'(1078);
			15605: out = 16'(-16332);
			15606: out = 16'(-24736);
			15607: out = 16'(-5792);
			15608: out = 16'(8814);
			15609: out = 16'(8315);
			15610: out = 16'(5215);
			15611: out = 16'(8918);
			15612: out = 16'(5486);
			15613: out = 16'(-11987);
			15614: out = 16'(-27788);
			15615: out = 16'(-12260);
			15616: out = 16'(3234);
			15617: out = 16'(6775);
			15618: out = 16'(5708);
			15619: out = 16'(11054);
			15620: out = 16'(7157);
			15621: out = 16'(-5176);
			15622: out = 16'(-14136);
			15623: out = 16'(-3905);
			15624: out = 16'(4600);
			15625: out = 16'(5564);
			15626: out = 16'(714);
			15627: out = 16'(472);
			15628: out = 16'(-426);
			15629: out = 16'(2498);
			15630: out = 16'(2940);
			15631: out = 16'(689);
			15632: out = 16'(145);
			15633: out = 16'(-2214);
			15634: out = 16'(-2562);
			15635: out = 16'(-2615);
			15636: out = 16'(253);
			15637: out = 16'(-924);
			15638: out = 16'(3494);
			15639: out = 16'(6559);
			15640: out = 16'(6650);
			15641: out = 16'(-2766);
			15642: out = 16'(-780);
			15643: out = 16'(765);
			15644: out = 16'(-5631);
			15645: out = 16'(-13823);
			15646: out = 16'(-2441);
			15647: out = 16'(8959);
			15648: out = 16'(4168);
			15649: out = 16'(4364);
			15650: out = 16'(3548);
			15651: out = 16'(3393);
			15652: out = 16'(-2777);
			15653: out = 16'(-13330);
			15654: out = 16'(-7033);
			15655: out = 16'(1473);
			15656: out = 16'(1676);
			15657: out = 16'(991);
			15658: out = 16'(6963);
			15659: out = 16'(9765);
			15660: out = 16'(1477);
			15661: out = 16'(-10036);
			15662: out = 16'(-17210);
			15663: out = 16'(-10714);
			15664: out = 16'(-1450);
			15665: out = 16'(3501);
			15666: out = 16'(8059);
			15667: out = 16'(11754);
			15668: out = 16'(9789);
			15669: out = 16'(2326);
			15670: out = 16'(-8012);
			15671: out = 16'(-10252);
			15672: out = 16'(-9797);
			15673: out = 16'(-6712);
			15674: out = 16'(1382);
			15675: out = 16'(7108);
			15676: out = 16'(4736);
			15677: out = 16'(-689);
			15678: out = 16'(595);
			15679: out = 16'(-90);
			15680: out = 16'(667);
			15681: out = 16'(-2037);
			15682: out = 16'(-7381);
			15683: out = 16'(-2733);
			15684: out = 16'(1469);
			15685: out = 16'(5155);
			15686: out = 16'(3647);
			15687: out = 16'(1553);
			15688: out = 16'(-3561);
			15689: out = 16'(1118);
			15690: out = 16'(6472);
			15691: out = 16'(3025);
			15692: out = 16'(-9585);
			15693: out = 16'(-6190);
			15694: out = 16'(8387);
			15695: out = 16'(9262);
			15696: out = 16'(4731);
			15697: out = 16'(158);
			15698: out = 16'(-670);
			15699: out = 16'(-5735);
			15700: out = 16'(-4655);
			15701: out = 16'(-1220);
			15702: out = 16'(4593);
			15703: out = 16'(3523);
			15704: out = 16'(5619);
			15705: out = 16'(-4370);
			15706: out = 16'(-5832);
			15707: out = 16'(1413);
			15708: out = 16'(5107);
			15709: out = 16'(1766);
			15710: out = 16'(-1988);
			15711: out = 16'(-2073);
			15712: out = 16'(136);
			15713: out = 16'(2640);
			15714: out = 16'(4729);
			15715: out = 16'(5882);
			15716: out = 16'(7257);
			15717: out = 16'(651);
			15718: out = 16'(-2905);
			15719: out = 16'(-8436);
			15720: out = 16'(-11949);
			15721: out = 16'(-2379);
			15722: out = 16'(11079);
			15723: out = 16'(11182);
			15724: out = 16'(380);
			15725: out = 16'(197);
			15726: out = 16'(3969);
			15727: out = 16'(4384);
			15728: out = 16'(-5649);
			15729: out = 16'(-14539);
			15730: out = 16'(-9728);
			15731: out = 16'(5426);
			15732: out = 16'(11807);
			15733: out = 16'(6759);
			15734: out = 16'(-5410);
			15735: out = 16'(-5163);
			15736: out = 16'(3033);
			15737: out = 16'(5133);
			15738: out = 16'(-3235);
			15739: out = 16'(-7568);
			15740: out = 16'(-1883);
			15741: out = 16'(5539);
			15742: out = 16'(1088);
			15743: out = 16'(-1816);
			15744: out = 16'(-2561);
			15745: out = 16'(-771);
			15746: out = 16'(1982);
			15747: out = 16'(-2851);
			15748: out = 16'(-9479);
			15749: out = 16'(-11519);
			15750: out = 16'(-137);
			15751: out = 16'(4639);
			15752: out = 16'(10266);
			15753: out = 16'(7775);
			15754: out = 16'(2098);
			15755: out = 16'(-7274);
			15756: out = 16'(-3564);
			15757: out = 16'(-3810);
			15758: out = 16'(-9690);
			15759: out = 16'(-3401);
			15760: out = 16'(9768);
			15761: out = 16'(12520);
			15762: out = 16'(4613);
			15763: out = 16'(176);
			15764: out = 16'(-1813);
			15765: out = 16'(-6903);
			15766: out = 16'(-10553);
			15767: out = 16'(-2240);
			15768: out = 16'(3045);
			15769: out = 16'(-452);
			15770: out = 16'(-3969);
			15771: out = 16'(3523);
			15772: out = 16'(7064);
			15773: out = 16'(3707);
			15774: out = 16'(-1082);
			15775: out = 16'(1050);
			15776: out = 16'(5957);
			15777: out = 16'(-1834);
			15778: out = 16'(-9847);
			15779: out = 16'(-4608);
			15780: out = 16'(6242);
			15781: out = 16'(1968);
			15782: out = 16'(-6860);
			15783: out = 16'(-3596);
			15784: out = 16'(9588);
			15785: out = 16'(8721);
			15786: out = 16'(853);
			15787: out = 16'(-1912);
			15788: out = 16'(861);
			15789: out = 16'(6442);
			15790: out = 16'(-900);
			15791: out = 16'(-6611);
			15792: out = 16'(-101);
			15793: out = 16'(7051);
			15794: out = 16'(5178);
			15795: out = 16'(145);
			15796: out = 16'(-324);
			15797: out = 16'(-3134);
			15798: out = 16'(-1038);
			15799: out = 16'(251);
			15800: out = 16'(719);
			15801: out = 16'(-2708);
			15802: out = 16'(5458);
			15803: out = 16'(8710);
			15804: out = 16'(1959);
			15805: out = 16'(-10257);
			15806: out = 16'(-17048);
			15807: out = 16'(-10425);
			15808: out = 16'(1959);
			15809: out = 16'(7589);
			15810: out = 16'(9533);
			15811: out = 16'(5349);
			15812: out = 16'(-1706);
			15813: out = 16'(-7567);
			15814: out = 16'(-2133);
			15815: out = 16'(226);
			15816: out = 16'(-3249);
			15817: out = 16'(-8540);
			15818: out = 16'(123);
			15819: out = 16'(1627);
			15820: out = 16'(3468);
			15821: out = 16'(2615);
			15822: out = 16'(259);
			15823: out = 16'(-3255);
			15824: out = 16'(-1992);
			15825: out = 16'(1147);
			15826: out = 16'(2129);
			15827: out = 16'(625);
			15828: out = 16'(-1584);
			15829: out = 16'(-2192);
			15830: out = 16'(556);
			15831: out = 16'(1662);
			15832: out = 16'(6430);
			15833: out = 16'(4017);
			15834: out = 16'(-5272);
			15835: out = 16'(-4329);
			15836: out = 16'(750);
			15837: out = 16'(8281);
			15838: out = 16'(7027);
			15839: out = 16'(367);
			15840: out = 16'(-5325);
			15841: out = 16'(-1167);
			15842: out = 16'(883);
			15843: out = 16'(-5349);
			15844: out = 16'(-14646);
			15845: out = 16'(-5757);
			15846: out = 16'(9366);
			15847: out = 16'(9674);
			15848: out = 16'(4267);
			15849: out = 16'(715);
			15850: out = 16'(4993);
			15851: out = 16'(6001);
			15852: out = 16'(783);
			15853: out = 16'(-8306);
			15854: out = 16'(-7077);
			15855: out = 16'(1705);
			15856: out = 16'(3750);
			15857: out = 16'(6209);
			15858: out = 16'(4899);
			15859: out = 16'(1942);
			15860: out = 16'(-386);
			15861: out = 16'(-4567);
			15862: out = 16'(-6886);
			15863: out = 16'(-8564);
			15864: out = 16'(-8245);
			15865: out = 16'(-4115);
			15866: out = 16'(5385);
			15867: out = 16'(9531);
			15868: out = 16'(5456);
			15869: out = 16'(2666);
			15870: out = 16'(415);
			15871: out = 16'(-3247);
			15872: out = 16'(-7701);
			15873: out = 16'(-219);
			15874: out = 16'(-256);
			15875: out = 16'(1046);
			15876: out = 16'(2659);
			15877: out = 16'(4230);
			15878: out = 16'(730);
			15879: out = 16'(-1176);
			15880: out = 16'(-2495);
			15881: out = 16'(-5593);
			15882: out = 16'(-6229);
			15883: out = 16'(-3409);
			15884: out = 16'(3370);
			15885: out = 16'(7099);
			15886: out = 16'(6215);
			15887: out = 16'(1195);
			15888: out = 16'(-63);
			15889: out = 16'(-1807);
			15890: out = 16'(-9019);
			15891: out = 16'(-19385);
			15892: out = 16'(-14023);
			15893: out = 16'(4900);
			15894: out = 16'(12220);
			15895: out = 16'(9309);
			15896: out = 16'(2860);
			15897: out = 16'(2028);
			15898: out = 16'(3541);
			15899: out = 16'(-10291);
			15900: out = 16'(-18306);
			15901: out = 16'(-11789);
			15902: out = 16'(2648);
			15903: out = 16'(10060);
			15904: out = 16'(8949);
			15905: out = 16'(4483);
			15906: out = 16'(736);
			15907: out = 16'(7);
			15908: out = 16'(714);
			15909: out = 16'(1282);
			15910: out = 16'(-1956);
			15911: out = 16'(-12101);
			15912: out = 16'(-6054);
			15913: out = 16'(3125);
			15914: out = 16'(4799);
			15915: out = 16'(862);
			15916: out = 16'(5056);
			15917: out = 16'(7722);
			15918: out = 16'(978);
			15919: out = 16'(-7980);
			15920: out = 16'(-4750);
			15921: out = 16'(9307);
			15922: out = 16'(10537);
			15923: out = 16'(-1779);
			15924: out = 16'(-7054);
			15925: out = 16'(-345);
			15926: out = 16'(1230);
			15927: out = 16'(-7691);
			15928: out = 16'(-2849);
			15929: out = 16'(-1668);
			15930: out = 16'(1727);
			15931: out = 16'(4262);
			15932: out = 16'(13594);
			15933: out = 16'(8992);
			15934: out = 16'(3128);
			15935: out = 16'(-7287);
			15936: out = 16'(-13704);
			15937: out = 16'(-10046);
			15938: out = 16'(1938);
			15939: out = 16'(6902);
			15940: out = 16'(4071);
			15941: out = 16'(1123);
			15942: out = 16'(3411);
			15943: out = 16'(3035);
			15944: out = 16'(-24);
			15945: out = 16'(4282);
			15946: out = 16'(5916);
			15947: out = 16'(3721);
			15948: out = 16'(-2047);
			15949: out = 16'(-2441);
			15950: out = 16'(-5485);
			15951: out = 16'(-916);
			15952: out = 16'(7647);
			15953: out = 16'(12717);
			15954: out = 16'(4289);
			15955: out = 16'(-8950);
			15956: out = 16'(-18755);
			15957: out = 16'(-16523);
			15958: out = 16'(-11886);
			15959: out = 16'(-1448);
			15960: out = 16'(5064);
			15961: out = 16'(6751);
			15962: out = 16'(4714);
			15963: out = 16'(4696);
			15964: out = 16'(3237);
			15965: out = 16'(-959);
			15966: out = 16'(-8568);
			15967: out = 16'(-10223);
			15968: out = 16'(-5140);
			15969: out = 16'(5770);
			15970: out = 16'(11281);
			15971: out = 16'(5649);
			15972: out = 16'(-9487);
			15973: out = 16'(-15608);
			15974: out = 16'(-2938);
			15975: out = 16'(3664);
			15976: out = 16'(856);
			15977: out = 16'(-4315);
			15978: out = 16'(1571);
			15979: out = 16'(7157);
			15980: out = 16'(6655);
			15981: out = 16'(-5096);
			15982: out = 16'(-10384);
			15983: out = 16'(1767);
			15984: out = 16'(9104);
			15985: out = 16'(268);
			15986: out = 16'(-10270);
			15987: out = 16'(-2273);
			15988: out = 16'(4939);
			15989: out = 16'(6870);
			15990: out = 16'(4101);
			15991: out = 16'(4955);
			15992: out = 16'(-637);
			15993: out = 16'(-2102);
			15994: out = 16'(-1644);
			15995: out = 16'(575);
			15996: out = 16'(49);
			15997: out = 16'(37);
			15998: out = 16'(2348);
			15999: out = 16'(5851);
			16000: out = 16'(2183);
			16001: out = 16'(3306);
			16002: out = 16'(2161);
			16003: out = 16'(-1865);
			16004: out = 16'(-8444);
			16005: out = 16'(-4338);
			16006: out = 16'(446);
			16007: out = 16'(695);
			16008: out = 16'(-790);
			16009: out = 16'(-1777);
			16010: out = 16'(5538);
			16011: out = 16'(9182);
			16012: out = 16'(2991);
			16013: out = 16'(-3593);
			16014: out = 16'(-4375);
			16015: out = 16'(-763);
			16016: out = 16'(61);
			16017: out = 16'(2769);
			16018: out = 16'(352);
			16019: out = 16'(-83);
			16020: out = 16'(-386);
			16021: out = 16'(209);
			16022: out = 16'(1377);
			16023: out = 16'(3324);
			16024: out = 16'(-1234);
			16025: out = 16'(-12050);
			16026: out = 16'(-1263);
			16027: out = 16'(11635);
			16028: out = 16'(12207);
			16029: out = 16'(1042);
			16030: out = 16'(-2122);
			16031: out = 16'(-1398);
			16032: out = 16'(-613);
			16033: out = 16'(-2586);
			16034: out = 16'(1947);
			16035: out = 16'(5256);
			16036: out = 16'(5005);
			16037: out = 16'(1912);
			16038: out = 16'(6383);
			16039: out = 16'(1155);
			16040: out = 16'(-4454);
			16041: out = 16'(-7869);
			16042: out = 16'(-2414);
			16043: out = 16'(-5196);
			16044: out = 16'(-2516);
			16045: out = 16'(1549);
			16046: out = 16'(4442);
			16047: out = 16'(3382);
			16048: out = 16'(2614);
			16049: out = 16'(1232);
			16050: out = 16'(-950);
			16051: out = 16'(-7186);
			16052: out = 16'(-8201);
			16053: out = 16'(-5899);
			16054: out = 16'(-1545);
			16055: out = 16'(-309);
			16056: out = 16'(2444);
			16057: out = 16'(501);
			16058: out = 16'(620);
			16059: out = 16'(10098);
			16060: out = 16'(2823);
			16061: out = 16'(-7523);
			16062: out = 16'(-11393);
			16063: out = 16'(1155);
			16064: out = 16'(4976);
			16065: out = 16'(8198);
			16066: out = 16'(4719);
			16067: out = 16'(-924);
			16068: out = 16'(-5084);
			16069: out = 16'(-5105);
			16070: out = 16'(-6640);
			16071: out = 16'(-8245);
			16072: out = 16'(-2807);
			16073: out = 16'(4372);
			16074: out = 16'(6889);
			16075: out = 16'(3158);
			16076: out = 16'(661);
			16077: out = 16'(-2415);
			16078: out = 16'(-1315);
			16079: out = 16'(30);
			16080: out = 16'(289);
			16081: out = 16'(-281);
			16082: out = 16'(1411);
			16083: out = 16'(2536);
			16084: out = 16'(2106);
			16085: out = 16'(-2125);
			16086: out = 16'(754);
			16087: out = 16'(5396);
			16088: out = 16'(5049);
			16089: out = 16'(-5281);
			16090: out = 16'(-8798);
			16091: out = 16'(-5650);
			16092: out = 16'(1747);
			16093: out = 16'(3944);
			16094: out = 16'(8345);
			16095: out = 16'(5413);
			16096: out = 16'(2208);
			16097: out = 16'(4074);
			16098: out = 16'(901);
			16099: out = 16'(-5200);
			16100: out = 16'(-5349);
			16101: out = 16'(4837);
			16102: out = 16'(48);
			16103: out = 16'(-1529);
			16104: out = 16'(758);
			16105: out = 16'(6776);
			16106: out = 16'(2875);
			16107: out = 16'(2577);
			16108: out = 16'(-25);
			16109: out = 16'(-4495);
			16110: out = 16'(-12440);
			16111: out = 16'(138);
			16112: out = 16'(10977);
			16113: out = 16'(6430);
			16114: out = 16'(-6855);
			16115: out = 16'(-9432);
			16116: out = 16'(-460);
			16117: out = 16'(2270);
			16118: out = 16'(-6255);
			16119: out = 16'(-5148);
			16120: out = 16'(7891);
			16121: out = 16'(13650);
			16122: out = 16'(2824);
			16123: out = 16'(-2590);
			16124: out = 16'(-1198);
			16125: out = 16'(2114);
			16126: out = 16'(-3620);
			16127: out = 16'(-3935);
			16128: out = 16'(-6628);
			16129: out = 16'(-371);
			16130: out = 16'(4915);
			16131: out = 16'(8238);
			16132: out = 16'(-3735);
			16133: out = 16'(-4689);
			16134: out = 16'(1543);
			16135: out = 16'(3209);
			16136: out = 16'(-7249);
			16137: out = 16'(-13212);
			16138: out = 16'(-9137);
			16139: out = 16'(1178);
			16140: out = 16'(3790);
			16141: out = 16'(4541);
			16142: out = 16'(1631);
			16143: out = 16'(700);
			16144: out = 16'(1415);
			16145: out = 16'(4946);
			16146: out = 16'(-2250);
			16147: out = 16'(-11088);
			16148: out = 16'(-1337);
			16149: out = 16'(2063);
			16150: out = 16'(-1947);
			16151: out = 16'(-6864);
			16152: out = 16'(1951);
			16153: out = 16'(2067);
			16154: out = 16'(-204);
			16155: out = 16'(-3710);
			16156: out = 16'(1717);
			16157: out = 16'(3062);
			16158: out = 16'(7654);
			16159: out = 16'(4216);
			16160: out = 16'(-1602);
			16161: out = 16'(-2891);
			16162: out = 16'(2501);
			16163: out = 16'(3530);
			16164: out = 16'(-63);
			16165: out = 16'(-2475);
			16166: out = 16'(-2587);
			16167: out = 16'(-2413);
			16168: out = 16'(532);
			16169: out = 16'(6147);
			16170: out = 16'(8459);
			16171: out = 16'(3862);
			16172: out = 16'(1192);
			16173: out = 16'(4836);
			16174: out = 16'(-1331);
			16175: out = 16'(-10343);
			16176: out = 16'(-11489);
			16177: out = 16'(2463);
			16178: out = 16'(8412);
			16179: out = 16'(6196);
			16180: out = 16'(-2003);
			16181: out = 16'(-2400);
			16182: out = 16'(712);
			16183: out = 16'(6547);
			16184: out = 16'(-342);
			16185: out = 16'(-7574);
			16186: out = 16'(-240);
			16187: out = 16'(8020);
			16188: out = 16'(5583);
			16189: out = 16'(-3479);
			16190: out = 16'(-4063);
			16191: out = 16'(2520);
			16192: out = 16'(7727);
			16193: out = 16'(3400);
			16194: out = 16'(-3228);
			16195: out = 16'(-6896);
			16196: out = 16'(-977);
			16197: out = 16'(1174);
			16198: out = 16'(-4856);
			16199: out = 16'(-14528);
			16200: out = 16'(-3187);
			16201: out = 16'(11338);
			16202: out = 16'(9418);
			16203: out = 16'(-6413);
			16204: out = 16'(-9436);
			16205: out = 16'(515);
			16206: out = 16'(6670);
			16207: out = 16'(-965);
			16208: out = 16'(-6496);
			16209: out = 16'(-3715);
			16210: out = 16'(2586);
			16211: out = 16'(1340);
			16212: out = 16'(-408);
			16213: out = 16'(-2864);
			16214: out = 16'(-1398);
			16215: out = 16'(111);
			16216: out = 16'(1331);
			16217: out = 16'(2308);
			16218: out = 16'(4267);
			16219: out = 16'(2896);
			16220: out = 16'(-2205);
			16221: out = 16'(-8756);
			16222: out = 16'(-6867);
			16223: out = 16'(694);
			16224: out = 16'(1748);
			16225: out = 16'(3834);
			16226: out = 16'(1167);
			16227: out = 16'(-299);
			16228: out = 16'(-178);
			16229: out = 16'(4060);
			16230: out = 16'(1782);
			16231: out = 16'(-557);
			16232: out = 16'(-168);
			16233: out = 16'(-139);
			16234: out = 16'(1242);
			16235: out = 16'(2470);
			16236: out = 16'(1872);
			16237: out = 16'(4458);
			16238: out = 16'(332);
			16239: out = 16'(-406);
			16240: out = 16'(-101);
			16241: out = 16'(3344);
			16242: out = 16'(-9082);
			16243: out = 16'(-8127);
			16244: out = 16'(85);
			16245: out = 16'(3892);
			16246: out = 16'(-7970);
			16247: out = 16'(-2940);
			16248: out = 16'(8405);
			16249: out = 16'(8513);
			16250: out = 16'(1352);
			16251: out = 16'(-2868);
			16252: out = 16'(-1406);
			16253: out = 16'(-464);
			16254: out = 16'(-3518);
			16255: out = 16'(-1568);
			16256: out = 16'(1138);
			16257: out = 16'(3019);
			16258: out = 16'(6058);
			16259: out = 16'(4336);
			16260: out = 16'(-3249);
			16261: out = 16'(-11642);
			16262: out = 16'(-8871);
			16263: out = 16'(-2747);
			16264: out = 16'(4898);
			16265: out = 16'(5832);
			16266: out = 16'(4300);
			16267: out = 16'(58);
			16268: out = 16'(229);
			16269: out = 16'(-1170);
			16270: out = 16'(-2932);
			16271: out = 16'(-9994);
			16272: out = 16'(-2156);
			16273: out = 16'(1694);
			16274: out = 16'(462);
			16275: out = 16'(4450);
			16276: out = 16'(8268);
			16277: out = 16'(6415);
			16278: out = 16'(-80);
			16279: out = 16'(-4926);
			16280: out = 16'(-4051);
			16281: out = 16'(-5771);
			16282: out = 16'(-5605);
			16283: out = 16'(3467);
			16284: out = 16'(7140);
			16285: out = 16'(6719);
			16286: out = 16'(1913);
			16287: out = 16'(-100);
			16288: out = 16'(-572);
			16289: out = 16'(298);
			16290: out = 16'(-1750);
			16291: out = 16'(-4106);
			16292: out = 16'(-5066);
			16293: out = 16'(-2384);
			16294: out = 16'(-638);
			16295: out = 16'(78);
			16296: out = 16'(1034);
			16297: out = 16'(5404);
			16298: out = 16'(4358);
			16299: out = 16'(-1237);
			16300: out = 16'(-3169);
			16301: out = 16'(-3451);
			16302: out = 16'(797);
			16303: out = 16'(2277);
			16304: out = 16'(2415);
			16305: out = 16'(-345);
			16306: out = 16'(3214);
			16307: out = 16'(2130);
			16308: out = 16'(-4078);
			16309: out = 16'(-12183);
			16310: out = 16'(-6050);
			16311: out = 16'(-420);
			16312: out = 16'(-14);
			16313: out = 16'(443);
			16314: out = 16'(8792);
			16315: out = 16'(7398);
			16316: out = 16'(-5003);
			16317: out = 16'(-15637);
			16318: out = 16'(-10417);
			16319: out = 16'(713);
			16320: out = 16'(5045);
			16321: out = 16'(3998);
			16322: out = 16'(7883);
			16323: out = 16'(7839);
			16324: out = 16'(4646);
			16325: out = 16'(2037);
			16326: out = 16'(-282);
			16327: out = 16'(-2480);
			16328: out = 16'(-4207);
			16329: out = 16'(-944);
			16330: out = 16'(3375);
			16331: out = 16'(3927);
			16332: out = 16'(-3172);
			16333: out = 16'(-6303);
			16334: out = 16'(616);
			16335: out = 16'(3728);
			16336: out = 16'(-2468);
			16337: out = 16'(-7460);
			16338: out = 16'(-3001);
			16339: out = 16'(3729);
			16340: out = 16'(1938);
			16341: out = 16'(2691);
			16342: out = 16'(11174);
			16343: out = 16'(12234);
			16344: out = 16'(8);
			16345: out = 16'(-11585);
			16346: out = 16'(-7139);
			16347: out = 16'(2537);
			16348: out = 16'(7143);
			16349: out = 16'(2993);
			16350: out = 16'(2303);
			16351: out = 16'(7288);
			16352: out = 16'(5609);
			16353: out = 16'(-3212);
			16354: out = 16'(-9983);
			16355: out = 16'(-7348);
			16356: out = 16'(-1767);
			16357: out = 16'(-1157);
			16358: out = 16'(-2757);
			16359: out = 16'(1084);
			16360: out = 16'(4073);
			16361: out = 16'(7360);
			16362: out = 16'(4895);
			16363: out = 16'(1286);
			16364: out = 16'(-3140);
			16365: out = 16'(-204);
			16366: out = 16'(-2639);
			16367: out = 16'(-9531);
			16368: out = 16'(-12250);
			16369: out = 16'(1043);
			16370: out = 16'(12713);
			16371: out = 16'(12255);
			16372: out = 16'(3284);
			16373: out = 16'(-5755);
			16374: out = 16'(-11517);
			16375: out = 16'(-13607);
			16376: out = 16'(-13436);
			16377: out = 16'(-1705);
			16378: out = 16'(3520);
			16379: out = 16'(5079);
			16380: out = 16'(3518);
			16381: out = 16'(-2631);
			16382: out = 16'(-7634);
			16383: out = 16'(-5236);
			16384: out = 16'(1386);
			16385: out = 16'(3);
			16386: out = 16'(712);
			16387: out = 16'(1075);
			16388: out = 16'(3936);
			16389: out = 16'(6272);
			16390: out = 16'(3624);
			16391: out = 16'(-648);
			16392: out = 16'(-2412);
			16393: out = 16'(-1455);
			16394: out = 16'(-6541);
			16395: out = 16'(-3729);
			16396: out = 16'(3547);
			16397: out = 16'(5685);
			16398: out = 16'(-25);
			16399: out = 16'(-1587);
			16400: out = 16'(3099);
			16401: out = 16'(4446);
			16402: out = 16'(964);
			16403: out = 16'(-6414);
			16404: out = 16'(-3615);
			16405: out = 16'(959);
			16406: out = 16'(-2066);
			16407: out = 16'(-1412);
			16408: out = 16'(8133);
			16409: out = 16'(12461);
			16410: out = 16'(2929);
			16411: out = 16'(-7931);
			16412: out = 16'(-5458);
			16413: out = 16'(2457);
			16414: out = 16'(639);
			16415: out = 16'(-8272);
			16416: out = 16'(-4156);
			16417: out = 16'(6726);
			16418: out = 16'(8649);
			16419: out = 16'(920);
			16420: out = 16'(2218);
			16421: out = 16'(5576);
			16422: out = 16'(790);
			16423: out = 16'(-10628);
			16424: out = 16'(-10719);
			16425: out = 16'(-1314);
			16426: out = 16'(5358);
			16427: out = 16'(4222);
			16428: out = 16'(2512);
			16429: out = 16'(3579);
			16430: out = 16'(2404);
			16431: out = 16'(-4630);
			16432: out = 16'(-5593);
			16433: out = 16'(-2325);
			16434: out = 16'(5580);
			16435: out = 16'(9747);
			16436: out = 16'(6655);
			16437: out = 16'(1249);
			16438: out = 16'(-406);
			16439: out = 16'(1034);
			16440: out = 16'(-579);
			16441: out = 16'(-3696);
			16442: out = 16'(-6110);
			16443: out = 16'(-2738);
			16444: out = 16'(3666);
			16445: out = 16'(-6820);
			16446: out = 16'(-10323);
			16447: out = 16'(902);
			16448: out = 16'(12859);
			16449: out = 16'(6451);
			16450: out = 16'(-7815);
			16451: out = 16'(-13161);
			16452: out = 16'(-4591);
			16453: out = 16'(-673);
			16454: out = 16'(1738);
			16455: out = 16'(5775);
			16456: out = 16'(10394);
			16457: out = 16'(7212);
			16458: out = 16'(-3);
			16459: out = 16'(-3490);
			16460: out = 16'(-2853);
			16461: out = 16'(-6530);
			16462: out = 16'(-9969);
			16463: out = 16'(-8773);
			16464: out = 16'(-431);
			16465: out = 16'(7869);
			16466: out = 16'(7913);
			16467: out = 16'(4096);
			16468: out = 16'(-1529);
			16469: out = 16'(-4772);
			16470: out = 16'(-7570);
			16471: out = 16'(-624);
			16472: out = 16'(2967);
			16473: out = 16'(125);
			16474: out = 16'(-5529);
			16475: out = 16'(3043);
			16476: out = 16'(7227);
			16477: out = 16'(2916);
			16478: out = 16'(720);
			16479: out = 16'(-165);
			16480: out = 16'(-1681);
			16481: out = 16'(-5896);
			16482: out = 16'(-3495);
			16483: out = 16'(1252);
			16484: out = 16'(9417);
			16485: out = 16'(8087);
			16486: out = 16'(-1176);
			16487: out = 16'(-6741);
			16488: out = 16'(-4043);
			16489: out = 16'(102);
			16490: out = 16'(-83);
			16491: out = 16'(408);
			16492: out = 16'(-760);
			16493: out = 16'(-1723);
			16494: out = 16'(-2171);
			16495: out = 16'(-992);
			16496: out = 16'(6141);
			16497: out = 16'(9445);
			16498: out = 16'(6500);
			16499: out = 16'(2063);
			16500: out = 16'(-8869);
			16501: out = 16'(-10053);
			16502: out = 16'(-1628);
			16503: out = 16'(6195);
			16504: out = 16'(1441);
			16505: out = 16'(-359);
			16506: out = 16'(5572);
			16507: out = 16'(10308);
			16508: out = 16'(-5657);
			16509: out = 16'(-14097);
			16510: out = 16'(-10792);
			16511: out = 16'(999);
			16512: out = 16'(1888);
			16513: out = 16'(8759);
			16514: out = 16'(10743);
			16515: out = 16'(8436);
			16516: out = 16'(1636);
			16517: out = 16'(-5352);
			16518: out = 16'(-10766);
			16519: out = 16'(-8847);
			16520: out = 16'(1184);
			16521: out = 16'(8574);
			16522: out = 16'(10020);
			16523: out = 16'(5139);
			16524: out = 16'(4);
			16525: out = 16'(-8410);
			16526: out = 16'(-5171);
			16527: out = 16'(-1191);
			16528: out = 16'(83);
			16529: out = 16'(-1566);
			16530: out = 16'(3732);
			16531: out = 16'(4119);
			16532: out = 16'(-1847);
			16533: out = 16'(-12369);
			16534: out = 16'(-3336);
			16535: out = 16'(2250);
			16536: out = 16'(1790);
			16537: out = 16'(74);
			16538: out = 16'(1404);
			16539: out = 16'(-2200);
			16540: out = 16'(-4789);
			16541: out = 16'(-1437);
			16542: out = 16'(5709);
			16543: out = 16'(4311);
			16544: out = 16'(1728);
			16545: out = 16'(2091);
			16546: out = 16'(-1244);
			16547: out = 16'(-4142);
			16548: out = 16'(-3424);
			16549: out = 16'(459);
			16550: out = 16'(-428);
			16551: out = 16'(171);
			16552: out = 16'(510);
			16553: out = 16'(895);
			16554: out = 16'(112);
			16555: out = 16'(-1215);
			16556: out = 16'(-576);
			16557: out = 16'(-1025);
			16558: out = 16'(-3556);
			16559: out = 16'(-2841);
			16560: out = 16'(3252);
			16561: out = 16'(7461);
			16562: out = 16'(5353);
			16563: out = 16'(-688);
			16564: out = 16'(-803);
			16565: out = 16'(-113);
			16566: out = 16'(-2204);
			16567: out = 16'(-4572);
			16568: out = 16'(21);
			16569: out = 16'(5107);
			16570: out = 16'(5268);
			16571: out = 16'(-174);
			16572: out = 16'(65);
			16573: out = 16'(-902);
			16574: out = 16'(-1033);
			16575: out = 16'(996);
			16576: out = 16'(4827);
			16577: out = 16'(2241);
			16578: out = 16'(-972);
			16579: out = 16'(262);
			16580: out = 16'(1555);
			16581: out = 16'(-679);
			16582: out = 16'(-3885);
			16583: out = 16'(-964);
			16584: out = 16'(5257);
			16585: out = 16'(9762);
			16586: out = 16'(5259);
			16587: out = 16'(-2154);
			16588: out = 16'(-2641);
			16589: out = 16'(-392);
			16590: out = 16'(662);
			16591: out = 16'(-1022);
			16592: out = 16'(-43);
			16593: out = 16'(1719);
			16594: out = 16'(4512);
			16595: out = 16'(-474);
			16596: out = 16'(-10381);
			16597: out = 16'(-3078);
			16598: out = 16'(6251);
			16599: out = 16'(7444);
			16600: out = 16'(-2723);
			16601: out = 16'(-4055);
			16602: out = 16'(-3431);
			16603: out = 16'(3233);
			16604: out = 16'(1098);
			16605: out = 16'(-6286);
			16606: out = 16'(-9195);
			16607: out = 16'(4056);
			16608: out = 16'(10004);
			16609: out = 16'(1609);
			16610: out = 16'(-19359);
			16611: out = 16'(-10255);
			16612: out = 16'(10293);
			16613: out = 16'(9994);
			16614: out = 16'(-8961);
			16615: out = 16'(-8738);
			16616: out = 16'(4538);
			16617: out = 16'(5559);
			16618: out = 16'(-7735);
			16619: out = 16'(-11141);
			16620: out = 16'(-3177);
			16621: out = 16'(2625);
			16622: out = 16'(2665);
			16623: out = 16'(431);
			16624: out = 16'(598);
			16625: out = 16'(1179);
			16626: out = 16'(2311);
			16627: out = 16'(-2519);
			16628: out = 16'(-5332);
			16629: out = 16'(-5438);
			16630: out = 16'(-1834);
			16631: out = 16'(-2578);
			16632: out = 16'(1970);
			16633: out = 16'(7095);
			16634: out = 16'(10049);
			16635: out = 16'(3613);
			16636: out = 16'(4104);
			16637: out = 16'(2776);
			16638: out = 16'(-2435);
			16639: out = 16'(-14857);
			16640: out = 16'(-3407);
			16641: out = 16'(6861);
			16642: out = 16'(5042);
			16643: out = 16'(-3219);
			16644: out = 16'(-2391);
			16645: out = 16'(541);
			16646: out = 16'(818);
			16647: out = 16'(-156);
			16648: out = 16'(-3436);
			16649: out = 16'(705);
			16650: out = 16'(5688);
			16651: out = 16'(2613);
			16652: out = 16'(-5271);
			16653: out = 16'(-11035);
			16654: out = 16'(-2164);
			16655: out = 16'(11841);
			16656: out = 16'(11460);
			16657: out = 16'(3656);
			16658: out = 16'(-4196);
			16659: out = 16'(-5867);
			16660: out = 16'(-2643);
			16661: out = 16'(172);
			16662: out = 16'(3134);
			16663: out = 16'(3662);
			16664: out = 16'(1006);
			16665: out = 16'(774);
			16666: out = 16'(769);
			16667: out = 16'(-2864);
			16668: out = 16'(-7607);
			16669: out = 16'(-11616);
			16670: out = 16'(2030);
			16671: out = 16'(13912);
			16672: out = 16'(11366);
			16673: out = 16'(1992);
			16674: out = 16'(-23);
			16675: out = 16'(1156);
			16676: out = 16'(-1936);
			16677: out = 16'(-6954);
			16678: out = 16'(-3034);
			16679: out = 16'(5075);
			16680: out = 16'(6159);
			16681: out = 16'(-2891);
			16682: out = 16'(68);
			16683: out = 16'(1814);
			16684: out = 16'(1190);
			16685: out = 16'(-114);
			16686: out = 16'(6786);
			16687: out = 16'(5129);
			16688: out = 16'(-2659);
			16689: out = 16'(-9719);
			16690: out = 16'(-14391);
			16691: out = 16'(-5513);
			16692: out = 16'(4577);
			16693: out = 16'(7523);
			16694: out = 16'(1175);
			16695: out = 16'(316);
			16696: out = 16'(-1340);
			16697: out = 16'(-2921);
			16698: out = 16'(-3863);
			16699: out = 16'(-357);
			16700: out = 16'(-2336);
			16701: out = 16'(-4444);
			16702: out = 16'(421);
			16703: out = 16'(-59);
			16704: out = 16'(842);
			16705: out = 16'(2261);
			16706: out = 16'(4089);
			16707: out = 16'(-3075);
			16708: out = 16'(-3902);
			16709: out = 16'(-4232);
			16710: out = 16'(-6473);
			16711: out = 16'(-5373);
			16712: out = 16'(-2259);
			16713: out = 16'(5978);
			16714: out = 16'(9359);
			16715: out = 16'(2448);
			16716: out = 16'(-11178);
			16717: out = 16'(-14364);
			16718: out = 16'(-6279);
			16719: out = 16'(-742);
			16720: out = 16'(9474);
			16721: out = 16'(9692);
			16722: out = 16'(5868);
			16723: out = 16'(2332);
			16724: out = 16'(458);
			16725: out = 16'(-2468);
			16726: out = 16'(-6415);
			16727: out = 16'(-5793);
			16728: out = 16'(-613);
			16729: out = 16'(5932);
			16730: out = 16'(4200);
			16731: out = 16'(448);
			16732: out = 16'(2282);
			16733: out = 16'(6329);
			16734: out = 16'(1621);
			16735: out = 16'(-6938);
			16736: out = 16'(-10621);
			16737: out = 16'(-1758);
			16738: out = 16'(1135);
			16739: out = 16'(1168);
			16740: out = 16'(3891);
			16741: out = 16'(4930);
			16742: out = 16'(1566);
			16743: out = 16'(1388);
			16744: out = 16'(4223);
			16745: out = 16'(1066);
			16746: out = 16'(-7108);
			16747: out = 16'(-5896);
			16748: out = 16'(4128);
			16749: out = 16'(4204);
			16750: out = 16'(1457);
			16751: out = 16'(1749);
			16752: out = 16'(4473);
			16753: out = 16'(551);
			16754: out = 16'(-7393);
			16755: out = 16'(-9748);
			16756: out = 16'(-4409);
			16757: out = 16'(3492);
			16758: out = 16'(10317);
			16759: out = 16'(13612);
			16760: out = 16'(5235);
			16761: out = 16'(-9077);
			16762: out = 16'(-8421);
			16763: out = 16'(4078);
			16764: out = 16'(6710);
			16765: out = 16'(-5221);
			16766: out = 16'(-12624);
			16767: out = 16'(-675);
			16768: out = 16'(10682);
			16769: out = 16'(6495);
			16770: out = 16'(1276);
			16771: out = 16'(542);
			16772: out = 16'(3666);
			16773: out = 16'(-1728);
			16774: out = 16'(-11965);
			16775: out = 16'(-10645);
			16776: out = 16'(592);
			16777: out = 16'(7746);
			16778: out = 16'(5870);
			16779: out = 16'(1906);
			16780: out = 16'(313);
			16781: out = 16'(-760);
			16782: out = 16'(-2606);
			16783: out = 16'(-2456);
			16784: out = 16'(-594);
			16785: out = 16'(315);
			16786: out = 16'(-603);
			16787: out = 16'(-3498);
			16788: out = 16'(-898);
			16789: out = 16'(960);
			16790: out = 16'(4582);
			16791: out = 16'(11218);
			16792: out = 16'(6109);
			16793: out = 16'(-3806);
			16794: out = 16'(-10603);
			16795: out = 16'(-6258);
			16796: out = 16'(-1221);
			16797: out = 16'(1583);
			16798: out = 16'(-361);
			16799: out = 16'(-2081);
			16800: out = 16'(-392);
			16801: out = 16'(1925);
			16802: out = 16'(962);
			16803: out = 16'(-3584);
			16804: out = 16'(-6317);
			16805: out = 16'(1213);
			16806: out = 16'(10607);
			16807: out = 16'(7684);
			16808: out = 16'(-6522);
			16809: out = 16'(-7675);
			16810: out = 16'(1643);
			16811: out = 16'(4409);
			16812: out = 16'(-5129);
			16813: out = 16'(-9412);
			16814: out = 16'(1244);
			16815: out = 16'(11753);
			16816: out = 16'(7833);
			16817: out = 16'(-2869);
			16818: out = 16'(-2895);
			16819: out = 16'(2556);
			16820: out = 16'(2312);
			16821: out = 16'(474);
			16822: out = 16'(-2430);
			16823: out = 16'(-1327);
			16824: out = 16'(-629);
			16825: out = 16'(-3427);
			16826: out = 16'(124);
			16827: out = 16'(3199);
			16828: out = 16'(4584);
			16829: out = 16'(3773);
			16830: out = 16'(-2953);
			16831: out = 16'(-6028);
			16832: out = 16'(-920);
			16833: out = 16'(6365);
			16834: out = 16'(4933);
			16835: out = 16'(-2575);
			16836: out = 16'(-5130);
			16837: out = 16'(1561);
			16838: out = 16'(5445);
			16839: out = 16'(4706);
			16840: out = 16'(1117);
			16841: out = 16'(-845);
			16842: out = 16'(-3945);
			16843: out = 16'(-843);
			16844: out = 16'(516);
			16845: out = 16'(632);
			16846: out = 16'(-305);
			16847: out = 16'(-3021);
			16848: out = 16'(-2628);
			16849: out = 16'(2682);
			16850: out = 16'(7685);
			16851: out = 16'(4772);
			16852: out = 16'(-636);
			16853: out = 16'(-1920);
			16854: out = 16'(2808);
			16855: out = 16'(3292);
			16856: out = 16'(4299);
			16857: out = 16'(1898);
			16858: out = 16'(-1677);
			16859: out = 16'(-7718);
			16860: out = 16'(-6864);
			16861: out = 16'(-5880);
			16862: out = 16'(-4108);
			16863: out = 16'(-1130);
			16864: out = 16'(9443);
			16865: out = 16'(8700);
			16866: out = 16'(-492);
			16867: out = 16'(-8076);
			16868: out = 16'(-990);
			16869: out = 16'(-118);
			16870: out = 16'(-5426);
			16871: out = 16'(-5673);
			16872: out = 16'(2494);
			16873: out = 16'(5915);
			16874: out = 16'(-1246);
			16875: out = 16'(-6452);
			16876: out = 16'(-1097);
			16877: out = 16'(7225);
			16878: out = 16'(2931);
			16879: out = 16'(-5200);
			16880: out = 16'(-8346);
			16881: out = 16'(2443);
			16882: out = 16'(876);
			16883: out = 16'(-4027);
			16884: out = 16'(-1850);
			16885: out = 16'(5726);
			16886: out = 16'(2585);
			16887: out = 16'(1167);
			16888: out = 16'(3367);
			16889: out = 16'(-2877);
			16890: out = 16'(-12293);
			16891: out = 16'(-5551);
			16892: out = 16'(9009);
			16893: out = 16'(4995);
			16894: out = 16'(-8311);
			16895: out = 16'(-4619);
			16896: out = 16'(10294);
			16897: out = 16'(5344);
			16898: out = 16'(-7672);
			16899: out = 16'(-8318);
			16900: out = 16'(4031);
			16901: out = 16'(5273);
			16902: out = 16'(1743);
			16903: out = 16'(2831);
			16904: out = 16'(6005);
			16905: out = 16'(-1878);
			16906: out = 16'(-8858);
			16907: out = 16'(-8649);
			16908: out = 16'(-1312);
			16909: out = 16'(229);
			16910: out = 16'(7059);
			16911: out = 16'(3679);
			16912: out = 16'(4837);
			16913: out = 16'(5865);
			16914: out = 16'(4411);
			16915: out = 16'(1220);
			16916: out = 16'(466);
			16917: out = 16'(-2675);
			16918: out = 16'(-10638);
			16919: out = 16'(-2942);
			16920: out = 16'(4713);
			16921: out = 16'(4059);
			16922: out = 16'(-2205);
			16923: out = 16'(2954);
			16924: out = 16'(7480);
			16925: out = 16'(3858);
			16926: out = 16'(-5477);
			16927: out = 16'(-699);
			16928: out = 16'(1565);
			16929: out = 16'(-397);
			16930: out = 16'(-5089);
			16931: out = 16'(179);
			16932: out = 16'(2742);
			16933: out = 16'(4731);
			16934: out = 16'(3211);
			16935: out = 16'(1905);
			16936: out = 16'(-8301);
			16937: out = 16'(-13224);
			16938: out = 16'(-8740);
			16939: out = 16'(3026);
			16940: out = 16'(5637);
			16941: out = 16'(6691);
			16942: out = 16'(4860);
			16943: out = 16'(1317);
			16944: out = 16'(-4088);
			16945: out = 16'(-6906);
			16946: out = 16'(-5841);
			16947: out = 16'(-1090);
			16948: out = 16'(2868);
			16949: out = 16'(8455);
			16950: out = 16'(8208);
			16951: out = 16'(1203);
			16952: out = 16'(-7936);
			16953: out = 16'(-13029);
			16954: out = 16'(-12669);
			16955: out = 16'(-8978);
			16956: out = 16'(-2496);
			16957: out = 16'(1451);
			16958: out = 16'(6674);
			16959: out = 16'(8238);
			16960: out = 16'(6109);
			16961: out = 16'(560);
			16962: out = 16'(-9);
			16963: out = 16'(-1982);
			16964: out = 16'(-5883);
			16965: out = 16'(-2427);
			16966: out = 16'(1182);
			16967: out = 16'(2875);
			16968: out = 16'(2211);
			16969: out = 16'(1207);
			16970: out = 16'(5128);
			16971: out = 16'(5961);
			16972: out = 16'(2546);
			16973: out = 16'(-2523);
			16974: out = 16'(-1562);
			16975: out = 16'(-2052);
			16976: out = 16'(-1406);
			16977: out = 16'(2863);
			16978: out = 16'(7210);
			16979: out = 16'(6154);
			16980: out = 16'(1776);
			16981: out = 16'(-1749);
			16982: out = 16'(-403);
			16983: out = 16'(-5735);
			16984: out = 16'(-8155);
			16985: out = 16'(-170);
			16986: out = 16'(12009);
			16987: out = 16'(10366);
			16988: out = 16'(2037);
			16989: out = 16'(-3242);
			16990: out = 16'(-2928);
			16991: out = 16'(-508);
			16992: out = 16'(-469);
			16993: out = 16'(-261);
			16994: out = 16'(-852);
			16995: out = 16'(1032);
			16996: out = 16'(-629);
			16997: out = 16'(3102);
			16998: out = 16'(8970);
			16999: out = 16'(2790);
			17000: out = 16'(-5095);
			17001: out = 16'(-6600);
			17002: out = 16'(-2978);
			17003: out = 16'(-7227);
			17004: out = 16'(-4959);
			17005: out = 16'(3649);
			17006: out = 16'(9325);
			17007: out = 16'(4005);
			17008: out = 16'(-146);
			17009: out = 16'(2823);
			17010: out = 16'(3746);
			17011: out = 16'(-6985);
			17012: out = 16'(-9798);
			17013: out = 16'(-2666);
			17014: out = 16'(6396);
			17015: out = 16'(4736);
			17016: out = 16'(911);
			17017: out = 16'(-1008);
			17018: out = 16'(120);
			17019: out = 16'(-1395);
			17020: out = 16'(-4607);
			17021: out = 16'(-3961);
			17022: out = 16'(-444);
			17023: out = 16'(2675);
			17024: out = 16'(3727);
			17025: out = 16'(1158);
			17026: out = 16'(-3463);
			17027: out = 16'(-3583);
			17028: out = 16'(1776);
			17029: out = 16'(2656);
			17030: out = 16'(-3932);
			17031: out = 16'(-8223);
			17032: out = 16'(-1544);
			17033: out = 16'(1257);
			17034: out = 16'(4279);
			17035: out = 16'(6230);
			17036: out = 16'(7077);
			17037: out = 16'(429);
			17038: out = 16'(-7673);
			17039: out = 16'(-12088);
			17040: out = 16'(-7198);
			17041: out = 16'(3532);
			17042: out = 16'(3427);
			17043: out = 16'(1560);
			17044: out = 16'(3044);
			17045: out = 16'(3523);
			17046: out = 16'(-1420);
			17047: out = 16'(-7287);
			17048: out = 16'(-7165);
			17049: out = 16'(-3737);
			17050: out = 16'(-2012);
			17051: out = 16'(-1551);
			17052: out = 16'(4087);
			17053: out = 16'(9592);
			17054: out = 16'(6210);
			17055: out = 16'(-1222);
			17056: out = 16'(-2799);
			17057: out = 16'(-534);
			17058: out = 16'(-3108);
			17059: out = 16'(-7054);
			17060: out = 16'(-1328);
			17061: out = 16'(7001);
			17062: out = 16'(1864);
			17063: out = 16'(2193);
			17064: out = 16'(4303);
			17065: out = 16'(5152);
			17066: out = 16'(-691);
			17067: out = 16'(-5148);
			17068: out = 16'(-4651);
			17069: out = 16'(-1315);
			17070: out = 16'(260);
			17071: out = 16'(476);
			17072: out = 16'(7936);
			17073: out = 16'(10678);
			17074: out = 16'(3694);
			17075: out = 16'(-4055);
			17076: out = 16'(-2599);
			17077: out = 16'(884);
			17078: out = 16'(-2213);
			17079: out = 16'(-7740);
			17080: out = 16'(-3166);
			17081: out = 16'(5970);
			17082: out = 16'(8811);
			17083: out = 16'(3594);
			17084: out = 16'(405);
			17085: out = 16'(-1277);
			17086: out = 16'(-2129);
			17087: out = 16'(-2990);
			17088: out = 16'(-4940);
			17089: out = 16'(-1663);
			17090: out = 16'(2099);
			17091: out = 16'(1876);
			17092: out = 16'(6163);
			17093: out = 16'(5568);
			17094: out = 16'(4212);
			17095: out = 16'(-3713);
			17096: out = 16'(-12345);
			17097: out = 16'(-19413);
			17098: out = 16'(-5887);
			17099: out = 16'(11094);
			17100: out = 16'(10483);
			17101: out = 16'(-486);
			17102: out = 16'(-3540);
			17103: out = 16'(1399);
			17104: out = 16'(929);
			17105: out = 16'(-6489);
			17106: out = 16'(-8532);
			17107: out = 16'(-1926);
			17108: out = 16'(4218);
			17109: out = 16'(-777);
			17110: out = 16'(3303);
			17111: out = 16'(7502);
			17112: out = 16'(3744);
			17113: out = 16'(-6209);
			17114: out = 16'(-4427);
			17115: out = 16'(3451);
			17116: out = 16'(3926);
			17117: out = 16'(-5753);
			17118: out = 16'(-9688);
			17119: out = 16'(-4888);
			17120: out = 16'(1960);
			17121: out = 16'(3092);
			17122: out = 16'(1737);
			17123: out = 16'(498);
			17124: out = 16'(-1775);
			17125: out = 16'(-5936);
			17126: out = 16'(-1473);
			17127: out = 16'(21);
			17128: out = 16'(336);
			17129: out = 16'(1046);
			17130: out = 16'(6140);
			17131: out = 16'(4052);
			17132: out = 16'(-1119);
			17133: out = 16'(-4404);
			17134: out = 16'(253);
			17135: out = 16'(-1627);
			17136: out = 16'(-3216);
			17137: out = 16'(-2451);
			17138: out = 16'(1240);
			17139: out = 16'(504);
			17140: out = 16'(607);
			17141: out = 16'(2501);
			17142: out = 16'(3891);
			17143: out = 16'(-1222);
			17144: out = 16'(-6071);
			17145: out = 16'(-4291);
			17146: out = 16'(3649);
			17147: out = 16'(3843);
			17148: out = 16'(4819);
			17149: out = 16'(3985);
			17150: out = 16'(4309);
			17151: out = 16'(1724);
			17152: out = 16'(967);
			17153: out = 16'(-3609);
			17154: out = 16'(-5075);
			17155: out = 16'(146);
			17156: out = 16'(2088);
			17157: out = 16'(957);
			17158: out = 16'(954);
			17159: out = 16'(4165);
			17160: out = 16'(1407);
			17161: out = 16'(-2251);
			17162: out = 16'(-2972);
			17163: out = 16'(494);
			17164: out = 16'(1888);
			17165: out = 16'(-1421);
			17166: out = 16'(-4106);
			17167: out = 16'(-1449);
			17168: out = 16'(-367);
			17169: out = 16'(3445);
			17170: out = 16'(5242);
			17171: out = 16'(5463);
			17172: out = 16'(-584);
			17173: out = 16'(1166);
			17174: out = 16'(-2949);
			17175: out = 16'(-6495);
			17176: out = 16'(-4019);
			17177: out = 16'(5889);
			17178: out = 16'(10809);
			17179: out = 16'(9643);
			17180: out = 16'(3195);
			17181: out = 16'(-5631);
			17182: out = 16'(-13729);
			17183: out = 16'(-11482);
			17184: out = 16'(-574);
			17185: out = 16'(3612);
			17186: out = 16'(4577);
			17187: out = 16'(4064);
			17188: out = 16'(3506);
			17189: out = 16'(-155);
			17190: out = 16'(-5715);
			17191: out = 16'(-5096);
			17192: out = 16'(2472);
			17193: out = 16'(5197);
			17194: out = 16'(1671);
			17195: out = 16'(-3611);
			17196: out = 16'(-678);
			17197: out = 16'(5390);
			17198: out = 16'(-4146);
			17199: out = 16'(-5858);
			17200: out = 16'(3597);
			17201: out = 16'(10125);
			17202: out = 16'(1300);
			17203: out = 16'(-11677);
			17204: out = 16'(-10625);
			17205: out = 16'(2062);
			17206: out = 16'(3713);
			17207: out = 16'(400);
			17208: out = 16'(479);
			17209: out = 16'(5281);
			17210: out = 16'(3361);
			17211: out = 16'(-1533);
			17212: out = 16'(-5996);
			17213: out = 16'(-4476);
			17214: out = 16'(-96);
			17215: out = 16'(-2180);
			17216: out = 16'(1304);
			17217: out = 16'(5828);
			17218: out = 16'(5312);
			17219: out = 16'(781);
			17220: out = 16'(-1461);
			17221: out = 16'(-577);
			17222: out = 16'(544);
			17223: out = 16'(-2563);
			17224: out = 16'(-894);
			17225: out = 16'(-246);
			17226: out = 16'(522);
			17227: out = 16'(4075);
			17228: out = 16'(5120);
			17229: out = 16'(2492);
			17230: out = 16'(-837);
			17231: out = 16'(-370);
			17232: out = 16'(-4522);
			17233: out = 16'(-3095);
			17234: out = 16'(2229);
			17235: out = 16'(5697);
			17236: out = 16'(4535);
			17237: out = 16'(1904);
			17238: out = 16'(4010);
			17239: out = 16'(7017);
			17240: out = 16'(2149);
			17241: out = 16'(-3728);
			17242: out = 16'(-4053);
			17243: out = 16'(-412);
			17244: out = 16'(-1986);
			17245: out = 16'(-3684);
			17246: out = 16'(-1573);
			17247: out = 16'(2842);
			17248: out = 16'(2402);
			17249: out = 16'(3041);
			17250: out = 16'(943);
			17251: out = 16'(-1509);
			17252: out = 16'(-3104);
			17253: out = 16'(-6389);
			17254: out = 16'(-2474);
			17255: out = 16'(2373);
			17256: out = 16'(3481);
			17257: out = 16'(-473);
			17258: out = 16'(1019);
			17259: out = 16'(256);
			17260: out = 16'(-4308);
			17261: out = 16'(-8399);
			17262: out = 16'(122);
			17263: out = 16'(6399);
			17264: out = 16'(3571);
			17265: out = 16'(-2507);
			17266: out = 16'(-776);
			17267: out = 16'(1872);
			17268: out = 16'(762);
			17269: out = 16'(-443);
			17270: out = 16'(-2232);
			17271: out = 16'(1912);
			17272: out = 16'(2862);
			17273: out = 16'(-1539);
			17274: out = 16'(-4829);
			17275: out = 16'(-1875);
			17276: out = 16'(1178);
			17277: out = 16'(-1321);
			17278: out = 16'(-2154);
			17279: out = 16'(-1683);
			17280: out = 16'(1561);
			17281: out = 16'(939);
			17282: out = 16'(253);
			17283: out = 16'(319);
			17284: out = 16'(6870);
			17285: out = 16'(7562);
			17286: out = 16'(1031);
			17287: out = 16'(-14739);
			17288: out = 16'(-10448);
			17289: out = 16'(1230);
			17290: out = 16'(2930);
			17291: out = 16'(-5063);
			17292: out = 16'(-510);
			17293: out = 16'(6512);
			17294: out = 16'(3904);
			17295: out = 16'(-3951);
			17296: out = 16'(-2792);
			17297: out = 16'(2834);
			17298: out = 16'(2124);
			17299: out = 16'(-4466);
			17300: out = 16'(-3393);
			17301: out = 16'(3934);
			17302: out = 16'(6862);
			17303: out = 16'(21);
			17304: out = 16'(-4915);
			17305: out = 16'(-5583);
			17306: out = 16'(1165);
			17307: out = 16'(7476);
			17308: out = 16'(4739);
			17309: out = 16'(-3019);
			17310: out = 16'(-5526);
			17311: out = 16'(837);
			17312: out = 16'(-1116);
			17313: out = 16'(4684);
			17314: out = 16'(3801);
			17315: out = 16'(-2991);
			17316: out = 16'(-13584);
			17317: out = 16'(-13589);
			17318: out = 16'(-8155);
			17319: out = 16'(1800);
			17320: out = 16'(11641);
			17321: out = 16'(14553);
			17322: out = 16'(7891);
			17323: out = 16'(-3101);
			17324: out = 16'(-12909);
			17325: out = 16'(-9227);
			17326: out = 16'(-7908);
			17327: out = 16'(-4660);
			17328: out = 16'(2934);
			17329: out = 16'(11731);
			17330: out = 16'(9968);
			17331: out = 16'(5077);
			17332: out = 16'(640);
			17333: out = 16'(-4826);
			17334: out = 16'(-9906);
			17335: out = 16'(-8570);
			17336: out = 16'(-1536);
			17337: out = 16'(-472);
			17338: out = 16'(2781);
			17339: out = 16'(-433);
			17340: out = 16'(-1347);
			17341: out = 16'(2703);
			17342: out = 16'(4243);
			17343: out = 16'(1889);
			17344: out = 16'(-763);
			17345: out = 16'(533);
			17346: out = 16'(3706);
			17347: out = 16'(2737);
			17348: out = 16'(-880);
			17349: out = 16'(-1782);
			17350: out = 16'(1683);
			17351: out = 16'(4088);
			17352: out = 16'(1002);
			17353: out = 16'(-6155);
			17354: out = 16'(-13177);
			17355: out = 16'(-7392);
			17356: out = 16'(-132);
			17357: out = 16'(3166);
			17358: out = 16'(4789);
			17359: out = 16'(7526);
			17360: out = 16'(4488);
			17361: out = 16'(-4340);
			17362: out = 16'(-10786);
			17363: out = 16'(-14139);
			17364: out = 16'(-4560);
			17365: out = 16'(3072);
			17366: out = 16'(4467);
			17367: out = 16'(460);
			17368: out = 16'(8622);
			17369: out = 16'(11783);
			17370: out = 16'(6857);
			17371: out = 16'(-94);
			17372: out = 16'(-3635);
			17373: out = 16'(-8797);
			17374: out = 16'(-11020);
			17375: out = 16'(-1527);
			17376: out = 16'(1522);
			17377: out = 16'(4930);
			17378: out = 16'(7840);
			17379: out = 16'(8986);
			17380: out = 16'(-2491);
			17381: out = 16'(-9791);
			17382: out = 16'(-7520);
			17383: out = 16'(884);
			17384: out = 16'(-2091);
			17385: out = 16'(-1066);
			17386: out = 16'(3704);
			17387: out = 16'(7797);
			17388: out = 16'(181);
			17389: out = 16'(678);
			17390: out = 16'(1829);
			17391: out = 16'(1573);
			17392: out = 16'(-1156);
			17393: out = 16'(-2584);
			17394: out = 16'(1105);
			17395: out = 16'(4962);
			17396: out = 16'(3723);
			17397: out = 16'(450);
			17398: out = 16'(176);
			17399: out = 16'(722);
			17400: out = 16'(-2806);
			17401: out = 16'(-13503);
			17402: out = 16'(-9989);
			17403: out = 16'(1893);
			17404: out = 16'(8211);
			17405: out = 16'(6766);
			17406: out = 16'(2908);
			17407: out = 16'(3838);
			17408: out = 16'(5891);
			17409: out = 16'(1588);
			17410: out = 16'(-6595);
			17411: out = 16'(-12571);
			17412: out = 16'(-9229);
			17413: out = 16'(407);
			17414: out = 16'(5747);
			17415: out = 16'(8488);
			17416: out = 16'(11018);
			17417: out = 16'(10184);
			17418: out = 16'(3632);
			17419: out = 16'(-8620);
			17420: out = 16'(-14630);
			17421: out = 16'(-9769);
			17422: out = 16'(-5526);
			17423: out = 16'(-1167);
			17424: out = 16'(2090);
			17425: out = 16'(4909);
			17426: out = 16'(4229);
			17427: out = 16'(2901);
			17428: out = 16'(2044);
			17429: out = 16'(1520);
			17430: out = 16'(-2949);
			17431: out = 16'(-6112);
			17432: out = 16'(-6767);
			17433: out = 16'(-1976);
			17434: out = 16'(2720);
			17435: out = 16'(9795);
			17436: out = 16'(4112);
			17437: out = 16'(-1145);
			17438: out = 16'(1082);
			17439: out = 16'(7190);
			17440: out = 16'(1797);
			17441: out = 16'(-7070);
			17442: out = 16'(-7848);
			17443: out = 16'(1364);
			17444: out = 16'(1584);
			17445: out = 16'(-4780);
			17446: out = 16'(-6542);
			17447: out = 16'(2472);
			17448: out = 16'(6168);
			17449: out = 16'(18);
			17450: out = 16'(-9911);
			17451: out = 16'(-10061);
			17452: out = 16'(1341);
			17453: out = 16'(10611);
			17454: out = 16'(9027);
			17455: out = 16'(3867);
			17456: out = 16'(-1);
			17457: out = 16'(3197);
			17458: out = 16'(1336);
			17459: out = 16'(-6766);
			17460: out = 16'(-15112);
			17461: out = 16'(-3685);
			17462: out = 16'(7352);
			17463: out = 16'(6644);
			17464: out = 16'(5140);
			17465: out = 16'(3291);
			17466: out = 16'(5353);
			17467: out = 16'(263);
			17468: out = 16'(-9259);
			17469: out = 16'(-14908);
			17470: out = 16'(-6036);
			17471: out = 16'(1808);
			17472: out = 16'(101);
			17473: out = 16'(283);
			17474: out = 16'(6360);
			17475: out = 16'(11011);
			17476: out = 16'(8108);
			17477: out = 16'(1514);
			17478: out = 16'(564);
			17479: out = 16'(808);
			17480: out = 16'(-1634);
			17481: out = 16'(-7048);
			17482: out = 16'(-5338);
			17483: out = 16'(-2547);
			17484: out = 16'(2994);
			17485: out = 16'(9180);
			17486: out = 16'(7473);
			17487: out = 16'(-2431);
			17488: out = 16'(-8047);
			17489: out = 16'(-1366);
			17490: out = 16'(1388);
			17491: out = 16'(1243);
			17492: out = 16'(-332);
			17493: out = 16'(-251);
			17494: out = 16'(-4279);
			17495: out = 16'(-5848);
			17496: out = 16'(-3346);
			17497: out = 16'(769);
			17498: out = 16'(278);
			17499: out = 16'(-141);
			17500: out = 16'(3676);
			17501: out = 16'(9193);
			17502: out = 16'(8874);
			17503: out = 16'(2007);
			17504: out = 16'(-2313);
			17505: out = 16'(-2352);
			17506: out = 16'(-3112);
			17507: out = 16'(-7250);
			17508: out = 16'(-7722);
			17509: out = 16'(-2321);
			17510: out = 16'(3658);
			17511: out = 16'(2385);
			17512: out = 16'(841);
			17513: out = 16'(-335);
			17514: out = 16'(1051);
			17515: out = 16'(3741);
			17516: out = 16'(2595);
			17517: out = 16'(-3640);
			17518: out = 16'(-7840);
			17519: out = 16'(-3107);
			17520: out = 16'(-310);
			17521: out = 16'(335);
			17522: out = 16'(1034);
			17523: out = 16'(4698);
			17524: out = 16'(6078);
			17525: out = 16'(603);
			17526: out = 16'(-7864);
			17527: out = 16'(-8836);
			17528: out = 16'(2385);
			17529: out = 16'(4859);
			17530: out = 16'(-2785);
			17531: out = 16'(-8151);
			17532: out = 16'(-723);
			17533: out = 16'(5629);
			17534: out = 16'(3914);
			17535: out = 16'(-391);
			17536: out = 16'(-2136);
			17537: out = 16'(3311);
			17538: out = 16'(2571);
			17539: out = 16'(268);
			17540: out = 16'(2246);
			17541: out = 16'(739);
			17542: out = 16'(-4454);
			17543: out = 16'(-4878);
			17544: out = 16'(3258);
			17545: out = 16'(4040);
			17546: out = 16'(2380);
			17547: out = 16'(1596);
			17548: out = 16'(5284);
			17549: out = 16'(9050);
			17550: out = 16'(4682);
			17551: out = 16'(-1503);
			17552: out = 16'(-5372);
			17553: out = 16'(-4558);
			17554: out = 16'(-7900);
			17555: out = 16'(-4608);
			17556: out = 16'(1040);
			17557: out = 16'(1311);
			17558: out = 16'(5101);
			17559: out = 16'(8725);
			17560: out = 16'(7018);
			17561: out = 16'(-1339);
			17562: out = 16'(-8506);
			17563: out = 16'(-6015);
			17564: out = 16'(57);
			17565: out = 16'(2215);
			17566: out = 16'(2133);
			17567: out = 16'(6749);
			17568: out = 16'(6898);
			17569: out = 16'(-387);
			17570: out = 16'(-6347);
			17571: out = 16'(-4659);
			17572: out = 16'(516);
			17573: out = 16'(1961);
			17574: out = 16'(2275);
			17575: out = 16'(22);
			17576: out = 16'(53);
			17577: out = 16'(-1126);
			17578: out = 16'(-3234);
			17579: out = 16'(2720);
			17580: out = 16'(4950);
			17581: out = 16'(-4);
			17582: out = 16'(-8946);
			17583: out = 16'(-7215);
			17584: out = 16'(-133);
			17585: out = 16'(7106);
			17586: out = 16'(6047);
			17587: out = 16'(853);
			17588: out = 16'(-6153);
			17589: out = 16'(-4939);
			17590: out = 16'(-719);
			17591: out = 16'(-40);
			17592: out = 16'(-6578);
			17593: out = 16'(-5684);
			17594: out = 16'(1993);
			17595: out = 16'(7489);
			17596: out = 16'(1432);
			17597: out = 16'(-658);
			17598: out = 16'(431);
			17599: out = 16'(116);
			17600: out = 16'(-8106);
			17601: out = 16'(-7842);
			17602: out = 16'(-2529);
			17603: out = 16'(2323);
			17604: out = 16'(6094);
			17605: out = 16'(5317);
			17606: out = 16'(2232);
			17607: out = 16'(-208);
			17608: out = 16'(153);
			17609: out = 16'(389);
			17610: out = 16'(-1985);
			17611: out = 16'(-5606);
			17612: out = 16'(-7521);
			17613: out = 16'(632);
			17614: out = 16'(2780);
			17615: out = 16'(605);
			17616: out = 16'(1042);
			17617: out = 16'(5407);
			17618: out = 16'(4002);
			17619: out = 16'(-919);
			17620: out = 16'(-1843);
			17621: out = 16'(-5042);
			17622: out = 16'(780);
			17623: out = 16'(1740);
			17624: out = 16'(544);
			17625: out = 16'(2004);
			17626: out = 16'(2951);
			17627: out = 16'(-1175);
			17628: out = 16'(-3582);
			17629: out = 16'(2358);
			17630: out = 16'(2607);
			17631: out = 16'(706);
			17632: out = 16'(638);
			17633: out = 16'(2167);
			17634: out = 16'(7717);
			17635: out = 16'(2820);
			17636: out = 16'(679);
			17637: out = 16'(3800);
			17638: out = 16'(2600);
			17639: out = 16'(-8529);
			17640: out = 16'(-10643);
			17641: out = 16'(3103);
			17642: out = 16'(9737);
			17643: out = 16'(5586);
			17644: out = 16'(-1204);
			17645: out = 16'(-325);
			17646: out = 16'(1148);
			17647: out = 16'(2598);
			17648: out = 16'(-1871);
			17649: out = 16'(-5205);
			17650: out = 16'(-3327);
			17651: out = 16'(992);
			17652: out = 16'(1388);
			17653: out = 16'(-906);
			17654: out = 16'(375);
			17655: out = 16'(-970);
			17656: out = 16'(5646);
			17657: out = 16'(4569);
			17658: out = 16'(-4174);
			17659: out = 16'(-9020);
			17660: out = 16'(-1984);
			17661: out = 16'(2784);
			17662: out = 16'(-2007);
			17663: out = 16'(-4759);
			17664: out = 16'(464);
			17665: out = 16'(9391);
			17666: out = 16'(7375);
			17667: out = 16'(-5887);
			17668: out = 16'(-6800);
			17669: out = 16'(-229);
			17670: out = 16'(3937);
			17671: out = 16'(-908);
			17672: out = 16'(-2728);
			17673: out = 16'(-2380);
			17674: out = 16'(2007);
			17675: out = 16'(3370);
			17676: out = 16'(733);
			17677: out = 16'(-2395);
			17678: out = 16'(-520);
			17679: out = 16'(1831);
			17680: out = 16'(188);
			17681: out = 16'(-5489);
			17682: out = 16'(-5818);
			17683: out = 16'(-228);
			17684: out = 16'(5912);
			17685: out = 16'(1908);
			17686: out = 16'(1062);
			17687: out = 16'(1912);
			17688: out = 16'(-955);
			17689: out = 16'(-9963);
			17690: out = 16'(-12107);
			17691: out = 16'(-4495);
			17692: out = 16'(5233);
			17693: out = 16'(7609);
			17694: out = 16'(4767);
			17695: out = 16'(-1101);
			17696: out = 16'(-4107);
			17697: out = 16'(459);
			17698: out = 16'(940);
			17699: out = 16'(-1985);
			17700: out = 16'(-1773);
			17701: out = 16'(5951);
			17702: out = 16'(7946);
			17703: out = 16'(3662);
			17704: out = 16'(-973);
			17705: out = 16'(628);
			17706: out = 16'(-4919);
			17707: out = 16'(-8000);
			17708: out = 16'(-5434);
			17709: out = 16'(3055);
			17710: out = 16'(3692);
			17711: out = 16'(4363);
			17712: out = 16'(3886);
			17713: out = 16'(4010);
			17714: out = 16'(3826);
			17715: out = 16'(897);
			17716: out = 16'(-1053);
			17717: out = 16'(-180);
			17718: out = 16'(-523);
			17719: out = 16'(-4448);
			17720: out = 16'(-5546);
			17721: out = 16'(-61);
			17722: out = 16'(3419);
			17723: out = 16'(6473);
			17724: out = 16'(1849);
			17725: out = 16'(7);
			17726: out = 16'(1528);
			17727: out = 16'(1613);
			17728: out = 16'(-6947);
			17729: out = 16'(-8857);
			17730: out = 16'(1850);
			17731: out = 16'(6577);
			17732: out = 16'(5879);
			17733: out = 16'(1380);
			17734: out = 16'(-1059);
			17735: out = 16'(-5158);
			17736: out = 16'(-2354);
			17737: out = 16'(-1760);
			17738: out = 16'(-3074);
			17739: out = 16'(-3220);
			17740: out = 16'(1471);
			17741: out = 16'(5540);
			17742: out = 16'(4079);
			17743: out = 16'(-426);
			17744: out = 16'(-951);
			17745: out = 16'(3724);
			17746: out = 16'(4333);
			17747: out = 16'(-1827);
			17748: out = 16'(-6687);
			17749: out = 16'(-3335);
			17750: out = 16'(2446);
			17751: out = 16'(3008);
			17752: out = 16'(-1179);
			17753: out = 16'(531);
			17754: out = 16'(2617);
			17755: out = 16'(-743);
			17756: out = 16'(-10613);
			17757: out = 16'(-2407);
			17758: out = 16'(3901);
			17759: out = 16'(1052);
			17760: out = 16'(-6867);
			17761: out = 16'(2095);
			17762: out = 16'(6172);
			17763: out = 16'(3699);
			17764: out = 16'(-334);
			17765: out = 16'(-471);
			17766: out = 16'(-555);
			17767: out = 16'(-4512);
			17768: out = 16'(-7184);
			17769: out = 16'(3509);
			17770: out = 16'(7877);
			17771: out = 16'(5157);
			17772: out = 16'(-1535);
			17773: out = 16'(213);
			17774: out = 16'(-3014);
			17775: out = 16'(-51);
			17776: out = 16'(1592);
			17777: out = 16'(-470);
			17778: out = 16'(-5283);
			17779: out = 16'(-4647);
			17780: out = 16'(-731);
			17781: out = 16'(2041);
			17782: out = 16'(126);
			17783: out = 16'(-659);
			17784: out = 16'(-3088);
			17785: out = 16'(-5594);
			17786: out = 16'(-1440);
			17787: out = 16'(1475);
			17788: out = 16'(2002);
			17789: out = 16'(930);
			17790: out = 16'(2220);
			17791: out = 16'(-1913);
			17792: out = 16'(-5295);
			17793: out = 16'(-3616);
			17794: out = 16'(4456);
			17795: out = 16'(2695);
			17796: out = 16'(912);
			17797: out = 16'(515);
			17798: out = 16'(2095);
			17799: out = 16'(-1801);
			17800: out = 16'(-3262);
			17801: out = 16'(-2755);
			17802: out = 16'(-460);
			17803: out = 16'(3907);
			17804: out = 16'(1811);
			17805: out = 16'(-1443);
			17806: out = 16'(-1093);
			17807: out = 16'(5813);
			17808: out = 16'(1932);
			17809: out = 16'(-1849);
			17810: out = 16'(-1060);
			17811: out = 16'(4094);
			17812: out = 16'(4162);
			17813: out = 16'(2951);
			17814: out = 16'(1415);
			17815: out = 16'(368);
			17816: out = 16'(-5183);
			17817: out = 16'(-4611);
			17818: out = 16'(-463);
			17819: out = 16'(1775);
			17820: out = 16'(-864);
			17821: out = 16'(-1023);
			17822: out = 16'(2612);
			17823: out = 16'(5370);
			17824: out = 16'(-1260);
			17825: out = 16'(-3179);
			17826: out = 16'(-2476);
			17827: out = 16'(1584);
			17828: out = 16'(5346);
			17829: out = 16'(1646);
			17830: out = 16'(-4223);
			17831: out = 16'(-4292);
			17832: out = 16'(2320);
			17833: out = 16'(5420);
			17834: out = 16'(3801);
			17835: out = 16'(809);
			17836: out = 16'(-603);
			17837: out = 16'(-4368);
			17838: out = 16'(-4274);
			17839: out = 16'(1437);
			17840: out = 16'(7306);
			17841: out = 16'(10);
			17842: out = 16'(-817);
			17843: out = 16'(2072);
			17844: out = 16'(5451);
			17845: out = 16'(-1152);
			17846: out = 16'(-2542);
			17847: out = 16'(-7770);
			17848: out = 16'(-10933);
			17849: out = 16'(-7728);
			17850: out = 16'(1936);
			17851: out = 16'(4185);
			17852: out = 16'(640);
			17853: out = 16'(618);
			17854: out = 16'(1006);
			17855: out = 16'(4503);
			17856: out = 16'(-919);
			17857: out = 16'(-10915);
			17858: out = 16'(-5184);
			17859: out = 16'(4109);
			17860: out = 16'(8498);
			17861: out = 16'(4309);
			17862: out = 16'(617);
			17863: out = 16'(-3218);
			17864: out = 16'(-2085);
			17865: out = 16'(438);
			17866: out = 16'(-337);
			17867: out = 16'(-764);
			17868: out = 16'(-2397);
			17869: out = 16'(-1587);
			17870: out = 16'(4);
			17871: out = 16'(3959);
			17872: out = 16'(1467);
			17873: out = 16'(613);
			17874: out = 16'(2777);
			17875: out = 16'(-852);
			17876: out = 16'(-7131);
			17877: out = 16'(-7944);
			17878: out = 16'(-309);
			17879: out = 16'(5292);
			17880: out = 16'(2975);
			17881: out = 16'(-630);
			17882: out = 16'(2177);
			17883: out = 16'(8798);
			17884: out = 16'(1610);
			17885: out = 16'(-6304);
			17886: out = 16'(-6538);
			17887: out = 16'(84);
			17888: out = 16'(187);
			17889: out = 16'(232);
			17890: out = 16'(2078);
			17891: out = 16'(3729);
			17892: out = 16'(569);
			17893: out = 16'(-778);
			17894: out = 16'(1529);
			17895: out = 16'(3329);
			17896: out = 16'(-2024);
			17897: out = 16'(-2567);
			17898: out = 16'(2093);
			17899: out = 16'(5289);
			17900: out = 16'(-445);
			17901: out = 16'(-3321);
			17902: out = 16'(-1260);
			17903: out = 16'(2238);
			17904: out = 16'(-821);
			17905: out = 16'(-2734);
			17906: out = 16'(-3855);
			17907: out = 16'(-788);
			17908: out = 16'(1857);
			17909: out = 16'(2317);
			17910: out = 16'(-250);
			17911: out = 16'(-1730);
			17912: out = 16'(-734);
			17913: out = 16'(5598);
			17914: out = 16'(-898);
			17915: out = 16'(-7307);
			17916: out = 16'(-4998);
			17917: out = 16'(3313);
			17918: out = 16'(2571);
			17919: out = 16'(-1817);
			17920: out = 16'(-10);
			17921: out = 16'(7217);
			17922: out = 16'(7168);
			17923: out = 16'(-2061);
			17924: out = 16'(-8870);
			17925: out = 16'(-3639);
			17926: out = 16'(5928);
			17927: out = 16'(2872);
			17928: out = 16'(-6011);
			17929: out = 16'(-4975);
			17930: out = 16'(5518);
			17931: out = 16'(9538);
			17932: out = 16'(1106);
			17933: out = 16'(-7371);
			17934: out = 16'(-4144);
			17935: out = 16'(6472);
			17936: out = 16'(6334);
			17937: out = 16'(-3457);
			17938: out = 16'(-7214);
			17939: out = 16'(200);
			17940: out = 16'(7946);
			17941: out = 16'(3190);
			17942: out = 16'(-8215);
			17943: out = 16'(-10497);
			17944: out = 16'(-424);
			17945: out = 16'(7495);
			17946: out = 16'(4960);
			17947: out = 16'(2657);
			17948: out = 16'(233);
			17949: out = 16'(-2768);
			17950: out = 16'(-7383);
			17951: out = 16'(-104);
			17952: out = 16'(792);
			17953: out = 16'(5088);
			17954: out = 16'(6458);
			17955: out = 16'(-358);
			17956: out = 16'(-3428);
			17957: out = 16'(-1224);
			17958: out = 16'(2662);
			17959: out = 16'(1198);
			17960: out = 16'(-3281);
			17961: out = 16'(-7154);
			17962: out = 16'(-5234);
			17963: out = 16'(152);
			17964: out = 16'(1891);
			17965: out = 16'(2757);
			17966: out = 16'(2866);
			17967: out = 16'(1874);
			17968: out = 16'(4049);
			17969: out = 16'(-1998);
			17970: out = 16'(-7237);
			17971: out = 16'(-6844);
			17972: out = 16'(1952);
			17973: out = 16'(2122);
			17974: out = 16'(2141);
			17975: out = 16'(1491);
			17976: out = 16'(34);
			17977: out = 16'(-466);
			17978: out = 16'(2289);
			17979: out = 16'(3473);
			17980: out = 16'(-32);
			17981: out = 16'(-6253);
			17982: out = 16'(-3833);
			17983: out = 16'(3093);
			17984: out = 16'(4852);
			17985: out = 16'(-2610);
			17986: out = 16'(-3765);
			17987: out = 16'(-518);
			17988: out = 16'(721);
			17989: out = 16'(345);
			17990: out = 16'(-508);
			17991: out = 16'(1335);
			17992: out = 16'(1409);
			17993: out = 16'(247);
			17994: out = 16'(-6305);
			17995: out = 16'(-1774);
			17996: out = 16'(6036);
			17997: out = 16'(4868);
			17998: out = 16'(-1615);
			17999: out = 16'(-6123);
			18000: out = 16'(-3977);
			18001: out = 16'(-1);
			18002: out = 16'(846);
			18003: out = 16'(2815);
			18004: out = 16'(5309);
			18005: out = 16'(4999);
			18006: out = 16'(257);
			18007: out = 16'(-839);
			18008: out = 16'(1610);
			18009: out = 16'(3653);
			18010: out = 16'(259);
			18011: out = 16'(900);
			18012: out = 16'(-1433);
			18013: out = 16'(-5464);
			18014: out = 16'(-7804);
			18015: out = 16'(1576);
			18016: out = 16'(7175);
			18017: out = 16'(5384);
			18018: out = 16'(0);
			18019: out = 16'(-2612);
			18020: out = 16'(-2052);
			18021: out = 16'(-3023);
			18022: out = 16'(-6327);
			18023: out = 16'(-2473);
			18024: out = 16'(-1075);
			18025: out = 16'(1942);
			18026: out = 16'(4455);
			18027: out = 16'(5695);
			18028: out = 16'(-2127);
			18029: out = 16'(-6727);
			18030: out = 16'(-4146);
			18031: out = 16'(691);
			18032: out = 16'(-482);
			18033: out = 16'(-3316);
			18034: out = 16'(-1441);
			18035: out = 16'(4434);
			18036: out = 16'(5882);
			18037: out = 16'(371);
			18038: out = 16'(-5791);
			18039: out = 16'(-4476);
			18040: out = 16'(2904);
			18041: out = 16'(6277);
			18042: out = 16'(2882);
			18043: out = 16'(-2801);
			18044: out = 16'(-7015);
			18045: out = 16'(-5655);
			18046: out = 16'(-2446);
			18047: out = 16'(495);
			18048: out = 16'(23);
			18049: out = 16'(5420);
			18050: out = 16'(3357);
			18051: out = 16'(-1883);
			18052: out = 16'(-4149);
			18053: out = 16'(1016);
			18054: out = 16'(2943);
			18055: out = 16'(-507);
			18056: out = 16'(-5664);
			18057: out = 16'(1727);
			18058: out = 16'(2385);
			18059: out = 16'(1059);
			18060: out = 16'(-1784);
			18061: out = 16'(371);
			18062: out = 16'(-2551);
			18063: out = 16'(1991);
			18064: out = 16'(7143);
			18065: out = 16'(3814);
			18066: out = 16'(-473);
			18067: out = 16'(888);
			18068: out = 16'(3805);
			18069: out = 16'(-832);
			18070: out = 16'(76);
			18071: out = 16'(76);
			18072: out = 16'(1404);
			18073: out = 16'(1576);
			18074: out = 16'(18);
			18075: out = 16'(-353);
			18076: out = 16'(-938);
			18077: out = 16'(-3129);
			18078: out = 16'(-4593);
			18079: out = 16'(-2783);
			18080: out = 16'(340);
			18081: out = 16'(2929);
			18082: out = 16'(6596);
			18083: out = 16'(837);
			18084: out = 16'(-4592);
			18085: out = 16'(-4860);
			18086: out = 16'(-147);
			18087: out = 16'(-2741);
			18088: out = 16'(-3137);
			18089: out = 16'(1370);
			18090: out = 16'(5844);
			18091: out = 16'(6423);
			18092: out = 16'(1645);
			18093: out = 16'(-692);
			18094: out = 16'(-854);
			18095: out = 16'(-990);
			18096: out = 16'(-3970);
			18097: out = 16'(1277);
			18098: out = 16'(8580);
			18099: out = 16'(3699);
			18100: out = 16'(-4610);
			18101: out = 16'(-5497);
			18102: out = 16'(2170);
			18103: out = 16'(4949);
			18104: out = 16'(3097);
			18105: out = 16'(-1113);
			18106: out = 16'(-3622);
			18107: out = 16'(-4942);
			18108: out = 16'(-3321);
			18109: out = 16'(1366);
			18110: out = 16'(3827);
			18111: out = 16'(1522);
			18112: out = 16'(3706);
			18113: out = 16'(1437);
			18114: out = 16'(-4512);
			18115: out = 16'(-11023);
			18116: out = 16'(-3718);
			18117: out = 16'(-1474);
			18118: out = 16'(1946);
			18119: out = 16'(4633);
			18120: out = 16'(5516);
			18121: out = 16'(420);
			18122: out = 16'(-3820);
			18123: out = 16'(-4095);
			18124: out = 16'(-2747);
			18125: out = 16'(-3780);
			18126: out = 16'(-5347);
			18127: out = 16'(-1012);
			18128: out = 16'(6195);
			18129: out = 16'(6244);
			18130: out = 16'(-1498);
			18131: out = 16'(-6402);
			18132: out = 16'(-1698);
			18133: out = 16'(4918);
			18134: out = 16'(5179);
			18135: out = 16'(1664);
			18136: out = 16'(54);
			18137: out = 16'(1729);
			18138: out = 16'(1952);
			18139: out = 16'(-513);
			18140: out = 16'(-5877);
			18141: out = 16'(-9854);
			18142: out = 16'(-2891);
			18143: out = 16'(5831);
			18144: out = 16'(3571);
			18145: out = 16'(-8089);
			18146: out = 16'(-1641);
			18147: out = 16'(7497);
			18148: out = 16'(8351);
			18149: out = 16'(-2193);
			18150: out = 16'(-4616);
			18151: out = 16'(-6229);
			18152: out = 16'(-1291);
			18153: out = 16'(1958);
			18154: out = 16'(241);
			18155: out = 16'(1977);
			18156: out = 16'(3268);
			18157: out = 16'(359);
			18158: out = 16'(-2931);
			18159: out = 16'(-1442);
			18160: out = 16'(3070);
			18161: out = 16'(2180);
			18162: out = 16'(-2604);
			18163: out = 16'(-10050);
			18164: out = 16'(-3301);
			18165: out = 16'(4180);
			18166: out = 16'(3721);
			18167: out = 16'(4151);
			18168: out = 16'(4269);
			18169: out = 16'(150);
			18170: out = 16'(-8161);
			18171: out = 16'(-6218);
			18172: out = 16'(-4948);
			18173: out = 16'(629);
			18174: out = 16'(5036);
			18175: out = 16'(5793);
			18176: out = 16'(3057);
			18177: out = 16'(207);
			18178: out = 16'(-3317);
			18179: out = 16'(-10714);
			18180: out = 16'(-3956);
			18181: out = 16'(-1421);
			18182: out = 16'(2825);
			18183: out = 16'(5772);
			18184: out = 16'(6868);
			18185: out = 16'(-2928);
			18186: out = 16'(-5366);
			18187: out = 16'(591);
			18188: out = 16'(-117);
			18189: out = 16'(-7422);
			18190: out = 16'(-7709);
			18191: out = 16'(2141);
			18192: out = 16'(7173);
			18193: out = 16'(7040);
			18194: out = 16'(4673);
			18195: out = 16'(3640);
			18196: out = 16'(1703);
			18197: out = 16'(-2643);
			18198: out = 16'(-2146);
			18199: out = 16'(385);
			18200: out = 16'(-622);
			18201: out = 16'(-950);
			18202: out = 16'(574);
			18203: out = 16'(3280);
			18204: out = 16'(4103);
			18205: out = 16'(6663);
			18206: out = 16'(3460);
			18207: out = 16'(-1088);
			18208: out = 16'(-6009);
			18209: out = 16'(-9036);
			18210: out = 16'(-7002);
			18211: out = 16'(-3178);
			18212: out = 16'(-152);
			18213: out = 16'(2512);
			18214: out = 16'(5306);
			18215: out = 16'(5459);
			18216: out = 16'(2426);
			18217: out = 16'(-96);
			18218: out = 16'(-5382);
			18219: out = 16'(-2500);
			18220: out = 16'(574);
			18221: out = 16'(-128);
			18222: out = 16'(58);
			18223: out = 16'(1293);
			18224: out = 16'(2522);
			18225: out = 16'(1550);
			18226: out = 16'(226);
			18227: out = 16'(-1903);
			18228: out = 16'(-2020);
			18229: out = 16'(-880);
			18230: out = 16'(-157);
			18231: out = 16'(972);
			18232: out = 16'(1800);
			18233: out = 16'(1074);
			18234: out = 16'(-3809);
			18235: out = 16'(-26);
			18236: out = 16'(-2927);
			18237: out = 16'(-3145);
			18238: out = 16'(1960);
			18239: out = 16'(5522);
			18240: out = 16'(2521);
			18241: out = 16'(-1679);
			18242: out = 16'(-1188);
			18243: out = 16'(3587);
			18244: out = 16'(5691);
			18245: out = 16'(3779);
			18246: out = 16'(-1246);
			18247: out = 16'(-6596);
			18248: out = 16'(-3878);
			18249: out = 16'(-306);
			18250: out = 16'(-972);
			18251: out = 16'(-2650);
			18252: out = 16'(2305);
			18253: out = 16'(7892);
			18254: out = 16'(4518);
			18255: out = 16'(-5118);
			18256: out = 16'(-4902);
			18257: out = 16'(-682);
			18258: out = 16'(-1045);
			18259: out = 16'(-5299);
			18260: out = 16'(2028);
			18261: out = 16'(10220);
			18262: out = 16'(12685);
			18263: out = 16'(6379);
			18264: out = 16'(291);
			18265: out = 16'(-1042);
			18266: out = 16'(-1637);
			18267: out = 16'(-4895);
			18268: out = 16'(-3931);
			18269: out = 16'(-159);
			18270: out = 16'(5709);
			18271: out = 16'(3822);
			18272: out = 16'(-3201);
			18273: out = 16'(-10148);
			18274: out = 16'(-4542);
			18275: out = 16'(1526);
			18276: out = 16'(509);
			18277: out = 16'(1251);
			18278: out = 16'(2761);
			18279: out = 16'(2914);
			18280: out = 16'(-1702);
			18281: out = 16'(-1641);
			18282: out = 16'(-1703);
			18283: out = 16'(4309);
			18284: out = 16'(6036);
			18285: out = 16'(-435);
			18286: out = 16'(-8810);
			18287: out = 16'(-7004);
			18288: out = 16'(2767);
			18289: out = 16'(8919);
			18290: out = 16'(9391);
			18291: out = 16'(3437);
			18292: out = 16'(-4315);
			18293: out = 16'(-9351);
			18294: out = 16'(-5460);
			18295: out = 16'(-2850);
			18296: out = 16'(-3311);
			18297: out = 16'(-4042);
			18298: out = 16'(-43);
			18299: out = 16'(5657);
			18300: out = 16'(7559);
			18301: out = 16'(4098);
			18302: out = 16'(56);
			18303: out = 16'(-2289);
			18304: out = 16'(-3048);
			18305: out = 16'(-3829);
			18306: out = 16'(-3476);
			18307: out = 16'(-7461);
			18308: out = 16'(-3969);
			18309: out = 16'(4040);
			18310: out = 16'(8772);
			18311: out = 16'(3017);
			18312: out = 16'(-4567);
			18313: out = 16'(-9007);
			18314: out = 16'(-6763);
			18315: out = 16'(-2837);
			18316: out = 16'(-2301);
			18317: out = 16'(-3496);
			18318: out = 16'(-229);
			18319: out = 16'(3588);
			18320: out = 16'(8146);
			18321: out = 16'(1361);
			18322: out = 16'(-7675);
			18323: out = 16'(-9430);
			18324: out = 16'(1850);
			18325: out = 16'(4430);
			18326: out = 16'(1583);
			18327: out = 16'(3120);
			18328: out = 16'(5343);
			18329: out = 16'(4265);
			18330: out = 16'(586);
			18331: out = 16'(548);
			18332: out = 16'(-500);
			18333: out = 16'(670);
			18334: out = 16'(-3567);
			18335: out = 16'(-7680);
			18336: out = 16'(-3161);
			18337: out = 16'(2346);
			18338: out = 16'(5843);
			18339: out = 16'(4794);
			18340: out = 16'(65);
			18341: out = 16'(1779);
			18342: out = 16'(-180);
			18343: out = 16'(-6752);
			18344: out = 16'(-13429);
			18345: out = 16'(-1971);
			18346: out = 16'(5973);
			18347: out = 16'(7119);
			18348: out = 16'(3588);
			18349: out = 16'(2547);
			18350: out = 16'(1224);
			18351: out = 16'(805);
			18352: out = 16'(-802);
			18353: out = 16'(-1971);
			18354: out = 16'(-2719);
			18355: out = 16'(-875);
			18356: out = 16'(-782);
			18357: out = 16'(-2868);
			18358: out = 16'(-3078);
			18359: out = 16'(3485);
			18360: out = 16'(7341);
			18361: out = 16'(1483);
			18362: out = 16'(449);
			18363: out = 16'(-421);
			18364: out = 16'(-612);
			18365: out = 16'(-2387);
			18366: out = 16'(-259);
			18367: out = 16'(1407);
			18368: out = 16'(1685);
			18369: out = 16'(-96);
			18370: out = 16'(2271);
			18371: out = 16'(411);
			18372: out = 16'(-415);
			18373: out = 16'(544);
			18374: out = 16'(4028);
			18375: out = 16'(3923);
			18376: out = 16'(3039);
			18377: out = 16'(1088);
			18378: out = 16'(-549);
			18379: out = 16'(-6079);
			18380: out = 16'(-5815);
			18381: out = 16'(-811);
			18382: out = 16'(4025);
			18383: out = 16'(2271);
			18384: out = 16'(502);
			18385: out = 16'(-440);
			18386: out = 16'(60);
			18387: out = 16'(-404);
			18388: out = 16'(-41);
			18389: out = 16'(554);
			18390: out = 16'(2638);
			18391: out = 16'(3303);
			18392: out = 16'(573);
			18393: out = 16'(-5675);
			18394: out = 16'(-5502);
			18395: out = 16'(6162);
			18396: out = 16'(10752);
			18397: out = 16'(6229);
			18398: out = 16'(-3309);
			18399: out = 16'(-7781);
			18400: out = 16'(-5871);
			18401: out = 16'(-1585);
			18402: out = 16'(1130);
			18403: out = 16'(4287);
			18404: out = 16'(3301);
			18405: out = 16'(2997);
			18406: out = 16'(-908);
			18407: out = 16'(-4006);
			18408: out = 16'(-6195);
			18409: out = 16'(1588);
			18410: out = 16'(3576);
			18411: out = 16'(1141);
			18412: out = 16'(-164);
			18413: out = 16'(3200);
			18414: out = 16'(264);
			18415: out = 16'(-5033);
			18416: out = 16'(-4116);
			18417: out = 16'(-1406);
			18418: out = 16'(1471);
			18419: out = 16'(1909);
			18420: out = 16'(1745);
			18421: out = 16'(-25);
			18422: out = 16'(-435);
			18423: out = 16'(-403);
			18424: out = 16'(-464);
			18425: out = 16'(751);
			18426: out = 16'(-516);
			18427: out = 16'(1555);
			18428: out = 16'(3339);
			18429: out = 16'(-437);
			18430: out = 16'(-6484);
			18431: out = 16'(-6394);
			18432: out = 16'(-304);
			18433: out = 16'(1721);
			18434: out = 16'(7208);
			18435: out = 16'(4330);
			18436: out = 16'(377);
			18437: out = 16'(-1506);
			18438: out = 16'(-321);
			18439: out = 16'(-2220);
			18440: out = 16'(-4540);
			18441: out = 16'(-3987);
			18442: out = 16'(-490);
			18443: out = 16'(898);
			18444: out = 16'(151);
			18445: out = 16'(1011);
			18446: out = 16'(5422);
			18447: out = 16'(6131);
			18448: out = 16'(305);
			18449: out = 16'(-8788);
			18450: out = 16'(-12202);
			18451: out = 16'(-3433);
			18452: out = 16'(4801);
			18453: out = 16'(4042);
			18454: out = 16'(523);
			18455: out = 16'(4572);
			18456: out = 16'(6902);
			18457: out = 16'(854);
			18458: out = 16'(-6832);
			18459: out = 16'(-960);
			18460: out = 16'(6954);
			18461: out = 16'(5993);
			18462: out = 16'(-2196);
			18463: out = 16'(-3135);
			18464: out = 16'(-59);
			18465: out = 16'(2586);
			18466: out = 16'(807);
			18467: out = 16'(-246);
			18468: out = 16'(-2654);
			18469: out = 16'(-1411);
			18470: out = 16'(476);
			18471: out = 16'(1538);
			18472: out = 16'(-1939);
			18473: out = 16'(-3074);
			18474: out = 16'(-1599);
			18475: out = 16'(-208);
			18476: out = 16'(31);
			18477: out = 16'(-457);
			18478: out = 16'(224);
			18479: out = 16'(-1790);
			18480: out = 16'(-7164);
			18481: out = 16'(-10045);
			18482: out = 16'(-2182);
			18483: out = 16'(7618);
			18484: out = 16'(7036);
			18485: out = 16'(775);
			18486: out = 16'(-1744);
			18487: out = 16'(815);
			18488: out = 16'(1475);
			18489: out = 16'(-3431);
			18490: out = 16'(-2952);
			18491: out = 16'(3433);
			18492: out = 16'(7733);
			18493: out = 16'(1603);
			18494: out = 16'(-4081);
			18495: out = 16'(-4796);
			18496: out = 16'(1484);
			18497: out = 16'(5558);
			18498: out = 16'(7039);
			18499: out = 16'(854);
			18500: out = 16'(-3496);
			18501: out = 16'(-1056);
			18502: out = 16'(792);
			18503: out = 16'(-6452);
			18504: out = 16'(-9710);
			18505: out = 16'(2987);
			18506: out = 16'(10334);
			18507: out = 16'(6211);
			18508: out = 16'(-1395);
			18509: out = 16'(695);
			18510: out = 16'(4326);
			18511: out = 16'(2267);
			18512: out = 16'(-6036);
			18513: out = 16'(-9623);
			18514: out = 16'(-2488);
			18515: out = 16'(1684);
			18516: out = 16'(998);
			18517: out = 16'(226);
			18518: out = 16'(1753);
			18519: out = 16'(2143);
			18520: out = 16'(785);
			18521: out = 16'(-276);
			18522: out = 16'(-329);
			18523: out = 16'(3123);
			18524: out = 16'(2065);
			18525: out = 16'(-1736);
			18526: out = 16'(-3036);
			18527: out = 16'(2499);
			18528: out = 16'(3450);
			18529: out = 16'(-412);
			18530: out = 16'(-2093);
			18531: out = 16'(-1363);
			18532: out = 16'(4936);
			18533: out = 16'(3829);
			18534: out = 16'(-3595);
			18535: out = 16'(-11307);
			18536: out = 16'(-2573);
			18537: out = 16'(5232);
			18538: out = 16'(3957);
			18539: out = 16'(-1177);
			18540: out = 16'(-820);
			18541: out = 16'(-285);
			18542: out = 16'(-3645);
			18543: out = 16'(-8850);
			18544: out = 16'(-880);
			18545: out = 16'(4536);
			18546: out = 16'(5343);
			18547: out = 16'(3612);
			18548: out = 16'(3798);
			18549: out = 16'(1185);
			18550: out = 16'(-2491);
			18551: out = 16'(-4771);
			18552: out = 16'(-2572);
			18553: out = 16'(394);
			18554: out = 16'(4034);
			18555: out = 16'(5062);
			18556: out = 16'(1779);
			18557: out = 16'(-3357);
			18558: out = 16'(-4036);
			18559: out = 16'(362);
			18560: out = 16'(3309);
			18561: out = 16'(683);
			18562: out = 16'(-2785);
			18563: out = 16'(-3601);
			18564: out = 16'(-4033);
			18565: out = 16'(-7151);
			18566: out = 16'(-4985);
			18567: out = 16'(4176);
			18568: out = 16'(10801);
			18569: out = 16'(10448);
			18570: out = 16'(225);
			18571: out = 16'(-4042);
			18572: out = 16'(-869);
			18573: out = 16'(-534);
			18574: out = 16'(-4352);
			18575: out = 16'(-5246);
			18576: out = 16'(-615);
			18577: out = 16'(3514);
			18578: out = 16'(1493);
			18579: out = 16'(-146);
			18580: out = 16'(-116);
			18581: out = 16'(-256);
			18582: out = 16'(-375);
			18583: out = 16'(-229);
			18584: out = 16'(-200);
			18585: out = 16'(-357);
			18586: out = 16'(-4535);
			18587: out = 16'(-1985);
			18588: out = 16'(30);
			18589: out = 16'(-357);
			18590: out = 16'(-149);
			18591: out = 16'(2965);
			18592: out = 16'(2401);
			18593: out = 16'(-103);
			18594: out = 16'(4071);
			18595: out = 16'(2049);
			18596: out = 16'(627);
			18597: out = 16'(-803);
			18598: out = 16'(-179);
			18599: out = 16'(-344);
			18600: out = 16'(-3170);
			18601: out = 16'(-7390);
			18602: out = 16'(-5405);
			18603: out = 16'(5446);
			18604: out = 16'(9958);
			18605: out = 16'(5090);
			18606: out = 16'(-1272);
			18607: out = 16'(-3959);
			18608: out = 16'(-4950);
			18609: out = 16'(-7811);
			18610: out = 16'(-6019);
			18611: out = 16'(1284);
			18612: out = 16'(7002);
			18613: out = 16'(-653);
			18614: out = 16'(-7547);
			18615: out = 16'(1814);
			18616: out = 16'(8521);
			18617: out = 16'(5759);
			18618: out = 16'(-1870);
			18619: out = 16'(-1839);
			18620: out = 16'(-2243);
			18621: out = 16'(-382);
			18622: out = 16'(9);
			18623: out = 16'(2620);
			18624: out = 16'(3189);
			18625: out = 16'(2299);
			18626: out = 16'(-1325);
			18627: out = 16'(-2518);
			18628: out = 16'(-4119);
			18629: out = 16'(2488);
			18630: out = 16'(2221);
			18631: out = 16'(-757);
			18632: out = 16'(-173);
			18633: out = 16'(4452);
			18634: out = 16'(4164);
			18635: out = 16'(-967);
			18636: out = 16'(-6172);
			18637: out = 16'(-5201);
			18638: out = 16'(-2357);
			18639: out = 16'(1458);
			18640: out = 16'(3971);
			18641: out = 16'(5684);
			18642: out = 16'(2803);
			18643: out = 16'(1519);
			18644: out = 16'(569);
			18645: out = 16'(-5791);
			18646: out = 16'(-5844);
			18647: out = 16'(-2232);
			18648: out = 16'(-1393);
			18649: out = 16'(-8008);
			18650: out = 16'(-8498);
			18651: out = 16'(-2651);
			18652: out = 16'(3780);
			18653: out = 16'(4045);
			18654: out = 16'(8020);
			18655: out = 16'(8240);
			18656: out = 16'(4348);
			18657: out = 16'(-4342);
			18658: out = 16'(-14293);
			18659: out = 16'(-13008);
			18660: out = 16'(-3816);
			18661: out = 16'(3568);
			18662: out = 16'(9385);
			18663: out = 16'(5642);
			18664: out = 16'(1956);
			18665: out = 16'(-424);
			18666: out = 16'(-117);
			18667: out = 16'(-4758);
			18668: out = 16'(-5387);
			18669: out = 16'(-4474);
			18670: out = 16'(-5405);
			18671: out = 16'(-538);
			18672: out = 16'(1848);
			18673: out = 16'(2413);
			18674: out = 16'(2100);
			18675: out = 16'(-1795);
			18676: out = 16'(-978);
			18677: out = 16'(1151);
			18678: out = 16'(1805);
			18679: out = 16'(-4154);
			18680: out = 16'(-1357);
			18681: out = 16'(964);
			18682: out = 16'(1829);
			18683: out = 16'(4227);
			18684: out = 16'(4258);
			18685: out = 16'(3189);
			18686: out = 16'(919);
			18687: out = 16'(-3561);
			18688: out = 16'(-383);
			18689: out = 16'(869);
			18690: out = 16'(4260);
			18691: out = 16'(7061);
			18692: out = 16'(5904);
			18693: out = 16'(-5036);
			18694: out = 16'(-10139);
			18695: out = 16'(-2166);
			18696: out = 16'(6491);
			18697: out = 16'(4530);
			18698: out = 16'(897);
			18699: out = 16'(2939);
			18700: out = 16'(3201);
			18701: out = 16'(1474);
			18702: out = 16'(-1680);
			18703: out = 16'(-223);
			18704: out = 16'(1355);
			18705: out = 16'(2593);
			18706: out = 16'(-1112);
			18707: out = 16'(-946);
			18708: out = 16'(3543);
			18709: out = 16'(793);
			18710: out = 16'(-6818);
			18711: out = 16'(-9287);
			18712: out = 16'(-180);
			18713: out = 16'(7740);
			18714: out = 16'(6830);
			18715: out = 16'(-632);
			18716: out = 16'(-4157);
			18717: out = 16'(-685);
			18718: out = 16'(3246);
			18719: out = 16'(1957);
			18720: out = 16'(-782);
			18721: out = 16'(-306);
			18722: out = 16'(-4507);
			18723: out = 16'(-7359);
			18724: out = 16'(-4614);
			18725: out = 16'(2386);
			18726: out = 16'(7009);
			18727: out = 16'(3383);
			18728: out = 16'(-1449);
			18729: out = 16'(-1196);
			18730: out = 16'(-3712);
			18731: out = 16'(-4076);
			18732: out = 16'(-4638);
			18733: out = 16'(-2721);
			18734: out = 16'(-2733);
			18735: out = 16'(5835);
			18736: out = 16'(6953);
			18737: out = 16'(-1206);
			18738: out = 16'(-10426);
			18739: out = 16'(-873);
			18740: out = 16'(8649);
			18741: out = 16'(1152);
			18742: out = 16'(-18338);
			18743: out = 16'(-17886);
			18744: out = 16'(-2308);
			18745: out = 16'(8068);
			18746: out = 16'(5707);
			18747: out = 16'(988);
			18748: out = 16'(4105);
			18749: out = 16'(4549);
			18750: out = 16'(-2661);
			18751: out = 16'(-10434);
			18752: out = 16'(-1462);
			18753: out = 16'(8281);
			18754: out = 16'(6849);
			18755: out = 16'(711);
			18756: out = 16'(103);
			18757: out = 16'(2172);
			18758: out = 16'(883);
			18759: out = 16'(-4348);
			18760: out = 16'(-2669);
			18761: out = 16'(126);
			18762: out = 16'(4371);
			18763: out = 16'(7023);
			18764: out = 16'(1757);
			18765: out = 16'(-6835);
			18766: out = 16'(-8692);
			18767: out = 16'(-443);
			18768: out = 16'(6935);
			18769: out = 16'(3364);
			18770: out = 16'(-1404);
			18771: out = 16'(-631);
			18772: out = 16'(-1545);
			18773: out = 16'(-2432);
			18774: out = 16'(-1713);
			18775: out = 16'(4829);
			18776: out = 16'(9164);
			18777: out = 16'(4780);
			18778: out = 16'(-4397);
			18779: out = 16'(-7105);
			18780: out = 16'(-2244);
			18781: out = 16'(1888);
			18782: out = 16'(1737);
			18783: out = 16'(4105);
			18784: out = 16'(6957);
			18785: out = 16'(4919);
			18786: out = 16'(-7453);
			18787: out = 16'(-12114);
			18788: out = 16'(-1594);
			18789: out = 16'(7191);
			18790: out = 16'(4890);
			18791: out = 16'(-371);
			18792: out = 16'(1546);
			18793: out = 16'(6504);
			18794: out = 16'(3754);
			18795: out = 16'(-2308);
			18796: out = 16'(-4003);
			18797: out = 16'(-434);
			18798: out = 16'(35);
			18799: out = 16'(-1593);
			18800: out = 16'(-2019);
			18801: out = 16'(483);
			18802: out = 16'(4881);
			18803: out = 16'(2582);
			18804: out = 16'(-2622);
			18805: out = 16'(-4209);
			18806: out = 16'(-4033);
			18807: out = 16'(794);
			18808: out = 16'(1304);
			18809: out = 16'(-106);
			18810: out = 16'(-282);
			18811: out = 16'(5590);
			18812: out = 16'(6251);
			18813: out = 16'(1219);
			18814: out = 16'(-5726);
			18815: out = 16'(-1185);
			18816: out = 16'(-2553);
			18817: out = 16'(-6756);
			18818: out = 16'(-4551);
			18819: out = 16'(439);
			18820: out = 16'(6047);
			18821: out = 16'(6851);
			18822: out = 16'(4741);
			18823: out = 16'(-2059);
			18824: out = 16'(-1446);
			18825: out = 16'(75);
			18826: out = 16'(-1702);
			18827: out = 16'(-11072);
			18828: out = 16'(-6962);
			18829: out = 16'(-804);
			18830: out = 16'(3378);
			18831: out = 16'(7462);
			18832: out = 16'(7282);
			18833: out = 16'(3833);
			18834: out = 16'(-3150);
			18835: out = 16'(-7671);
			18836: out = 16'(-12765);
			18837: out = 16'(-6744);
			18838: out = 16'(168);
			18839: out = 16'(2636);
			18840: out = 16'(5462);
			18841: out = 16'(8887);
			18842: out = 16'(8077);
			18843: out = 16'(1209);
			18844: out = 16'(-11641);
			18845: out = 16'(-9486);
			18846: out = 16'(-2771);
			18847: out = 16'(117);
			18848: out = 16'(-2016);
			18849: out = 16'(-236);
			18850: out = 16'(1315);
			18851: out = 16'(2941);
			18852: out = 16'(4032);
			18853: out = 16'(7218);
			18854: out = 16'(3447);
			18855: out = 16'(-3161);
			18856: out = 16'(-7777);
			18857: out = 16'(-5791);
			18858: out = 16'(-2400);
			18859: out = 16'(2880);
			18860: out = 16'(5172);
			18861: out = 16'(833);
			18862: out = 16'(-3096);
			18863: out = 16'(1226);
			18864: out = 16'(7831);
			18865: out = 16'(3396);
			18866: out = 16'(-6376);
			18867: out = 16'(-10827);
			18868: out = 16'(-4516);
			18869: out = 16'(698);
			18870: out = 16'(1199);
			18871: out = 16'(480);
			18872: out = 16'(4708);
			18873: out = 16'(6329);
			18874: out = 16'(17);
			18875: out = 16'(-9107);
			18876: out = 16'(-7522);
			18877: out = 16'(1999);
			18878: out = 16'(2324);
			18879: out = 16'(532);
			18880: out = 16'(2374);
			18881: out = 16'(6101);
			18882: out = 16'(3987);
			18883: out = 16'(-2327);
			18884: out = 16'(-3025);
			18885: out = 16'(1011);
			18886: out = 16'(-343);
			18887: out = 16'(-2198);
			18888: out = 16'(-2111);
			18889: out = 16'(2628);
			18890: out = 16'(6514);
			18891: out = 16'(5356);
			18892: out = 16'(681);
			18893: out = 16'(-4754);
			18894: out = 16'(-7302);
			18895: out = 16'(-3935);
			18896: out = 16'(838);
			18897: out = 16'(2041);
			18898: out = 16'(650);
			18899: out = 16'(-1126);
			18900: out = 16'(1487);
			18901: out = 16'(2083);
			18902: out = 16'(2962);
			18903: out = 16'(5353);
			18904: out = 16'(7775);
			18905: out = 16'(-776);
			18906: out = 16'(-11695);
			18907: out = 16'(-11320);
			18908: out = 16'(-627);
			18909: out = 16'(4692);
			18910: out = 16'(2912);
			18911: out = 16'(2460);
			18912: out = 16'(648);
			18913: out = 16'(-1264);
			18914: out = 16'(-4650);
			18915: out = 16'(-2808);
			18916: out = 16'(1183);
			18917: out = 16'(6024);
			18918: out = 16'(1375);
			18919: out = 16'(-4790);
			18920: out = 16'(-2976);
			18921: out = 16'(5395);
			18922: out = 16'(5024);
			18923: out = 16'(-3297);
			18924: out = 16'(-9000);
			18925: out = 16'(2614);
			18926: out = 16'(9434);
			18927: out = 16'(6079);
			18928: out = 16'(-1069);
			18929: out = 16'(-9125);
			18930: out = 16'(-9233);
			18931: out = 16'(-5355);
			18932: out = 16'(-1180);
			18933: out = 16'(2132);
			18934: out = 16'(8843);
			18935: out = 16'(12232);
			18936: out = 16'(6667);
			18937: out = 16'(-3463);
			18938: out = 16'(-8358);
			18939: out = 16'(-1914);
			18940: out = 16'(3997);
			18941: out = 16'(-644);
			18942: out = 16'(-6401);
			18943: out = 16'(-4365);
			18944: out = 16'(1808);
			18945: out = 16'(1578);
			18946: out = 16'(832);
			18947: out = 16'(3367);
			18948: out = 16'(9585);
			18949: out = 16'(9388);
			18950: out = 16'(-881);
			18951: out = 16'(-7366);
			18952: out = 16'(-4782);
			18953: out = 16'(463);
			18954: out = 16'(-162);
			18955: out = 16'(-2710);
			18956: out = 16'(-1114);
			18957: out = 16'(2763);
			18958: out = 16'(1641);
			18959: out = 16'(516);
			18960: out = 16'(-522);
			18961: out = 16'(777);
			18962: out = 16'(1672);
			18963: out = 16'(271);
			18964: out = 16'(-720);
			18965: out = 16'(738);
			18966: out = 16'(1640);
			18967: out = 16'(386);
			18968: out = 16'(-2533);
			18969: out = 16'(-2336);
			18970: out = 16'(596);
			18971: out = 16'(1759);
			18972: out = 16'(531);
			18973: out = 16'(-486);
			18974: out = 16'(560);
			18975: out = 16'(1670);
			18976: out = 16'(-212);
			18977: out = 16'(-3781);
			18978: out = 16'(-5121);
			18979: out = 16'(-1832);
			18980: out = 16'(-349);
			18981: out = 16'(1455);
			18982: out = 16'(2663);
			18983: out = 16'(4096);
			18984: out = 16'(3699);
			18985: out = 16'(1803);
			18986: out = 16'(-2288);
			18987: out = 16'(-4067);
			18988: out = 16'(-2878);
			18989: out = 16'(2590);
			18990: out = 16'(2484);
			18991: out = 16'(-881);
			18992: out = 16'(-2342);
			18993: out = 16'(1360);
			18994: out = 16'(-1187);
			18995: out = 16'(-6064);
			18996: out = 16'(-2241);
			18997: out = 16'(7212);
			18998: out = 16'(9999);
			18999: out = 16'(3382);
			19000: out = 16'(-3251);
			19001: out = 16'(-3080);
			19002: out = 16'(-19);
			19003: out = 16'(-286);
			19004: out = 16'(-2469);
			19005: out = 16'(-2420);
			19006: out = 16'(-812);
			19007: out = 16'(-92);
			19008: out = 16'(-244);
			19009: out = 16'(-1160);
			19010: out = 16'(6271);
			19011: out = 16'(10081);
			19012: out = 16'(5632);
			19013: out = 16'(-5830);
			19014: out = 16'(-9448);
			19015: out = 16'(-10758);
			19016: out = 16'(-7939);
			19017: out = 16'(-21);
			19018: out = 16'(8226);
			19019: out = 16'(12507);
			19020: out = 16'(10460);
			19021: out = 16'(4000);
			19022: out = 16'(-3572);
			19023: out = 16'(-4977);
			19024: out = 16'(-1043);
			19025: out = 16'(1026);
			19026: out = 16'(-4130);
			19027: out = 16'(-5325);
			19028: out = 16'(-800);
			19029: out = 16'(4577);
			19030: out = 16'(4421);
			19031: out = 16'(3839);
			19032: out = 16'(3951);
			19033: out = 16'(3708);
			19034: out = 16'(-203);
			19035: out = 16'(-6520);
			19036: out = 16'(-9030);
			19037: out = 16'(-6137);
			19038: out = 16'(-2133);
			19039: out = 16'(-234);
			19040: out = 16'(3365);
			19041: out = 16'(6802);
			19042: out = 16'(4500);
			19043: out = 16'(-5610);
			19044: out = 16'(-7518);
			19045: out = 16'(-339);
			19046: out = 16'(5300);
			19047: out = 16'(-293);
			19048: out = 16'(-588);
			19049: out = 16'(2740);
			19050: out = 16'(4815);
			19051: out = 16'(-1080);
			19052: out = 16'(-3804);
			19053: out = 16'(-4699);
			19054: out = 16'(-2825);
			19055: out = 16'(-2783);
			19056: out = 16'(-2997);
			19057: out = 16'(-2668);
			19058: out = 16'(1001);
			19059: out = 16'(3894);
			19060: out = 16'(4053);
			19061: out = 16'(1460);
			19062: out = 16'(453);
			19063: out = 16'(-1354);
			19064: out = 16'(-7351);
			19065: out = 16'(-12841);
			19066: out = 16'(-9392);
			19067: out = 16'(1426);
			19068: out = 16'(6214);
			19069: out = 16'(6858);
			19070: out = 16'(4224);
			19071: out = 16'(4627);
			19072: out = 16'(3880);
			19073: out = 16'(1347);
			19074: out = 16'(-9669);
			19075: out = 16'(-15231);
			19076: out = 16'(-7687);
			19077: out = 16'(4420);
			19078: out = 16'(5952);
			19079: out = 16'(1894);
			19080: out = 16'(1049);
			19081: out = 16'(6416);
			19082: out = 16'(5153);
			19083: out = 16'(1382);
			19084: out = 16'(-2139);
			19085: out = 16'(-4288);
			19086: out = 16'(-3699);
			19087: out = 16'(-1553);
			19088: out = 16'(712);
			19089: out = 16'(2645);
			19090: out = 16'(8718);
			19091: out = 16'(9633);
			19092: out = 16'(5009);
			19093: out = 16'(-687);
			19094: out = 16'(-3522);
			19095: out = 16'(-2257);
			19096: out = 16'(-1400);
			19097: out = 16'(-1506);
			19098: out = 16'(-3631);
			19099: out = 16'(1921);
			19100: out = 16'(3606);
			19101: out = 16'(372);
			19102: out = 16'(-5546);
			19103: out = 16'(270);
			19104: out = 16'(1555);
			19105: out = 16'(-781);
			19106: out = 16'(-1074);
			19107: out = 16'(1425);
			19108: out = 16'(963);
			19109: out = 16'(91);
			19110: out = 16'(2352);
			19111: out = 16'(5082);
			19112: out = 16'(2279);
			19113: out = 16'(-2545);
			19114: out = 16'(-4334);
			19115: out = 16'(-682);
			19116: out = 16'(1068);
			19117: out = 16'(4168);
			19118: out = 16'(7238);
			19119: out = 16'(4972);
			19120: out = 16'(265);
			19121: out = 16'(-4865);
			19122: out = 16'(-8101);
			19123: out = 16'(-10236);
			19124: out = 16'(-5943);
			19125: out = 16'(471);
			19126: out = 16'(5179);
			19127: out = 16'(5385);
			19128: out = 16'(5779);
			19129: out = 16'(1963);
			19130: out = 16'(-2559);
			19131: out = 16'(-4239);
			19132: out = 16'(-956);
			19133: out = 16'(2822);
			19134: out = 16'(2419);
			19135: out = 16'(-893);
			19136: out = 16'(-1154);
			19137: out = 16'(-715);
			19138: out = 16'(971);
			19139: out = 16'(1517);
			19140: out = 16'(-270);
			19141: out = 16'(-252);
			19142: out = 16'(-981);
			19143: out = 16'(-1957);
			19144: out = 16'(-3711);
			19145: out = 16'(-4238);
			19146: out = 16'(-1372);
			19147: out = 16'(6118);
			19148: out = 16'(10056);
			19149: out = 16'(995);
			19150: out = 16'(-7855);
			19151: out = 16'(-8505);
			19152: out = 16'(-2550);
			19153: out = 16'(-2421);
			19154: out = 16'(-773);
			19155: out = 16'(4584);
			19156: out = 16'(10339);
			19157: out = 16'(6410);
			19158: out = 16'(1825);
			19159: out = 16'(-3166);
			19160: out = 16'(-5804);
			19161: out = 16'(-10406);
			19162: out = 16'(-2395);
			19163: out = 16'(815);
			19164: out = 16'(3007);
			19165: out = 16'(3805);
			19166: out = 16'(7428);
			19167: out = 16'(343);
			19168: out = 16'(-4331);
			19169: out = 16'(-1339);
			19170: out = 16'(1287);
			19171: out = 16'(-2703);
			19172: out = 16'(-7491);
			19173: out = 16'(-4462);
			19174: out = 16'(1309);
			19175: out = 16'(5889);
			19176: out = 16'(2575);
			19177: out = 16'(628);
			19178: out = 16'(3613);
			19179: out = 16'(4380);
			19180: out = 16'(-2715);
			19181: out = 16'(-8430);
			19182: out = 16'(-4602);
			19183: out = 16'(-101);
			19184: out = 16'(-466);
			19185: out = 16'(-2234);
			19186: out = 16'(1542);
			19187: out = 16'(5639);
			19188: out = 16'(6242);
			19189: out = 16'(1001);
			19190: out = 16'(-4118);
			19191: out = 16'(-5589);
			19192: out = 16'(-3197);
			19193: out = 16'(-1087);
			19194: out = 16'(125);
			19195: out = 16'(303);
			19196: out = 16'(7470);
			19197: out = 16'(7322);
			19198: out = 16'(-544);
			19199: out = 16'(-9821);
			19200: out = 16'(-2017);
			19201: out = 16'(2124);
			19202: out = 16'(709);
			19203: out = 16'(-758);
			19204: out = 16'(1353);
			19205: out = 16'(4995);
			19206: out = 16'(3574);
			19207: out = 16'(-908);
			19208: out = 16'(-3230);
			19209: out = 16'(2854);
			19210: out = 16'(6605);
			19211: out = 16'(3040);
			19212: out = 16'(-5501);
			19213: out = 16'(-2853);
			19214: out = 16'(-298);
			19215: out = 16'(-1364);
			19216: out = 16'(-3139);
			19217: out = 16'(806);
			19218: out = 16'(4022);
			19219: out = 16'(3355);
			19220: out = 16'(-786);
			19221: out = 16'(-3069);
			19222: out = 16'(-2697);
			19223: out = 16'(-530);
			19224: out = 16'(-798);
			19225: out = 16'(103);
			19226: out = 16'(464);
			19227: out = 16'(4892);
			19228: out = 16'(6032);
			19229: out = 16'(2162);
			19230: out = 16'(-5833);
			19231: out = 16'(-2249);
			19232: out = 16'(4389);
			19233: out = 16'(696);
			19234: out = 16'(-12047);
			19235: out = 16'(-12328);
			19236: out = 16'(-741);
			19237: out = 16'(2889);
			19238: out = 16'(1643);
			19239: out = 16'(-331);
			19240: out = 16'(7114);
			19241: out = 16'(11190);
			19242: out = 16'(3443);
			19243: out = 16'(-14089);
			19244: out = 16'(-16627);
			19245: out = 16'(-779);
			19246: out = 16'(624);
			19247: out = 16'(3657);
			19248: out = 16'(-6);
			19249: out = 16'(2555);
			19250: out = 16'(6440);
			19251: out = 16'(8253);
			19252: out = 16'(-3154);
			19253: out = 16'(-8952);
			19254: out = 16'(691);
			19255: out = 16'(3497);
			19256: out = 16'(-182);
			19257: out = 16'(-2690);
			19258: out = 16'(3636);
			19259: out = 16'(8665);
			19260: out = 16'(7109);
			19261: out = 16'(1075);
			19262: out = 16'(-3190);
			19263: out = 16'(-5728);
			19264: out = 16'(-7493);
			19265: out = 16'(-5930);
			19266: out = 16'(-374);
			19267: out = 16'(3614);
			19268: out = 16'(4191);
			19269: out = 16'(2700);
			19270: out = 16'(1358);
			19271: out = 16'(-253);
			19272: out = 16'(-142);
			19273: out = 16'(-183);
			19274: out = 16'(-756);
			19275: out = 16'(-2543);
			19276: out = 16'(-423);
			19277: out = 16'(-174);
			19278: out = 16'(-82);
			19279: out = 16'(31);
			19280: out = 16'(3744);
			19281: out = 16'(1044);
			19282: out = 16'(-1375);
			19283: out = 16'(-2492);
			19284: out = 16'(-1192);
			19285: out = 16'(-2396);
			19286: out = 16'(-266);
			19287: out = 16'(2807);
			19288: out = 16'(3822);
			19289: out = 16'(6675);
			19290: out = 16'(4751);
			19291: out = 16'(-1777);
			19292: out = 16'(-7830);
			19293: out = 16'(-6544);
			19294: out = 16'(-1644);
			19295: out = 16'(-866);
			19296: out = 16'(-3651);
			19297: out = 16'(-5553);
			19298: out = 16'(2924);
			19299: out = 16'(6977);
			19300: out = 16'(1033);
			19301: out = 16'(-9225);
			19302: out = 16'(-3550);
			19303: out = 16'(2615);
			19304: out = 16'(-53);
			19305: out = 16'(-4799);
			19306: out = 16'(-7177);
			19307: out = 16'(-1418);
			19308: out = 16'(3033);
			19309: out = 16'(1845);
			19310: out = 16'(-2269);
			19311: out = 16'(-3350);
			19312: out = 16'(-2568);
			19313: out = 16'(-1593);
			19314: out = 16'(277);
			19315: out = 16'(1931);
			19316: out = 16'(2484);
			19317: out = 16'(2650);
			19318: out = 16'(4021);
			19319: out = 16'(2990);
			19320: out = 16'(448);
			19321: out = 16'(-846);
			19322: out = 16'(895);
			19323: out = 16'(553);
			19324: out = 16'(-264);
			19325: out = 16'(767);
			19326: out = 16'(2166);
			19327: out = 16'(7140);
			19328: out = 16'(3055);
			19329: out = 16'(-1649);
			19330: out = 16'(-2357);
			19331: out = 16'(-2188);
			19332: out = 16'(-4755);
			19333: out = 16'(-2490);
			19334: out = 16'(5584);
			19335: out = 16'(7537);
			19336: out = 16'(6709);
			19337: out = 16'(4539);
			19338: out = 16'(4263);
			19339: out = 16'(1201);
			19340: out = 16'(-1430);
			19341: out = 16'(-3482);
			19342: out = 16'(-1494);
			19343: out = 16'(60);
			19344: out = 16'(65);
			19345: out = 16'(857);
			19346: out = 16'(7283);
			19347: out = 16'(11116);
			19348: out = 16'(3366);
			19349: out = 16'(-9527);
			19350: out = 16'(-13452);
			19351: out = 16'(-5235);
			19352: out = 16'(997);
			19353: out = 16'(588);
			19354: out = 16'(1556);
			19355: out = 16'(6517);
			19356: out = 16'(6296);
			19357: out = 16'(1783);
			19358: out = 16'(-2990);
			19359: out = 16'(-3989);
			19360: out = 16'(-6376);
			19361: out = 16'(-3717);
			19362: out = 16'(-3359);
			19363: out = 16'(-946);
			19364: out = 16'(2025);
			19365: out = 16'(6146);
			19366: out = 16'(3553);
			19367: out = 16'(576);
			19368: out = 16'(-986);
			19369: out = 16'(-3374);
			19370: out = 16'(-6751);
			19371: out = 16'(-7932);
			19372: out = 16'(-5973);
			19373: out = 16'(-2253);
			19374: out = 16'(-598);
			19375: out = 16'(3406);
			19376: out = 16'(6793);
			19377: out = 16'(3327);
			19378: out = 16'(15);
			19379: out = 16'(-3032);
			19380: out = 16'(-3259);
			19381: out = 16'(-3505);
			19382: out = 16'(-1147);
			19383: out = 16'(-805);
			19384: out = 16'(3138);
			19385: out = 16'(9726);
			19386: out = 16'(10831);
			19387: out = 16'(975);
			19388: out = 16'(-12807);
			19389: out = 16'(-17133);
			19390: out = 16'(-5736);
			19391: out = 16'(473);
			19392: out = 16'(-4830);
			19393: out = 16'(-10360);
			19394: out = 16'(-1288);
			19395: out = 16'(6570);
			19396: out = 16'(8435);
			19397: out = 16'(3911);
			19398: out = 16'(176);
			19399: out = 16'(-6501);
			19400: out = 16'(-6156);
			19401: out = 16'(-1173);
			19402: out = 16'(3575);
			19403: out = 16'(2753);
			19404: out = 16'(946);
			19405: out = 16'(1760);
			19406: out = 16'(4216);
			19407: out = 16'(221);
			19408: out = 16'(1517);
			19409: out = 16'(3462);
			19410: out = 16'(2984);
			19411: out = 16'(-2963);
			19412: out = 16'(-5897);
			19413: out = 16'(-3594);
			19414: out = 16'(2568);
			19415: out = 16'(5629);
			19416: out = 16'(5515);
			19417: out = 16'(4550);
			19418: out = 16'(5014);
			19419: out = 16'(2702);
			19420: out = 16'(-5642);
			19421: out = 16'(-7945);
			19422: out = 16'(-249);
			19423: out = 16'(6423);
			19424: out = 16'(4754);
			19425: out = 16'(-1136);
			19426: out = 16'(1098);
			19427: out = 16'(7451);
			19428: out = 16'(9531);
			19429: out = 16'(-2715);
			19430: out = 16'(-6557);
			19431: out = 16'(90);
			19432: out = 16'(4948);
			19433: out = 16'(-1473);
			19434: out = 16'(-2914);
			19435: out = 16'(1017);
			19436: out = 16'(1232);
			19437: out = 16'(-1556);
			19438: out = 16'(-1731);
			19439: out = 16'(1546);
			19440: out = 16'(3417);
			19441: out = 16'(1974);
			19442: out = 16'(298);
			19443: out = 16'(-1882);
			19444: out = 16'(-3525);
			19445: out = 16'(-1598);
			19446: out = 16'(2259);
			19447: out = 16'(4033);
			19448: out = 16'(2759);
			19449: out = 16'(-606);
			19450: out = 16'(-370);
			19451: out = 16'(-2722);
			19452: out = 16'(-4242);
			19453: out = 16'(44);
			19454: out = 16'(4439);
			19455: out = 16'(2958);
			19456: out = 16'(-2783);
			19457: out = 16'(-5147);
			19458: out = 16'(-1240);
			19459: out = 16'(1697);
			19460: out = 16'(917);
			19461: out = 16'(-532);
			19462: out = 16'(-2401);
			19463: out = 16'(-4910);
			19464: out = 16'(-7084);
			19465: out = 16'(-2868);
			19466: out = 16'(4701);
			19467: out = 16'(9602);
			19468: out = 16'(4205);
			19469: out = 16'(-2686);
			19470: out = 16'(-4348);
			19471: out = 16'(1033);
			19472: out = 16'(-2216);
			19473: out = 16'(-7103);
			19474: out = 16'(-3132);
			19475: out = 16'(4855);
			19476: out = 16'(4048);
			19477: out = 16'(-532);
			19478: out = 16'(647);
			19479: out = 16'(-647);
			19480: out = 16'(-745);
			19481: out = 16'(-4579);
			19482: out = 16'(-5621);
			19483: out = 16'(-2756);
			19484: out = 16'(794);
			19485: out = 16'(-2364);
			19486: out = 16'(-6127);
			19487: out = 16'(-517);
			19488: out = 16'(6010);
			19489: out = 16'(9126);
			19490: out = 16'(5479);
			19491: out = 16'(-454);
			19492: out = 16'(-5018);
			19493: out = 16'(-3386);
			19494: out = 16'(-328);
			19495: out = 16'(-22);
			19496: out = 16'(1871);
			19497: out = 16'(3465);
			19498: out = 16'(4833);
			19499: out = 16'(2126);
			19500: out = 16'(-3527);
			19501: out = 16'(-8499);
			19502: out = 16'(-3799);
			19503: out = 16'(5943);
			19504: out = 16'(7851);
			19505: out = 16'(2407);
			19506: out = 16'(-4659);
			19507: out = 16'(-5404);
			19508: out = 16'(-224);
			19509: out = 16'(36);
			19510: out = 16'(786);
			19511: out = 16'(2790);
			19512: out = 16'(3145);
			19513: out = 16'(514);
			19514: out = 16'(248);
			19515: out = 16'(3956);
			19516: out = 16'(5269);
			19517: out = 16'(2334);
			19518: out = 16'(-4213);
			19519: out = 16'(-3901);
			19520: out = 16'(106);
			19521: out = 16'(-474);
			19522: out = 16'(-4787);
			19523: out = 16'(-1810);
			19524: out = 16'(5024);
			19525: out = 16'(3543);
			19526: out = 16'(121);
			19527: out = 16'(-3958);
			19528: out = 16'(-3968);
			19529: out = 16'(-2292);
			19530: out = 16'(-289);
			19531: out = 16'(-36);
			19532: out = 16'(-183);
			19533: out = 16'(145);
			19534: out = 16'(1551);
			19535: out = 16'(4820);
			19536: out = 16'(6806);
			19537: out = 16'(5925);
			19538: out = 16'(1333);
			19539: out = 16'(-5068);
			19540: out = 16'(-11989);
			19541: out = 16'(-11307);
			19542: out = 16'(-128);
			19543: out = 16'(2100);
			19544: out = 16'(-995);
			19545: out = 16'(-2371);
			19546: out = 16'(2320);
			19547: out = 16'(3724);
			19548: out = 16'(-2528);
			19549: out = 16'(-8638);
			19550: out = 16'(-3321);
			19551: out = 16'(2236);
			19552: out = 16'(8027);
			19553: out = 16'(4665);
			19554: out = 16'(-486);
			19555: out = 16'(-1471);
			19556: out = 16'(-738);
			19557: out = 16'(-4754);
			19558: out = 16'(-7815);
			19559: out = 16'(198);
			19560: out = 16'(269);
			19561: out = 16'(-917);
			19562: out = 16'(-1351);
			19563: out = 16'(2571);
			19564: out = 16'(1939);
			19565: out = 16'(1662);
			19566: out = 16'(360);
			19567: out = 16'(353);
			19568: out = 16'(-236);
			19569: out = 16'(643);
			19570: out = 16'(-3355);
			19571: out = 16'(-10204);
			19572: out = 16'(-5881);
			19573: out = 16'(3450);
			19574: out = 16'(13096);
			19575: out = 16'(11965);
			19576: out = 16'(5165);
			19577: out = 16'(-9289);
			19578: out = 16'(-10091);
			19579: out = 16'(-3313);
			19580: out = 16'(-13);
			19581: out = 16'(-1216);
			19582: out = 16'(6901);
			19583: out = 16'(14516);
			19584: out = 16'(10384);
			19585: out = 16'(1705);
			19586: out = 16'(-4644);
			19587: out = 16'(-5647);
			19588: out = 16'(-5611);
			19589: out = 16'(-4299);
			19590: out = 16'(-3004);
			19591: out = 16'(-1449);
			19592: out = 16'(-938);
			19593: out = 16'(422);
			19594: out = 16'(6593);
			19595: out = 16'(9454);
			19596: out = 16'(5359);
			19597: out = 16'(-150);
			19598: out = 16'(-3563);
			19599: out = 16'(-1575);
			19600: out = 16'(-1398);
			19601: out = 16'(-4440);
			19602: out = 16'(-2818);
			19603: out = 16'(1646);
			19604: out = 16'(3617);
			19605: out = 16'(1272);
			19606: out = 16'(141);
			19607: out = 16'(-859);
			19608: out = 16'(-3028);
			19609: out = 16'(-5007);
			19610: out = 16'(1024);
			19611: out = 16'(1671);
			19612: out = 16'(1201);
			19613: out = 16'(-136);
			19614: out = 16'(2156);
			19615: out = 16'(14);
			19616: out = 16'(41);
			19617: out = 16'(-332);
			19618: out = 16'(-214);
			19619: out = 16'(-5074);
			19620: out = 16'(-2424);
			19621: out = 16'(1234);
			19622: out = 16'(1747);
			19623: out = 16'(35);
			19624: out = 16'(298);
			19625: out = 16'(1322);
			19626: out = 16'(1880);
			19627: out = 16'(-227);
			19628: out = 16'(412);
			19629: out = 16'(-2974);
			19630: out = 16'(-5839);
			19631: out = 16'(1108);
			19632: out = 16'(3179);
			19633: out = 16'(3191);
			19634: out = 16'(1524);
			19635: out = 16'(1662);
			19636: out = 16'(-7809);
			19637: out = 16'(-10955);
			19638: out = 16'(-6512);
			19639: out = 16'(824);
			19640: out = 16'(3083);
			19641: out = 16'(42);
			19642: out = 16'(-1225);
			19643: out = 16'(3559);
			19644: out = 16'(6578);
			19645: out = 16'(4381);
			19646: out = 16'(33);
			19647: out = 16'(1118);
			19648: out = 16'(2787);
			19649: out = 16'(-748);
			19650: out = 16'(-12841);
			19651: out = 16'(-15908);
			19652: out = 16'(2985);
			19653: out = 16'(8960);
			19654: out = 16'(4712);
			19655: out = 16'(-3259);
			19656: out = 16'(-3122);
			19657: out = 16'(-1020);
			19658: out = 16'(1430);
			19659: out = 16'(292);
			19660: out = 16'(910);
			19661: out = 16'(4206);
			19662: out = 16'(6588);
			19663: out = 16'(4612);
			19664: out = 16'(1355);
			19665: out = 16'(-1097);
			19666: out = 16'(3681);
			19667: out = 16'(5460);
			19668: out = 16'(1415);
			19669: out = 16'(-5006);
			19670: out = 16'(1195);
			19671: out = 16'(6165);
			19672: out = 16'(3643);
			19673: out = 16'(-2364);
			19674: out = 16'(-1183);
			19675: out = 16'(4910);
			19676: out = 16'(5944);
			19677: out = 16'(-2109);
			19678: out = 16'(-8744);
			19679: out = 16'(-5241);
			19680: out = 16'(5361);
			19681: out = 16'(7716);
			19682: out = 16'(2762);
			19683: out = 16'(-7903);
			19684: out = 16'(-6631);
			19685: out = 16'(626);
			19686: out = 16'(-509);
			19687: out = 16'(-5195);
			19688: out = 16'(-4225);
			19689: out = 16'(2332);
			19690: out = 16'(5116);
			19691: out = 16'(7050);
			19692: out = 16'(4153);
			19693: out = 16'(-1523);
			19694: out = 16'(-7853);
			19695: out = 16'(-4089);
			19696: out = 16'(-1051);
			19697: out = 16'(-1919);
			19698: out = 16'(-5551);
			19699: out = 16'(-1248);
			19700: out = 16'(-1764);
			19701: out = 16'(-3197);
			19702: out = 16'(-3360);
			19703: out = 16'(2116);
			19704: out = 16'(738);
			19705: out = 16'(-541);
			19706: out = 16'(-757);
			19707: out = 16'(188);
			19708: out = 16'(114);
			19709: out = 16'(272);
			19710: out = 16'(1618);
			19711: out = 16'(1707);
			19712: out = 16'(871);
			19713: out = 16'(-3640);
			19714: out = 16'(-3767);
			19715: out = 16'(698);
			19716: out = 16'(177);
			19717: out = 16'(-3255);
			19718: out = 16'(-4739);
			19719: out = 16'(421);
			19720: out = 16'(8400);
			19721: out = 16'(4617);
			19722: out = 16'(-2118);
			19723: out = 16'(-4465);
			19724: out = 16'(293);
			19725: out = 16'(-3956);
			19726: out = 16'(-5211);
			19727: out = 16'(-1157);
			19728: out = 16'(6167);
			19729: out = 16'(2507);
			19730: out = 16'(2239);
			19731: out = 16'(1495);
			19732: out = 16'(-284);
			19733: out = 16'(-2937);
			19734: out = 16'(-857);
			19735: out = 16'(512);
			19736: out = 16'(31);
			19737: out = 16'(261);
			19738: out = 16'(4357);
			19739: out = 16'(4721);
			19740: out = 16'(778);
			19741: out = 16'(-714);
			19742: out = 16'(-1501);
			19743: out = 16'(-218);
			19744: out = 16'(461);
			19745: out = 16'(2078);
			19746: out = 16'(-3433);
			19747: out = 16'(-3830);
			19748: out = 16'(-2394);
			19749: out = 16'(-265);
			19750: out = 16'(4962);
			19751: out = 16'(8650);
			19752: out = 16'(8650);
			19753: out = 16'(5218);
			19754: out = 16'(2099);
			19755: out = 16'(-2900);
			19756: out = 16'(-4476);
			19757: out = 16'(-1052);
			19758: out = 16'(1270);
			19759: out = 16'(5811);
			19760: out = 16'(3019);
			19761: out = 16'(-948);
			19762: out = 16'(-295);
			19763: out = 16'(1331);
			19764: out = 16'(532);
			19765: out = 16'(395);
			19766: out = 16'(4044);
			19767: out = 16'(8447);
			19768: out = 16'(1828);
			19769: out = 16'(-7987);
			19770: out = 16'(-8434);
			19771: out = 16'(897);
			19772: out = 16'(7270);
			19773: out = 16'(3979);
			19774: out = 16'(-1267);
			19775: out = 16'(-766);
			19776: out = 16'(2496);
			19777: out = 16'(861);
			19778: out = 16'(-4599);
			19779: out = 16'(-7558);
			19780: out = 16'(-2308);
			19781: out = 16'(1292);
			19782: out = 16'(1623);
			19783: out = 16'(2421);
			19784: out = 16'(-2155);
			19785: out = 16'(-3366);
			19786: out = 16'(-3450);
			19787: out = 16'(-2424);
			19788: out = 16'(-4657);
			19789: out = 16'(-998);
			19790: out = 16'(748);
			19791: out = 16'(-589);
			19792: out = 16'(834);
			19793: out = 16'(427);
			19794: out = 16'(377);
			19795: out = 16'(-578);
			19796: out = 16'(919);
			19797: out = 16'(-1344);
			19798: out = 16'(-1065);
			19799: out = 16'(-2177);
			19800: out = 16'(-2622);
			19801: out = 16'(400);
			19802: out = 16'(8227);
			19803: out = 16'(8542);
			19804: out = 16'(345);
			19805: out = 16'(-3928);
			19806: out = 16'(-6100);
			19807: out = 16'(-8241);
			19808: out = 16'(-8544);
			19809: out = 16'(1375);
			19810: out = 16'(5291);
			19811: out = 16'(3034);
			19812: out = 16'(-309);
			19813: out = 16'(1993);
			19814: out = 16'(5497);
			19815: out = 16'(4214);
			19816: out = 16'(751);
			19817: out = 16'(-379);
			19818: out = 16'(-1843);
			19819: out = 16'(-4894);
			19820: out = 16'(-3014);
			19821: out = 16'(4203);
			19822: out = 16'(5329);
			19823: out = 16'(-213);
			19824: out = 16'(-4043);
			19825: out = 16'(-2052);
			19826: out = 16'(-2450);
			19827: out = 16'(-6087);
			19828: out = 16'(-4601);
			19829: out = 16'(5028);
			19830: out = 16'(10715);
			19831: out = 16'(8206);
			19832: out = 16'(2019);
			19833: out = 16'(-948);
			19834: out = 16'(-1791);
			19835: out = 16'(-546);
			19836: out = 16'(-881);
			19837: out = 16'(638);
			19838: out = 16'(3447);
			19839: out = 16'(3391);
			19840: out = 16'(239);
			19841: out = 16'(-2116);
			19842: out = 16'(38);
			19843: out = 16'(841);
			19844: out = 16'(2001);
			19845: out = 16'(-302);
			19846: out = 16'(-1107);
			19847: out = 16'(1046);
			19848: out = 16'(7146);
			19849: out = 16'(4450);
			19850: out = 16'(-2911);
			19851: out = 16'(-5391);
			19852: out = 16'(1230);
			19853: out = 16'(2341);
			19854: out = 16'(-3353);
			19855: out = 16'(-7436);
			19856: out = 16'(-3838);
			19857: out = 16'(-531);
			19858: out = 16'(-79);
			19859: out = 16'(2663);
			19860: out = 16'(4932);
			19861: out = 16'(8012);
			19862: out = 16'(2259);
			19863: out = 16'(-7522);
			19864: out = 16'(-10964);
			19865: out = 16'(-3812);
			19866: out = 16'(2534);
			19867: out = 16'(3607);
			19868: out = 16'(6131);
			19869: out = 16'(724);
			19870: out = 16'(-3955);
			19871: out = 16'(-7415);
			19872: out = 16'(-4950);
			19873: out = 16'(-4388);
			19874: out = 16'(297);
			19875: out = 16'(1400);
			19876: out = 16'(94);
			19877: out = 16'(263);
			19878: out = 16'(4614);
			19879: out = 16'(5031);
			19880: out = 16'(763);
			19881: out = 16'(-2175);
			19882: out = 16'(-1755);
			19883: out = 16'(-3309);
			19884: out = 16'(-7170);
			19885: out = 16'(-5030);
			19886: out = 16'(-4127);
			19887: out = 16'(261);
			19888: out = 16'(6054);
			19889: out = 16'(10435);
			19890: out = 16'(5303);
			19891: out = 16'(-2886);
			19892: out = 16'(-9510);
			19893: out = 16'(-10314);
			19894: out = 16'(-2596);
			19895: out = 16'(2477);
			19896: out = 16'(4755);
			19897: out = 16'(4985);
			19898: out = 16'(260);
			19899: out = 16'(-1988);
			19900: out = 16'(-1356);
			19901: out = 16'(-284);
			19902: out = 16'(-3059);
			19903: out = 16'(-6503);
			19904: out = 16'(-4636);
			19905: out = 16'(2578);
			19906: out = 16'(5794);
			19907: out = 16'(3608);
			19908: out = 16'(-19);
			19909: out = 16'(1689);
			19910: out = 16'(4057);
			19911: out = 16'(4706);
			19912: out = 16'(-5076);
			19913: out = 16'(-11537);
			19914: out = 16'(-5557);
			19915: out = 16'(2405);
			19916: out = 16'(7476);
			19917: out = 16'(6873);
			19918: out = 16'(3565);
			19919: out = 16'(-830);
			19920: out = 16'(-5913);
			19921: out = 16'(-6887);
			19922: out = 16'(-2812);
			19923: out = 16'(-133);
			19924: out = 16'(4741);
			19925: out = 16'(4972);
			19926: out = 16'(3366);
			19927: out = 16'(3875);
			19928: out = 16'(3320);
			19929: out = 16'(3834);
			19930: out = 16'(2215);
			19931: out = 16'(-1035);
			19932: out = 16'(-8134);
			19933: out = 16'(-6086);
			19934: out = 16'(-2247);
			19935: out = 16'(-2447);
			19936: out = 16'(205);
			19937: out = 16'(3870);
			19938: out = 16'(8580);
			19939: out = 16'(7780);
			19940: out = 16'(2950);
			19941: out = 16'(-2747);
			19942: out = 16'(-2930);
			19943: out = 16'(-1580);
			19944: out = 16'(-1372);
			19945: out = 16'(-985);
			19946: out = 16'(3002);
			19947: out = 16'(4555);
			19948: out = 16'(979);
			19949: out = 16'(-3083);
			19950: out = 16'(-3870);
			19951: out = 16'(-3450);
			19952: out = 16'(-1942);
			19953: out = 16'(-917);
			19954: out = 16'(3076);
			19955: out = 16'(102);
			19956: out = 16'(-6797);
			19957: out = 16'(-9846);
			19958: out = 16'(648);
			19959: out = 16'(6654);
			19960: out = 16'(5520);
			19961: out = 16'(3256);
			19962: out = 16'(-1372);
			19963: out = 16'(-10300);
			19964: out = 16'(-12491);
			19965: out = 16'(1228);
			19966: out = 16'(7471);
			19967: out = 16'(6586);
			19968: out = 16'(2179);
			19969: out = 16'(2083);
			19970: out = 16'(1530);
			19971: out = 16'(-1988);
			19972: out = 16'(-5214);
			19973: out = 16'(-1652);
			19974: out = 16'(3669);
			19975: out = 16'(5906);
			19976: out = 16'(2150);
			19977: out = 16'(-2026);
			19978: out = 16'(-1313);
			19979: out = 16'(-2424);
			19980: out = 16'(-1985);
			19981: out = 16'(-650);
			19982: out = 16'(1788);
			19983: out = 16'(-4597);
			19984: out = 16'(-3048);
			19985: out = 16'(2376);
			19986: out = 16'(5014);
			19987: out = 16'(509);
			19988: out = 16'(-550);
			19989: out = 16'(683);
			19990: out = 16'(1595);
			19991: out = 16'(-148);
			19992: out = 16'(-1014);
			19993: out = 16'(-2037);
			19994: out = 16'(-2660);
			19995: out = 16'(-4551);
			19996: out = 16'(-352);
			19997: out = 16'(685);
			19998: out = 16'(-171);
			19999: out = 16'(15);
			20000: out = 16'(93);
			20001: out = 16'(719);
			20002: out = 16'(3981);
			20003: out = 16'(7681);
			20004: out = 16'(5813);
			20005: out = 16'(877);
			20006: out = 16'(-2986);
			20007: out = 16'(-4979);
			20008: out = 16'(-5205);
			20009: out = 16'(-5590);
			20010: out = 16'(423);
			20011: out = 16'(6124);
			20012: out = 16'(-128);
			20013: out = 16'(-1994);
			20014: out = 16'(-415);
			20015: out = 16'(1520);
			20016: out = 16'(-2464);
			20017: out = 16'(-583);
			20018: out = 16'(2305);
			20019: out = 16'(1974);
			20020: out = 16'(-5154);
			20021: out = 16'(-7103);
			20022: out = 16'(-2431);
			20023: out = 16'(4371);
			20024: out = 16'(3922);
			20025: out = 16'(6239);
			20026: out = 16'(-992);
			20027: out = 16'(-3546);
			20028: out = 16'(-1342);
			20029: out = 16'(4551);
			20030: out = 16'(-582);
			20031: out = 16'(-2560);
			20032: out = 16'(73);
			20033: out = 16'(4503);
			20034: out = 16'(575);
			20035: out = 16'(-603);
			20036: out = 16'(766);
			20037: out = 16'(3546);
			20038: out = 16'(-2732);
			20039: out = 16'(-1920);
			20040: out = 16'(559);
			20041: out = 16'(1374);
			20042: out = 16'(-7148);
			20043: out = 16'(-2988);
			20044: out = 16'(534);
			20045: out = 16'(210);
			20046: out = 16'(1626);
			20047: out = 16'(5137);
			20048: out = 16'(197);
			20049: out = 16'(-8827);
			20050: out = 16'(-5661);
			20051: out = 16'(2559);
			20052: out = 16'(5800);
			20053: out = 16'(537);
			20054: out = 16'(-1298);
			20055: out = 16'(-1278);
			20056: out = 16'(3597);
			20057: out = 16'(2644);
			20058: out = 16'(-2646);
			20059: out = 16'(-5337);
			20060: out = 16'(-2230);
			20061: out = 16'(648);
			20062: out = 16'(669);
			20063: out = 16'(177);
			20064: out = 16'(4244);
			20065: out = 16'(8280);
			20066: out = 16'(8745);
			20067: out = 16'(5871);
			20068: out = 16'(1251);
			20069: out = 16'(-5149);
			20070: out = 16'(-8739);
			20071: out = 16'(-2968);
			20072: out = 16'(-3819);
			20073: out = 16'(-524);
			20074: out = 16'(3815);
			20075: out = 16'(7539);
			20076: out = 16'(533);
			20077: out = 16'(-633);
			20078: out = 16'(-1027);
			20079: out = 16'(-2899);
			20080: out = 16'(-4277);
			20081: out = 16'(-1960);
			20082: out = 16'(2258);
			20083: out = 16'(3958);
			20084: out = 16'(-291);
			20085: out = 16'(929);
			20086: out = 16'(2745);
			20087: out = 16'(2939);
			20088: out = 16'(316);
			20089: out = 16'(439);
			20090: out = 16'(-1055);
			20091: out = 16'(-3694);
			20092: out = 16'(-5399);
			20093: out = 16'(-1286);
			20094: out = 16'(-8);
			20095: out = 16'(-142);
			20096: out = 16'(2665);
			20097: out = 16'(5192);
			20098: out = 16'(5306);
			20099: out = 16'(-706);
			20100: out = 16'(-5881);
			20101: out = 16'(-6095);
			20102: out = 16'(2611);
			20103: out = 16'(4480);
			20104: out = 16'(366);
			20105: out = 16'(-2358);
			20106: out = 16'(-692);
			20107: out = 16'(-2142);
			20108: out = 16'(-5280);
			20109: out = 16'(-4990);
			20110: out = 16'(3700);
			20111: out = 16'(4242);
			20112: out = 16'(-120);
			20113: out = 16'(-1845);
			20114: out = 16'(2870);
			20115: out = 16'(2749);
			20116: out = 16'(1269);
			20117: out = 16'(1968);
			20118: out = 16'(3222);
			20119: out = 16'(-5942);
			20120: out = 16'(-16090);
			20121: out = 16'(-15471);
			20122: out = 16'(-670);
			20123: out = 16'(5095);
			20124: out = 16'(5096);
			20125: out = 16'(3355);
			20126: out = 16'(2053);
			20127: out = 16'(3489);
			20128: out = 16'(2089);
			20129: out = 16'(-2024);
			20130: out = 16'(-4915);
			20131: out = 16'(-1046);
			20132: out = 16'(3087);
			20133: out = 16'(698);
			20134: out = 16'(-6913);
			20135: out = 16'(-3829);
			20136: out = 16'(-450);
			20137: out = 16'(5877);
			20138: out = 16'(8705);
			20139: out = 16'(3602);
			20140: out = 16'(-2766);
			20141: out = 16'(-8574);
			20142: out = 16'(-9625);
			20143: out = 16'(-2533);
			20144: out = 16'(849);
			20145: out = 16'(5302);
			20146: out = 16'(7110);
			20147: out = 16'(5752);
			20148: out = 16'(-1027);
			20149: out = 16'(-2647);
			20150: out = 16'(-1316);
			20151: out = 16'(204);
			20152: out = 16'(-245);
			20153: out = 16'(1294);
			20154: out = 16'(2091);
			20155: out = 16'(1123);
			20156: out = 16'(-5037);
			20157: out = 16'(-2388);
			20158: out = 16'(1130);
			20159: out = 16'(5090);
			20160: out = 16'(6960);
			20161: out = 16'(5316);
			20162: out = 16'(-3347);
			20163: out = 16'(-7772);
			20164: out = 16'(-565);
			20165: out = 16'(5146);
			20166: out = 16'(3003);
			20167: out = 16'(-1528);
			20168: out = 16'(-2116);
			20169: out = 16'(-1291);
			20170: out = 16'(-6323);
			20171: out = 16'(-9642);
			20172: out = 16'(-4092);
			20173: out = 16'(2897);
			20174: out = 16'(7358);
			20175: out = 16'(6910);
			20176: out = 16'(4376);
			20177: out = 16'(689);
			20178: out = 16'(-3156);
			20179: out = 16'(-5092);
			20180: out = 16'(-4610);
			20181: out = 16'(-1791);
			20182: out = 16'(-1479);
			20183: out = 16'(955);
			20184: out = 16'(2108);
			20185: out = 16'(1961);
			20186: out = 16'(-1915);
			20187: out = 16'(535);
			20188: out = 16'(1716);
			20189: out = 16'(-833);
			20190: out = 16'(-8868);
			20191: out = 16'(-4036);
			20192: out = 16'(1219);
			20193: out = 16'(1939);
			20194: out = 16'(53);
			20195: out = 16'(7317);
			20196: out = 16'(6928);
			20197: out = 16'(-1400);
			20198: out = 16'(-8910);
			20199: out = 16'(-4813);
			20200: out = 16'(-635);
			20201: out = 16'(1283);
			20202: out = 16'(5370);
			20203: out = 16'(8552);
			20204: out = 16'(5624);
			20205: out = 16'(-2201);
			20206: out = 16'(-7116);
			20207: out = 16'(-5831);
			20208: out = 16'(979);
			20209: out = 16'(5107);
			20210: out = 16'(4785);
			20211: out = 16'(2001);
			20212: out = 16'(2987);
			20213: out = 16'(2355);
			20214: out = 16'(-1788);
			20215: out = 16'(-4863);
			20216: out = 16'(-5979);
			20217: out = 16'(-2114);
			20218: out = 16'(67);
			20219: out = 16'(-1259);
			20220: out = 16'(-8463);
			20221: out = 16'(-2142);
			20222: out = 16'(9765);
			20223: out = 16'(13521);
			20224: out = 16'(8520);
			20225: out = 16'(1985);
			20226: out = 16'(-3271);
			20227: out = 16'(-9148);
			20228: out = 16'(-15511);
			20229: out = 16'(-10660);
			20230: out = 16'(2137);
			20231: out = 16'(10118);
			20232: out = 16'(9151);
			20233: out = 16'(4690);
			20234: out = 16'(1696);
			20235: out = 16'(-2497);
			20236: out = 16'(-7271);
			20237: out = 16'(-12827);
			20238: out = 16'(-5692);
			20239: out = 16'(4135);
			20240: out = 16'(6068);
			20241: out = 16'(6528);
			20242: out = 16'(4585);
			20243: out = 16'(2089);
			20244: out = 16'(-552);
			20245: out = 16'(-3179);
			20246: out = 16'(-2391);
			20247: out = 16'(-3397);
			20248: out = 16'(-6012);
			20249: out = 16'(-10497);
			20250: out = 16'(-2181);
			20251: out = 16'(1180);
			20252: out = 16'(202);
			20253: out = 16'(778);
			20254: out = 16'(9439);
			20255: out = 16'(6140);
			20256: out = 16'(-5159);
			20257: out = 16'(-13317);
			20258: out = 16'(-1715);
			20259: out = 16'(1363);
			20260: out = 16'(-411);
			20261: out = 16'(941);
			20262: out = 16'(1867);
			20263: out = 16'(1350);
			20264: out = 16'(-417);
			20265: out = 16'(964);
			20266: out = 16'(1746);
			20267: out = 16'(1568);
			20268: out = 16'(-3463);
			20269: out = 16'(-6128);
			20270: out = 16'(688);
			20271: out = 16'(4560);
			20272: out = 16'(7016);
			20273: out = 16'(6810);
			20274: out = 16'(5660);
			20275: out = 16'(-6341);
			20276: out = 16'(-7627);
			20277: out = 16'(-1461);
			20278: out = 16'(4165);
			20279: out = 16'(4758);
			20280: out = 16'(1695);
			20281: out = 16'(-434);
			20282: out = 16'(478);
			20283: out = 16'(2562);
			20284: out = 16'(1192);
			20285: out = 16'(-2188);
			20286: out = 16'(-3979);
			20287: out = 16'(-1909);
			20288: out = 16'(2597);
			20289: out = 16'(2947);
			20290: out = 16'(-876);
			20291: out = 16'(-2279);
			20292: out = 16'(3538);
			20293: out = 16'(9188);
			20294: out = 16'(7380);
			20295: out = 16'(818);
			20296: out = 16'(-4874);
			20297: out = 16'(-3664);
			20298: out = 16'(-1872);
			20299: out = 16'(-2311);
			20300: out = 16'(-3045);
			20301: out = 16'(3344);
			20302: out = 16'(8305);
			20303: out = 16'(8289);
			20304: out = 16'(4809);
			20305: out = 16'(-323);
			20306: out = 16'(-7354);
			20307: out = 16'(-9983);
			20308: out = 16'(-2743);
			20309: out = 16'(967);
			20310: out = 16'(1305);
			20311: out = 16'(-970);
			20312: out = 16'(-1995);
			20313: out = 16'(-1348);
			20314: out = 16'(-500);
			20315: out = 16'(27);
			20316: out = 16'(271);
			20317: out = 16'(3601);
			20318: out = 16'(1568);
			20319: out = 16'(304);
			20320: out = 16'(-284);
			20321: out = 16'(231);
			20322: out = 16'(-3549);
			20323: out = 16'(-1672);
			20324: out = 16'(2986);
			20325: out = 16'(4175);
			20326: out = 16'(686);
			20327: out = 16'(-1582);
			20328: out = 16'(-2122);
			20329: out = 16'(249);
			20330: out = 16'(-726);
			20331: out = 16'(2335);
			20332: out = 16'(617);
			20333: out = 16'(-3796);
			20334: out = 16'(-15878);
			20335: out = 16'(-3451);
			20336: out = 16'(5943);
			20337: out = 16'(2028);
			20338: out = 16'(-5321);
			20339: out = 16'(2580);
			20340: out = 16'(6769);
			20341: out = 16'(1312);
			20342: out = 16'(-5652);
			20343: out = 16'(-2358);
			20344: out = 16'(-952);
			20345: out = 16'(-1707);
			20346: out = 16'(20);
			20347: out = 16'(587);
			20348: out = 16'(-5319);
			20349: out = 16'(-7646);
			20350: out = 16'(2020);
			20351: out = 16'(9573);
			20352: out = 16'(9853);
			20353: out = 16'(4635);
			20354: out = 16'(-591);
			20355: out = 16'(386);
			20356: out = 16'(-9229);
			20357: out = 16'(-11272);
			20358: out = 16'(-1428);
			20359: out = 16'(8769);
			20360: out = 16'(4469);
			20361: out = 16'(268);
			20362: out = 16'(266);
			20363: out = 16'(125);
			20364: out = 16'(-160);
			20365: out = 16'(4045);
			20366: out = 16'(8382);
			20367: out = 16'(4842);
			20368: out = 16'(-1431);
			20369: out = 16'(-5598);
			20370: out = 16'(-3252);
			20371: out = 16'(12);
			20372: out = 16'(-847);
			20373: out = 16'(-560);
			20374: out = 16'(1122);
			20375: out = 16'(1590);
			20376: out = 16'(77);
			20377: out = 16'(-264);
			20378: out = 16'(989);
			20379: out = 16'(2280);
			20380: out = 16'(4509);
			20381: out = 16'(658);
			20382: out = 16'(-1258);
			20383: out = 16'(-3386);
			20384: out = 16'(-5041);
			20385: out = 16'(-3158);
			20386: out = 16'(2076);
			20387: out = 16'(5262);
			20388: out = 16'(5786);
			20389: out = 16'(-59);
			20390: out = 16'(3373);
			20391: out = 16'(3638);
			20392: out = 16'(-1405);
			20393: out = 16'(-4216);
			20394: out = 16'(-3748);
			20395: out = 16'(-5033);
			20396: out = 16'(-7120);
			20397: out = 16'(-1946);
			20398: out = 16'(3031);
			20399: out = 16'(4946);
			20400: out = 16'(4842);
			20401: out = 16'(7701);
			20402: out = 16'(7415);
			20403: out = 16'(762);
			20404: out = 16'(-10197);
			20405: out = 16'(-14955);
			20406: out = 16'(-9201);
			20407: out = 16'(-581);
			20408: out = 16'(3168);
			20409: out = 16'(5412);
			20410: out = 16'(7004);
			20411: out = 16'(5864);
			20412: out = 16'(-3079);
			20413: out = 16'(-10600);
			20414: out = 16'(-3041);
			20415: out = 16'(3635);
			20416: out = 16'(4507);
			20417: out = 16'(697);
			20418: out = 16'(154);
			20419: out = 16'(-6225);
			20420: out = 16'(-5373);
			20421: out = 16'(1556);
			20422: out = 16'(7307);
			20423: out = 16'(1329);
			20424: out = 16'(-3449);
			20425: out = 16'(-2084);
			20426: out = 16'(1163);
			20427: out = 16'(-8432);
			20428: out = 16'(-7842);
			20429: out = 16'(2355);
			20430: out = 16'(11178);
			20431: out = 16'(6033);
			20432: out = 16'(-3666);
			20433: out = 16'(-8556);
			20434: out = 16'(-6690);
			20435: out = 16'(-8469);
			20436: out = 16'(-5400);
			20437: out = 16'(1684);
			20438: out = 16'(11776);
			20439: out = 16'(12416);
			20440: out = 16'(6399);
			20441: out = 16'(-7482);
			20442: out = 16'(-11872);
			20443: out = 16'(-3498);
			20444: out = 16'(1480);
			20445: out = 16'(-576);
			20446: out = 16'(-2738);
			20447: out = 16'(2012);
			20448: out = 16'(5658);
			20449: out = 16'(6740);
			20450: out = 16'(2449);
			20451: out = 16'(774);
			20452: out = 16'(3396);
			20453: out = 16'(2835);
			20454: out = 16'(-2547);
			20455: out = 16'(-7595);
			20456: out = 16'(-9186);
			20457: out = 16'(-2883);
			20458: out = 16'(504);
			20459: out = 16'(5019);
			20460: out = 16'(9486);
			20461: out = 16'(9745);
			20462: out = 16'(-248);
			20463: out = 16'(-6458);
			20464: out = 16'(-2280);
			20465: out = 16'(3800);
			20466: out = 16'(2517);
			20467: out = 16'(-1565);
			20468: out = 16'(-2994);
			20469: out = 16'(-2091);
			20470: out = 16'(-1386);
			20471: out = 16'(929);
			20472: out = 16'(4062);
			20473: out = 16'(6154);
			20474: out = 16'(5426);
			20475: out = 16'(2486);
			20476: out = 16'(-2482);
			20477: out = 16'(-5097);
			20478: out = 16'(-7035);
			20479: out = 16'(542);
			20480: out = 16'(3124);
			20481: out = 16'(-535);
			20482: out = 16'(-1052);
			20483: out = 16'(73);
			20484: out = 16'(-2515);
			20485: out = 16'(-6115);
			20486: out = 16'(-2773);
			20487: out = 16'(7444);
			20488: out = 16'(7442);
			20489: out = 16'(-1060);
			20490: out = 16'(-4260);
			20491: out = 16'(-1522);
			20492: out = 16'(2074);
			20493: out = 16'(1010);
			20494: out = 16'(447);
			20495: out = 16'(-421);
			20496: out = 16'(2769);
			20497: out = 16'(2288);
			20498: out = 16'(-2136);
			20499: out = 16'(-6703);
			20500: out = 16'(-1602);
			20501: out = 16'(5361);
			20502: out = 16'(5628);
			20503: out = 16'(474);
			20504: out = 16'(-4336);
			20505: out = 16'(-4393);
			20506: out = 16'(-2592);
			20507: out = 16'(-743);
			20508: out = 16'(-515);
			20509: out = 16'(5380);
			20510: out = 16'(9188);
			20511: out = 16'(4189);
			20512: out = 16'(-1709);
			20513: out = 16'(-2522);
			20514: out = 16'(1439);
			20515: out = 16'(499);
			20516: out = 16'(-3918);
			20517: out = 16'(-9243);
			20518: out = 16'(-5855);
			20519: out = 16'(1230);
			20520: out = 16'(3670);
			20521: out = 16'(965);
			20522: out = 16'(-226);
			20523: out = 16'(401);
			20524: out = 16'(2029);
			20525: out = 16'(-3902);
			20526: out = 16'(-3064);
			20527: out = 16'(757);
			20528: out = 16'(-139);
			20529: out = 16'(-1521);
			20530: out = 16'(406);
			20531: out = 16'(5102);
			20532: out = 16'(7243);
			20533: out = 16'(2435);
			20534: out = 16'(321);
			20535: out = 16'(-1164);
			20536: out = 16'(-1961);
			20537: out = 16'(431);
			20538: out = 16'(5754);
			20539: out = 16'(6602);
			20540: out = 16'(1207);
			20541: out = 16'(-4930);
			20542: out = 16'(-4464);
			20543: out = 16'(-1289);
			20544: out = 16'(-119);
			20545: out = 16'(38);
			20546: out = 16'(4765);
			20547: out = 16'(5519);
			20548: out = 16'(-197);
			20549: out = 16'(-7338);
			20550: out = 16'(-3282);
			20551: out = 16'(789);
			20552: out = 16'(1174);
			20553: out = 16'(-672);
			20554: out = 16'(-3204);
			20555: out = 16'(-1154);
			20556: out = 16'(-94);
			20557: out = 16'(1099);
			20558: out = 16'(7286);
			20559: out = 16'(6713);
			20560: out = 16'(2682);
			20561: out = 16'(-1273);
			20562: out = 16'(-1562);
			20563: out = 16'(-3747);
			20564: out = 16'(-5663);
			20565: out = 16'(-2466);
			20566: out = 16'(6475);
			20567: out = 16'(5842);
			20568: out = 16'(2271);
			20569: out = 16'(-2341);
			20570: out = 16'(-3589);
			20571: out = 16'(-7548);
			20572: out = 16'(-2964);
			20573: out = 16'(2707);
			20574: out = 16'(4601);
			20575: out = 16'(14);
			20576: out = 16'(-440);
			20577: out = 16'(21);
			20578: out = 16'(-813);
			20579: out = 16'(-2180);
			20580: out = 16'(-7559);
			20581: out = 16'(-5524);
			20582: out = 16'(1674);
			20583: out = 16'(5719);
			20584: out = 16'(1050);
			20585: out = 16'(-1651);
			20586: out = 16'(700);
			20587: out = 16'(4528);
			20588: out = 16'(3534);
			20589: out = 16'(2288);
			20590: out = 16'(806);
			20591: out = 16'(-1461);
			20592: out = 16'(-8168);
			20593: out = 16'(-3226);
			20594: out = 16'(3625);
			20595: out = 16'(5367);
			20596: out = 16'(1758);
			20597: out = 16'(-52);
			20598: out = 16'(676);
			20599: out = 16'(1237);
			20600: out = 16'(-1779);
			20601: out = 16'(-2051);
			20602: out = 16'(-3262);
			20603: out = 16'(-2001);
			20604: out = 16'(2205);
			20605: out = 16'(3057);
			20606: out = 16'(4202);
			20607: out = 16'(3286);
			20608: out = 16'(1130);
			20609: out = 16'(-425);
			20610: out = 16'(-629);
			20611: out = 16'(-1559);
			20612: out = 16'(-4176);
			20613: out = 16'(-5106);
			20614: out = 16'(-1401);
			20615: out = 16'(2929);
			20616: out = 16'(2422);
			20617: out = 16'(196);
			20618: out = 16'(-884);
			20619: out = 16'(3630);
			20620: out = 16'(4627);
			20621: out = 16'(-777);
			20622: out = 16'(-2319);
			20623: out = 16'(418);
			20624: out = 16'(2373);
			20625: out = 16'(-188);
			20626: out = 16'(-322);
			20627: out = 16'(2686);
			20628: out = 16'(7201);
			20629: out = 16'(7545);
			20630: out = 16'(1339);
			20631: out = 16'(-1087);
			20632: out = 16'(-3488);
			20633: out = 16'(-4885);
			20634: out = 16'(-3516);
			20635: out = 16'(1713);
			20636: out = 16'(3665);
			20637: out = 16'(2290);
			20638: out = 16'(1174);
			20639: out = 16'(-1457);
			20640: out = 16'(-2527);
			20641: out = 16'(-2547);
			20642: out = 16'(-1640);
			20643: out = 16'(-1763);
			20644: out = 16'(-1722);
			20645: out = 16'(-611);
			20646: out = 16'(1789);
			20647: out = 16'(1113);
			20648: out = 16'(-1141);
			20649: out = 16'(-3537);
			20650: out = 16'(-876);
			20651: out = 16'(3395);
			20652: out = 16'(1390);
			20653: out = 16'(-5022);
			20654: out = 16'(-6921);
			20655: out = 16'(-3351);
			20656: out = 16'(5104);
			20657: out = 16'(2459);
			20658: out = 16'(-317);
			20659: out = 16'(1564);
			20660: out = 16'(1876);
			20661: out = 16'(-5852);
			20662: out = 16'(-9322);
			20663: out = 16'(-2979);
			20664: out = 16'(-692);
			20665: out = 16'(-1907);
			20666: out = 16'(-2619);
			20667: out = 16'(803);
			20668: out = 16'(1490);
			20669: out = 16'(621);
			20670: out = 16'(-1050);
			20671: out = 16'(-923);
			20672: out = 16'(-41);
			20673: out = 16'(2888);
			20674: out = 16'(4554);
			20675: out = 16'(2995);
			20676: out = 16'(-419);
			20677: out = 16'(-5036);
			20678: out = 16'(-178);
			20679: out = 16'(5483);
			20680: out = 16'(4481);
			20681: out = 16'(-6457);
			20682: out = 16'(-5350);
			20683: out = 16'(-1267);
			20684: out = 16'(-156);
			20685: out = 16'(-1054);
			20686: out = 16'(5334);
			20687: out = 16'(7896);
			20688: out = 16'(3619);
			20689: out = 16'(-2216);
			20690: out = 16'(-1037);
			20691: out = 16'(-837);
			20692: out = 16'(-3968);
			20693: out = 16'(-4126);
			20694: out = 16'(7778);
			20695: out = 16'(12713);
			20696: out = 16'(3454);
			20697: out = 16'(-11923);
			20698: out = 16'(-6077);
			20699: out = 16'(442);
			20700: out = 16'(3684);
			20701: out = 16'(730);
			20702: out = 16'(2163);
			20703: out = 16'(7);
			20704: out = 16'(2090);
			20705: out = 16'(2444);
			20706: out = 16'(-227);
			20707: out = 16'(-4241);
			20708: out = 16'(-1558);
			20709: out = 16'(1737);
			20710: out = 16'(-895);
			20711: out = 16'(-4691);
			20712: out = 16'(-2191);
			20713: out = 16'(4568);
			20714: out = 16'(6410);
			20715: out = 16'(686);
			20716: out = 16'(-1317);
			20717: out = 16'(28);
			20718: out = 16'(-2134);
			20719: out = 16'(-7660);
			20720: out = 16'(-9227);
			20721: out = 16'(-774);
			20722: out = 16'(8449);
			20723: out = 16'(10745);
			20724: out = 16'(560);
			20725: out = 16'(-4177);
			20726: out = 16'(-2499);
			20727: out = 16'(-679);
			20728: out = 16'(-8166);
			20729: out = 16'(-8367);
			20730: out = 16'(-2420);
			20731: out = 16'(1535);
			20732: out = 16'(-3376);
			20733: out = 16'(-2092);
			20734: out = 16'(2386);
			20735: out = 16'(4237);
			20736: out = 16'(2090);
			20737: out = 16'(426);
			20738: out = 16'(-1896);
			20739: out = 16'(-4726);
			20740: out = 16'(-4891);
			20741: out = 16'(-5313);
			20742: out = 16'(-2695);
			20743: out = 16'(2510);
			20744: out = 16'(7604);
			20745: out = 16'(4168);
			20746: out = 16'(-1228);
			20747: out = 16'(-4864);
			20748: out = 16'(-5017);
			20749: out = 16'(-4982);
			20750: out = 16'(-3445);
			20751: out = 16'(1357);
			20752: out = 16'(7056);
			20753: out = 16'(7772);
			20754: out = 16'(946);
			20755: out = 16'(-5232);
			20756: out = 16'(-3258);
			20757: out = 16'(2235);
			20758: out = 16'(5659);
			20759: out = 16'(2760);
			20760: out = 16'(-343);
			20761: out = 16'(39);
			20762: out = 16'(381);
			20763: out = 16'(-1750);
			20764: out = 16'(-1606);
			20765: out = 16'(4109);
			20766: out = 16'(2916);
			20767: out = 16'(-294);
			20768: out = 16'(-5076);
			20769: out = 16'(-6597);
			20770: out = 16'(-3619);
			20771: out = 16'(2830);
			20772: out = 16'(7632);
			20773: out = 16'(8936);
			20774: out = 16'(6110);
			20775: out = 16'(4904);
			20776: out = 16'(870);
			20777: out = 16'(-7183);
			20778: out = 16'(-14609);
			20779: out = 16'(-7423);
			20780: out = 16'(5754);
			20781: out = 16'(9171);
			20782: out = 16'(1725);
			20783: out = 16'(465);
			20784: out = 16'(4786);
			20785: out = 16'(6491);
			20786: out = 16'(762);
			20787: out = 16'(-876);
			20788: out = 16'(-2782);
			20789: out = 16'(-4238);
			20790: out = 16'(-5101);
			20791: out = 16'(-3565);
			20792: out = 16'(3377);
			20793: out = 16'(7128);
			20794: out = 16'(5612);
			20795: out = 16'(484);
			20796: out = 16'(182);
			20797: out = 16'(-2809);
			20798: out = 16'(-5766);
			20799: out = 16'(-5144);
			20800: out = 16'(1979);
			20801: out = 16'(4713);
			20802: out = 16'(5059);
			20803: out = 16'(3064);
			20804: out = 16'(-1356);
			20805: out = 16'(-10285);
			20806: out = 16'(-8769);
			20807: out = 16'(3263);
			20808: out = 16'(8387);
			20809: out = 16'(1045);
			20810: out = 16'(-4053);
			20811: out = 16'(-1485);
			20812: out = 16'(-414);
			20813: out = 16'(-5299);
			20814: out = 16'(-4681);
			20815: out = 16'(1407);
			20816: out = 16'(1394);
			20817: out = 16'(-1742);
			20818: out = 16'(-1953);
			20819: out = 16'(1022);
			20820: out = 16'(1655);
			20821: out = 16'(-2369);
			20822: out = 16'(1824);
			20823: out = 16'(6570);
			20824: out = 16'(2016);
			20825: out = 16'(-2626);
			20826: out = 16'(-5660);
			20827: out = 16'(-2985);
			20828: out = 16'(123);
			20829: out = 16'(147);
			20830: out = 16'(3022);
			20831: out = 16'(4683);
			20832: out = 16'(1807);
			20833: out = 16'(-4649);
			20834: out = 16'(-5477);
			20835: out = 16'(-2288);
			20836: out = 16'(2262);
			20837: out = 16'(4188);
			20838: out = 16'(6130);
			20839: out = 16'(1182);
			20840: out = 16'(-5227);
			20841: out = 16'(-6317);
			20842: out = 16'(1245);
			20843: out = 16'(1918);
			20844: out = 16'(-2194);
			20845: out = 16'(-1441);
			20846: out = 16'(6796);
			20847: out = 16'(7926);
			20848: out = 16'(161);
			20849: out = 16'(-5682);
			20850: out = 16'(1257);
			20851: out = 16'(4159);
			20852: out = 16'(697);
			20853: out = 16'(-3558);
			20854: out = 16'(-982);
			20855: out = 16'(3845);
			20856: out = 16'(4066);
			20857: out = 16'(1722);
			20858: out = 16'(1741);
			20859: out = 16'(4385);
			20860: out = 16'(480);
			20861: out = 16'(-6757);
			20862: out = 16'(-9864);
			20863: out = 16'(-1233);
			20864: out = 16'(1567);
			20865: out = 16'(1529);
			20866: out = 16'(2111);
			20867: out = 16'(4816);
			20868: out = 16'(3736);
			20869: out = 16'(1627);
			20870: out = 16'(-984);
			20871: out = 16'(-71);
			20872: out = 16'(-3557);
			20873: out = 16'(-502);
			20874: out = 16'(171);
			20875: out = 16'(-5604);
			20876: out = 16'(-10262);
			20877: out = 16'(-2961);
			20878: out = 16'(5777);
			20879: out = 16'(3852);
			20880: out = 16'(727);
			20881: out = 16'(-1001);
			20882: out = 16'(418);
			20883: out = 16'(-1016);
			20884: out = 16'(-2581);
			20885: out = 16'(-1725);
			20886: out = 16'(2285);
			20887: out = 16'(2223);
			20888: out = 16'(-1804);
			20889: out = 16'(-4358);
			20890: out = 16'(-1763);
			20891: out = 16'(-153);
			20892: out = 16'(-782);
			20893: out = 16'(-650);
			20894: out = 16'(4031);
			20895: out = 16'(4276);
			20896: out = 16'(-1904);
			20897: out = 16'(-5744);
			20898: out = 16'(-2606);
			20899: out = 16'(576);
			20900: out = 16'(111);
			20901: out = 16'(1669);
			20902: out = 16'(3449);
			20903: out = 16'(209);
			20904: out = 16'(-6100);
			20905: out = 16'(-5731);
			20906: out = 16'(-3083);
			20907: out = 16'(-1562);
			20908: out = 16'(-891);
			20909: out = 16'(3958);
			20910: out = 16'(-70);
			20911: out = 16'(-1063);
			20912: out = 16'(2848);
			20913: out = 16'(8925);
			20914: out = 16'(4348);
			20915: out = 16'(-2024);
			20916: out = 16'(-5631);
			20917: out = 16'(-3532);
			20918: out = 16'(-3201);
			20919: out = 16'(-2914);
			20920: out = 16'(-815);
			20921: out = 16'(4163);
			20922: out = 16'(5613);
			20923: out = 16'(3445);
			20924: out = 16'(-177);
			20925: out = 16'(-700);
			20926: out = 16'(-297);
			20927: out = 16'(-2772);
			20928: out = 16'(-4532);
			20929: out = 16'(944);
			20930: out = 16'(9906);
			20931: out = 16'(10438);
			20932: out = 16'(3905);
			20933: out = 16'(-3118);
			20934: out = 16'(-4757);
			20935: out = 16'(-105);
			20936: out = 16'(478);
			20937: out = 16'(-834);
			20938: out = 16'(-1156);
			20939: out = 16'(-334);
			20940: out = 16'(-199);
			20941: out = 16'(1402);
			20942: out = 16'(3745);
			20943: out = 16'(2950);
			20944: out = 16'(-157);
			20945: out = 16'(-2879);
			20946: out = 16'(-3175);
			20947: out = 16'(-3055);
			20948: out = 16'(2533);
			20949: out = 16'(4137);
			20950: out = 16'(3134);
			20951: out = 16'(97);
			20952: out = 16'(1710);
			20953: out = 16'(45);
			20954: out = 16'(-268);
			20955: out = 16'(-1143);
			20956: out = 16'(-2842);
			20957: out = 16'(-6137);
			20958: out = 16'(-2419);
			20959: out = 16'(4970);
			20960: out = 16'(6688);
			20961: out = 16'(1558);
			20962: out = 16'(-1521);
			20963: out = 16'(965);
			20964: out = 16'(3387);
			20965: out = 16'(-3305);
			20966: out = 16'(-8599);
			20967: out = 16'(-8318);
			20968: out = 16'(-4469);
			20969: out = 16'(2730);
			20970: out = 16'(2922);
			20971: out = 16'(520);
			20972: out = 16'(-1102);
			20973: out = 16'(-41);
			20974: out = 16'(4);
			20975: out = 16'(26);
			20976: out = 16'(-536);
			20977: out = 16'(-3948);
			20978: out = 16'(267);
			20979: out = 16'(1840);
			20980: out = 16'(-1982);
			20981: out = 16'(-6312);
			20982: out = 16'(-2046);
			20983: out = 16'(5270);
			20984: out = 16'(5765);
			20985: out = 16'(-772);
			20986: out = 16'(-6326);
			20987: out = 16'(-3352);
			20988: out = 16'(1479);
			20989: out = 16'(1480);
			20990: out = 16'(-619);
			20991: out = 16'(2229);
			20992: out = 16'(5900);
			20993: out = 16'(4417);
			20994: out = 16'(-2597);
			20995: out = 16'(-5721);
			20996: out = 16'(-5044);
			20997: out = 16'(-1685);
			20998: out = 16'(1838);
			20999: out = 16'(3477);
			21000: out = 16'(2704);
			21001: out = 16'(1295);
			21002: out = 16'(-620);
			21003: out = 16'(-3972);
			21004: out = 16'(-6882);
			21005: out = 16'(-4254);
			21006: out = 16'(2832);
			21007: out = 16'(5730);
			21008: out = 16'(4200);
			21009: out = 16'(1445);
			21010: out = 16'(-183);
			21011: out = 16'(203);
			21012: out = 16'(-3752);
			21013: out = 16'(-3400);
			21014: out = 16'(1437);
			21015: out = 16'(3011);
			21016: out = 16'(-4625);
			21017: out = 16'(-10642);
			21018: out = 16'(-7223);
			21019: out = 16'(1203);
			21020: out = 16'(5759);
			21021: out = 16'(8574);
			21022: out = 16'(11072);
			21023: out = 16'(8016);
			21024: out = 16'(1883);
			21025: out = 16'(-7192);
			21026: out = 16'(-6808);
			21027: out = 16'(634);
			21028: out = 16'(3368);
			21029: out = 16'(1922);
			21030: out = 16'(3554);
			21031: out = 16'(4933);
			21032: out = 16'(-129);
			21033: out = 16'(-7848);
			21034: out = 16'(-5087);
			21035: out = 16'(3849);
			21036: out = 16'(4297);
			21037: out = 16'(1123);
			21038: out = 16'(61);
			21039: out = 16'(2584);
			21040: out = 16'(2930);
			21041: out = 16'(2644);
			21042: out = 16'(744);
			21043: out = 16'(-2470);
			21044: out = 16'(-4495);
			21045: out = 16'(4680);
			21046: out = 16'(6572);
			21047: out = 16'(1044);
			21048: out = 16'(-5315);
			21049: out = 16'(1330);
			21050: out = 16'(527);
			21051: out = 16'(-4157);
			21052: out = 16'(-8337);
			21053: out = 16'(-2864);
			21054: out = 16'(-828);
			21055: out = 16'(-275);
			21056: out = 16'(-1820);
			21057: out = 16'(-1702);
			21058: out = 16'(2456);
			21059: out = 16'(4090);
			21060: out = 16'(1037);
			21061: out = 16'(-4672);
			21062: out = 16'(-2973);
			21063: out = 16'(-5748);
			21064: out = 16'(-7391);
			21065: out = 16'(-6112);
			21066: out = 16'(-126);
			21067: out = 16'(0);
			21068: out = 16'(1751);
			21069: out = 16'(4046);
			21070: out = 16'(3647);
			21071: out = 16'(2880);
			21072: out = 16'(1810);
			21073: out = 16'(-3287);
			21074: out = 16'(-12300);
			21075: out = 16'(-11368);
			21076: out = 16'(276);
			21077: out = 16'(10270);
			21078: out = 16'(7508);
			21079: out = 16'(-2619);
			21080: out = 16'(-4422);
			21081: out = 16'(1424);
			21082: out = 16'(2726);
			21083: out = 16'(-1653);
			21084: out = 16'(-3952);
			21085: out = 16'(2246);
			21086: out = 16'(7855);
			21087: out = 16'(5372);
			21088: out = 16'(-474);
			21089: out = 16'(-659);
			21090: out = 16'(2346);
			21091: out = 16'(314);
			21092: out = 16'(-2124);
			21093: out = 16'(-1948);
			21094: out = 16'(1975);
			21095: out = 16'(3727);
			21096: out = 16'(-3534);
			21097: out = 16'(-3303);
			21098: out = 16'(4134);
			21099: out = 16'(8414);
			21100: out = 16'(5838);
			21101: out = 16'(-2294);
			21102: out = 16'(-5230);
			21103: out = 16'(-2312);
			21104: out = 16'(-419);
			21105: out = 16'(-2289);
			21106: out = 16'(-331);
			21107: out = 16'(7352);
			21108: out = 16'(12354);
			21109: out = 16'(7875);
			21110: out = 16'(-1858);
			21111: out = 16'(-8746);
			21112: out = 16'(-8298);
			21113: out = 16'(-12460);
			21114: out = 16'(-7315);
			21115: out = 16'(3655);
			21116: out = 16'(10871);
			21117: out = 16'(6568);
			21118: out = 16'(1515);
			21119: out = 16'(649);
			21120: out = 16'(3966);
			21121: out = 16'(3605);
			21122: out = 16'(-621);
			21123: out = 16'(-7578);
			21124: out = 16'(-9561);
			21125: out = 16'(-3134);
			21126: out = 16'(974);
			21127: out = 16'(1208);
			21128: out = 16'(-377);
			21129: out = 16'(-34);
			21130: out = 16'(-138);
			21131: out = 16'(4);
			21132: out = 16'(-151);
			21133: out = 16'(983);
			21134: out = 16'(1528);
			21135: out = 16'(871);
			21136: out = 16'(-341);
			21137: out = 16'(1491);
			21138: out = 16'(2733);
			21139: out = 16'(3133);
			21140: out = 16'(-3007);
			21141: out = 16'(-8891);
			21142: out = 16'(-9248);
			21143: out = 16'(-333);
			21144: out = 16'(1909);
			21145: out = 16'(-597);
			21146: out = 16'(-1479);
			21147: out = 16'(6227);
			21148: out = 16'(5176);
			21149: out = 16'(-550);
			21150: out = 16'(-3767);
			21151: out = 16'(-471);
			21152: out = 16'(-2796);
			21153: out = 16'(-5656);
			21154: out = 16'(-3629);
			21155: out = 16'(3262);
			21156: out = 16'(2882);
			21157: out = 16'(1796);
			21158: out = 16'(2014);
			21159: out = 16'(1919);
			21160: out = 16'(-7011);
			21161: out = 16'(-10490);
			21162: out = 16'(-5342);
			21163: out = 16'(-10);
			21164: out = 16'(874);
			21165: out = 16'(1194);
			21166: out = 16'(2851);
			21167: out = 16'(1863);
			21168: out = 16'(2616);
			21169: out = 16'(784);
			21170: out = 16'(421);
			21171: out = 16'(-162);
			21172: out = 16'(429);
			21173: out = 16'(-1557);
			21174: out = 16'(-609);
			21175: out = 16'(977);
			21176: out = 16'(356);
			21177: out = 16'(1189);
			21178: out = 16'(4644);
			21179: out = 16'(4599);
			21180: out = 16'(-2768);
			21181: out = 16'(-5033);
			21182: out = 16'(867);
			21183: out = 16'(7140);
			21184: out = 16'(3716);
			21185: out = 16'(5692);
			21186: out = 16'(1557);
			21187: out = 16'(-4300);
			21188: out = 16'(-10111);
			21189: out = 16'(-1610);
			21190: out = 16'(2754);
			21191: out = 16'(5759);
			21192: out = 16'(5691);
			21193: out = 16'(6249);
			21194: out = 16'(-841);
			21195: out = 16'(-3237);
			21196: out = 16'(1011);
			21197: out = 16'(8445);
			21198: out = 16'(1088);
			21199: out = 16'(-3891);
			21200: out = 16'(-3134);
			21201: out = 16'(-268);
			21202: out = 16'(-823);
			21203: out = 16'(-3545);
			21204: out = 16'(-4977);
			21205: out = 16'(-1874);
			21206: out = 16'(4111);
			21207: out = 16'(6572);
			21208: out = 16'(2799);
			21209: out = 16'(-2498);
			21210: out = 16'(-1248);
			21211: out = 16'(-3526);
			21212: out = 16'(-7005);
			21213: out = 16'(-6105);
			21214: out = 16'(2562);
			21215: out = 16'(7112);
			21216: out = 16'(4082);
			21217: out = 16'(-1411);
			21218: out = 16'(-1689);
			21219: out = 16'(-1414);
			21220: out = 16'(-346);
			21221: out = 16'(1160);
			21222: out = 16'(3376);
			21223: out = 16'(593);
			21224: out = 16'(-6348);
			21225: out = 16'(-10193);
			21226: out = 16'(-3743);
			21227: out = 16'(2398);
			21228: out = 16'(6644);
			21229: out = 16'(3334);
			21230: out = 16'(191);
			21231: out = 16'(1660);
			21232: out = 16'(3793);
			21233: out = 16'(130);
			21234: out = 16'(-4092);
			21235: out = 16'(-631);
			21236: out = 16'(1988);
			21237: out = 16'(2727);
			21238: out = 16'(1197);
			21239: out = 16'(-66);
			21240: out = 16'(-3327);
			21241: out = 16'(-3309);
			21242: out = 16'(216);
			21243: out = 16'(3833);
			21244: out = 16'(5266);
			21245: out = 16'(2850);
			21246: out = 16'(1510);
			21247: out = 16'(2053);
			21248: out = 16'(5773);
			21249: out = 16'(-1283);
			21250: out = 16'(-6383);
			21251: out = 16'(-6234);
			21252: out = 16'(-69);
			21253: out = 16'(-2892);
			21254: out = 16'(1298);
			21255: out = 16'(6827);
			21256: out = 16'(5199);
			21257: out = 16'(719);
			21258: out = 16'(208);
			21259: out = 16'(1573);
			21260: out = 16'(-1384);
			21261: out = 16'(-8162);
			21262: out = 16'(-4838);
			21263: out = 16'(3233);
			21264: out = 16'(4014);
			21265: out = 16'(1640);
			21266: out = 16'(-2948);
			21267: out = 16'(-327);
			21268: out = 16'(3475);
			21269: out = 16'(1675);
			21270: out = 16'(-1431);
			21271: out = 16'(-1461);
			21272: out = 16'(-215);
			21273: out = 16'(-2370);
			21274: out = 16'(-2968);
			21275: out = 16'(-85);
			21276: out = 16'(6271);
			21277: out = 16'(10215);
			21278: out = 16'(5806);
			21279: out = 16'(-261);
			21280: out = 16'(-6285);
			21281: out = 16'(-10788);
			21282: out = 16'(-8440);
			21283: out = 16'(-2065);
			21284: out = 16'(5776);
			21285: out = 16'(7727);
			21286: out = 16'(2177);
			21287: out = 16'(-3252);
			21288: out = 16'(-2811);
			21289: out = 16'(-920);
			21290: out = 16'(-6362);
			21291: out = 16'(-3239);
			21292: out = 16'(1385);
			21293: out = 16'(4952);
			21294: out = 16'(3774);
			21295: out = 16'(2253);
			21296: out = 16'(202);
			21297: out = 16'(-1198);
			21298: out = 16'(-3775);
			21299: out = 16'(-4728);
			21300: out = 16'(-4515);
			21301: out = 16'(-219);
			21302: out = 16'(3663);
			21303: out = 16'(3583);
			21304: out = 16'(-1409);
			21305: out = 16'(-1950);
			21306: out = 16'(3867);
			21307: out = 16'(8755);
			21308: out = 16'(5264);
			21309: out = 16'(-1241);
			21310: out = 16'(-4980);
			21311: out = 16'(-5569);
			21312: out = 16'(-6703);
			21313: out = 16'(-7843);
			21314: out = 16'(-3751);
			21315: out = 16'(5454);
			21316: out = 16'(8956);
			21317: out = 16'(5319);
			21318: out = 16'(-1249);
			21319: out = 16'(-2435);
			21320: out = 16'(-953);
			21321: out = 16'(843);
			21322: out = 16'(-3630);
			21323: out = 16'(-5807);
			21324: out = 16'(2253);
			21325: out = 16'(7060);
			21326: out = 16'(2527);
			21327: out = 16'(-4358);
			21328: out = 16'(-2490);
			21329: out = 16'(4086);
			21330: out = 16'(3786);
			21331: out = 16'(-3543);
			21332: out = 16'(-7253);
			21333: out = 16'(-216);
			21334: out = 16'(7239);
			21335: out = 16'(6662);
			21336: out = 16'(721);
			21337: out = 16'(-77);
			21338: out = 16'(-610);
			21339: out = 16'(196);
			21340: out = 16'(654);
			21341: out = 16'(3395);
			21342: out = 16'(912);
			21343: out = 16'(-33);
			21344: out = 16'(-1392);
			21345: out = 16'(-3195);
			21346: out = 16'(-5443);
			21347: out = 16'(-2467);
			21348: out = 16'(0);
			21349: out = 16'(-1502);
			21350: out = 16'(-5826);
			21351: out = 16'(-1127);
			21352: out = 16'(3060);
			21353: out = 16'(-1110);
			21354: out = 16'(-2243);
			21355: out = 16'(386);
			21356: out = 16'(6371);
			21357: out = 16'(5895);
			21358: out = 16'(2434);
			21359: out = 16'(-4260);
			21360: out = 16'(-4398);
			21361: out = 16'(-3590);
			21362: out = 16'(-3577);
			21363: out = 16'(-5855);
			21364: out = 16'(2333);
			21365: out = 16'(7942);
			21366: out = 16'(821);
			21367: out = 16'(-3868);
			21368: out = 16'(-2442);
			21369: out = 16'(1689);
			21370: out = 16'(-551);
			21371: out = 16'(2252);
			21372: out = 16'(299);
			21373: out = 16'(-834);
			21374: out = 16'(-2001);
			21375: out = 16'(1989);
			21376: out = 16'(371);
			21377: out = 16'(-399);
			21378: out = 16'(-1489);
			21379: out = 16'(-862);
			21380: out = 16'(-4525);
			21381: out = 16'(-2706);
			21382: out = 16'(1370);
			21383: out = 16'(2627);
			21384: out = 16'(2163);
			21385: out = 16'(2664);
			21386: out = 16'(3889);
			21387: out = 16'(2877);
			21388: out = 16'(620);
			21389: out = 16'(-4105);
			21390: out = 16'(-6399);
			21391: out = 16'(-4044);
			21392: out = 16'(-381);
			21393: out = 16'(530);
			21394: out = 16'(-903);
			21395: out = 16'(594);
			21396: out = 16'(7086);
			21397: out = 16'(4502);
			21398: out = 16'(-1754);
			21399: out = 16'(-4080);
			21400: out = 16'(2051);
			21401: out = 16'(3343);
			21402: out = 16'(1605);
			21403: out = 16'(-48);
			21404: out = 16'(2333);
			21405: out = 16'(6475);
			21406: out = 16'(3906);
			21407: out = 16'(-3330);
			21408: out = 16'(-8160);
			21409: out = 16'(-5613);
			21410: out = 16'(-4695);
			21411: out = 16'(-5405);
			21412: out = 16'(-3085);
			21413: out = 16'(5648);
			21414: out = 16'(7706);
			21415: out = 16'(4110);
			21416: out = 16'(-912);
			21417: out = 16'(427);
			21418: out = 16'(59);
			21419: out = 16'(1625);
			21420: out = 16'(1148);
			21421: out = 16'(841);
			21422: out = 16'(-1593);
			21423: out = 16'(2718);
			21424: out = 16'(4470);
			21425: out = 16'(439);
			21426: out = 16'(-8353);
			21427: out = 16'(-3781);
			21428: out = 16'(3308);
			21429: out = 16'(1491);
			21430: out = 16'(-6957);
			21431: out = 16'(-4487);
			21432: out = 16'(4652);
			21433: out = 16'(8217);
			21434: out = 16'(4378);
			21435: out = 16'(367);
			21436: out = 16'(-16);
			21437: out = 16'(-2699);
			21438: out = 16'(-10578);
			21439: out = 16'(-12625);
			21440: out = 16'(-7376);
			21441: out = 16'(-1001);
			21442: out = 16'(-828);
			21443: out = 16'(3787);
			21444: out = 16'(5272);
			21445: out = 16'(6165);
			21446: out = 16'(3522);
			21447: out = 16'(2563);
			21448: out = 16'(-5943);
			21449: out = 16'(-10154);
			21450: out = 16'(-7013);
			21451: out = 16'(2000);
			21452: out = 16'(5442);
			21453: out = 16'(5980);
			21454: out = 16'(3043);
			21455: out = 16'(194);
			21456: out = 16'(-4605);
			21457: out = 16'(-2076);
			21458: out = 16'(-89);
			21459: out = 16'(-3064);
			21460: out = 16'(-4670);
			21461: out = 16'(1650);
			21462: out = 16'(8830);
			21463: out = 16'(8462);
			21464: out = 16'(1057);
			21465: out = 16'(-48);
			21466: out = 16'(923);
			21467: out = 16'(-1054);
			21468: out = 16'(-2436);
			21469: out = 16'(-2246);
			21470: out = 16'(1986);
			21471: out = 16'(4144);
			21472: out = 16'(1783);
			21473: out = 16'(-2248);
			21474: out = 16'(-2157);
			21475: out = 16'(508);
			21476: out = 16'(-519);
			21477: out = 16'(-1324);
			21478: out = 16'(-4502);
			21479: out = 16'(-3791);
			21480: out = 16'(699);
			21481: out = 16'(5093);
			21482: out = 16'(5550);
			21483: out = 16'(5622);
			21484: out = 16'(6282);
			21485: out = 16'(8172);
			21486: out = 16'(-3269);
			21487: out = 16'(-14408);
			21488: out = 16'(-16170);
			21489: out = 16'(-5155);
			21490: out = 16'(1282);
			21491: out = 16'(6087);
			21492: out = 16'(7808);
			21493: out = 16'(5936);
			21494: out = 16'(2493);
			21495: out = 16'(618);
			21496: out = 16'(-1641);
			21497: out = 16'(-5329);
			21498: out = 16'(59);
			21499: out = 16'(465);
			21500: out = 16'(-1612);
			21501: out = 16'(-2237);
			21502: out = 16'(5694);
			21503: out = 16'(2469);
			21504: out = 16'(-3204);
			21505: out = 16'(-3726);
			21506: out = 16'(4068);
			21507: out = 16'(3141);
			21508: out = 16'(-2103);
			21509: out = 16'(-4921);
			21510: out = 16'(-809);
			21511: out = 16'(4974);
			21512: out = 16'(6631);
			21513: out = 16'(4835);
			21514: out = 16'(1079);
			21515: out = 16'(413);
			21516: out = 16'(-3985);
			21517: out = 16'(-4116);
			21518: out = 16'(530);
			21519: out = 16'(3257);
			21520: out = 16'(208);
			21521: out = 16'(-1434);
			21522: out = 16'(-897);
			21523: out = 16'(-5314);
			21524: out = 16'(-5788);
			21525: out = 16'(-2013);
			21526: out = 16'(3075);
			21527: out = 16'(4293);
			21528: out = 16'(2362);
			21529: out = 16'(845);
			21530: out = 16'(-1662);
			21531: out = 16'(-4896);
			21532: out = 16'(282);
			21533: out = 16'(5608);
			21534: out = 16'(1711);
			21535: out = 16'(-9155);
			21536: out = 16'(-5685);
			21537: out = 16'(-189);
			21538: out = 16'(772);
			21539: out = 16'(-3353);
			21540: out = 16'(393);
			21541: out = 16'(3879);
			21542: out = 16'(5391);
			21543: out = 16'(2735);
			21544: out = 16'(2108);
			21545: out = 16'(55);
			21546: out = 16'(-666);
			21547: out = 16'(-1319);
			21548: out = 16'(-116);
			21549: out = 16'(-281);
			21550: out = 16'(1036);
			21551: out = 16'(1427);
			21552: out = 16'(-747);
			21553: out = 16'(-13);
			21554: out = 16'(-717);
			21555: out = 16'(2062);
			21556: out = 16'(5371);
			21557: out = 16'(6054);
			21558: out = 16'(1103);
			21559: out = 16'(-1359);
			21560: out = 16'(-2238);
			21561: out = 16'(-4234);
			21562: out = 16'(-6883);
			21563: out = 16'(-523);
			21564: out = 16'(7750);
			21565: out = 16'(6336);
			21566: out = 16'(-5332);
			21567: out = 16'(-11195);
			21568: out = 16'(-6066);
			21569: out = 16'(2478);
			21570: out = 16'(4901);
			21571: out = 16'(7104);
			21572: out = 16'(5307);
			21573: out = 16'(-1501);
			21574: out = 16'(-2709);
			21575: out = 16'(-4106);
			21576: out = 16'(-1673);
			21577: out = 16'(35);
			21578: out = 16'(1952);
			21579: out = 16'(-155);
			21580: out = 16'(678);
			21581: out = 16'(1872);
			21582: out = 16'(2629);
			21583: out = 16'(-3398);
			21584: out = 16'(-2655);
			21585: out = 16'(-260);
			21586: out = 16'(-2794);
			21587: out = 16'(-2938);
			21588: out = 16'(-2352);
			21589: out = 16'(-477);
			21590: out = 16'(688);
			21591: out = 16'(8738);
			21592: out = 16'(4628);
			21593: out = 16'(-1956);
			21594: out = 16'(-5064);
			21595: out = 16'(-414);
			21596: out = 16'(-696);
			21597: out = 16'(-3370);
			21598: out = 16'(-5293);
			21599: out = 16'(-2980);
			21600: out = 16'(-652);
			21601: out = 16'(800);
			21602: out = 16'(530);
			21603: out = 16'(-36);
			21604: out = 16'(1687);
			21605: out = 16'(8);
			21606: out = 16'(-4285);
			21607: out = 16'(-6281);
			21608: out = 16'(3530);
			21609: out = 16'(3953);
			21610: out = 16'(-1233);
			21611: out = 16'(-4605);
			21612: out = 16'(-74);
			21613: out = 16'(5973);
			21614: out = 16'(7456);
			21615: out = 16'(1072);
			21616: out = 16'(-12600);
			21617: out = 16'(-11115);
			21618: out = 16'(-4218);
			21619: out = 16'(2665);
			21620: out = 16'(6533);
			21621: out = 16'(6713);
			21622: out = 16'(3209);
			21623: out = 16'(-2762);
			21624: out = 16'(-8225);
			21625: out = 16'(-5381);
			21626: out = 16'(-441);
			21627: out = 16'(4663);
			21628: out = 16'(6027);
			21629: out = 16'(2590);
			21630: out = 16'(471);
			21631: out = 16'(313);
			21632: out = 16'(-19);
			21633: out = 16'(574);
			21634: out = 16'(1034);
			21635: out = 16'(4776);
			21636: out = 16'(4961);
			21637: out = 16'(-69);
			21638: out = 16'(-4781);
			21639: out = 16'(-1146);
			21640: out = 16'(4422);
			21641: out = 16'(4834);
			21642: out = 16'(532);
			21643: out = 16'(-355);
			21644: out = 16'(-1641);
			21645: out = 16'(-4501);
			21646: out = 16'(-3379);
			21647: out = 16'(461);
			21648: out = 16'(1567);
			21649: out = 16'(-28);
			21650: out = 16'(1915);
			21651: out = 16'(4016);
			21652: out = 16'(2635);
			21653: out = 16'(-648);
			21654: out = 16'(139);
			21655: out = 16'(-1058);
			21656: out = 16'(-874);
			21657: out = 16'(1778);
			21658: out = 16'(5777);
			21659: out = 16'(1059);
			21660: out = 16'(-5534);
			21661: out = 16'(-8354);
			21662: out = 16'(-4147);
			21663: out = 16'(1212);
			21664: out = 16'(2920);
			21665: out = 16'(2556);
			21666: out = 16'(1099);
			21667: out = 16'(-2671);
			21668: out = 16'(-5112);
			21669: out = 16'(-2126);
			21670: out = 16'(3434);
			21671: out = 16'(6002);
			21672: out = 16'(1483);
			21673: out = 16'(-1338);
			21674: out = 16'(-3580);
			21675: out = 16'(-8263);
			21676: out = 16'(-4178);
			21677: out = 16'(1980);
			21678: out = 16'(3859);
			21679: out = 16'(-1565);
			21680: out = 16'(1129);
			21681: out = 16'(423);
			21682: out = 16'(-179);
			21683: out = 16'(-123);
			21684: out = 16'(8276);
			21685: out = 16'(3179);
			21686: out = 16'(-4271);
			21687: out = 16'(-7600);
			21688: out = 16'(-84);
			21689: out = 16'(50);
			21690: out = 16'(-464);
			21691: out = 16'(-992);
			21692: out = 16'(273);
			21693: out = 16'(1452);
			21694: out = 16'(3493);
			21695: out = 16'(1866);
			21696: out = 16'(-4273);
			21697: out = 16'(-519);
			21698: out = 16'(1372);
			21699: out = 16'(1364);
			21700: out = 16'(-1651);
			21701: out = 16'(-1570);
			21702: out = 16'(-1978);
			21703: out = 16'(1322);
			21704: out = 16'(3122);
			21705: out = 16'(-1649);
			21706: out = 16'(-3364);
			21707: out = 16'(230);
			21708: out = 16'(3696);
			21709: out = 16'(-254);
			21710: out = 16'(0);
			21711: out = 16'(2003);
			21712: out = 16'(3314);
			21713: out = 16'(-382);
			21714: out = 16'(846);
			21715: out = 16'(1285);
			21716: out = 16'(1342);
			21717: out = 16'(-2079);
			21718: out = 16'(-4408);
			21719: out = 16'(-3676);
			21720: out = 16'(3525);
			21721: out = 16'(9693);
			21722: out = 16'(11318);
			21723: out = 16'(2961);
			21724: out = 16'(-2148);
			21725: out = 16'(-2284);
			21726: out = 16'(-1493);
			21727: out = 16'(-726);
			21728: out = 16'(1715);
			21729: out = 16'(2827);
			21730: out = 16'(-420);
			21731: out = 16'(-629);
			21732: out = 16'(1187);
			21733: out = 16'(1909);
			21734: out = 16'(-796);
			21735: out = 16'(178);
			21736: out = 16'(229);
			21737: out = 16'(-3279);
			21738: out = 16'(-8701);
			21739: out = 16'(-968);
			21740: out = 16'(3533);
			21741: out = 16'(5003);
			21742: out = 16'(2472);
			21743: out = 16'(1809);
			21744: out = 16'(-1065);
			21745: out = 16'(-2667);
			21746: out = 16'(-3464);
			21747: out = 16'(-176);
			21748: out = 16'(694);
			21749: out = 16'(3005);
			21750: out = 16'(2081);
			21751: out = 16'(-582);
			21752: out = 16'(-6355);
			21753: out = 16'(-3303);
			21754: out = 16'(218);
			21755: out = 16'(-498);
			21756: out = 16'(-429);
			21757: out = 16'(959);
			21758: out = 16'(1119);
			21759: out = 16'(-884);
			21760: out = 16'(-3304);
			21761: out = 16'(223);
			21762: out = 16'(1442);
			21763: out = 16'(-1617);
			21764: out = 16'(-5194);
			21765: out = 16'(-1695);
			21766: out = 16'(696);
			21767: out = 16'(219);
			21768: out = 16'(176);
			21769: out = 16'(1250);
			21770: out = 16'(3507);
			21771: out = 16'(3819);
			21772: out = 16'(946);
			21773: out = 16'(-793);
			21774: out = 16'(-5766);
			21775: out = 16'(-7345);
			21776: out = 16'(-4429);
			21777: out = 16'(-217);
			21778: out = 16'(-8);
			21779: out = 16'(2205);
			21780: out = 16'(6083);
			21781: out = 16'(4712);
			21782: out = 16'(1549);
			21783: out = 16'(-4326);
			21784: out = 16'(-8040);
			21785: out = 16'(-6945);
			21786: out = 16'(-1352);
			21787: out = 16'(2753);
			21788: out = 16'(3562);
			21789: out = 16'(3014);
			21790: out = 16'(5764);
			21791: out = 16'(2756);
			21792: out = 16'(-3698);
			21793: out = 16'(-6549);
			21794: out = 16'(992);
			21795: out = 16'(1315);
			21796: out = 16'(-3721);
			21797: out = 16'(-4383);
			21798: out = 16'(5904);
			21799: out = 16'(8758);
			21800: out = 16'(2782);
			21801: out = 16'(-5007);
			21802: out = 16'(-4823);
			21803: out = 16'(392);
			21804: out = 16'(1493);
			21805: out = 16'(-772);
			21806: out = 16'(405);
			21807: out = 16'(2743);
			21808: out = 16'(4667);
			21809: out = 16'(2296);
			21810: out = 16'(-1950);
			21811: out = 16'(-2220);
			21812: out = 16'(-2008);
			21813: out = 16'(-641);
			21814: out = 16'(-997);
			21815: out = 16'(-2865);
			21816: out = 16'(-1746);
			21817: out = 16'(4105);
			21818: out = 16'(7385);
			21819: out = 16'(4088);
			21820: out = 16'(137);
			21821: out = 16'(502);
			21822: out = 16'(537);
			21823: out = 16'(-4170);
			21824: out = 16'(-9215);
			21825: out = 16'(-4893);
			21826: out = 16'(1829);
			21827: out = 16'(1503);
			21828: out = 16'(6495);
			21829: out = 16'(2021);
			21830: out = 16'(-91);
			21831: out = 16'(-272);
			21832: out = 16'(2769);
			21833: out = 16'(-1397);
			21834: out = 16'(-961);
			21835: out = 16'(2396);
			21836: out = 16'(2181);
			21837: out = 16'(530);
			21838: out = 16'(-712);
			21839: out = 16'(271);
			21840: out = 16'(96);
			21841: out = 16'(-767);
			21842: out = 16'(-4259);
			21843: out = 16'(-3993);
			21844: out = 16'(1476);
			21845: out = 16'(3037);
			21846: out = 16'(2762);
			21847: out = 16'(402);
			21848: out = 16'(45);
			21849: out = 16'(1252);
			21850: out = 16'(3926);
			21851: out = 16'(2592);
			21852: out = 16'(-128);
			21853: out = 16'(-517);
			21854: out = 16'(3122);
			21855: out = 16'(3590);
			21856: out = 16'(1046);
			21857: out = 16'(-1796);
			21858: out = 16'(-851);
			21859: out = 16'(-2379);
			21860: out = 16'(-3205);
			21861: out = 16'(357);
			21862: out = 16'(2507);
			21863: out = 16'(2787);
			21864: out = 16'(-1552);
			21865: out = 16'(-5467);
			21866: out = 16'(-720);
			21867: out = 16'(1136);
			21868: out = 16'(779);
			21869: out = 16'(-136);
			21870: out = 16'(3318);
			21871: out = 16'(-427);
			21872: out = 16'(-3817);
			21873: out = 16'(-5711);
			21874: out = 16'(-3076);
			21875: out = 16'(-5653);
			21876: out = 16'(-223);
			21877: out = 16'(6956);
			21878: out = 16'(8926);
			21879: out = 16'(1040);
			21880: out = 16'(-4493);
			21881: out = 16'(-8281);
			21882: out = 16'(-8814);
			21883: out = 16'(-1014);
			21884: out = 16'(5896);
			21885: out = 16'(5389);
			21886: out = 16'(-2074);
			21887: out = 16'(-5548);
			21888: out = 16'(-3594);
			21889: out = 16'(2568);
			21890: out = 16'(3295);
			21891: out = 16'(-909);
			21892: out = 16'(-1902);
			21893: out = 16'(2262);
			21894: out = 16'(3378);
			21895: out = 16'(-1751);
			21896: out = 16'(-4967);
			21897: out = 16'(-2158);
			21898: out = 16'(1860);
			21899: out = 16'(1515);
			21900: out = 16'(1900);
			21901: out = 16'(1815);
			21902: out = 16'(-507);
			21903: out = 16'(-6811);
			21904: out = 16'(-8797);
			21905: out = 16'(-5987);
			21906: out = 16'(3262);
			21907: out = 16'(9074);
			21908: out = 16'(7572);
			21909: out = 16'(652);
			21910: out = 16'(-1936);
			21911: out = 16'(-1152);
			21912: out = 16'(-2470);
			21913: out = 16'(-2952);
			21914: out = 16'(-164);
			21915: out = 16'(4386);
			21916: out = 16'(3662);
			21917: out = 16'(2761);
			21918: out = 16'(115);
			21919: out = 16'(2574);
			21920: out = 16'(3253);
			21921: out = 16'(-333);
			21922: out = 16'(-9169);
			21923: out = 16'(-7077);
			21924: out = 16'(1567);
			21925: out = 16'(3384);
			21926: out = 16'(592);
			21927: out = 16'(2368);
			21928: out = 16'(4489);
			21929: out = 16'(-1913);
			21930: out = 16'(-6514);
			21931: out = 16'(-3158);
			21932: out = 16'(3974);
			21933: out = 16'(3759);
			21934: out = 16'(4900);
			21935: out = 16'(2372);
			21936: out = 16'(622);
			21937: out = 16'(-1433);
			21938: out = 16'(3329);
			21939: out = 16'(1366);
			21940: out = 16'(-659);
			21941: out = 16'(-1490);
			21942: out = 16'(-314);
			21943: out = 16'(-484);
			21944: out = 16'(-617);
			21945: out = 16'(916);
			21946: out = 16'(5963);
			21947: out = 16'(5776);
			21948: out = 16'(3592);
			21949: out = 16'(-287);
			21950: out = 16'(-2920);
			21951: out = 16'(-8288);
			21952: out = 16'(-8679);
			21953: out = 16'(-5381);
			21954: out = 16'(990);
			21955: out = 16'(2609);
			21956: out = 16'(8022);
			21957: out = 16'(5810);
			21958: out = 16'(-1826);
			21959: out = 16'(-4086);
			21960: out = 16'(-5597);
			21961: out = 16'(-4828);
			21962: out = 16'(-1115);
			21963: out = 16'(7524);
			21964: out = 16'(5941);
			21965: out = 16'(1079);
			21966: out = 16'(-2931);
			21967: out = 16'(-259);
			21968: out = 16'(-6087);
			21969: out = 16'(-5114);
			21970: out = 16'(-1445);
			21971: out = 16'(2045);
			21972: out = 16'(1604);
			21973: out = 16'(1931);
			21974: out = 16'(540);
			21975: out = 16'(-1458);
			21976: out = 16'(-174);
			21977: out = 16'(2388);
			21978: out = 16'(2480);
			21979: out = 16'(-1640);
			21980: out = 16'(-2794);
			21981: out = 16'(-7348);
			21982: out = 16'(-4035);
			21983: out = 16'(1959);
			21984: out = 16'(6170);
			21985: out = 16'(3740);
			21986: out = 16'(1787);
			21987: out = 16'(-3194);
			21988: out = 16'(-8694);
			21989: out = 16'(-11368);
			21990: out = 16'(-2605);
			21991: out = 16'(2572);
			21992: out = 16'(-689);
			21993: out = 16'(-2608);
			21994: out = 16'(2081);
			21995: out = 16'(5399);
			21996: out = 16'(2007);
			21997: out = 16'(-3724);
			21998: out = 16'(-5212);
			21999: out = 16'(-4732);
			22000: out = 16'(-2778);
			22001: out = 16'(1007);
			22002: out = 16'(2472);
			22003: out = 16'(-1683);
			22004: out = 16'(-4521);
			22005: out = 16'(1573);
			22006: out = 16'(10093);
			22007: out = 16'(7378);
			22008: out = 16'(-4737);
			22009: out = 16'(-13206);
			22010: out = 16'(-1258);
			22011: out = 16'(4555);
			22012: out = 16'(1875);
			22013: out = 16'(-2860);
			22014: out = 16'(2426);
			22015: out = 16'(681);
			22016: out = 16'(188);
			22017: out = 16'(37);
			22018: out = 16'(469);
			22019: out = 16'(-23);
			22020: out = 16'(2330);
			22021: out = 16'(3291);
			22022: out = 16'(-400);
			22023: out = 16'(20);
			22024: out = 16'(1087);
			22025: out = 16'(1808);
			22026: out = 16'(-651);
			22027: out = 16'(541);
			22028: out = 16'(-1169);
			22029: out = 16'(242);
			22030: out = 16'(2116);
			22031: out = 16'(3893);
			22032: out = 16'(460);
			22033: out = 16'(1706);
			22034: out = 16'(4478);
			22035: out = 16'(1373);
			22036: out = 16'(-4479);
			22037: out = 16'(-6952);
			22038: out = 16'(-3122);
			22039: out = 16'(1916);
			22040: out = 16'(2058);
			22041: out = 16'(1764);
			22042: out = 16'(2182);
			22043: out = 16'(2722);
			22044: out = 16'(1794);
			22045: out = 16'(1826);
			22046: out = 16'(1003);
			22047: out = 16'(-629);
			22048: out = 16'(-1347);
			22049: out = 16'(-1917);
			22050: out = 16'(-3047);
			22051: out = 16'(-1624);
			22052: out = 16'(5935);
			22053: out = 16'(4011);
			22054: out = 16'(-2172);
			22055: out = 16'(-5515);
			22056: out = 16'(3432);
			22057: out = 16'(-73);
			22058: out = 16'(-1344);
			22059: out = 16'(-4930);
			22060: out = 16'(-5380);
			22061: out = 16'(-1738);
			22062: out = 16'(6914);
			22063: out = 16'(7246);
			22064: out = 16'(367);
			22065: out = 16'(-6822);
			22066: out = 16'(-2215);
			22067: out = 16'(1435);
			22068: out = 16'(-491);
			22069: out = 16'(362);
			22070: out = 16'(4483);
			22071: out = 16'(5172);
			22072: out = 16'(-1469);
			22073: out = 16'(-9261);
			22074: out = 16'(-9486);
			22075: out = 16'(-3724);
			22076: out = 16'(2515);
			22077: out = 16'(6389);
			22078: out = 16'(4847);
			22079: out = 16'(2428);
			22080: out = 16'(-1240);
			22081: out = 16'(-4265);
			22082: out = 16'(-2310);
			22083: out = 16'(-600);
			22084: out = 16'(353);
			22085: out = 16'(-90);
			22086: out = 16'(286);
			22087: out = 16'(-240);
			22088: out = 16'(95);
			22089: out = 16'(-568);
			22090: out = 16'(-729);
			22091: out = 16'(-612);
			22092: out = 16'(2968);
			22093: out = 16'(3685);
			22094: out = 16'(-393);
			22095: out = 16'(-7339);
			22096: out = 16'(-4829);
			22097: out = 16'(1013);
			22098: out = 16'(1672);
			22099: out = 16'(583);
			22100: out = 16'(2740);
			22101: out = 16'(5428);
			22102: out = 16'(3734);
			22103: out = 16'(3307);
			22104: out = 16'(23);
			22105: out = 16'(656);
			22106: out = 16'(1877);
			22107: out = 16'(2674);
			22108: out = 16'(-3800);
			22109: out = 16'(-4402);
			22110: out = 16'(-1943);
			22111: out = 16'(-4655);
			22112: out = 16'(-4638);
			22113: out = 16'(-1910);
			22114: out = 16'(6206);
			22115: out = 16'(10637);
			22116: out = 16'(5860);
			22117: out = 16'(-1346);
			22118: out = 16'(-2054);
			22119: out = 16'(167);
			22120: out = 16'(-3603);
			22121: out = 16'(-9345);
			22122: out = 16'(-7064);
			22123: out = 16'(2744);
			22124: out = 16'(9614);
			22125: out = 16'(6180);
			22126: out = 16'(2675);
			22127: out = 16'(1624);
			22128: out = 16'(1687);
			22129: out = 16'(-3449);
			22130: out = 16'(-3465);
			22131: out = 16'(-2555);
			22132: out = 16'(-3853);
			22133: out = 16'(780);
			22134: out = 16'(6223);
			22135: out = 16'(4876);
			22136: out = 16'(-3407);
			22137: out = 16'(-5981);
			22138: out = 16'(-1287);
			22139: out = 16'(3248);
			22140: out = 16'(2167);
			22141: out = 16'(2047);
			22142: out = 16'(1674);
			22143: out = 16'(-268);
			22144: out = 16'(-3358);
			22145: out = 16'(398);
			22146: out = 16'(-501);
			22147: out = 16'(-162);
			22148: out = 16'(-2807);
			22149: out = 16'(-5758);
			22150: out = 16'(-2342);
			22151: out = 16'(2731);
			22152: out = 16'(3937);
			22153: out = 16'(1651);
			22154: out = 16'(2566);
			22155: out = 16'(3754);
			22156: out = 16'(3065);
			22157: out = 16'(-1600);
			22158: out = 16'(-6350);
			22159: out = 16'(-10122);
			22160: out = 16'(-7234);
			22161: out = 16'(729);
			22162: out = 16'(8097);
			22163: out = 16'(12152);
			22164: out = 16'(9819);
			22165: out = 16'(2808);
			22166: out = 16'(-3348);
			22167: out = 16'(-13532);
			22168: out = 16'(-13728);
			22169: out = 16'(-6835);
			22170: out = 16'(957);
			22171: out = 16'(3190);
			22172: out = 16'(7044);
			22173: out = 16'(7437);
			22174: out = 16'(3422);
			22175: out = 16'(471);
			22176: out = 16'(-1751);
			22177: out = 16'(-1596);
			22178: out = 16'(-30);
			22179: out = 16'(-1488);
			22180: out = 16'(-23);
			22181: out = 16'(-1428);
			22182: out = 16'(-898);
			22183: out = 16'(3346);
			22184: out = 16'(3964);
			22185: out = 16'(1071);
			22186: out = 16'(1354);
			22187: out = 16'(5403);
			22188: out = 16'(1070);
			22189: out = 16'(-7279);
			22190: out = 16'(-7783);
			22191: out = 16'(3223);
			22192: out = 16'(5141);
			22193: out = 16'(2295);
			22194: out = 16'(-2174);
			22195: out = 16'(-1861);
			22196: out = 16'(-1769);
			22197: out = 16'(-346);
			22198: out = 16'(-946);
			22199: out = 16'(-722);
			22200: out = 16'(2770);
			22201: out = 16'(3557);
			22202: out = 16'(5440);
			22203: out = 16'(3979);
			22204: out = 16'(-1995);
			22205: out = 16'(-11333);
			22206: out = 16'(-11411);
			22207: out = 16'(-5999);
			22208: out = 16'(-2724);
			22209: out = 16'(-73);
			22210: out = 16'(3139);
			22211: out = 16'(4136);
			22212: out = 16'(1699);
			22213: out = 16'(4590);
			22214: out = 16'(2531);
			22215: out = 16'(-224);
			22216: out = 16'(-4048);
			22217: out = 16'(-4683);
			22218: out = 16'(-6378);
			22219: out = 16'(-2210);
			22220: out = 16'(3494);
			22221: out = 16'(4035);
			22222: out = 16'(2798);
			22223: out = 16'(-203);
			22224: out = 16'(-1075);
			22225: out = 16'(-1273);
			22226: out = 16'(915);
			22227: out = 16'(-1856);
			22228: out = 16'(-2266);
			22229: out = 16'(53);
			22230: out = 16'(0);
			22231: out = 16'(-290);
			22232: out = 16'(2725);
			22233: out = 16'(6216);
			22234: out = 16'(4242);
			22235: out = 16'(1464);
			22236: out = 16'(13);
			22237: out = 16'(-1255);
			22238: out = 16'(-4138);
			22239: out = 16'(-7013);
			22240: out = 16'(-2587);
			22241: out = 16'(4030);
			22242: out = 16'(5508);
			22243: out = 16'(797);
			22244: out = 16'(-396);
			22245: out = 16'(-1621);
			22246: out = 16'(-5230);
			22247: out = 16'(-307);
			22248: out = 16'(2339);
			22249: out = 16'(3757);
			22250: out = 16'(1923);
			22251: out = 16'(330);
			22252: out = 16'(2744);
			22253: out = 16'(5129);
			22254: out = 16'(2221);
			22255: out = 16'(-2971);
			22256: out = 16'(-7125);
			22257: out = 16'(-3744);
			22258: out = 16'(1717);
			22259: out = 16'(4264);
			22260: out = 16'(3423);
			22261: out = 16'(4788);
			22262: out = 16'(5281);
			22263: out = 16'(2321);
			22264: out = 16'(-1838);
			22265: out = 16'(-3529);
			22266: out = 16'(-3296);
			22267: out = 16'(-4037);
			22268: out = 16'(-8071);
			22269: out = 16'(-387);
			22270: out = 16'(7399);
			22271: out = 16'(7010);
			22272: out = 16'(-45);
			22273: out = 16'(-1573);
			22274: out = 16'(-1067);
			22275: out = 16'(-3003);
			22276: out = 16'(-7128);
			22277: out = 16'(-6035);
			22278: out = 16'(1324);
			22279: out = 16'(8204);
			22280: out = 16'(8595);
			22281: out = 16'(2484);
			22282: out = 16'(-224);
			22283: out = 16'(-272);
			22284: out = 16'(-1131);
			22285: out = 16'(-4178);
			22286: out = 16'(-3804);
			22287: out = 16'(-4300);
			22288: out = 16'(-6211);
			22289: out = 16'(-555);
			22290: out = 16'(1076);
			22291: out = 16'(6324);
			22292: out = 16'(6808);
			22293: out = 16'(2247);
			22294: out = 16'(-7889);
			22295: out = 16'(-5707);
			22296: out = 16'(362);
			22297: out = 16'(-755);
			22298: out = 16'(-3276);
			22299: out = 16'(-1095);
			22300: out = 16'(3955);
			22301: out = 16'(3041);
			22302: out = 16'(-1977);
			22303: out = 16'(-8034);
			22304: out = 16'(-7778);
			22305: out = 16'(-3950);
			22306: out = 16'(-879);
			22307: out = 16'(-4524);
			22308: out = 16'(-2891);
			22309: out = 16'(5937);
			22310: out = 16'(12347);
			22311: out = 16'(9506);
			22312: out = 16'(697);
			22313: out = 16'(-4593);
			22314: out = 16'(-2508);
			22315: out = 16'(1325);
			22316: out = 16'(15);
			22317: out = 16'(-2684);
			22318: out = 16'(-802);
			22319: out = 16'(5212);
			22320: out = 16'(3109);
			22321: out = 16'(-4754);
			22322: out = 16'(-9600);
			22323: out = 16'(-2229);
			22324: out = 16'(219);
			22325: out = 16'(-991);
			22326: out = 16'(-2483);
			22327: out = 16'(652);
			22328: out = 16'(2967);
			22329: out = 16'(4308);
			22330: out = 16'(3042);
			22331: out = 16'(2059);
			22332: out = 16'(-830);
			22333: out = 16'(-1279);
			22334: out = 16'(-3927);
			22335: out = 16'(-7641);
			22336: out = 16'(-2574);
			22337: out = 16'(2841);
			22338: out = 16'(5108);
			22339: out = 16'(4520);
			22340: out = 16'(4528);
			22341: out = 16'(8250);
			22342: out = 16'(8218);
			22343: out = 16'(660);
			22344: out = 16'(-11982);
			22345: out = 16'(-7346);
			22346: out = 16'(2240);
			22347: out = 16'(5230);
			22348: out = 16'(-152);
			22349: out = 16'(1503);
			22350: out = 16'(1072);
			22351: out = 16'(-2431);
			22352: out = 16'(-6644);
			22353: out = 16'(1557);
			22354: out = 16'(4442);
			22355: out = 16'(2831);
			22356: out = 16'(-128);
			22357: out = 16'(1780);
			22358: out = 16'(468);
			22359: out = 16'(-464);
			22360: out = 16'(718);
			22361: out = 16'(3169);
			22362: out = 16'(4395);
			22363: out = 16'(2131);
			22364: out = 16'(-604);
			22365: out = 16'(-149);
			22366: out = 16'(-2593);
			22367: out = 16'(-4572);
			22368: out = 16'(-4069);
			22369: out = 16'(483);
			22370: out = 16'(-282);
			22371: out = 16'(2682);
			22372: out = 16'(4813);
			22373: out = 16'(3111);
			22374: out = 16'(-5139);
			22375: out = 16'(-5240);
			22376: out = 16'(1539);
			22377: out = 16'(7949);
			22378: out = 16'(6980);
			22379: out = 16'(1945);
			22380: out = 16'(-2633);
			22381: out = 16'(-2471);
			22382: out = 16'(1073);
			22383: out = 16'(-2618);
			22384: out = 16'(-8962);
			22385: out = 16'(-9835);
			22386: out = 16'(897);
			22387: out = 16'(-517);
			22388: out = 16'(1987);
			22389: out = 16'(2577);
			22390: out = 16'(2735);
			22391: out = 16'(-490);
			22392: out = 16'(2461);
			22393: out = 16'(2302);
			22394: out = 16'(-1052);
			22395: out = 16'(-7139);
			22396: out = 16'(-4098);
			22397: out = 16'(-4548);
			22398: out = 16'(-6151);
			22399: out = 16'(329);
			22400: out = 16'(3886);
			22401: out = 16'(2583);
			22402: out = 16'(-186);
			22403: out = 16'(2199);
			22404: out = 16'(2007);
			22405: out = 16'(-1772);
			22406: out = 16'(-5641);
			22407: out = 16'(-3075);
			22408: out = 16'(22);
			22409: out = 16'(2086);
			22410: out = 16'(1851);
			22411: out = 16'(1889);
			22412: out = 16'(148);
			22413: out = 16'(-3112);
			22414: out = 16'(-6331);
			22415: out = 16'(-6101);
			22416: out = 16'(-2797);
			22417: out = 16'(-142);
			22418: out = 16'(1499);
			22419: out = 16'(2447);
			22420: out = 16'(2124);
			22421: out = 16'(781);
			22422: out = 16'(171);
			22423: out = 16'(895);
			22424: out = 16'(2316);
			22425: out = 16'(2722);
			22426: out = 16'(4973);
			22427: out = 16'(6055);
			22428: out = 16'(3081);
			22429: out = 16'(-5050);
			22430: out = 16'(-5004);
			22431: out = 16'(-240);
			22432: out = 16'(1404);
			22433: out = 16'(-531);
			22434: out = 16'(-889);
			22435: out = 16'(3445);
			22436: out = 16'(5071);
			22437: out = 16'(138);
			22438: out = 16'(782);
			22439: out = 16'(6351);
			22440: out = 16'(8126);
			22441: out = 16'(701);
			22442: out = 16'(-929);
			22443: out = 16'(-2156);
			22444: out = 16'(-4161);
			22445: out = 16'(-8501);
			22446: out = 16'(-3566);
			22447: out = 16'(148);
			22448: out = 16'(2841);
			22449: out = 16'(3919);
			22450: out = 16'(7206);
			22451: out = 16'(5227);
			22452: out = 16'(1063);
			22453: out = 16'(-3713);
			22454: out = 16'(-6217);
			22455: out = 16'(-2812);
			22456: out = 16'(709);
			22457: out = 16'(1314);
			22458: out = 16'(-304);
			22459: out = 16'(-128);
			22460: out = 16'(-194);
			22461: out = 16'(-599);
			22462: out = 16'(-2312);
			22463: out = 16'(1670);
			22464: out = 16'(-804);
			22465: out = 16'(-3199);
			22466: out = 16'(-3859);
			22467: out = 16'(1871);
			22468: out = 16'(2);
			22469: out = 16'(2531);
			22470: out = 16'(6146);
			22471: out = 16'(5620);
			22472: out = 16'(-8347);
			22473: out = 16'(-13949);
			22474: out = 16'(-6518);
			22475: out = 16'(3452);
			22476: out = 16'(990);
			22477: out = 16'(1016);
			22478: out = 16'(4282);
			22479: out = 16'(5228);
			22480: out = 16'(-3679);
			22481: out = 16'(-4891);
			22482: out = 16'(-714);
			22483: out = 16'(1087);
			22484: out = 16'(-6257);
			22485: out = 16'(-6231);
			22486: out = 16'(-1835);
			22487: out = 16'(3332);
			22488: out = 16'(5915);
			22489: out = 16'(9354);
			22490: out = 16'(6102);
			22491: out = 16'(-3327);
			22492: out = 16'(-14790);
			22493: out = 16'(-10157);
			22494: out = 16'(-4504);
			22495: out = 16'(-1850);
			22496: out = 16'(836);
			22497: out = 16'(3331);
			22498: out = 16'(5898);
			22499: out = 16'(5649);
			22500: out = 16'(3150);
			22501: out = 16'(-1396);
			22502: out = 16'(-4487);
			22503: out = 16'(-7853);
			22504: out = 16'(-9352);
			22505: out = 16'(-2629);
			22506: out = 16'(2339);
			22507: out = 16'(5943);
			22508: out = 16'(5610);
			22509: out = 16'(2198);
			22510: out = 16'(-2489);
			22511: out = 16'(-4657);
			22512: out = 16'(-3972);
			22513: out = 16'(-1196);
			22514: out = 16'(1598);
			22515: out = 16'(5018);
			22516: out = 16'(6733);
			22517: out = 16'(5683);
			22518: out = 16'(802);
			22519: out = 16'(-797);
			22520: out = 16'(-656);
			22521: out = 16'(926);
			22522: out = 16'(4132);
			22523: out = 16'(2039);
			22524: out = 16'(-4061);
			22525: out = 16'(-6853);
			22526: out = 16'(2364);
			22527: out = 16'(10144);
			22528: out = 16'(10369);
			22529: out = 16'(2279);
			22530: out = 16'(-3583);
			22531: out = 16'(-6058);
			22532: out = 16'(-202);
			22533: out = 16'(2262);
			22534: out = 16'(-515);
			22535: out = 16'(-3100);
			22536: out = 16'(1629);
			22537: out = 16'(4762);
			22538: out = 16'(2980);
			22539: out = 16'(2629);
			22540: out = 16'(2678);
			22541: out = 16'(-861);
			22542: out = 16'(-7697);
			22543: out = 16'(-7607);
			22544: out = 16'(-2922);
			22545: out = 16'(3975);
			22546: out = 16'(5286);
			22547: out = 16'(2704);
			22548: out = 16'(0);
			22549: out = 16'(1794);
			22550: out = 16'(2810);
			22551: out = 16'(-893);
			22552: out = 16'(-3522);
			22553: out = 16'(-4334);
			22554: out = 16'(-1179);
			22555: out = 16'(1624);
			22556: out = 16'(30);
			22557: out = 16'(-1891);
			22558: out = 16'(-582);
			22559: out = 16'(1960);
			22560: out = 16'(-76);
			22561: out = 16'(-2148);
			22562: out = 16'(-2243);
			22563: out = 16'(927);
			22564: out = 16'(1413);
			22565: out = 16'(2421);
			22566: out = 16'(-995);
			22567: out = 16'(-3073);
			22568: out = 16'(-1934);
			22569: out = 16'(616);
			22570: out = 16'(-882);
			22571: out = 16'(-1450);
			22572: out = 16'(1122);
			22573: out = 16'(136);
			22574: out = 16'(-14);
			22575: out = 16'(1718);
			22576: out = 16'(4392);
			22577: out = 16'(-26);
			22578: out = 16'(4196);
			22579: out = 16'(6728);
			22580: out = 16'(3153);
			22581: out = 16'(-8015);
			22582: out = 16'(-8843);
			22583: out = 16'(-4049);
			22584: out = 16'(1397);
			22585: out = 16'(1496);
			22586: out = 16'(627);
			22587: out = 16'(-1155);
			22588: out = 16'(199);
			22589: out = 16'(2868);
			22590: out = 16'(3598);
			22591: out = 16'(-853);
			22592: out = 16'(-6724);
			22593: out = 16'(-7961);
			22594: out = 16'(1223);
			22595: out = 16'(4353);
			22596: out = 16'(3531);
			22597: out = 16'(1466);
			22598: out = 16'(101);
			22599: out = 16'(-670);
			22600: out = 16'(-2515);
			22601: out = 16'(-4086);
			22602: out = 16'(-2598);
			22603: out = 16'(-539);
			22604: out = 16'(1538);
			22605: out = 16'(1571);
			22606: out = 16'(269);
			22607: out = 16'(1664);
			22608: out = 16'(2694);
			22609: out = 16'(1951);
			22610: out = 16'(30);
			22611: out = 16'(1797);
			22612: out = 16'(849);
			22613: out = 16'(-1327);
			22614: out = 16'(-2563);
			22615: out = 16'(1827);
			22616: out = 16'(1927);
			22617: out = 16'(1073);
			22618: out = 16'(-717);
			22619: out = 16'(-857);
			22620: out = 16'(-1447);
			22621: out = 16'(118);
			22622: out = 16'(301);
			22623: out = 16'(-1252);
			22624: out = 16'(-7223);
			22625: out = 16'(-3060);
			22626: out = 16'(5774);
			22627: out = 16'(8922);
			22628: out = 16'(3719);
			22629: out = 16'(-3185);
			22630: out = 16'(-7944);
			22631: out = 16'(-8468);
			22632: out = 16'(-3229);
			22633: out = 16'(1463);
			22634: out = 16'(4197);
			22635: out = 16'(4280);
			22636: out = 16'(2902);
			22637: out = 16'(-95);
			22638: out = 16'(-1340);
			22639: out = 16'(-763);
			22640: out = 16'(-1199);
			22641: out = 16'(-1577);
			22642: out = 16'(-1483);
			22643: out = 16'(2146);
			22644: out = 16'(5930);
			22645: out = 16'(4919);
			22646: out = 16'(580);
			22647: out = 16'(-1193);
			22648: out = 16'(-831);
			22649: out = 16'(-5592);
			22650: out = 16'(-8184);
			22651: out = 16'(-4200);
			22652: out = 16'(3076);
			22653: out = 16'(1619);
			22654: out = 16'(2170);
			22655: out = 16'(2899);
			22656: out = 16'(4601);
			22657: out = 16'(2216);
			22658: out = 16'(1409);
			22659: out = 16'(-274);
			22660: out = 16'(712);
			22661: out = 16'(1287);
			22662: out = 16'(480);
			22663: out = 16'(-3981);
			22664: out = 16'(-2559);
			22665: out = 16'(5329);
			22666: out = 16'(5372);
			22667: out = 16'(2352);
			22668: out = 16'(-2405);
			22669: out = 16'(-2459);
			22670: out = 16'(-740);
			22671: out = 16'(1051);
			22672: out = 16'(-914);
			22673: out = 16'(360);
			22674: out = 16'(5481);
			22675: out = 16'(7005);
			22676: out = 16'(1878);
			22677: out = 16'(-1313);
			22678: out = 16'(1326);
			22679: out = 16'(266);
			22680: out = 16'(-6791);
			22681: out = 16'(-9586);
			22682: out = 16'(-754);
			22683: out = 16'(727);
			22684: out = 16'(2372);
			22685: out = 16'(576);
			22686: out = 16'(26);
			22687: out = 16'(-387);
			22688: out = 16'(35);
			22689: out = 16'(259);
			22690: out = 16'(2586);
			22691: out = 16'(3637);
			22692: out = 16'(2725);
			22693: out = 16'(-2938);
			22694: out = 16'(-6610);
			22695: out = 16'(-3771);
			22696: out = 16'(1430);
			22697: out = 16'(2096);
			22698: out = 16'(-1038);
			22699: out = 16'(-3148);
			22700: out = 16'(-3388);
			22701: out = 16'(-1057);
			22702: out = 16'(539);
			22703: out = 16'(564);
			22704: out = 16'(-105);
			22705: out = 16'(2177);
			22706: out = 16'(5053);
			22707: out = 16'(5178);
			22708: out = 16'(2416);
			22709: out = 16'(-7492);
			22710: out = 16'(-12143);
			22711: out = 16'(-7634);
			22712: out = 16'(54);
			22713: out = 16'(579);
			22714: out = 16'(-751);
			22715: out = 16'(219);
			22716: out = 16'(3128);
			22717: out = 16'(4428);
			22718: out = 16'(1942);
			22719: out = 16'(-1425);
			22720: out = 16'(-3044);
			22721: out = 16'(-3073);
			22722: out = 16'(-1639);
			22723: out = 16'(-354);
			22724: out = 16'(599);
			22725: out = 16'(2830);
			22726: out = 16'(2169);
			22727: out = 16'(630);
			22728: out = 16'(-1976);
			22729: out = 16'(-2527);
			22730: out = 16'(-941);
			22731: out = 16'(3191);
			22732: out = 16'(3342);
			22733: out = 16'(-202);
			22734: out = 16'(-1338);
			22735: out = 16'(3894);
			22736: out = 16'(6738);
			22737: out = 16'(3138);
			22738: out = 16'(-1585);
			22739: out = 16'(-129);
			22740: out = 16'(2810);
			22741: out = 16'(495);
			22742: out = 16'(-9924);
			22743: out = 16'(-3837);
			22744: out = 16'(4995);
			22745: out = 16'(7316);
			22746: out = 16'(2302);
			22747: out = 16'(217);
			22748: out = 16'(-829);
			22749: out = 16'(18);
			22750: out = 16'(405);
			22751: out = 16'(4018);
			22752: out = 16'(2332);
			22753: out = 16'(2630);
			22754: out = 16'(5518);
			22755: out = 16'(2516);
			22756: out = 16'(-1769);
			22757: out = 16'(-3107);
			22758: out = 16'(-267);
			22759: out = 16'(-1874);
			22760: out = 16'(-2778);
			22761: out = 16'(-2760);
			22762: out = 16'(931);
			22763: out = 16'(3582);
			22764: out = 16'(4439);
			22765: out = 16'(1482);
			22766: out = 16'(-1148);
			22767: out = 16'(-2830);
			22768: out = 16'(-4868);
			22769: out = 16'(-5992);
			22770: out = 16'(-3717);
			22771: out = 16'(-324);
			22772: out = 16'(33);
			22773: out = 16'(-494);
			22774: out = 16'(39);
			22775: out = 16'(-114);
			22776: out = 16'(4593);
			22777: out = 16'(-2791);
			22778: out = 16'(-3809);
			22779: out = 16'(585);
			22780: out = 16'(-356);
			22781: out = 16'(-2403);
			22782: out = 16'(-1247);
			22783: out = 16'(3335);
			22784: out = 16'(5486);
			22785: out = 16'(1062);
			22786: out = 16'(-2112);
			22787: out = 16'(-4464);
			22788: out = 16'(-6800);
			22789: out = 16'(-1073);
			22790: out = 16'(4285);
			22791: out = 16'(5277);
			22792: out = 16'(1643);
			22793: out = 16'(-3663);
			22794: out = 16'(-1254);
			22795: out = 16'(1317);
			22796: out = 16'(-531);
			22797: out = 16'(-5869);
			22798: out = 16'(1385);
			22799: out = 16'(4978);
			22800: out = 16'(-382);
			22801: out = 16'(-8445);
			22802: out = 16'(2805);
			22803: out = 16'(9279);
			22804: out = 16'(2010);
			22805: out = 16'(-10188);
			22806: out = 16'(-6847);
			22807: out = 16'(671);
			22808: out = 16'(401);
			22809: out = 16'(-6321);
			22810: out = 16'(-4212);
			22811: out = 16'(3714);
			22812: out = 16'(9119);
			22813: out = 16'(6730);
			22814: out = 16'(3056);
			22815: out = 16'(1445);
			22816: out = 16'(1174);
			22817: out = 16'(-1433);
			22818: out = 16'(-4777);
			22819: out = 16'(-7693);
			22820: out = 16'(-4961);
			22821: out = 16'(1980);
			22822: out = 16'(7767);
			22823: out = 16'(5043);
			22824: out = 16'(1226);
			22825: out = 16'(-357);
			22826: out = 16'(492);
			22827: out = 16'(-1075);
			22828: out = 16'(-1563);
			22829: out = 16'(163);
			22830: out = 16'(2411);
			22831: out = 16'(-92);
			22832: out = 16'(-1054);
			22833: out = 16'(-263);
			22834: out = 16'(2125);
			22835: out = 16'(2061);
			22836: out = 16'(643);
			22837: out = 16'(-3039);
			22838: out = 16'(-5222);
			22839: out = 16'(-3693);
			22840: out = 16'(646);
			22841: out = 16'(3077);
			22842: out = 16'(3451);
			22843: out = 16'(4090);
			22844: out = 16'(1631);
			22845: out = 16'(640);
			22846: out = 16'(-1528);
			22847: out = 16'(-3122);
			22848: out = 16'(-3410);
			22849: out = 16'(-761);
			22850: out = 16'(-490);
			22851: out = 16'(-734);
			22852: out = 16'(1459);
			22853: out = 16'(2043);
			22854: out = 16'(-694);
			22855: out = 16'(-3664);
			22856: out = 16'(-5002);
			22857: out = 16'(-145);
			22858: out = 16'(328);
			22859: out = 16'(348);
			22860: out = 16'(1842);
			22861: out = 16'(5654);
			22862: out = 16'(1445);
			22863: out = 16'(-1280);
			22864: out = 16'(622);
			22865: out = 16'(142);
			22866: out = 16'(-7561);
			22867: out = 16'(-10701);
			22868: out = 16'(-3474);
			22869: out = 16'(2780);
			22870: out = 16'(1704);
			22871: out = 16'(-330);
			22872: out = 16'(2116);
			22873: out = 16'(3855);
			22874: out = 16'(3463);
			22875: out = 16'(343);
			22876: out = 16'(-1278);
			22877: out = 16'(-1086);
			22878: out = 16'(488);
			22879: out = 16'(400);
			22880: out = 16'(-167);
			22881: out = 16'(212);
			22882: out = 16'(2984);
			22883: out = 16'(2783);
			22884: out = 16'(-982);
			22885: out = 16'(-5174);
			22886: out = 16'(-2941);
			22887: out = 16'(-771);
			22888: out = 16'(44);
			22889: out = 16'(-1559);
			22890: out = 16'(-1496);
			22891: out = 16'(1273);
			22892: out = 16'(5070);
			22893: out = 16'(4424);
			22894: out = 16'(-61);
			22895: out = 16'(-1257);
			22896: out = 16'(574);
			22897: out = 16'(1597);
			22898: out = 16'(414);
			22899: out = 16'(-1127);
			22900: out = 16'(-451);
			22901: out = 16'(-99);
			22902: out = 16'(59);
			22903: out = 16'(-337);
			22904: out = 16'(2067);
			22905: out = 16'(1402);
			22906: out = 16'(-200);
			22907: out = 16'(-212);
			22908: out = 16'(7252);
			22909: out = 16'(7076);
			22910: out = 16'(-59);
			22911: out = 16'(-8052);
			22912: out = 16'(-4323);
			22913: out = 16'(-2407);
			22914: out = 16'(-1484);
			22915: out = 16'(959);
			22916: out = 16'(5289);
			22917: out = 16'(2624);
			22918: out = 16'(-317);
			22919: out = 16'(-106);
			22920: out = 16'(490);
			22921: out = 16'(-2875);
			22922: out = 16'(-2857);
			22923: out = 16'(1258);
			22924: out = 16'(1356);
			22925: out = 16'(245);
			22926: out = 16'(1475);
			22927: out = 16'(4262);
			22928: out = 16'(1683);
			22929: out = 16'(-4203);
			22930: out = 16'(-6855);
			22931: out = 16'(-3000);
			22932: out = 16'(254);
			22933: out = 16'(497);
			22934: out = 16'(-1189);
			22935: out = 16'(-486);
			22936: out = 16'(-592);
			22937: out = 16'(-2314);
			22938: out = 16'(-3865);
			22939: out = 16'(803);
			22940: out = 16'(5981);
			22941: out = 16'(4259);
			22942: out = 16'(-1301);
			22943: out = 16'(-2319);
			22944: out = 16'(463);
			22945: out = 16'(-334);
			22946: out = 16'(-862);
			22947: out = 16'(-699);
			22948: out = 16'(-479);
			22949: out = 16'(-3312);
			22950: out = 16'(-4553);
			22951: out = 16'(-4000);
			22952: out = 16'(-1983);
			22953: out = 16'(-480);
			22954: out = 16'(3895);
			22955: out = 16'(5694);
			22956: out = 16'(3900);
			22957: out = 16'(-1351);
			22958: out = 16'(-3392);
			22959: out = 16'(-5087);
			22960: out = 16'(-3206);
			22961: out = 16'(-417);
			22962: out = 16'(148);
			22963: out = 16'(1597);
			22964: out = 16'(2071);
			22965: out = 16'(1485);
			22966: out = 16'(75);
			22967: out = 16'(1690);
			22968: out = 16'(2);
			22969: out = 16'(-2871);
			22970: out = 16'(-1737);
			22971: out = 16'(6489);
			22972: out = 16'(9130);
			22973: out = 16'(3134);
			22974: out = 16'(-5982);
			22975: out = 16'(-5791);
			22976: out = 16'(-4175);
			22977: out = 16'(-1799);
			22978: out = 16'(-887);
			22979: out = 16'(324);
			22980: out = 16'(3027);
			22981: out = 16'(5739);
			22982: out = 16'(3508);
			22983: out = 16'(-4963);
			22984: out = 16'(-1079);
			22985: out = 16'(1386);
			22986: out = 16'(1143);
			22987: out = 16'(-79);
			22988: out = 16'(1374);
			22989: out = 16'(1961);
			22990: out = 16'(875);
			22991: out = 16'(247);
			22992: out = 16'(2090);
			22993: out = 16'(3926);
			22994: out = 16'(2378);
			22995: out = 16'(-607);
			22996: out = 16'(-378);
			22997: out = 16'(-2473);
			22998: out = 16'(-3264);
			22999: out = 16'(-1011);
			23000: out = 16'(1509);
			23001: out = 16'(9891);
			23002: out = 16'(6948);
			23003: out = 16'(-139);
			23004: out = 16'(-2156);
			23005: out = 16'(-844);
			23006: out = 16'(-4273);
			23007: out = 16'(-10605);
			23008: out = 16'(-9537);
			23009: out = 16'(-204);
			23010: out = 16'(8030);
			23011: out = 16'(7045);
			23012: out = 16'(2502);
			23013: out = 16'(412);
			23014: out = 16'(232);
			23015: out = 16'(-2606);
			23016: out = 16'(-4850);
			23017: out = 16'(-1271);
			23018: out = 16'(242);
			23019: out = 16'(883);
			23020: out = 16'(2776);
			23021: out = 16'(5040);
			23022: out = 16'(1107);
			23023: out = 16'(-5662);
			23024: out = 16'(-6327);
			23025: out = 16'(448);
			23026: out = 16'(1536);
			23027: out = 16'(-791);
			23028: out = 16'(-1185);
			23029: out = 16'(1992);
			23030: out = 16'(1638);
			23031: out = 16'(-1815);
			23032: out = 16'(-1263);
			23033: out = 16'(2877);
			23034: out = 16'(-566);
			23035: out = 16'(-6400);
			23036: out = 16'(-8958);
			23037: out = 16'(-3293);
			23038: out = 16'(339);
			23039: out = 16'(6454);
			23040: out = 16'(3852);
			23041: out = 16'(1585);
			23042: out = 16'(1454);
			23043: out = 16'(577);
			23044: out = 16'(-4920);
			23045: out = 16'(-8013);
			23046: out = 16'(-4797);
			23047: out = 16'(-359);
			23048: out = 16'(447);
			23049: out = 16'(846);
			23050: out = 16'(3543);
			23051: out = 16'(3961);
			23052: out = 16'(1755);
			23053: out = 16'(-2507);
			23054: out = 16'(-5814);
			23055: out = 16'(-10947);
			23056: out = 16'(-4283);
			23057: out = 16'(-543);
			23058: out = 16'(1505);
			23059: out = 16'(3959);
			23060: out = 16'(6061);
			23061: out = 16'(2946);
			23062: out = 16'(-512);
			23063: out = 16'(520);
			23064: out = 16'(-107);
			23065: out = 16'(672);
			23066: out = 16'(-1021);
			23067: out = 16'(-2090);
			23068: out = 16'(2525);
			23069: out = 16'(1884);
			23070: out = 16'(-48);
			23071: out = 16'(1293);
			23072: out = 16'(5517);
			23073: out = 16'(6412);
			23074: out = 16'(1429);
			23075: out = 16'(-3824);
			23076: out = 16'(-2272);
			23077: out = 16'(4023);
			23078: out = 16'(6666);
			23079: out = 16'(3355);
			23080: out = 16'(-1206);
			23081: out = 16'(255);
			23082: out = 16'(2977);
			23083: out = 16'(2944);
			23084: out = 16'(-1084);
			23085: out = 16'(-1669);
			23086: out = 16'(-2399);
			23087: out = 16'(1761);
			23088: out = 16'(5813);
			23089: out = 16'(6094);
			23090: out = 16'(2218);
			23091: out = 16'(1498);
			23092: out = 16'(739);
			23093: out = 16'(-5507);
			23094: out = 16'(-5072);
			23095: out = 16'(-361);
			23096: out = 16'(2945);
			23097: out = 16'(-1013);
			23098: out = 16'(-269);
			23099: out = 16'(-776);
			23100: out = 16'(-173);
			23101: out = 16'(-856);
			23102: out = 16'(-2885);
			23103: out = 16'(-4904);
			23104: out = 16'(-4639);
			23105: out = 16'(-2518);
			23106: out = 16'(304);
			23107: out = 16'(96);
			23108: out = 16'(110);
			23109: out = 16'(3203);
			23110: out = 16'(7293);
			23111: out = 16'(6488);
			23112: out = 16'(278);
			23113: out = 16'(-6539);
			23114: out = 16'(-10163);
			23115: out = 16'(-2811);
			23116: out = 16'(-663);
			23117: out = 16'(-1983);
			23118: out = 16'(-2917);
			23119: out = 16'(-379);
			23120: out = 16'(-240);
			23121: out = 16'(1630);
			23122: out = 16'(3888);
			23123: out = 16'(-13);
			23124: out = 16'(-4681);
			23125: out = 16'(-3850);
			23126: out = 16'(1691);
			23127: out = 16'(-616);
			23128: out = 16'(614);
			23129: out = 16'(-1697);
			23130: out = 16'(-3630);
			23131: out = 16'(-6859);
			23132: out = 16'(-58);
			23133: out = 16'(1200);
			23134: out = 16'(1911);
			23135: out = 16'(3369);
			23136: out = 16'(764);
			23137: out = 16'(-2162);
			23138: out = 16'(-1350);
			23139: out = 16'(2497);
			23140: out = 16'(4136);
			23141: out = 16'(-438);
			23142: out = 16'(-4537);
			23143: out = 16'(-4336);
			23144: out = 16'(-2874);
			23145: out = 16'(827);
			23146: out = 16'(4267);
			23147: out = 16'(5916);
			23148: out = 16'(3965);
			23149: out = 16'(912);
			23150: out = 16'(-1873);
			23151: out = 16'(-3262);
			23152: out = 16'(-2515);
			23153: out = 16'(1106);
			23154: out = 16'(1277);
			23155: out = 16'(-1789);
			23156: out = 16'(-1622);
			23157: out = 16'(4661);
			23158: out = 16'(10355);
			23159: out = 16'(5512);
			23160: out = 16'(-3105);
			23161: out = 16'(-254);
			23162: out = 16'(-61);
			23163: out = 16'(-2908);
			23164: out = 16'(-5892);
			23165: out = 16'(-691);
			23166: out = 16'(4320);
			23167: out = 16'(4297);
			23168: out = 16'(-144);
			23169: out = 16'(-525);
			23170: out = 16'(2671);
			23171: out = 16'(6611);
			23172: out = 16'(4489);
			23173: out = 16'(-1296);
			23174: out = 16'(-4887);
			23175: out = 16'(-4429);
			23176: out = 16'(-1905);
			23177: out = 16'(371);
			23178: out = 16'(3805);
			23179: out = 16'(3432);
			23180: out = 16'(1097);
			23181: out = 16'(-2364);
			23182: out = 16'(-2047);
			23183: out = 16'(-3680);
			23184: out = 16'(-1456);
			23185: out = 16'(-318);
			23186: out = 16'(131);
			23187: out = 16'(704);
			23188: out = 16'(4642);
			23189: out = 16'(2456);
			23190: out = 16'(-6220);
			23191: out = 16'(-9832);
			23192: out = 16'(-5956);
			23193: out = 16'(-1511);
			23194: out = 16'(-551);
			23195: out = 16'(4207);
			23196: out = 16'(6552);
			23197: out = 16'(5175);
			23198: out = 16'(311);
			23199: out = 16'(-980);
			23200: out = 16'(-4432);
			23201: out = 16'(-5852);
			23202: out = 16'(-4459);
			23203: out = 16'(2325);
			23204: out = 16'(3600);
			23205: out = 16'(3749);
			23206: out = 16'(1226);
			23207: out = 16'(215);
			23208: out = 16'(-672);
			23209: out = 16'(5195);
			23210: out = 16'(6764);
			23211: out = 16'(155);
			23212: out = 16'(-7871);
			23213: out = 16'(-13335);
			23214: out = 16'(-9646);
			23215: out = 16'(-715);
			23216: out = 16'(3089);
			23217: out = 16'(2771);
			23218: out = 16'(2028);
			23219: out = 16'(4739);
			23220: out = 16'(4837);
			23221: out = 16'(-340);
			23222: out = 16'(-8407);
			23223: out = 16'(-6833);
			23224: out = 16'(2026);
			23225: out = 16'(4823);
			23226: out = 16'(-2343);
			23227: out = 16'(-3900);
			23228: out = 16'(3635);
			23229: out = 16'(4180);
			23230: out = 16'(-2476);
			23231: out = 16'(-4899);
			23232: out = 16'(2366);
			23233: out = 16'(7160);
			23234: out = 16'(3950);
			23235: out = 16'(-33);
			23236: out = 16'(105);
			23237: out = 16'(-1557);
			23238: out = 16'(-975);
			23239: out = 16'(-765);
			23240: out = 16'(21);
			23241: out = 16'(-1162);
			23242: out = 16'(3647);
			23243: out = 16'(3079);
			23244: out = 16'(-127);
			23245: out = 16'(-3155);
			23246: out = 16'(-3153);
			23247: out = 16'(62);
			23248: out = 16'(2515);
			23249: out = 16'(2005);
			23250: out = 16'(-971);
			23251: out = 16'(692);
			23252: out = 16'(1661);
			23253: out = 16'(-695);
			23254: out = 16'(-4740);
			23255: out = 16'(-1464);
			23256: out = 16'(1446);
			23257: out = 16'(1140);
			23258: out = 16'(106);
			23259: out = 16'(-315);
			23260: out = 16'(1129);
			23261: out = 16'(1253);
			23262: out = 16'(-853);
			23263: out = 16'(-7112);
			23264: out = 16'(-6065);
			23265: out = 16'(-1282);
			23266: out = 16'(2505);
			23267: out = 16'(5651);
			23268: out = 16'(6412);
			23269: out = 16'(4701);
			23270: out = 16'(173);
			23271: out = 16'(-2625);
			23272: out = 16'(-5150);
			23273: out = 16'(-3100);
			23274: out = 16'(-927);
			23275: out = 16'(-1098);
			23276: out = 16'(-4383);
			23277: out = 16'(-2563);
			23278: out = 16'(1837);
			23279: out = 16'(4284);
			23280: out = 16'(3485);
			23281: out = 16'(3997);
			23282: out = 16'(2109);
			23283: out = 16'(-4249);
			23284: out = 16'(-7192);
			23285: out = 16'(-5372);
			23286: out = 16'(-409);
			23287: out = 16'(597);
			23288: out = 16'(2546);
			23289: out = 16'(-234);
			23290: out = 16'(3808);
			23291: out = 16'(7273);
			23292: out = 16'(5530);
			23293: out = 16'(-3997);
			23294: out = 16'(-4049);
			23295: out = 16'(2838);
			23296: out = 16'(7459);
			23297: out = 16'(2397);
			23298: out = 16'(160);
			23299: out = 16'(-1518);
			23300: out = 16'(-3097);
			23301: out = 16'(-1790);
			23302: out = 16'(402);
			23303: out = 16'(-1157);
			23304: out = 16'(-1916);
			23305: out = 16'(5594);
			23306: out = 16'(7821);
			23307: out = 16'(871);
			23308: out = 16'(-6905);
			23309: out = 16'(-4135);
			23310: out = 16'(-1462);
			23311: out = 16'(-5657);
			23312: out = 16'(-9586);
			23313: out = 16'(-2015);
			23314: out = 16'(2509);
			23315: out = 16'(2042);
			23316: out = 16'(552);
			23317: out = 16'(5368);
			23318: out = 16'(8409);
			23319: out = 16'(5271);
			23320: out = 16'(-3210);
			23321: out = 16'(-9090);
			23322: out = 16'(-5243);
			23323: out = 16'(-3498);
			23324: out = 16'(-1594);
			23325: out = 16'(1320);
			23326: out = 16'(6597);
			23327: out = 16'(4549);
			23328: out = 16'(4285);
			23329: out = 16'(2768);
			23330: out = 16'(-1449);
			23331: out = 16'(-9089);
			23332: out = 16'(-5560);
			23333: out = 16'(2434);
			23334: out = 16'(3522);
			23335: out = 16'(674);
			23336: out = 16'(-1381);
			23337: out = 16'(-368);
			23338: out = 16'(625);
			23339: out = 16'(30);
			23340: out = 16'(21);
			23341: out = 16'(-1092);
			23342: out = 16'(-3646);
			23343: out = 16'(-5640);
			23344: out = 16'(-277);
			23345: out = 16'(3219);
			23346: out = 16'(1618);
			23347: out = 16'(-689);
			23348: out = 16'(1029);
			23349: out = 16'(1085);
			23350: out = 16'(-3282);
			23351: out = 16'(-6026);
			23352: out = 16'(-2407);
			23353: out = 16'(4612);
			23354: out = 16'(6135);
			23355: out = 16'(4171);
			23356: out = 16'(2378);
			23357: out = 16'(3670);
			23358: out = 16'(84);
			23359: out = 16'(-6188);
			23360: out = 16'(-11060);
			23361: out = 16'(-3083);
			23362: out = 16'(904);
			23363: out = 16'(742);
			23364: out = 16'(4657);
			23365: out = 16'(10264);
			23366: out = 16'(7434);
			23367: out = 16'(-335);
			23368: out = 16'(-3911);
			23369: out = 16'(-5115);
			23370: out = 16'(-5662);
			23371: out = 16'(-4405);
			23372: out = 16'(1147);
			23373: out = 16'(5186);
			23374: out = 16'(5145);
			23375: out = 16'(3773);
			23376: out = 16'(4160);
			23377: out = 16'(3068);
			23378: out = 16'(829);
			23379: out = 16'(-1102);
			23380: out = 16'(-1598);
			23381: out = 16'(-3245);
			23382: out = 16'(-1042);
			23383: out = 16'(762);
			23384: out = 16'(2151);
			23385: out = 16'(4097);
			23386: out = 16'(2359);
			23387: out = 16'(2806);
			23388: out = 16'(2756);
			23389: out = 16'(1996);
			23390: out = 16'(-1429);
			23391: out = 16'(-1350);
			23392: out = 16'(-3004);
			23393: out = 16'(-5277);
			23394: out = 16'(-5496);
			23395: out = 16'(5053);
			23396: out = 16'(9100);
			23397: out = 16'(2533);
			23398: out = 16'(-5652);
			23399: out = 16'(-8453);
			23400: out = 16'(-6826);
			23401: out = 16'(-3522);
			23402: out = 16'(1912);
			23403: out = 16'(2319);
			23404: out = 16'(2548);
			23405: out = 16'(2777);
			23406: out = 16'(3893);
			23407: out = 16'(-16);
			23408: out = 16'(-2220);
			23409: out = 16'(-4124);
			23410: out = 16'(-4857);
			23411: out = 16'(-2329);
			23412: out = 16'(510);
			23413: out = 16'(3056);
			23414: out = 16'(4118);
			23415: out = 16'(4113);
			23416: out = 16'(578);
			23417: out = 16'(387);
			23418: out = 16'(3187);
			23419: out = 16'(3356);
			23420: out = 16'(3);
			23421: out = 16'(-3761);
			23422: out = 16'(-3125);
			23423: out = 16'(-243);
			23424: out = 16'(2262);
			23425: out = 16'(652);
			23426: out = 16'(-202);
			23427: out = 16'(429);
			23428: out = 16'(1564);
			23429: out = 16'(-2924);
			23430: out = 16'(-6246);
			23431: out = 16'(-5407);
			23432: out = 16'(-1335);
			23433: out = 16'(-621);
			23434: out = 16'(1756);
			23435: out = 16'(4790);
			23436: out = 16'(5366);
			23437: out = 16'(1119);
			23438: out = 16'(-2965);
			23439: out = 16'(-6356);
			23440: out = 16'(-7535);
			23441: out = 16'(-4279);
			23442: out = 16'(1137);
			23443: out = 16'(1940);
			23444: out = 16'(-178);
			23445: out = 16'(-3206);
			23446: out = 16'(4543);
			23447: out = 16'(6785);
			23448: out = 16'(-318);
			23449: out = 16'(-7166);
			23450: out = 16'(-1719);
			23451: out = 16'(3314);
			23452: out = 16'(-666);
			23453: out = 16'(-8252);
			23454: out = 16'(-3503);
			23455: out = 16'(1796);
			23456: out = 16'(921);
			23457: out = 16'(-339);
			23458: out = 16'(-489);
			23459: out = 16'(3138);
			23460: out = 16'(3336);
			23461: out = 16'(-64);
			23462: out = 16'(-118);
			23463: out = 16'(1700);
			23464: out = 16'(2690);
			23465: out = 16'(1580);
			23466: out = 16'(2687);
			23467: out = 16'(625);
			23468: out = 16'(-563);
			23469: out = 16'(46);
			23470: out = 16'(450);
			23471: out = 16'(1598);
			23472: out = 16'(1538);
			23473: out = 16'(1943);
			23474: out = 16'(2241);
			23475: out = 16'(2592);
			23476: out = 16'(1147);
			23477: out = 16'(426);
			23478: out = 16'(101);
			23479: out = 16'(-25);
			23480: out = 16'(-2674);
			23481: out = 16'(-1019);
			23482: out = 16'(4220);
			23483: out = 16'(2327);
			23484: out = 16'(213);
			23485: out = 16'(1032);
			23486: out = 16'(3502);
			23487: out = 16'(-484);
			23488: out = 16'(-3874);
			23489: out = 16'(-5158);
			23490: out = 16'(-3922);
			23491: out = 16'(-5060);
			23492: out = 16'(-3451);
			23493: out = 16'(474);
			23494: out = 16'(5727);
			23495: out = 16'(6568);
			23496: out = 16'(-871);
			23497: out = 16'(-6892);
			23498: out = 16'(-5369);
			23499: out = 16'(987);
			23500: out = 16'(-963);
			23501: out = 16'(-1137);
			23502: out = 16'(-159);
			23503: out = 16'(2697);
			23504: out = 16'(7063);
			23505: out = 16'(3914);
			23506: out = 16'(-2344);
			23507: out = 16'(-5263);
			23508: out = 16'(-438);
			23509: out = 16'(242);
			23510: out = 16'(-2427);
			23511: out = 16'(-4324);
			23512: out = 16'(321);
			23513: out = 16'(3138);
			23514: out = 16'(2552);
			23515: out = 16'(-2240);
			23516: out = 16'(-4313);
			23517: out = 16'(-6354);
			23518: out = 16'(-152);
			23519: out = 16'(2374);
			23520: out = 16'(-566);
			23521: out = 16'(-4321);
			23522: out = 16'(92);
			23523: out = 16'(3493);
			23524: out = 16'(1723);
			23525: out = 16'(-705);
			23526: out = 16'(189);
			23527: out = 16'(-1103);
			23528: out = 16'(-6388);
			23529: out = 16'(-8568);
			23530: out = 16'(-2446);
			23531: out = 16'(6360);
			23532: out = 16'(8654);
			23533: out = 16'(5414);
			23534: out = 16'(1300);
			23535: out = 16'(657);
			23536: out = 16'(-308);
			23537: out = 16'(-3393);
			23538: out = 16'(-7998);
			23539: out = 16'(-3574);
			23540: out = 16'(3952);
			23541: out = 16'(6709);
			23542: out = 16'(4431);
			23543: out = 16'(3619);
			23544: out = 16'(5172);
			23545: out = 16'(5026);
			23546: out = 16'(-437);
			23547: out = 16'(-2423);
			23548: out = 16'(-4813);
			23549: out = 16'(-5657);
			23550: out = 16'(-2466);
			23551: out = 16'(1304);
			23552: out = 16'(3951);
			23553: out = 16'(2985);
			23554: out = 16'(1738);
			23555: out = 16'(2558);
			23556: out = 16'(4950);
			23557: out = 16'(3304);
			23558: out = 16'(-1576);
			23559: out = 16'(-7608);
			23560: out = 16'(-4981);
			23561: out = 16'(-1398);
			23562: out = 16'(-32);
			23563: out = 16'(-365);
			23564: out = 16'(3102);
			23565: out = 16'(3441);
			23566: out = 16'(1356);
			23567: out = 16'(-1452);
			23568: out = 16'(-384);
			23569: out = 16'(-696);
			23570: out = 16'(1621);
			23571: out = 16'(5096);
			23572: out = 16'(4467);
			23573: out = 16'(-3375);
			23574: out = 16'(-5643);
			23575: out = 16'(1658);
			23576: out = 16'(2388);
			23577: out = 16'(-1833);
			23578: out = 16'(-7466);
			23579: out = 16'(-6479);
			23580: out = 16'(-1662);
			23581: out = 16'(2014);
			23582: out = 16'(2779);
			23583: out = 16'(3248);
			23584: out = 16'(1938);
			23585: out = 16'(-224);
			23586: out = 16'(-3819);
			23587: out = 16'(-4198);
			23588: out = 16'(-792);
			23589: out = 16'(1972);
			23590: out = 16'(2113);
			23591: out = 16'(1034);
			23592: out = 16'(676);
			23593: out = 16'(2125);
			23594: out = 16'(1256);
			23595: out = 16'(-1187);
			23596: out = 16'(-3359);
			23597: out = 16'(-2968);
			23598: out = 16'(-3085);
			23599: out = 16'(-2865);
			23600: out = 16'(-3103);
			23601: out = 16'(-3324);
			23602: out = 16'(4642);
			23603: out = 16'(9617);
			23604: out = 16'(6802);
			23605: out = 16'(-977);
			23606: out = 16'(-6961);
			23607: out = 16'(-6991);
			23608: out = 16'(-5674);
			23609: out = 16'(-6208);
			23610: out = 16'(-428);
			23611: out = 16'(1611);
			23612: out = 16'(1089);
			23613: out = 16'(-1009);
			23614: out = 16'(440);
			23615: out = 16'(2938);
			23616: out = 16'(4955);
			23617: out = 16'(2552);
			23618: out = 16'(-2521);
			23619: out = 16'(-5519);
			23620: out = 16'(-2850);
			23621: out = 16'(1576);
			23622: out = 16'(3218);
			23623: out = 16'(768);
			23624: out = 16'(-259);
			23625: out = 16'(158);
			23626: out = 16'(4);
			23627: out = 16'(208);
			23628: out = 16'(-119);
			23629: out = 16'(554);
			23630: out = 16'(2223);
			23631: out = 16'(3892);
			23632: out = 16'(6636);
			23633: out = 16'(7323);
			23634: out = 16'(4490);
			23635: out = 16'(-388);
			23636: out = 16'(-2888);
			23637: out = 16'(-2867);
			23638: out = 16'(-2042);
			23639: out = 16'(-1133);
			23640: out = 16'(885);
			23641: out = 16'(3846);
			23642: out = 16'(5230);
			23643: out = 16'(3002);
			23644: out = 16'(-1479);
			23645: out = 16'(-3461);
			23646: out = 16'(-2071);
			23647: out = 16'(-210);
			23648: out = 16'(-220);
			23649: out = 16'(590);
			23650: out = 16'(3473);
			23651: out = 16'(5611);
			23652: out = 16'(1837);
			23653: out = 16'(315);
			23654: out = 16'(-1707);
			23655: out = 16'(-2603);
			23656: out = 16'(-3490);
			23657: out = 16'(-4540);
			23658: out = 16'(-5553);
			23659: out = 16'(-3022);
			23660: out = 16'(1793);
			23661: out = 16'(3807);
			23662: out = 16'(935);
			23663: out = 16'(-2381);
			23664: out = 16'(-3093);
			23665: out = 16'(-4734);
			23666: out = 16'(-3853);
			23667: out = 16'(36);
			23668: out = 16'(4386);
			23669: out = 16'(1414);
			23670: out = 16'(-1414);
			23671: out = 16'(-2959);
			23672: out = 16'(293);
			23673: out = 16'(942);
			23674: out = 16'(2715);
			23675: out = 16'(-4992);
			23676: out = 16'(-11338);
			23677: out = 16'(-7429);
			23678: out = 16'(2355);
			23679: out = 16'(5284);
			23680: out = 16'(3308);
			23681: out = 16'(3002);
			23682: out = 16'(3816);
			23683: out = 16'(1824);
			23684: out = 16'(-2523);
			23685: out = 16'(-4452);
			23686: out = 16'(-3015);
			23687: out = 16'(2331);
			23688: out = 16'(4956);
			23689: out = 16'(2039);
			23690: out = 16'(-7184);
			23691: out = 16'(-2252);
			23692: out = 16'(3044);
			23693: out = 16'(3123);
			23694: out = 16'(-977);
			23695: out = 16'(-407);
			23696: out = 16'(1108);
			23697: out = 16'(2001);
			23698: out = 16'(2801);
			23699: out = 16'(3640);
			23700: out = 16'(4413);
			23701: out = 16'(1711);
			23702: out = 16'(-2711);
			23703: out = 16'(-4772);
			23704: out = 16'(-1778);
			23705: out = 16'(-78);
			23706: out = 16'(-1924);
			23707: out = 16'(-4449);
			23708: out = 16'(-1409);
			23709: out = 16'(2421);
			23710: out = 16'(4195);
			23711: out = 16'(3149);
			23712: out = 16'(7001);
			23713: out = 16'(4166);
			23714: out = 16'(-2590);
			23715: out = 16'(-7313);
			23716: out = 16'(885);
			23717: out = 16'(3167);
			23718: out = 16'(315);
			23719: out = 16'(-3242);
			23720: out = 16'(-2988);
			23721: out = 16'(1379);
			23722: out = 16'(6269);
			23723: out = 16'(6263);
			23724: out = 16'(1923);
			23725: out = 16'(-695);
			23726: out = 16'(2153);
			23727: out = 16'(3420);
			23728: out = 16'(-1569);
			23729: out = 16'(-8950);
			23730: out = 16'(-4378);
			23731: out = 16'(6335);
			23732: out = 16'(7219);
			23733: out = 16'(70);
			23734: out = 16'(-7139);
			23735: out = 16'(-5654);
			23736: out = 16'(-287);
			23737: out = 16'(-3519);
			23738: out = 16'(-5659);
			23739: out = 16'(-3991);
			23740: out = 16'(456);
			23741: out = 16'(325);
			23742: out = 16'(2246);
			23743: out = 16'(2138);
			23744: out = 16'(1306);
			23745: out = 16'(-270);
			23746: out = 16'(-2032);
			23747: out = 16'(-4409);
			23748: out = 16'(-3558);
			23749: out = 16'(74);
			23750: out = 16'(1846);
			23751: out = 16'(-2241);
			23752: out = 16'(-7005);
			23753: out = 16'(-6733);
			23754: out = 16'(-1731);
			23755: out = 16'(2373);
			23756: out = 16'(4195);
			23757: out = 16'(3659);
			23758: out = 16'(-427);
			23759: out = 16'(-2508);
			23760: out = 16'(-1477);
			23761: out = 16'(444);
			23762: out = 16'(258);
			23763: out = 16'(-5);
			23764: out = 16'(661);
			23765: out = 16'(-224);
			23766: out = 16'(-4470);
			23767: out = 16'(-4816);
			23768: out = 16'(48);
			23769: out = 16'(4204);
			23770: out = 16'(1259);
			23771: out = 16'(6);
			23772: out = 16'(661);
			23773: out = 16'(5004);
			23774: out = 16'(5201);
			23775: out = 16'(250);
			23776: out = 16'(-8389);
			23777: out = 16'(-7282);
			23778: out = 16'(2637);
			23779: out = 16'(5633);
			23780: out = 16'(4479);
			23781: out = 16'(98);
			23782: out = 16'(27);
			23783: out = 16'(2254);
			23784: out = 16'(4468);
			23785: out = 16'(-181);
			23786: out = 16'(-4276);
			23787: out = 16'(-2169);
			23788: out = 16'(3169);
			23789: out = 16'(3269);
			23790: out = 16'(341);
			23791: out = 16'(-846);
			23792: out = 16'(-221);
			23793: out = 16'(2621);
			23794: out = 16'(5268);
			23795: out = 16'(5515);
			23796: out = 16'(2451);
			23797: out = 16'(-1732);
			23798: out = 16'(-4289);
			23799: out = 16'(-5062);
			23800: out = 16'(-4584);
			23801: out = 16'(-1625);
			23802: out = 16'(4302);
			23803: out = 16'(7707);
			23804: out = 16'(4740);
			23805: out = 16'(-133);
			23806: out = 16'(-1463);
			23807: out = 16'(1353);
			23808: out = 16'(3376);
			23809: out = 16'(-816);
			23810: out = 16'(-285);
			23811: out = 16'(3632);
			23812: out = 16'(4588);
			23813: out = 16'(-4576);
			23814: out = 16'(-9113);
			23815: out = 16'(-8558);
			23816: out = 16'(-3261);
			23817: out = 16'(-395);
			23818: out = 16'(7019);
			23819: out = 16'(6304);
			23820: out = 16'(1078);
			23821: out = 16'(-2766);
			23822: out = 16'(607);
			23823: out = 16'(1157);
			23824: out = 16'(-1883);
			23825: out = 16'(-4600);
			23826: out = 16'(-700);
			23827: out = 16'(-268);
			23828: out = 16'(-2136);
			23829: out = 16'(-2420);
			23830: out = 16'(-359);
			23831: out = 16'(2113);
			23832: out = 16'(1209);
			23833: out = 16'(-1766);
			23834: out = 16'(-2697);
			23835: out = 16'(-351);
			23836: out = 16'(472);
			23837: out = 16'(-2355);
			23838: out = 16'(-4129);
			23839: out = 16'(-2303);
			23840: out = 16'(4073);
			23841: out = 16'(6812);
			23842: out = 16'(3420);
			23843: out = 16'(-419);
			23844: out = 16'(-2347);
			23845: out = 16'(-4435);
			23846: out = 16'(-7950);
			23847: out = 16'(-7372);
			23848: out = 16'(-2640);
			23849: out = 16'(3516);
			23850: out = 16'(5398);
			23851: out = 16'(2939);
			23852: out = 16'(498);
			23853: out = 16'(1450);
			23854: out = 16'(3899);
			23855: out = 16'(3638);
			23856: out = 16'(-1142);
			23857: out = 16'(-4765);
			23858: out = 16'(-3240);
			23859: out = 16'(280);
			23860: out = 16'(5897);
			23861: out = 16'(1417);
			23862: out = 16'(-5635);
			23863: out = 16'(-7766);
			23864: out = 16'(-639);
			23865: out = 16'(605);
			23866: out = 16'(1332);
			23867: out = 16'(5302);
			23868: out = 16'(5694);
			23869: out = 16'(6892);
			23870: out = 16'(2723);
			23871: out = 16'(-2756);
			23872: out = 16'(-7604);
			23873: out = 16'(-1893);
			23874: out = 16'(571);
			23875: out = 16'(-256);
			23876: out = 16'(53);
			23877: out = 16'(-279);
			23878: out = 16'(911);
			23879: out = 16'(2986);
			23880: out = 16'(5873);
			23881: out = 16'(7248);
			23882: out = 16'(3469);
			23883: out = 16'(-3459);
			23884: out = 16'(-7400);
			23885: out = 16'(-803);
			23886: out = 16'(55);
			23887: out = 16'(230);
			23888: out = 16'(2541);
			23889: out = 16'(4976);
			23890: out = 16'(6237);
			23891: out = 16'(2654);
			23892: out = 16'(-1835);
			23893: out = 16'(-3114);
			23894: out = 16'(-1952);
			23895: out = 16'(-789);
			23896: out = 16'(-506);
			23897: out = 16'(-30);
			23898: out = 16'(3186);
			23899: out = 16'(5239);
			23900: out = 16'(4602);
			23901: out = 16'(-387);
			23902: out = 16'(-5162);
			23903: out = 16'(-9124);
			23904: out = 16'(-5365);
			23905: out = 16'(421);
			23906: out = 16'(-180);
			23907: out = 16'(1436);
			23908: out = 16'(3756);
			23909: out = 16'(864);
			23910: out = 16'(-10635);
			23911: out = 16'(-5389);
			23912: out = 16'(3953);
			23913: out = 16'(5319);
			23914: out = 16'(-4598);
			23915: out = 16'(-4734);
			23916: out = 16'(-59);
			23917: out = 16'(3355);
			23918: out = 16'(-935);
			23919: out = 16'(456);
			23920: out = 16'(-3003);
			23921: out = 16'(-3500);
			23922: out = 16'(-2479);
			23923: out = 16'(-942);
			23924: out = 16'(-73);
			23925: out = 16'(280);
			23926: out = 16'(122);
			23927: out = 16'(33);
			23928: out = 16'(-745);
			23929: out = 16'(-482);
			23930: out = 16'(802);
			23931: out = 16'(1434);
			23932: out = 16'(-3228);
			23933: out = 16'(-6005);
			23934: out = 16'(-2964);
			23935: out = 16'(2002);
			23936: out = 16'(751);
			23937: out = 16'(-2439);
			23938: out = 16'(-2350);
			23939: out = 16'(811);
			23940: out = 16'(1990);
			23941: out = 16'(-630);
			23942: out = 16'(-477);
			23943: out = 16'(2533);
			23944: out = 16'(1706);
			23945: out = 16'(700);
			23946: out = 16'(-194);
			23947: out = 16'(225);
			23948: out = 16'(261);
			23949: out = 16'(122);
			23950: out = 16'(2349);
			23951: out = 16'(5105);
			23952: out = 16'(5109);
			23953: out = 16'(-94);
			23954: out = 16'(-3086);
			23955: out = 16'(-3651);
			23956: out = 16'(-2333);
			23957: out = 16'(-1304);
			23958: out = 16'(2855);
			23959: out = 16'(3651);
			23960: out = 16'(1154);
			23961: out = 16'(303);
			23962: out = 16'(1664);
			23963: out = 16'(3457);
			23964: out = 16'(3762);
			23965: out = 16'(2120);
			23966: out = 16'(656);
			23967: out = 16'(-3321);
			23968: out = 16'(-5856);
			23969: out = 16'(-3331);
			23970: out = 16'(-588);
			23971: out = 16'(796);
			23972: out = 16'(1094);
			23973: out = 16'(2151);
			23974: out = 16'(5797);
			23975: out = 16'(3942);
			23976: out = 16'(1453);
			23977: out = 16'(1964);
			23978: out = 16'(3402);
			23979: out = 16'(2406);
			23980: out = 16'(-930);
			23981: out = 16'(-3696);
			23982: out = 16'(-4935);
			23983: out = 16'(-857);
			23984: out = 16'(1088);
			23985: out = 16'(155);
			23986: out = 16'(179);
			23987: out = 16'(2810);
			23988: out = 16'(4499);
			23989: out = 16'(967);
			23990: out = 16'(-5435);
			23991: out = 16'(-6231);
			23992: out = 16'(-2068);
			23993: out = 16'(890);
			23994: out = 16'(-1443);
			23995: out = 16'(-6122);
			23996: out = 16'(-1801);
			23997: out = 16'(4750);
			23998: out = 16'(2792);
			23999: out = 16'(-8963);
			24000: out = 16'(-9489);
			24001: out = 16'(-1258);
			24002: out = 16'(4198);
			24003: out = 16'(-220);
			24004: out = 16'(-2255);
			24005: out = 16'(-518);
			24006: out = 16'(2358);
			24007: out = 16'(120);
			24008: out = 16'(-1139);
			24009: out = 16'(-1281);
			24010: out = 16'(2172);
			24011: out = 16'(3450);
			24012: out = 16'(-163);
			24013: out = 16'(-7330);
			24014: out = 16'(-8230);
			24015: out = 16'(-1523);
			24016: out = 16'(3692);
			24017: out = 16'(114);
			24018: out = 16'(-6337);
			24019: out = 16'(-6568);
			24020: out = 16'(1191);
			24021: out = 16'(4203);
			24022: out = 16'(3773);
			24023: out = 16'(2782);
			24024: out = 16'(2867);
			24025: out = 16'(4332);
			24026: out = 16'(-9);
			24027: out = 16'(-5807);
			24028: out = 16'(-6101);
			24029: out = 16'(3213);
			24030: out = 16'(2901);
			24031: out = 16'(-3552);
			24032: out = 16'(-5765);
			24033: out = 16'(3914);
			24034: out = 16'(8204);
			24035: out = 16'(6790);
			24036: out = 16'(3402);
			24037: out = 16'(1766);
			24038: out = 16'(1797);
			24039: out = 16'(723);
			24040: out = 16'(-68);
			24041: out = 16'(-197);
			24042: out = 16'(-665);
			24043: out = 16'(-1659);
			24044: out = 16'(1201);
			24045: out = 16'(5445);
			24046: out = 16'(2875);
			24047: out = 16'(-431);
			24048: out = 16'(-4);
			24049: out = 16'(2191);
			24050: out = 16'(20);
			24051: out = 16'(-876);
			24052: out = 16'(2650);
			24053: out = 16'(5704);
			24054: out = 16'(2086);
			24055: out = 16'(-3013);
			24056: out = 16'(-2624);
			24057: out = 16'(-23);
			24058: out = 16'(-1416);
			24059: out = 16'(-882);
			24060: out = 16'(3471);
			24061: out = 16'(4888);
			24062: out = 16'(-1573);
			24063: out = 16'(-6835);
			24064: out = 16'(-6913);
			24065: out = 16'(-3097);
			24066: out = 16'(-525);
			24067: out = 16'(4578);
			24068: out = 16'(5420);
			24069: out = 16'(3214);
			24070: out = 16'(-1032);
			24071: out = 16'(136);
			24072: out = 16'(-703);
			24073: out = 16'(856);
			24074: out = 16'(821);
			24075: out = 16'(-1417);
			24076: out = 16'(-2924);
			24077: out = 16'(-3493);
			24078: out = 16'(-5055);
			24079: out = 16'(-7669);
			24080: out = 16'(-5942);
			24081: out = 16'(-1059);
			24082: out = 16'(3734);
			24083: out = 16'(3346);
			24084: out = 16'(-61);
			24085: out = 16'(-1769);
			24086: out = 16'(1775);
			24087: out = 16'(3384);
			24088: out = 16'(-1405);
			24089: out = 16'(-4549);
			24090: out = 16'(-1423);
			24091: out = 16'(2179);
			24092: out = 16'(705);
			24093: out = 16'(-4523);
			24094: out = 16'(-2958);
			24095: out = 16'(901);
			24096: out = 16'(249);
			24097: out = 16'(3826);
			24098: out = 16'(5611);
			24099: out = 16'(3164);
			24100: out = 16'(-3524);
			24101: out = 16'(-3430);
			24102: out = 16'(-204);
			24103: out = 16'(2557);
			24104: out = 16'(1608);
			24105: out = 16'(4459);
			24106: out = 16'(809);
			24107: out = 16'(511);
			24108: out = 16'(1913);
			24109: out = 16'(1228);
			24110: out = 16'(-3009);
			24111: out = 16'(-8160);
			24112: out = 16'(-7894);
			24113: out = 16'(-209);
			24114: out = 16'(3491);
			24115: out = 16'(4621);
			24116: out = 16'(3562);
			24117: out = 16'(2536);
			24118: out = 16'(2528);
			24119: out = 16'(888);
			24120: out = 16'(-336);
			24121: out = 16'(-95);
			24122: out = 16'(-352);
			24123: out = 16'(72);
			24124: out = 16'(-755);
			24125: out = 16'(-2348);
			24126: out = 16'(-2609);
			24127: out = 16'(-3042);
			24128: out = 16'(-530);
			24129: out = 16'(3208);
			24130: out = 16'(6140);
			24131: out = 16'(2393);
			24132: out = 16'(1714);
			24133: out = 16'(3062);
			24134: out = 16'(3527);
			24135: out = 16'(-689);
			24136: out = 16'(-957);
			24137: out = 16'(692);
			24138: out = 16'(1000);
			24139: out = 16'(-2721);
			24140: out = 16'(-5089);
			24141: out = 16'(-6150);
			24142: out = 16'(-4689);
			24143: out = 16'(-11);
			24144: out = 16'(4927);
			24145: out = 16'(6796);
			24146: out = 16'(4810);
			24147: out = 16'(361);
			24148: out = 16'(-901);
			24149: out = 16'(-2295);
			24150: out = 16'(-3378);
			24151: out = 16'(-3350);
			24152: out = 16'(4371);
			24153: out = 16'(5961);
			24154: out = 16'(3388);
			24155: out = 16'(-1027);
			24156: out = 16'(-3203);
			24157: out = 16'(-6819);
			24158: out = 16'(-4767);
			24159: out = 16'(2264);
			24160: out = 16'(5388);
			24161: out = 16'(4795);
			24162: out = 16'(1864);
			24163: out = 16'(26);
			24164: out = 16'(-1308);
			24165: out = 16'(1527);
			24166: out = 16'(2427);
			24167: out = 16'(1290);
			24168: out = 16'(-1601);
			24169: out = 16'(-2701);
			24170: out = 16'(-3286);
			24171: out = 16'(-2064);
			24172: out = 16'(-268);
			24173: out = 16'(-113);
			24174: out = 16'(-862);
			24175: out = 16'(-1265);
			24176: out = 16'(-1082);
			24177: out = 16'(-104);
			24178: out = 16'(-1477);
			24179: out = 16'(-1890);
			24180: out = 16'(-77);
			24181: out = 16'(3896);
			24182: out = 16'(3787);
			24183: out = 16'(3221);
			24184: out = 16'(976);
			24185: out = 16'(-2095);
			24186: out = 16'(-3810);
			24187: out = 16'(-3087);
			24188: out = 16'(-3910);
			24189: out = 16'(-5979);
			24190: out = 16'(-839);
			24191: out = 16'(4460);
			24192: out = 16'(4433);
			24193: out = 16'(-1382);
			24194: out = 16'(-3106);
			24195: out = 16'(-1613);
			24196: out = 16'(1821);
			24197: out = 16'(1286);
			24198: out = 16'(-3246);
			24199: out = 16'(-3446);
			24200: out = 16'(130);
			24201: out = 16'(2668);
			24202: out = 16'(1577);
			24203: out = 16'(1620);
			24204: out = 16'(1684);
			24205: out = 16'(906);
			24206: out = 16'(-1489);
			24207: out = 16'(-4994);
			24208: out = 16'(-4254);
			24209: out = 16'(-982);
			24210: out = 16'(1239);
			24211: out = 16'(4029);
			24212: out = 16'(1179);
			24213: out = 16'(269);
			24214: out = 16'(4161);
			24215: out = 16'(9730);
			24216: out = 16'(3283);
			24217: out = 16'(-6302);
			24218: out = 16'(-9302);
			24219: out = 16'(-987);
			24220: out = 16'(-206);
			24221: out = 16'(-848);
			24222: out = 16'(212);
			24223: out = 16'(4131);
			24224: out = 16'(4608);
			24225: out = 16'(335);
			24226: out = 16'(-3787);
			24227: out = 16'(-399);
			24228: out = 16'(5898);
			24229: out = 16'(8325);
			24230: out = 16'(2962);
			24231: out = 16'(-2532);
			24232: out = 16'(-1604);
			24233: out = 16'(2028);
			24234: out = 16'(1248);
			24235: out = 16'(-2609);
			24236: out = 16'(-5742);
			24237: out = 16'(-900);
			24238: out = 16'(-1);
			24239: out = 16'(-1497);
			24240: out = 16'(205);
			24241: out = 16'(5947);
			24242: out = 16'(5779);
			24243: out = 16'(1336);
			24244: out = 16'(-1359);
			24245: out = 16'(-1707);
			24246: out = 16'(-754);
			24247: out = 16'(-515);
			24248: out = 16'(-538);
			24249: out = 16'(-3105);
			24250: out = 16'(-1891);
			24251: out = 16'(-791);
			24252: out = 16'(440);
			24253: out = 16'(3512);
			24254: out = 16'(763);
			24255: out = 16'(-3143);
			24256: out = 16'(-6941);
			24257: out = 16'(-8088);
			24258: out = 16'(-4186);
			24259: out = 16'(1559);
			24260: out = 16'(4394);
			24261: out = 16'(3475);
			24262: out = 16'(366);
			24263: out = 16'(-1258);
			24264: out = 16'(-3412);
			24265: out = 16'(-5309);
			24266: out = 16'(-1234);
			24267: out = 16'(2656);
			24268: out = 16'(3109);
			24269: out = 16'(-1980);
			24270: out = 16'(-7417);
			24271: out = 16'(-2936);
			24272: out = 16'(6104);
			24273: out = 16'(7952);
			24274: out = 16'(1510);
			24275: out = 16'(-2383);
			24276: out = 16'(712);
			24277: out = 16'(4329);
			24278: out = 16'(1366);
			24279: out = 16'(-3519);
			24280: out = 16'(-4451);
			24281: out = 16'(-738);
			24282: out = 16'(1510);
			24283: out = 16'(1851);
			24284: out = 16'(-421);
			24285: out = 16'(-903);
			24286: out = 16'(84);
			24287: out = 16'(1583);
			24288: out = 16'(284);
			24289: out = 16'(466);
			24290: out = 16'(1808);
			24291: out = 16'(1213);
			24292: out = 16'(293);
			24293: out = 16'(-2470);
			24294: out = 16'(-3467);
			24295: out = 16'(-822);
			24296: out = 16'(-508);
			24297: out = 16'(368);
			24298: out = 16'(838);
			24299: out = 16'(2093);
			24300: out = 16'(4790);
			24301: out = 16'(3831);
			24302: out = 16'(-665);
			24303: out = 16'(-3209);
			24304: out = 16'(1883);
			24305: out = 16'(4372);
			24306: out = 16'(977);
			24307: out = 16'(-5080);
			24308: out = 16'(-4193);
			24309: out = 16'(-3852);
			24310: out = 16'(-144);
			24311: out = 16'(1705);
			24312: out = 16'(1659);
			24313: out = 16'(1899);
			24314: out = 16'(4570);
			24315: out = 16'(4422);
			24316: out = 16'(-1491);
			24317: out = 16'(-5566);
			24318: out = 16'(-7517);
			24319: out = 16'(-3898);
			24320: out = 16'(235);
			24321: out = 16'(2527);
			24322: out = 16'(437);
			24323: out = 16'(674);
			24324: out = 16'(1311);
			24325: out = 16'(45);
			24326: out = 16'(-3861);
			24327: out = 16'(-3178);
			24328: out = 16'(-366);
			24329: out = 16'(50);
			24330: out = 16'(-138);
			24331: out = 16'(2385);
			24332: out = 16'(3230);
			24333: out = 16'(-748);
			24334: out = 16'(-1611);
			24335: out = 16'(-597);
			24336: out = 16'(1368);
			24337: out = 16'(1700);
			24338: out = 16'(3793);
			24339: out = 16'(1757);
			24340: out = 16'(-1610);
			24341: out = 16'(-3651);
			24342: out = 16'(-1089);
			24343: out = 16'(420);
			24344: out = 16'(502);
			24345: out = 16'(-137);
			24346: out = 16'(-159);
			24347: out = 16'(-2066);
			24348: out = 16'(-4651);
			24349: out = 16'(-4195);
			24350: out = 16'(794);
			24351: out = 16'(4759);
			24352: out = 16'(3637);
			24353: out = 16'(-380);
			24354: out = 16'(-3069);
			24355: out = 16'(-5459);
			24356: out = 16'(-3746);
			24357: out = 16'(-1279);
			24358: out = 16'(538);
			24359: out = 16'(1841);
			24360: out = 16'(4943);
			24361: out = 16'(6768);
			24362: out = 16'(4145);
			24363: out = 16'(-1824);
			24364: out = 16'(-6540);
			24365: out = 16'(-6194);
			24366: out = 16'(-3052);
			24367: out = 16'(405);
			24368: out = 16'(2042);
			24369: out = 16'(5119);
			24370: out = 16'(5188);
			24371: out = 16'(1701);
			24372: out = 16'(-3970);
			24373: out = 16'(-2007);
			24374: out = 16'(588);
			24375: out = 16'(-493);
			24376: out = 16'(-2393);
			24377: out = 16'(-985);
			24378: out = 16'(392);
			24379: out = 16'(-5);
			24380: out = 16'(291);
			24381: out = 16'(3050);
			24382: out = 16'(4380);
			24383: out = 16'(3059);
			24384: out = 16'(684);
			24385: out = 16'(751);
			24386: out = 16'(-1334);
			24387: out = 16'(-2756);
			24388: out = 16'(-463);
			24389: out = 16'(1835);
			24390: out = 16'(2294);
			24391: out = 16'(408);
			24392: out = 16'(-993);
			24393: out = 16'(-191);
			24394: out = 16'(-574);
			24395: out = 16'(-1395);
			24396: out = 16'(-154);
			24397: out = 16'(3635);
			24398: out = 16'(2945);
			24399: out = 16'(1419);
			24400: out = 16'(2732);
			24401: out = 16'(6673);
			24402: out = 16'(-660);
			24403: out = 16'(-8091);
			24404: out = 16'(-8736);
			24405: out = 16'(-546);
			24406: out = 16'(-2019);
			24407: out = 16'(-1334);
			24408: out = 16'(-163);
			24409: out = 16'(2038);
			24410: out = 16'(2869);
			24411: out = 16'(1335);
			24412: out = 16'(-1060);
			24413: out = 16'(-341);
			24414: out = 16'(998);
			24415: out = 16'(456);
			24416: out = 16'(-5297);
			24417: out = 16'(-8716);
			24418: out = 16'(-3382);
			24419: out = 16'(3394);
			24420: out = 16'(3097);
			24421: out = 16'(-882);
			24422: out = 16'(-147);
			24423: out = 16'(4210);
			24424: out = 16'(4674);
			24425: out = 16'(-592);
			24426: out = 16'(-5082);
			24427: out = 16'(-1788);
			24428: out = 16'(1853);
			24429: out = 16'(1353);
			24430: out = 16'(-1034);
			24431: out = 16'(34);
			24432: out = 16'(4174);
			24433: out = 16'(5924);
			24434: out = 16'(1685);
			24435: out = 16'(-4999);
			24436: out = 16'(-5644);
			24437: out = 16'(-1176);
			24438: out = 16'(2230);
			24439: out = 16'(3280);
			24440: out = 16'(1544);
			24441: out = 16'(3429);
			24442: out = 16'(3474);
			24443: out = 16'(-657);
			24444: out = 16'(-5105);
			24445: out = 16'(-1349);
			24446: out = 16'(3982);
			24447: out = 16'(2536);
			24448: out = 16'(-1952);
			24449: out = 16'(-2784);
			24450: out = 16'(2255);
			24451: out = 16'(5623);
			24452: out = 16'(3745);
			24453: out = 16'(-2180);
			24454: out = 16'(-4272);
			24455: out = 16'(-2343);
			24456: out = 16'(-1484);
			24457: out = 16'(-1056);
			24458: out = 16'(-963);
			24459: out = 16'(1077);
			24460: out = 16'(3484);
			24461: out = 16'(498);
			24462: out = 16'(-3254);
			24463: out = 16'(-4748);
			24464: out = 16'(-2191);
			24465: out = 16'(1678);
			24466: out = 16'(1044);
			24467: out = 16'(-1422);
			24468: out = 16'(-103);
			24469: out = 16'(3102);
			24470: out = 16'(4472);
			24471: out = 16'(295);
			24472: out = 16'(-3310);
			24473: out = 16'(-3178);
			24474: out = 16'(-285);
			24475: out = 16'(-2675);
			24476: out = 16'(-3426);
			24477: out = 16'(2722);
			24478: out = 16'(3753);
			24479: out = 16'(1336);
			24480: out = 16'(446);
			24481: out = 16'(4080);
			24482: out = 16'(3630);
			24483: out = 16'(-2159);
			24484: out = 16'(-7114);
			24485: out = 16'(-4380);
			24486: out = 16'(-856);
			24487: out = 16'(982);
			24488: out = 16'(430);
			24489: out = 16'(3142);
			24490: out = 16'(7199);
			24491: out = 16'(4303);
			24492: out = 16'(-4809);
			24493: out = 16'(-11137);
			24494: out = 16'(-6567);
			24495: out = 16'(1732);
			24496: out = 16'(5148);
			24497: out = 16'(1340);
			24498: out = 16'(-2600);
			24499: out = 16'(-1759);
			24500: out = 16'(1614);
			24501: out = 16'(1445);
			24502: out = 16'(-228);
			24503: out = 16'(-414);
			24504: out = 16'(4534);
			24505: out = 16'(3181);
			24506: out = 16'(-3715);
			24507: out = 16'(-5058);
			24508: out = 16'(-162);
			24509: out = 16'(3899);
			24510: out = 16'(1442);
			24511: out = 16'(-589);
			24512: out = 16'(-1128);
			24513: out = 16'(3524);
			24514: out = 16'(3817);
			24515: out = 16'(-369);
			24516: out = 16'(-690);
			24517: out = 16'(2401);
			24518: out = 16'(2303);
			24519: out = 16'(-2246);
			24520: out = 16'(-5472);
			24521: out = 16'(-2238);
			24522: out = 16'(534);
			24523: out = 16'(-574);
			24524: out = 16'(122);
			24525: out = 16'(811);
			24526: out = 16'(2090);
			24527: out = 16'(2314);
			24528: out = 16'(3694);
			24529: out = 16'(-534);
			24530: out = 16'(-1338);
			24531: out = 16'(443);
			24532: out = 16'(1883);
			24533: out = 16'(16);
			24534: out = 16'(-2911);
			24535: out = 16'(-3493);
			24536: out = 16'(-401);
			24537: out = 16'(4540);
			24538: out = 16'(3490);
			24539: out = 16'(564);
			24540: out = 16'(-91);
			24541: out = 16'(932);
			24542: out = 16'(380);
			24543: out = 16'(-3053);
			24544: out = 16'(-6374);
			24545: out = 16'(-5438);
			24546: out = 16'(-1488);
			24547: out = 16'(1804);
			24548: out = 16'(1677);
			24549: out = 16'(-23);
			24550: out = 16'(-268);
			24551: out = 16'(947);
			24552: out = 16'(1566);
			24553: out = 16'(1381);
			24554: out = 16'(-264);
			24555: out = 16'(-2328);
			24556: out = 16'(-5093);
			24557: out = 16'(-4540);
			24558: out = 16'(-871);
			24559: out = 16'(4143);
			24560: out = 16'(1590);
			24561: out = 16'(-3091);
			24562: out = 16'(-766);
			24563: out = 16'(4022);
			24564: out = 16'(5063);
			24565: out = 16'(3406);
			24566: out = 16'(3578);
			24567: out = 16'(-1070);
			24568: out = 16'(-4224);
			24569: out = 16'(-3445);
			24570: out = 16'(-64);
			24571: out = 16'(69);
			24572: out = 16'(-5082);
			24573: out = 16'(-5530);
			24574: out = 16'(1958);
			24575: out = 16'(1750);
			24576: out = 16'(2321);
			24577: out = 16'(1084);
			24578: out = 16'(1940);
			24579: out = 16'(1111);
			24580: out = 16'(2545);
			24581: out = 16'(-224);
			24582: out = 16'(-3891);
			24583: out = 16'(-5509);
			24584: out = 16'(-4892);
			24585: out = 16'(-2207);
			24586: out = 16'(2123);
			24587: out = 16'(5285);
			24588: out = 16'(4358);
			24589: out = 16'(1277);
			24590: out = 16'(-300);
			24591: out = 16'(-301);
			24592: out = 16'(-2521);
			24593: out = 16'(-4294);
			24594: out = 16'(-2987);
			24595: out = 16'(839);
			24596: out = 16'(1393);
			24597: out = 16'(2516);
			24598: out = 16'(1309);
			24599: out = 16'(-452);
			24600: out = 16'(-841);
			24601: out = 16'(894);
			24602: out = 16'(2390);
			24603: out = 16'(1529);
			24604: out = 16'(-324);
			24605: out = 16'(-3524);
			24606: out = 16'(-1781);
			24607: out = 16'(341);
			24608: out = 16'(790);
			24609: out = 16'(2126);
			24610: out = 16'(4855);
			24611: out = 16'(5424);
			24612: out = 16'(2848);
			24613: out = 16'(-49);
			24614: out = 16'(-4646);
			24615: out = 16'(-7994);
			24616: out = 16'(-5077);
			24617: out = 16'(3427);
			24618: out = 16'(5848);
			24619: out = 16'(-278);
			24620: out = 16'(-5901);
			24621: out = 16'(-1298);
			24622: out = 16'(1513);
			24623: out = 16'(1455);
			24624: out = 16'(-675);
			24625: out = 16'(549);
			24626: out = 16'(3122);
			24627: out = 16'(2935);
			24628: out = 16'(-1118);
			24629: out = 16'(-5056);
			24630: out = 16'(-5536);
			24631: out = 16'(-2034);
			24632: out = 16'(2278);
			24633: out = 16'(3247);
			24634: out = 16'(99);
			24635: out = 16'(-1220);
			24636: out = 16'(553);
			24637: out = 16'(2416);
			24638: out = 16'(1334);
			24639: out = 16'(-59);
			24640: out = 16'(-295);
			24641: out = 16'(-422);
			24642: out = 16'(-1425);
			24643: out = 16'(-5315);
			24644: out = 16'(-2630);
			24645: out = 16'(613);
			24646: out = 16'(-828);
			24647: out = 16'(-4821);
			24648: out = 16'(-951);
			24649: out = 16'(7003);
			24650: out = 16'(9276);
			24651: out = 16'(1744);
			24652: out = 16'(-3971);
			24653: out = 16'(-6187);
			24654: out = 16'(-5590);
			24655: out = 16'(-7482);
			24656: out = 16'(-5571);
			24657: out = 16'(-2728);
			24658: out = 16'(3141);
			24659: out = 16'(7263);
			24660: out = 16'(6525);
			24661: out = 16'(-831);
			24662: out = 16'(-4464);
			24663: out = 16'(-1133);
			24664: out = 16'(515);
			24665: out = 16'(-1352);
			24666: out = 16'(-1847);
			24667: out = 16'(1546);
			24668: out = 16'(1497);
			24669: out = 16'(145);
			24670: out = 16'(-1063);
			24671: out = 16'(530);
			24672: out = 16'(-181);
			24673: out = 16'(1847);
			24674: out = 16'(740);
			24675: out = 16'(539);
			24676: out = 16'(1602);
			24677: out = 16'(2020);
			24678: out = 16'(-1878);
			24679: out = 16'(-5006);
			24680: out = 16'(-2678);
			24681: out = 16'(921);
			24682: out = 16'(2517);
			24683: out = 16'(-646);
			24684: out = 16'(-4394);
			24685: out = 16'(-896);
			24686: out = 16'(1565);
			24687: out = 16'(4395);
			24688: out = 16'(6093);
			24689: out = 16'(3578);
			24690: out = 16'(2568);
			24691: out = 16'(-2961);
			24692: out = 16'(-7875);
			24693: out = 16'(-3704);
			24694: out = 16'(-1254);
			24695: out = 16'(4142);
			24696: out = 16'(6611);
			24697: out = 16'(7583);
			24698: out = 16'(6778);
			24699: out = 16'(3182);
			24700: out = 16'(-9484);
			24701: out = 16'(-22152);
			24702: out = 16'(-6013);
			24703: out = 16'(6359);
			24704: out = 16'(8338);
			24705: out = 16'(2589);
			24706: out = 16'(554);
			24707: out = 16'(1599);
			24708: out = 16'(1804);
			24709: out = 16'(-1116);
			24710: out = 16'(-2366);
			24711: out = 16'(-1011);
			24712: out = 16'(1653);
			24713: out = 16'(2077);
			24714: out = 16'(393);
			24715: out = 16'(-761);
			24716: out = 16'(-822);
			24717: out = 16'(1766);
			24718: out = 16'(4002);
			24719: out = 16'(-3071);
			24720: out = 16'(-4409);
			24721: out = 16'(-1369);
			24722: out = 16'(1588);
			24723: out = 16'(-901);
			24724: out = 16'(-708);
			24725: out = 16'(1987);
			24726: out = 16'(3586);
			24727: out = 16'(402);
			24728: out = 16'(-2227);
			24729: out = 16'(-2177);
			24730: out = 16'(-737);
			24731: out = 16'(-1142);
			24732: out = 16'(-957);
			24733: out = 16'(852);
			24734: out = 16'(4385);
			24735: out = 16'(7126);
			24736: out = 16'(1741);
			24737: out = 16'(444);
			24738: out = 16'(-2569);
			24739: out = 16'(-5964);
			24740: out = 16'(-5642);
			24741: out = 16'(-1638);
			24742: out = 16'(353);
			24743: out = 16'(238);
			24744: out = 16'(1652);
			24745: out = 16'(2505);
			24746: out = 16'(-515);
			24747: out = 16'(-4418);
			24748: out = 16'(-3160);
			24749: out = 16'(-1574);
			24750: out = 16'(-531);
			24751: out = 16'(-822);
			24752: out = 16'(649);
			24753: out = 16'(1361);
			24754: out = 16'(2626);
			24755: out = 16'(1605);
			24756: out = 16'(-382);
			24757: out = 16'(-3396);
			24758: out = 16'(-3067);
			24759: out = 16'(-1371);
			24760: out = 16'(610);
			24761: out = 16'(21);
			24762: out = 16'(3499);
			24763: out = 16'(3194);
			24764: out = 16'(1102);
			24765: out = 16'(32);
			24766: out = 16'(2077);
			24767: out = 16'(1787);
			24768: out = 16'(112);
			24769: out = 16'(-864);
			24770: out = 16'(2177);
			24771: out = 16'(-1021);
			24772: out = 16'(-4935);
			24773: out = 16'(-3146);
			24774: out = 16'(3083);
			24775: out = 16'(3354);
			24776: out = 16'(-1845);
			24777: out = 16'(-4983);
			24778: out = 16'(-1058);
			24779: out = 16'(4757);
			24780: out = 16'(4984);
			24781: out = 16'(1119);
			24782: out = 16'(-744);
			24783: out = 16'(-429);
			24784: out = 16'(-111);
			24785: out = 16'(-2667);
			24786: out = 16'(-6101);
			24787: out = 16'(-2563);
			24788: out = 16'(1991);
			24789: out = 16'(5283);
			24790: out = 16'(5432);
			24791: out = 16'(522);
			24792: out = 16'(-1031);
			24793: out = 16'(-946);
			24794: out = 16'(-1520);
			24795: out = 16'(-3403);
			24796: out = 16'(-3316);
			24797: out = 16'(-427);
			24798: out = 16'(2061);
			24799: out = 16'(1617);
			24800: out = 16'(-382);
			24801: out = 16'(102);
			24802: out = 16'(2746);
			24803: out = 16'(3621);
			24804: out = 16'(2193);
			24805: out = 16'(-260);
			24806: out = 16'(-1191);
			24807: out = 16'(-1420);
			24808: out = 16'(-4192);
			24809: out = 16'(-3669);
			24810: out = 16'(-1189);
			24811: out = 16'(185);
			24812: out = 16'(380);
			24813: out = 16'(1609);
			24814: out = 16'(4078);
			24815: out = 16'(3765);
			24816: out = 16'(135);
			24817: out = 16'(-489);
			24818: out = 16'(2345);
			24819: out = 16'(3277);
			24820: out = 16'(489);
			24821: out = 16'(-2602);
			24822: out = 16'(-1685);
			24823: out = 16'(-2295);
			24824: out = 16'(-4812);
			24825: out = 16'(1278);
			24826: out = 16'(7392);
			24827: out = 16'(6073);
			24828: out = 16'(-809);
			24829: out = 16'(1545);
			24830: out = 16'(2981);
			24831: out = 16'(1670);
			24832: out = 16'(-3215);
			24833: out = 16'(-4102);
			24834: out = 16'(-2395);
			24835: out = 16'(1006);
			24836: out = 16'(1870);
			24837: out = 16'(-278);
			24838: out = 16'(-73);
			24839: out = 16'(-1018);
			24840: out = 16'(-129);
			24841: out = 16'(2143);
			24842: out = 16'(1769);
			24843: out = 16'(-1347);
			24844: out = 16'(-2513);
			24845: out = 16'(-923);
			24846: out = 16'(695);
			24847: out = 16'(-5340);
			24848: out = 16'(-5892);
			24849: out = 16'(3275);
			24850: out = 16'(7801);
			24851: out = 16'(3416);
			24852: out = 16'(-4762);
			24853: out = 16'(-5533);
			24854: out = 16'(-536);
			24855: out = 16'(232);
			24856: out = 16'(-5711);
			24857: out = 16'(-7093);
			24858: out = 16'(1411);
			24859: out = 16'(3627);
			24860: out = 16'(2661);
			24861: out = 16'(2643);
			24862: out = 16'(5737);
			24863: out = 16'(418);
			24864: out = 16'(-1007);
			24865: out = 16'(884);
			24866: out = 16'(4359);
			24867: out = 16'(-1142);
			24868: out = 16'(-2149);
			24869: out = 16'(-2986);
			24870: out = 16'(-2645);
			24871: out = 16'(-4426);
			24872: out = 16'(1030);
			24873: out = 16'(3559);
			24874: out = 16'(3517);
			24875: out = 16'(2266);
			24876: out = 16'(3536);
			24877: out = 16'(1874);
			24878: out = 16'(-2179);
			24879: out = 16'(-6060);
			24880: out = 16'(-3135);
			24881: out = 16'(-752);
			24882: out = 16'(275);
			24883: out = 16'(183);
			24884: out = 16'(2360);
			24885: out = 16'(795);
			24886: out = 16'(-249);
			24887: out = 16'(587);
			24888: out = 16'(3619);
			24889: out = 16'(962);
			24890: out = 16'(-477);
			24891: out = 16'(-479);
			24892: out = 16'(-2990);
			24893: out = 16'(-1764);
			24894: out = 16'(-2943);
			24895: out = 16'(-2868);
			24896: out = 16'(177);
			24897: out = 16'(1964);
			24898: out = 16'(2477);
			24899: out = 16'(2172);
			24900: out = 16'(2055);
			24901: out = 16'(-947);
			24902: out = 16'(465);
			24903: out = 16'(1888);
			24904: out = 16'(180);
			24905: out = 16'(-6673);
			24906: out = 16'(-2670);
			24907: out = 16'(2938);
			24908: out = 16'(1443);
			24909: out = 16'(-7590);
			24910: out = 16'(-6047);
			24911: out = 16'(2298);
			24912: out = 16'(7348);
			24913: out = 16'(3064);
			24914: out = 16'(-87);
			24915: out = 16'(-1089);
			24916: out = 16'(210);
			24917: out = 16'(-838);
			24918: out = 16'(-3742);
			24919: out = 16'(-2353);
			24920: out = 16'(2764);
			24921: out = 16'(4908);
			24922: out = 16'(4143);
			24923: out = 16'(470);
			24924: out = 16'(1470);
			24925: out = 16'(3500);
			24926: out = 16'(1169);
			24927: out = 16'(-6839);
			24928: out = 16'(-7817);
			24929: out = 16'(-572);
			24930: out = 16'(3157);
			24931: out = 16'(5266);
			24932: out = 16'(-1550);
			24933: out = 16'(-5146);
			24934: out = 16'(67);
			24935: out = 16'(4741);
			24936: out = 16'(3802);
			24937: out = 16'(-1567);
			24938: out = 16'(-3955);
			24939: out = 16'(-166);
			24940: out = 16'(137);
			24941: out = 16'(-4235);
			24942: out = 16'(-5848);
			24943: out = 16'(2192);
			24944: out = 16'(4927);
			24945: out = 16'(2735);
			24946: out = 16'(-834);
			24947: out = 16'(-765);
			24948: out = 16'(2890);
			24949: out = 16'(2070);
			24950: out = 16'(-1341);
			24951: out = 16'(-1441);
			24952: out = 16'(-699);
			24953: out = 16'(2629);
			24954: out = 16'(2887);
			24955: out = 16'(-578);
			24956: out = 16'(-5662);
			24957: out = 16'(-2252);
			24958: out = 16'(4437);
			24959: out = 16'(6113);
			24960: out = 16'(2499);
			24961: out = 16'(867);
			24962: out = 16'(2866);
			24963: out = 16'(1454);
			24964: out = 16'(-5456);
			24965: out = 16'(-7811);
			24966: out = 16'(-1252);
			24967: out = 16'(4128);
			24968: out = 16'(771);
			24969: out = 16'(174);
			24970: out = 16'(1023);
			24971: out = 16'(1935);
			24972: out = 16'(348);
			24973: out = 16'(1254);
			24974: out = 16'(2838);
			24975: out = 16'(1982);
			24976: out = 16'(-2961);
			24977: out = 16'(-8883);
			24978: out = 16'(-6958);
			24979: out = 16'(-3768);
			24980: out = 16'(-2148);
			24981: out = 16'(370);
			24982: out = 16'(4614);
			24983: out = 16'(6086);
			24984: out = 16'(3430);
			24985: out = 16'(-673);
			24986: out = 16'(-3946);
			24987: out = 16'(-5006);
			24988: out = 16'(-2869);
			24989: out = 16'(1032);
			24990: out = 16'(2183);
			24991: out = 16'(862);
			24992: out = 16'(-661);
			24993: out = 16'(-1376);
			24994: out = 16'(-4265);
			24995: out = 16'(-1486);
			24996: out = 16'(1596);
			24997: out = 16'(2078);
			24998: out = 16'(886);
			24999: out = 16'(-292);
			25000: out = 16'(2042);
			25001: out = 16'(3449);
			25002: out = 16'(386);
			25003: out = 16'(-2025);
			25004: out = 16'(-2928);
			25005: out = 16'(-2479);
			25006: out = 16'(-2269);
			25007: out = 16'(2008);
			25008: out = 16'(1337);
			25009: out = 16'(-1622);
			25010: out = 16'(-2595);
			25011: out = 16'(3331);
			25012: out = 16'(4404);
			25013: out = 16'(932);
			25014: out = 16'(-2890);
			25015: out = 16'(-775);
			25016: out = 16'(2683);
			25017: out = 16'(3284);
			25018: out = 16'(85);
			25019: out = 16'(-2300);
			25020: out = 16'(410);
			25021: out = 16'(3367);
			25022: out = 16'(1953);
			25023: out = 16'(-3153);
			25024: out = 16'(-3408);
			25025: out = 16'(-3164);
			25026: out = 16'(-2433);
			25027: out = 16'(-2340);
			25028: out = 16'(1714);
			25029: out = 16'(355);
			25030: out = 16'(1980);
			25031: out = 16'(5993);
			25032: out = 16'(6580);
			25033: out = 16'(1964);
			25034: out = 16'(-2606);
			25035: out = 16'(-3285);
			25036: out = 16'(-2226);
			25037: out = 16'(-4403);
			25038: out = 16'(-5250);
			25039: out = 16'(-133);
			25040: out = 16'(7168);
			25041: out = 16'(6178);
			25042: out = 16'(2001);
			25043: out = 16'(-596);
			25044: out = 16'(-196);
			25045: out = 16'(-1781);
			25046: out = 16'(-2247);
			25047: out = 16'(214);
			25048: out = 16'(3926);
			25049: out = 16'(1978);
			25050: out = 16'(-703);
			25051: out = 16'(-1990);
			25052: out = 16'(961);
			25053: out = 16'(2968);
			25054: out = 16'(1296);
			25055: out = 16'(-4916);
			25056: out = 16'(-7241);
			25057: out = 16'(-291);
			25058: out = 16'(4502);
			25059: out = 16'(4522);
			25060: out = 16'(-603);
			25061: out = 16'(-4124);
			25062: out = 16'(-978);
			25063: out = 16'(1598);
			25064: out = 16'(-839);
			25065: out = 16'(-4868);
			25066: out = 16'(-5398);
			25067: out = 16'(32);
			25068: out = 16'(4213);
			25069: out = 16'(4444);
			25070: out = 16'(-282);
			25071: out = 16'(234);
			25072: out = 16'(-3998);
			25073: out = 16'(-9266);
			25074: out = 16'(-10372);
			25075: out = 16'(-1840);
			25076: out = 16'(1920);
			25077: out = 16'(2009);
			25078: out = 16'(2973);
			25079: out = 16'(5683);
			25080: out = 16'(3598);
			25081: out = 16'(107);
			25082: out = 16'(-1936);
			25083: out = 16'(-2338);
			25084: out = 16'(-3384);
			25085: out = 16'(-1850);
			25086: out = 16'(349);
			25087: out = 16'(-577);
			25088: out = 16'(-375);
			25089: out = 16'(3362);
			25090: out = 16'(5040);
			25091: out = 16'(-1202);
			25092: out = 16'(-4461);
			25093: out = 16'(-3244);
			25094: out = 16'(143);
			25095: out = 16'(121);
			25096: out = 16'(1650);
			25097: out = 16'(3967);
			25098: out = 16'(4701);
			25099: out = 16'(516);
			25100: out = 16'(-2634);
			25101: out = 16'(-3570);
			25102: out = 16'(-452);
			25103: out = 16'(1580);
			25104: out = 16'(286);
			25105: out = 16'(358);
			25106: out = 16'(1412);
			25107: out = 16'(1229);
			25108: out = 16'(235);
			25109: out = 16'(-251);
			25110: out = 16'(1454);
			25111: out = 16'(1842);
			25112: out = 16'(-19);
			25113: out = 16'(-364);
			25114: out = 16'(3294);
			25115: out = 16'(5813);
			25116: out = 16'(2661);
			25117: out = 16'(1215);
			25118: out = 16'(-4972);
			25119: out = 16'(-7106);
			25120: out = 16'(-2732);
			25121: out = 16'(4408);
			25122: out = 16'(2205);
			25123: out = 16'(-3028);
			25124: out = 16'(-2280);
			25125: out = 16'(6727);
			25126: out = 16'(6566);
			25127: out = 16'(1711);
			25128: out = 16'(-540);
			25129: out = 16'(3527);
			25130: out = 16'(531);
			25131: out = 16'(-4066);
			25132: out = 16'(-5571);
			25133: out = 16'(-391);
			25134: out = 16'(214);
			25135: out = 16'(416);
			25136: out = 16'(-981);
			25137: out = 16'(-667);
			25138: out = 16'(1132);
			25139: out = 16'(2195);
			25140: out = 16'(1176);
			25141: out = 16'(-446);
			25142: out = 16'(-76);
			25143: out = 16'(-1085);
			25144: out = 16'(-692);
			25145: out = 16'(-273);
			25146: out = 16'(-1142);
			25147: out = 16'(-508);
			25148: out = 16'(-577);
			25149: out = 16'(-1768);
			25150: out = 16'(-2427);
			25151: out = 16'(-853);
			25152: out = 16'(2624);
			25153: out = 16'(2658);
			25154: out = 16'(-897);
			25155: out = 16'(-2529);
			25156: out = 16'(-1629);
			25157: out = 16'(-2051);
			25158: out = 16'(-4727);
			25159: out = 16'(-2134);
			25160: out = 16'(1759);
			25161: out = 16'(6394);
			25162: out = 16'(5388);
			25163: out = 16'(-295);
			25164: out = 16'(-6146);
			25165: out = 16'(-6631);
			25166: out = 16'(-4213);
			25167: out = 16'(-1254);
			25168: out = 16'(1704);
			25169: out = 16'(5094);
			25170: out = 16'(4207);
			25171: out = 16'(-390);
			25172: out = 16'(707);
			25173: out = 16'(104);
			25174: out = 16'(-655);
			25175: out = 16'(-840);
			25176: out = 16'(-376);
			25177: out = 16'(2993);
			25178: out = 16'(2348);
			25179: out = 16'(-1004);
			25180: out = 16'(-2458);
			25181: out = 16'(555);
			25182: out = 16'(1261);
			25183: out = 16'(-1233);
			25184: out = 16'(-3275);
			25185: out = 16'(-610);
			25186: out = 16'(448);
			25187: out = 16'(-866);
			25188: out = 16'(-2410);
			25189: out = 16'(-129);
			25190: out = 16'(2513);
			25191: out = 16'(4335);
			25192: out = 16'(3255);
			25193: out = 16'(4128);
			25194: out = 16'(-5551);
			25195: out = 16'(-9948);
			25196: out = 16'(-6147);
			25197: out = 16'(66);
			25198: out = 16'(1961);
			25199: out = 16'(5299);
			25200: out = 16'(7505);
			25201: out = 16'(2866);
			25202: out = 16'(-2714);
			25203: out = 16'(-5541);
			25204: out = 16'(-2540);
			25205: out = 16'(-227);
			25206: out = 16'(454);
			25207: out = 16'(-2326);
			25208: out = 16'(272);
			25209: out = 16'(6964);
			25210: out = 16'(9901);
			25211: out = 16'(3496);
			25212: out = 16'(-3968);
			25213: out = 16'(-5533);
			25214: out = 16'(-1422);
			25215: out = 16'(-782);
			25216: out = 16'(-1357);
			25217: out = 16'(-247);
			25218: out = 16'(1461);
			25219: out = 16'(4165);
			25220: out = 16'(2088);
			25221: out = 16'(-954);
			25222: out = 16'(-719);
			25223: out = 16'(1613);
			25224: out = 16'(1237);
			25225: out = 16'(-1625);
			25226: out = 16'(-2071);
			25227: out = 16'(1463);
			25228: out = 16'(5155);
			25229: out = 16'(2787);
			25230: out = 16'(-3314);
			25231: out = 16'(-5115);
			25232: out = 16'(-1949);
			25233: out = 16'(1107);
			25234: out = 16'(-995);
			25235: out = 16'(-5783);
			25236: out = 16'(-2050);
			25237: out = 16'(4414);
			25238: out = 16'(6866);
			25239: out = 16'(4523);
			25240: out = 16'(-456);
			25241: out = 16'(-1081);
			25242: out = 16'(-884);
			25243: out = 16'(-3757);
			25244: out = 16'(-8383);
			25245: out = 16'(-6853);
			25246: out = 16'(-1009);
			25247: out = 16'(2968);
			25248: out = 16'(5916);
			25249: out = 16'(2603);
			25250: out = 16'(373);
			25251: out = 16'(-2154);
			25252: out = 16'(-5053);
			25253: out = 16'(-5836);
			25254: out = 16'(-1199);
			25255: out = 16'(3631);
			25256: out = 16'(4164);
			25257: out = 16'(-762);
			25258: out = 16'(-1147);
			25259: out = 16'(960);
			25260: out = 16'(1439);
			25261: out = 16'(845);
			25262: out = 16'(282);
			25263: out = 16'(-362);
			25264: out = 16'(-551);
			25265: out = 16'(2123);
			25266: out = 16'(3620);
			25267: out = 16'(2125);
			25268: out = 16'(-391);
			25269: out = 16'(1563);
			25270: out = 16'(317);
			25271: out = 16'(-2168);
			25272: out = 16'(-4857);
			25273: out = 16'(-3016);
			25274: out = 16'(-1021);
			25275: out = 16'(1348);
			25276: out = 16'(1617);
			25277: out = 16'(2797);
			25278: out = 16'(3121);
			25279: out = 16'(4829);
			25280: out = 16'(1028);
			25281: out = 16'(-6029);
			25282: out = 16'(-6029);
			25283: out = 16'(-2155);
			25284: out = 16'(2119);
			25285: out = 16'(4363);
			25286: out = 16'(6849);
			25287: out = 16'(3681);
			25288: out = 16'(-589);
			25289: out = 16'(-2697);
			25290: out = 16'(-1173);
			25291: out = 16'(-54);
			25292: out = 16'(-1979);
			25293: out = 16'(-3202);
			25294: out = 16'(362);
			25295: out = 16'(3526);
			25296: out = 16'(6193);
			25297: out = 16'(6032);
			25298: out = 16'(2331);
			25299: out = 16'(-2800);
			25300: out = 16'(-5831);
			25301: out = 16'(-3681);
			25302: out = 16'(-1325);
			25303: out = 16'(-1496);
			25304: out = 16'(-3322);
			25305: out = 16'(1833);
			25306: out = 16'(7090);
			25307: out = 16'(4015);
			25308: out = 16'(-4162);
			25309: out = 16'(-4269);
			25310: out = 16'(1317);
			25311: out = 16'(666);
			25312: out = 16'(-2444);
			25313: out = 16'(-2993);
			25314: out = 16'(51);
			25315: out = 16'(-623);
			25316: out = 16'(-477);
			25317: out = 16'(-668);
			25318: out = 16'(1871);
			25319: out = 16'(1138);
			25320: out = 16'(-2628);
			25321: out = 16'(-6982);
			25322: out = 16'(-2705);
			25323: out = 16'(5307);
			25324: out = 16'(7192);
			25325: out = 16'(812);
			25326: out = 16'(-3782);
			25327: out = 16'(-2482);
			25328: out = 16'(-462);
			25329: out = 16'(391);
			25330: out = 16'(-1627);
			25331: out = 16'(-2167);
			25332: out = 16'(373);
			25333: out = 16'(4998);
			25334: out = 16'(3101);
			25335: out = 16'(-3729);
			25336: out = 16'(-8239);
			25337: out = 16'(-1138);
			25338: out = 16'(3377);
			25339: out = 16'(1747);
			25340: out = 16'(-1685);
			25341: out = 16'(1523);
			25342: out = 16'(3371);
			25343: out = 16'(1197);
			25344: out = 16'(-3953);
			25345: out = 16'(-3819);
			25346: out = 16'(298);
			25347: out = 16'(5120);
			25348: out = 16'(3914);
			25349: out = 16'(-1288);
			25350: out = 16'(-3557);
			25351: out = 16'(-2108);
			25352: out = 16'(-1368);
			25353: out = 16'(-2441);
			25354: out = 16'(1849);
			25355: out = 16'(4811);
			25356: out = 16'(4564);
			25357: out = 16'(539);
			25358: out = 16'(303);
			25359: out = 16'(-316);
			25360: out = 16'(2462);
			25361: out = 16'(4144);
			25362: out = 16'(3490);
			25363: out = 16'(-447);
			25364: out = 16'(-1967);
			25365: out = 16'(-2645);
			25366: out = 16'(-3692);
			25367: out = 16'(-3365);
			25368: out = 16'(845);
			25369: out = 16'(4685);
			25370: out = 16'(5262);
			25371: out = 16'(3536);
			25372: out = 16'(1557);
			25373: out = 16'(-2320);
			25374: out = 16'(-5685);
			25375: out = 16'(-3381);
			25376: out = 16'(1777);
			25377: out = 16'(3046);
			25378: out = 16'(524);
			25379: out = 16'(-262);
			25380: out = 16'(-1068);
			25381: out = 16'(-3083);
			25382: out = 16'(-4725);
			25383: out = 16'(-2624);
			25384: out = 16'(-224);
			25385: out = 16'(1150);
			25386: out = 16'(2014);
			25387: out = 16'(3372);
			25388: out = 16'(215);
			25389: out = 16'(-766);
			25390: out = 16'(343);
			25391: out = 16'(1163);
			25392: out = 16'(2255);
			25393: out = 16'(-672);
			25394: out = 16'(-404);
			25395: out = 16'(1494);
			25396: out = 16'(3536);
			25397: out = 16'(-5751);
			25398: out = 16'(-7096);
			25399: out = 16'(-1061);
			25400: out = 16'(804);
			25401: out = 16'(-3886);
			25402: out = 16'(-5027);
			25403: out = 16'(-620);
			25404: out = 16'(1953);
			25405: out = 16'(1143);
			25406: out = 16'(-327);
			25407: out = 16'(495);
			25408: out = 16'(1322);
			25409: out = 16'(66);
			25410: out = 16'(-1776);
			25411: out = 16'(-4248);
			25412: out = 16'(-6034);
			25413: out = 16'(-3397);
			25414: out = 16'(-786);
			25415: out = 16'(239);
			25416: out = 16'(-1421);
			25417: out = 16'(-973);
			25418: out = 16'(4940);
			25419: out = 16'(9690);
			25420: out = 16'(4566);
			25421: out = 16'(-7268);
			25422: out = 16'(-6239);
			25423: out = 16'(589);
			25424: out = 16'(3011);
			25425: out = 16'(-2638);
			25426: out = 16'(-2982);
			25427: out = 16'(-2528);
			25428: out = 16'(-1909);
			25429: out = 16'(-3124);
			25430: out = 16'(2026);
			25431: out = 16'(1673);
			25432: out = 16'(1319);
			25433: out = 16'(-507);
			25434: out = 16'(494);
			25435: out = 16'(24);
			25436: out = 16'(3120);
			25437: out = 16'(2190);
			25438: out = 16'(-3372);
			25439: out = 16'(-3135);
			25440: out = 16'(3405);
			25441: out = 16'(7299);
			25442: out = 16'(2289);
			25443: out = 16'(-4577);
			25444: out = 16'(-6660);
			25445: out = 16'(-2129);
			25446: out = 16'(2160);
			25447: out = 16'(3997);
			25448: out = 16'(1086);
			25449: out = 16'(697);
			25450: out = 16'(3115);
			25451: out = 16'(4108);
			25452: out = 16'(598);
			25453: out = 16'(-3070);
			25454: out = 16'(-2263);
			25455: out = 16'(1697);
			25456: out = 16'(6994);
			25457: out = 16'(4601);
			25458: out = 16'(-574);
			25459: out = 16'(-2599);
			25460: out = 16'(-1563);
			25461: out = 16'(-882);
			25462: out = 16'(-1301);
			25463: out = 16'(-780);
			25464: out = 16'(-310);
			25465: out = 16'(2717);
			25466: out = 16'(3109);
			25467: out = 16'(1235);
			25468: out = 16'(3791);
			25469: out = 16'(-209);
			25470: out = 16'(-2215);
			25471: out = 16'(-2695);
			25472: out = 16'(-179);
			25473: out = 16'(-7079);
			25474: out = 16'(-4535);
			25475: out = 16'(2601);
			25476: out = 16'(5372);
			25477: out = 16'(4116);
			25478: out = 16'(3286);
			25479: out = 16'(3134);
			25480: out = 16'(102);
			25481: out = 16'(-6309);
			25482: out = 16'(-6989);
			25483: out = 16'(-2773);
			25484: out = 16'(-36);
			25485: out = 16'(137);
			25486: out = 16'(522);
			25487: out = 16'(4569);
			25488: out = 16'(5870);
			25489: out = 16'(-456);
			25490: out = 16'(-8108);
			25491: out = 16'(-9301);
			25492: out = 16'(-3762);
			25493: out = 16'(-493);
			25494: out = 16'(-834);
			25495: out = 16'(-2651);
			25496: out = 16'(-180);
			25497: out = 16'(4104);
			25498: out = 16'(3904);
			25499: out = 16'(23);
			25500: out = 16'(-4814);
			25501: out = 16'(-7381);
			25502: out = 16'(-4784);
			25503: out = 16'(-173);
			25504: out = 16'(4246);
			25505: out = 16'(4596);
			25506: out = 16'(2041);
			25507: out = 16'(176);
			25508: out = 16'(967);
			25509: out = 16'(-1151);
			25510: out = 16'(-7473);
			25511: out = 16'(-11078);
			25512: out = 16'(-4734);
			25513: out = 16'(3945);
			25514: out = 16'(5217);
			25515: out = 16'(7469);
			25516: out = 16'(5121);
			25517: out = 16'(2252);
			25518: out = 16'(-1145);
			25519: out = 16'(-487);
			25520: out = 16'(-2442);
			25521: out = 16'(-3272);
			25522: out = 16'(-2425);
			25523: out = 16'(451);
			25524: out = 16'(3051);
			25525: out = 16'(5177);
			25526: out = 16'(5438);
			25527: out = 16'(3484);
			25528: out = 16'(897);
			25529: out = 16'(-2433);
			25530: out = 16'(-4795);
			25531: out = 16'(-4428);
			25532: out = 16'(1394);
			25533: out = 16'(4834);
			25534: out = 16'(5627);
			25535: out = 16'(4721);
			25536: out = 16'(4360);
			25537: out = 16'(-239);
			25538: out = 16'(-5115);
			25539: out = 16'(-6038);
			25540: out = 16'(-375);
			25541: out = 16'(2875);
			25542: out = 16'(3295);
			25543: out = 16'(1771);
			25544: out = 16'(2538);
			25545: out = 16'(4330);
			25546: out = 16'(6114);
			25547: out = 16'(2424);
			25548: out = 16'(-4771);
			25549: out = 16'(-7916);
			25550: out = 16'(-3477);
			25551: out = 16'(1189);
			25552: out = 16'(1080);
			25553: out = 16'(139);
			25554: out = 16'(835);
			25555: out = 16'(835);
			25556: out = 16'(-1768);
			25557: out = 16'(-3996);
			25558: out = 16'(-1582);
			25559: out = 16'(504);
			25560: out = 16'(-113);
			25561: out = 16'(1884);
			25562: out = 16'(375);
			25563: out = 16'(2267);
			25564: out = 16'(3274);
			25565: out = 16'(980);
			25566: out = 16'(-2606);
			25567: out = 16'(-4883);
			25568: out = 16'(-4532);
			25569: out = 16'(-1943);
			25570: out = 16'(1691);
			25571: out = 16'(4651);
			25572: out = 16'(5116);
			25573: out = 16'(2677);
			25574: out = 16'(52);
			25575: out = 16'(-2300);
			25576: out = 16'(-2786);
			25577: out = 16'(-2537);
			25578: out = 16'(-932);
			25579: out = 16'(-3016);
			25580: out = 16'(-2491);
			25581: out = 16'(735);
			25582: out = 16'(5638);
			25583: out = 16'(1995);
			25584: out = 16'(545);
			25585: out = 16'(-570);
			25586: out = 16'(-1208);
			25587: out = 16'(-7372);
			25588: out = 16'(-4701);
			25589: out = 16'(-1100);
			25590: out = 16'(730);
			25591: out = 16'(3310);
			25592: out = 16'(6891);
			25593: out = 16'(4600);
			25594: out = 16'(-963);
			25595: out = 16'(-742);
			25596: out = 16'(-337);
			25597: out = 16'(-1019);
			25598: out = 16'(-2956);
			25599: out = 16'(-2333);
			25600: out = 16'(-382);
			25601: out = 16'(-314);
			25602: out = 16'(-269);
			25603: out = 16'(2735);
			25604: out = 16'(5096);
			25605: out = 16'(1703);
			25606: out = 16'(-4802);
			25607: out = 16'(-6741);
			25608: out = 16'(631);
			25609: out = 16'(2777);
			25610: out = 16'(1076);
			25611: out = 16'(442);
			25612: out = 16'(1948);
			25613: out = 16'(2099);
			25614: out = 16'(-936);
			25615: out = 16'(-3706);
			25616: out = 16'(-3199);
			25617: out = 16'(644);
			25618: out = 16'(1222);
			25619: out = 16'(-382);
			25620: out = 16'(560);
			25621: out = 16'(2844);
			25622: out = 16'(4212);
			25623: out = 16'(1651);
			25624: out = 16'(-2359);
			25625: out = 16'(-6579);
			25626: out = 16'(-2651);
			25627: out = 16'(1729);
			25628: out = 16'(1741);
			25629: out = 16'(392);
			25630: out = 16'(1141);
			25631: out = 16'(3939);
			25632: out = 16'(3898);
			25633: out = 16'(-88);
			25634: out = 16'(-3667);
			25635: out = 16'(-3743);
			25636: out = 16'(-2363);
			25637: out = 16'(-2639);
			25638: out = 16'(-3949);
			25639: out = 16'(-832);
			25640: out = 16'(4682);
			25641: out = 16'(6067);
			25642: out = 16'(1082);
			25643: out = 16'(-3345);
			25644: out = 16'(-3242);
			25645: out = 16'(-535);
			25646: out = 16'(29);
			25647: out = 16'(-9);
			25648: out = 16'(752);
			25649: out = 16'(1288);
			25650: out = 16'(-960);
			25651: out = 16'(-4651);
			25652: out = 16'(-5620);
			25653: out = 16'(-2550);
			25654: out = 16'(239);
			25655: out = 16'(4162);
			25656: out = 16'(3503);
			25657: out = 16'(2147);
			25658: out = 16'(2565);
			25659: out = 16'(4101);
			25660: out = 16'(2036);
			25661: out = 16'(-2495);
			25662: out = 16'(-5825);
			25663: out = 16'(-3463);
			25664: out = 16'(-1532);
			25665: out = 16'(-170);
			25666: out = 16'(396);
			25667: out = 16'(1763);
			25668: out = 16'(3133);
			25669: out = 16'(4077);
			25670: out = 16'(2655);
			25671: out = 16'(-8);
			25672: out = 16'(-3708);
			25673: out = 16'(-2822);
			25674: out = 16'(172);
			25675: out = 16'(1304);
			25676: out = 16'(-1926);
			25677: out = 16'(-1344);
			25678: out = 16'(1295);
			25679: out = 16'(1799);
			25680: out = 16'(-1175);
			25681: out = 16'(-3685);
			25682: out = 16'(-3109);
			25683: out = 16'(227);
			25684: out = 16'(3440);
			25685: out = 16'(2510);
			25686: out = 16'(45);
			25687: out = 16'(-385);
			25688: out = 16'(1409);
			25689: out = 16'(1836);
			25690: out = 16'(-713);
			25691: out = 16'(-2268);
			25692: out = 16'(373);
			25693: out = 16'(1245);
			25694: out = 16'(349);
			25695: out = 16'(-1417);
			25696: out = 16'(-353);
			25697: out = 16'(1036);
			25698: out = 16'(3310);
			25699: out = 16'(2548);
			25700: out = 16'(133);
			25701: out = 16'(-141);
			25702: out = 16'(-2019);
			25703: out = 16'(-1942);
			25704: out = 16'(1694);
			25705: out = 16'(6301);
			25706: out = 16'(4739);
			25707: out = 16'(-825);
			25708: out = 16'(-5146);
			25709: out = 16'(-4929);
			25710: out = 16'(-2347);
			25711: out = 16'(-704);
			25712: out = 16'(533);
			25713: out = 16'(1439);
			25714: out = 16'(325);
			25715: out = 16'(554);
			25716: out = 16'(3435);
			25717: out = 16'(4262);
			25718: out = 16'(-4988);
			25719: out = 16'(-6877);
			25720: out = 16'(-1174);
			25721: out = 16'(4428);
			25722: out = 16'(-114);
			25723: out = 16'(-3124);
			25724: out = 16'(-3426);
			25725: out = 16'(-781);
			25726: out = 16'(8);
			25727: out = 16'(889);
			25728: out = 16'(575);
			25729: out = 16'(-72);
			25730: out = 16'(98);
			25731: out = 16'(-1695);
			25732: out = 16'(-705);
			25733: out = 16'(-2298);
			25734: out = 16'(-4085);
			25735: out = 16'(1644);
			25736: out = 16'(6421);
			25737: out = 16'(3267);
			25738: out = 16'(-4379);
			25739: out = 16'(-5318);
			25740: out = 16'(-1423);
			25741: out = 16'(790);
			25742: out = 16'(826);
			25743: out = 16'(4659);
			25744: out = 16'(4635);
			25745: out = 16'(691);
			25746: out = 16'(-4411);
			25747: out = 16'(-3321);
			25748: out = 16'(-800);
			25749: out = 16'(2089);
			25750: out = 16'(1872);
			25751: out = 16'(714);
			25752: out = 16'(177);
			25753: out = 16'(1442);
			25754: out = 16'(3137);
			25755: out = 16'(3102);
			25756: out = 16'(334);
			25757: out = 16'(-1630);
			25758: out = 16'(494);
			25759: out = 16'(3933);
			25760: out = 16'(1820);
			25761: out = 16'(486);
			25762: out = 16'(-427);
			25763: out = 16'(1531);
			25764: out = 16'(2970);
			25765: out = 16'(-1148);
			25766: out = 16'(-5864);
			25767: out = 16'(-4546);
			25768: out = 16'(2747);
			25769: out = 16'(2017);
			25770: out = 16'(969);
			25771: out = 16'(-477);
			25772: out = 16'(240);
			25773: out = 16'(-406);
			25774: out = 16'(1794);
			25775: out = 16'(914);
			25776: out = 16'(-1170);
			25777: out = 16'(-85);
			25778: out = 16'(-15);
			25779: out = 16'(-1245);
			25780: out = 16'(-2618);
			25781: out = 16'(-629);
			25782: out = 16'(3082);
			25783: out = 16'(4816);
			25784: out = 16'(2720);
			25785: out = 16'(-121);
			25786: out = 16'(-411);
			25787: out = 16'(71);
			25788: out = 16'(-2041);
			25789: out = 16'(-4957);
			25790: out = 16'(-56);
			25791: out = 16'(1889);
			25792: out = 16'(1239);
			25793: out = 16'(-106);
			25794: out = 16'(1989);
			25795: out = 16'(523);
			25796: out = 16'(-1276);
			25797: out = 16'(-1706);
			25798: out = 16'(-229);
			25799: out = 16'(1083);
			25800: out = 16'(527);
			25801: out = 16'(-559);
			25802: out = 16'(-100);
			25803: out = 16'(-362);
			25804: out = 16'(-861);
			25805: out = 16'(-545);
			25806: out = 16'(1734);
			25807: out = 16'(3037);
			25808: out = 16'(1824);
			25809: out = 16'(-1668);
			25810: out = 16'(-3300);
			25811: out = 16'(-510);
			25812: out = 16'(1119);
			25813: out = 16'(573);
			25814: out = 16'(-308);
			25815: out = 16'(-369);
			25816: out = 16'(-41);
			25817: out = 16'(-3650);
			25818: out = 16'(-7119);
			25819: out = 16'(-2470);
			25820: out = 16'(3443);
			25821: out = 16'(8734);
			25822: out = 16'(6117);
			25823: out = 16'(-900);
			25824: out = 16'(-5054);
			25825: out = 16'(-2904);
			25826: out = 16'(-1390);
			25827: out = 16'(-4201);
			25828: out = 16'(-4772);
			25829: out = 16'(-2021);
			25830: out = 16'(2370);
			25831: out = 16'(2961);
			25832: out = 16'(309);
			25833: out = 16'(741);
			25834: out = 16'(2429);
			25835: out = 16'(107);
			25836: out = 16'(-6710);
			25837: out = 16'(-6566);
			25838: out = 16'(-1165);
			25839: out = 16'(3162);
			25840: out = 16'(1932);
			25841: out = 16'(1870);
			25842: out = 16'(1309);
			25843: out = 16'(1887);
			25844: out = 16'(1893);
			25845: out = 16'(118);
			25846: out = 16'(-2857);
			25847: out = 16'(-5235);
			25848: out = 16'(-3769);
			25849: out = 16'(2025);
			25850: out = 16'(4293);
			25851: out = 16'(2674);
			25852: out = 16'(-327);
			25853: out = 16'(-2604);
			25854: out = 16'(-2427);
			25855: out = 16'(-2378);
			25856: out = 16'(332);
			25857: out = 16'(5081);
			25858: out = 16'(4014);
			25859: out = 16'(648);
			25860: out = 16'(-1008);
			25861: out = 16'(-146);
			25862: out = 16'(-2301);
			25863: out = 16'(-6702);
			25864: out = 16'(-8093);
			25865: out = 16'(-3009);
			25866: out = 16'(3324);
			25867: out = 16'(6643);
			25868: out = 16'(6190);
			25869: out = 16'(4242);
			25870: out = 16'(2221);
			25871: out = 16'(1995);
			25872: out = 16'(1282);
			25873: out = 16'(-2342);
			25874: out = 16'(-7909);
			25875: out = 16'(-8881);
			25876: out = 16'(-3795);
			25877: out = 16'(2543);
			25878: out = 16'(5203);
			25879: out = 16'(5620);
			25880: out = 16'(4484);
			25881: out = 16'(1417);
			25882: out = 16'(-2071);
			25883: out = 16'(-134);
			25884: out = 16'(-154);
			25885: out = 16'(-41);
			25886: out = 16'(188);
			25887: out = 16'(1413);
			25888: out = 16'(327);
			25889: out = 16'(-718);
			25890: out = 16'(-780);
			25891: out = 16'(-83);
			25892: out = 16'(-648);
			25893: out = 16'(-2066);
			25894: out = 16'(-1884);
			25895: out = 16'(324);
			25896: out = 16'(702);
			25897: out = 16'(1705);
			25898: out = 16'(2537);
			25899: out = 16'(1157);
			25900: out = 16'(-5203);
			25901: out = 16'(-5909);
			25902: out = 16'(-3089);
			25903: out = 16'(-2145);
			25904: out = 16'(-4336);
			25905: out = 16'(-2461);
			25906: out = 16'(5072);
			25907: out = 16'(9086);
			25908: out = 16'(5121);
			25909: out = 16'(-3305);
			25910: out = 16'(-4006);
			25911: out = 16'(-747);
			25912: out = 16'(-1254);
			25913: out = 16'(-3569);
			25914: out = 16'(-2359);
			25915: out = 16'(357);
			25916: out = 16'(1262);
			25917: out = 16'(3636);
			25918: out = 16'(4098);
			25919: out = 16'(1605);
			25920: out = 16'(-1832);
			25921: out = 16'(191);
			25922: out = 16'(223);
			25923: out = 16'(-1067);
			25924: out = 16'(-2128);
			25925: out = 16'(310);
			25926: out = 16'(2008);
			25927: out = 16'(1595);
			25928: out = 16'(889);
			25929: out = 16'(2465);
			25930: out = 16'(3501);
			25931: out = 16'(208);
			25932: out = 16'(-3719);
			25933: out = 16'(-2340);
			25934: out = 16'(2752);
			25935: out = 16'(3436);
			25936: out = 16'(187);
			25937: out = 16'(-1490);
			25938: out = 16'(-356);
			25939: out = 16'(865);
			25940: out = 16'(-1991);
			25941: out = 16'(-5336);
			25942: out = 16'(-2927);
			25943: out = 16'(934);
			25944: out = 16'(3996);
			25945: out = 16'(3707);
			25946: out = 16'(2110);
			25947: out = 16'(-2721);
			25948: out = 16'(-1922);
			25949: out = 16'(437);
			25950: out = 16'(-518);
			25951: out = 16'(-2665);
			25952: out = 16'(-2578);
			25953: out = 16'(2495);
			25954: out = 16'(6692);
			25955: out = 16'(3730);
			25956: out = 16'(93);
			25957: out = 16'(-979);
			25958: out = 16'(-413);
			25959: out = 16'(-3601);
			25960: out = 16'(-6023);
			25961: out = 16'(-5378);
			25962: out = 16'(-535);
			25963: out = 16'(1976);
			25964: out = 16'(4096);
			25965: out = 16'(856);
			25966: out = 16'(-519);
			25967: out = 16'(1832);
			25968: out = 16'(4047);
			25969: out = 16'(2106);
			25970: out = 16'(-389);
			25971: out = 16'(-1252);
			25972: out = 16'(-3223);
			25973: out = 16'(-4231);
			25974: out = 16'(-2064);
			25975: out = 16'(2576);
			25976: out = 16'(3294);
			25977: out = 16'(3852);
			25978: out = 16'(2782);
			25979: out = 16'(1373);
			25980: out = 16'(-2123);
			25981: out = 16'(-2411);
			25982: out = 16'(-1753);
			25983: out = 16'(1895);
			25984: out = 16'(5096);
			25985: out = 16'(2835);
			25986: out = 16'(-2504);
			25987: out = 16'(-6608);
			25988: out = 16'(-7398);
			25989: out = 16'(-2820);
			25990: out = 16'(567);
			25991: out = 16'(4738);
			25992: out = 16'(6274);
			25993: out = 16'(3910);
			25994: out = 16'(-948);
			25995: out = 16'(260);
			25996: out = 16'(3731);
			25997: out = 16'(1659);
			25998: out = 16'(-2998);
			25999: out = 16'(-4649);
			26000: out = 16'(-2407);
			26001: out = 16'(-84);
			26002: out = 16'(-119);
			26003: out = 16'(-437);
			26004: out = 16'(-1449);
			26005: out = 16'(-155);
			26006: out = 16'(2474);
			26007: out = 16'(6694);
			26008: out = 16'(1972);
			26009: out = 16'(-7328);
			26010: out = 16'(-10588);
			26011: out = 16'(-543);
			26012: out = 16'(4439);
			26013: out = 16'(1102);
			26014: out = 16'(387);
			26015: out = 16'(3208);
			26016: out = 16'(2258);
			26017: out = 16'(-2512);
			26018: out = 16'(-2843);
			26019: out = 16'(1012);
			26020: out = 16'(1231);
			26021: out = 16'(-2566);
			26022: out = 16'(-2247);
			26023: out = 16'(4098);
			26024: out = 16'(6618);
			26025: out = 16'(1581);
			26026: out = 16'(-4630);
			26027: out = 16'(-2760);
			26028: out = 16'(-803);
			26029: out = 16'(-954);
			26030: out = 16'(-2576);
			26031: out = 16'(111);
			26032: out = 16'(-4061);
			26033: out = 16'(-3138);
			26034: out = 16'(2406);
			26035: out = 16'(6218);
			26036: out = 16'(-2252);
			26037: out = 16'(-8000);
			26038: out = 16'(-3734);
			26039: out = 16'(5255);
			26040: out = 16'(2356);
			26041: out = 16'(37);
			26042: out = 16'(1636);
			26043: out = 16'(3898);
			26044: out = 16'(-226);
			26045: out = 16'(-5444);
			26046: out = 16'(-4277);
			26047: out = 16'(1543);
			26048: out = 16'(-115);
			26049: out = 16'(256);
			26050: out = 16'(773);
			26051: out = 16'(1292);
			26052: out = 16'(-1769);
			26053: out = 16'(-141);
			26054: out = 16'(282);
			26055: out = 16'(-227);
			26056: out = 16'(-478);
			26057: out = 16'(1642);
			26058: out = 16'(4830);
			26059: out = 16'(3739);
			26060: out = 16'(-1777);
			26061: out = 16'(-4659);
			26062: out = 16'(-2722);
			26063: out = 16'(647);
			26064: out = 16'(1384);
			26065: out = 16'(163);
			26066: out = 16'(125);
			26067: out = 16'(-672);
			26068: out = 16'(-1763);
			26069: out = 16'(-1501);
			26070: out = 16'(2718);
			26071: out = 16'(3188);
			26072: out = 16'(38);
			26073: out = 16'(-3238);
			26074: out = 16'(-1984);
			26075: out = 16'(-209);
			26076: out = 16'(2029);
			26077: out = 16'(3662);
			26078: out = 16'(3835);
			26079: out = 16'(1103);
			26080: out = 16'(-252);
			26081: out = 16'(-225);
			26082: out = 16'(-770);
			26083: out = 16'(-3650);
			26084: out = 16'(-2070);
			26085: out = 16'(2662);
			26086: out = 16'(3980);
			26087: out = 16'(2821);
			26088: out = 16'(909);
			26089: out = 16'(-1014);
			26090: out = 16'(-3318);
			26091: out = 16'(-879);
			26092: out = 16'(1703);
			26093: out = 16'(802);
			26094: out = 16'(-2604);
			26095: out = 16'(-1453);
			26096: out = 16'(2221);
			26097: out = 16'(2641);
			26098: out = 16'(-912);
			26099: out = 16'(-4854);
			26100: out = 16'(-1958);
			26101: out = 16'(450);
			26102: out = 16'(-176);
			26103: out = 16'(82);
			26104: out = 16'(2791);
			26105: out = 16'(2851);
			26106: out = 16'(1028);
			26107: out = 16'(1409);
			26108: out = 16'(244);
			26109: out = 16'(-2946);
			26110: out = 16'(-5011);
			26111: out = 16'(-1120);
			26112: out = 16'(-747);
			26113: out = 16'(1629);
			26114: out = 16'(2314);
			26115: out = 16'(1856);
			26116: out = 16'(-1534);
			26117: out = 16'(-1985);
			26118: out = 16'(-869);
			26119: out = 16'(972);
			26120: out = 16'(1364);
			26121: out = 16'(891);
			26122: out = 16'(971);
			26123: out = 16'(3056);
			26124: out = 16'(4282);
			26125: out = 16'(-706);
			26126: out = 16'(-6865);
			26127: out = 16'(-7559);
			26128: out = 16'(-2290);
			26129: out = 16'(-1039);
			26130: out = 16'(-1392);
			26131: out = 16'(-963);
			26132: out = 16'(920);
			26133: out = 16'(1642);
			26134: out = 16'(1416);
			26135: out = 16'(2529);
			26136: out = 16'(3057);
			26137: out = 16'(-653);
			26138: out = 16'(-6117);
			26139: out = 16'(-6171);
			26140: out = 16'(-764);
			26141: out = 16'(1271);
			26142: out = 16'(2676);
			26143: out = 16'(691);
			26144: out = 16'(-1455);
			26145: out = 16'(-2079);
			26146: out = 16'(2685);
			26147: out = 16'(4710);
			26148: out = 16'(2817);
			26149: out = 16'(-184);
			26150: out = 16'(490);
			26151: out = 16'(2789);
			26152: out = 16'(2545);
			26153: out = 16'(-1067);
			26154: out = 16'(-4724);
			26155: out = 16'(-3117);
			26156: out = 16'(-60);
			26157: out = 16'(375);
			26158: out = 16'(-2305);
			26159: out = 16'(-529);
			26160: out = 16'(1363);
			26161: out = 16'(3191);
			26162: out = 16'(5454);
			26163: out = 16'(2878);
			26164: out = 16'(-935);
			26165: out = 16'(-4504);
			26166: out = 16'(-5271);
			26167: out = 16'(-2899);
			26168: out = 16'(-502);
			26169: out = 16'(686);
			26170: out = 16'(1974);
			26171: out = 16'(3288);
			26172: out = 16'(3801);
			26173: out = 16'(2032);
			26174: out = 16'(-773);
			26175: out = 16'(-3861);
			26176: out = 16'(-756);
			26177: out = 16'(1577);
			26178: out = 16'(577);
			26179: out = 16'(-2156);
			26180: out = 16'(1033);
			26181: out = 16'(4018);
			26182: out = 16'(3569);
			26183: out = 16'(-312);
			26184: out = 16'(1223);
			26185: out = 16'(863);
			26186: out = 16'(334);
			26187: out = 16'(-388);
			26188: out = 16'(-736);
			26189: out = 16'(-5360);
			26190: out = 16'(-6559);
			26191: out = 16'(-549);
			26192: out = 16'(2560);
			26193: out = 16'(5741);
			26194: out = 16'(2158);
			26195: out = 16'(-1317);
			26196: out = 16'(-1976);
			26197: out = 16'(1178);
			26198: out = 16'(-1045);
			26199: out = 16'(-3031);
			26200: out = 16'(-983);
			26201: out = 16'(-426);
			26202: out = 16'(-4442);
			26203: out = 16'(-4023);
			26204: out = 16'(4538);
			26205: out = 16'(5652);
			26206: out = 16'(1029);
			26207: out = 16'(-2914);
			26208: out = 16'(1433);
			26209: out = 16'(4277);
			26210: out = 16'(4027);
			26211: out = 16'(-2179);
			26212: out = 16'(-6799);
			26213: out = 16'(-6447);
			26214: out = 16'(185);
			26215: out = 16'(3068);
			26216: out = 16'(950);
			26217: out = 16'(-2057);
			26218: out = 16'(-834);
			26219: out = 16'(2246);
			26220: out = 16'(3354);
			26221: out = 16'(1786);
			26222: out = 16'(-1866);
			26223: out = 16'(-1848);
			26224: out = 16'(-223);
			26225: out = 16'(-489);
			26226: out = 16'(-5000);
			26227: out = 16'(-3403);
			26228: out = 16'(437);
			26229: out = 16'(1059);
			26230: out = 16'(-1042);
			26231: out = 16'(641);
			26232: out = 16'(5742);
			26233: out = 16'(7168);
			26234: out = 16'(1191);
			26235: out = 16'(-2426);
			26236: out = 16'(-3514);
			26237: out = 16'(-3510);
			26238: out = 16'(-4870);
			26239: out = 16'(-4911);
			26240: out = 16'(-1248);
			26241: out = 16'(3582);
			26242: out = 16'(5202);
			26243: out = 16'(4520);
			26244: out = 16'(1357);
			26245: out = 16'(-475);
			26246: out = 16'(77);
			26247: out = 16'(-273);
			26248: out = 16'(-222);
			26249: out = 16'(-3222);
			26250: out = 16'(-5139);
			26251: out = 16'(-736);
			26252: out = 16'(1252);
			26253: out = 16'(582);
			26254: out = 16'(-632);
			26255: out = 16'(1880);
			26256: out = 16'(1379);
			26257: out = 16'(874);
			26258: out = 16'(-919);
			26259: out = 16'(-1135);
			26260: out = 16'(2816);
			26261: out = 16'(3265);
			26262: out = 16'(-375);
			26263: out = 16'(-4343);
			26264: out = 16'(-4101);
			26265: out = 16'(-1258);
			26266: out = 16'(378);
			26267: out = 16'(457);
			26268: out = 16'(3763);
			26269: out = 16'(4349);
			26270: out = 16'(4515);
			26271: out = 16'(2032);
			26272: out = 16'(-771);
			26273: out = 16'(-719);
			26274: out = 16'(1558);
			26275: out = 16'(303);
			26276: out = 16'(-4211);
			26277: out = 16'(-2254);
			26278: out = 16'(2465);
			26279: out = 16'(5232);
			26280: out = 16'(3922);
			26281: out = 16'(64);
			26282: out = 16'(-272);
			26283: out = 16'(-1393);
			26284: out = 16'(-4218);
			26285: out = 16'(-6448);
			26286: out = 16'(-1831);
			26287: out = 16'(1624);
			26288: out = 16'(1735);
			26289: out = 16'(573);
			26290: out = 16'(1214);
			26291: out = 16'(1702);
			26292: out = 16'(2183);
			26293: out = 16'(1497);
			26294: out = 16'(-959);
			26295: out = 16'(-5331);
			26296: out = 16'(-5173);
			26297: out = 16'(-454);
			26298: out = 16'(-267);
			26299: out = 16'(-2177);
			26300: out = 16'(-2957);
			26301: out = 16'(-1034);
			26302: out = 16'(613);
			26303: out = 16'(186);
			26304: out = 16'(2191);
			26305: out = 16'(5157);
			26306: out = 16'(2899);
			26307: out = 16'(-3476);
			26308: out = 16'(-6456);
			26309: out = 16'(-2718);
			26310: out = 16'(188);
			26311: out = 16'(-1950);
			26312: out = 16'(-4423);
			26313: out = 16'(-1345);
			26314: out = 16'(2180);
			26315: out = 16'(997);
			26316: out = 16'(-3125);
			26317: out = 16'(-362);
			26318: out = 16'(6372);
			26319: out = 16'(5280);
			26320: out = 16'(1537);
			26321: out = 16'(-280);
			26322: out = 16'(493);
			26323: out = 16'(-2525);
			26324: out = 16'(-1143);
			26325: out = 16'(842);
			26326: out = 16'(2269);
			26327: out = 16'(565);
			26328: out = 16'(3197);
			26329: out = 16'(2669);
			26330: out = 16'(-535);
			26331: out = 16'(-3550);
			26332: out = 16'(3250);
			26333: out = 16'(4449);
			26334: out = 16'(12);
			26335: out = 16'(-4818);
			26336: out = 16'(254);
			26337: out = 16'(2947);
			26338: out = 16'(1721);
			26339: out = 16'(-1441);
			26340: out = 16'(83);
			26341: out = 16'(2388);
			26342: out = 16'(3870);
			26343: out = 16'(1813);
			26344: out = 16'(-2821);
			26345: out = 16'(-3858);
			26346: out = 16'(-4853);
			26347: out = 16'(-3881);
			26348: out = 16'(-296);
			26349: out = 16'(3034);
			26350: out = 16'(2978);
			26351: out = 16'(1115);
			26352: out = 16'(-435);
			26353: out = 16'(-1576);
			26354: out = 16'(208);
			26355: out = 16'(3007);
			26356: out = 16'(3179);
			26357: out = 16'(-757);
			26358: out = 16'(-3197);
			26359: out = 16'(-1114);
			26360: out = 16'(1558);
			26361: out = 16'(-327);
			26362: out = 16'(-2607);
			26363: out = 16'(-1961);
			26364: out = 16'(1546);
			26365: out = 16'(3024);
			26366: out = 16'(-136);
			26367: out = 16'(-2292);
			26368: out = 16'(-1596);
			26369: out = 16'(330);
			26370: out = 16'(1984);
			26371: out = 16'(856);
			26372: out = 16'(-668);
			26373: out = 16'(-635);
			26374: out = 16'(-231);
			26375: out = 16'(1365);
			26376: out = 16'(-293);
			26377: out = 16'(-2728);
			26378: out = 16'(-1452);
			26379: out = 16'(-396);
			26380: out = 16'(203);
			26381: out = 16'(-456);
			26382: out = 16'(-748);
			26383: out = 16'(283);
			26384: out = 16'(1688);
			26385: out = 16'(2062);
			26386: out = 16'(1155);
			26387: out = 16'(246);
			26388: out = 16'(-818);
			26389: out = 16'(-295);
			26390: out = 16'(694);
			26391: out = 16'(30);
			26392: out = 16'(-2343);
			26393: out = 16'(-2645);
			26394: out = 16'(-186);
			26395: out = 16'(-281);
			26396: out = 16'(458);
			26397: out = 16'(-1427);
			26398: out = 16'(-1603);
			26399: out = 16'(1968);
			26400: out = 16'(7605);
			26401: out = 16'(7443);
			26402: out = 16'(1886);
			26403: out = 16'(-4595);
			26404: out = 16'(-5006);
			26405: out = 16'(-3616);
			26406: out = 16'(-1299);
			26407: out = 16'(-17);
			26408: out = 16'(-787);
			26409: out = 16'(-1530);
			26410: out = 16'(-999);
			26411: out = 16'(597);
			26412: out = 16'(2090);
			26413: out = 16'(3170);
			26414: out = 16'(2718);
			26415: out = 16'(-229);
			26416: out = 16'(-4778);
			26417: out = 16'(-1123);
			26418: out = 16'(695);
			26419: out = 16'(-1664);
			26420: out = 16'(-4269);
			26421: out = 16'(885);
			26422: out = 16'(5102);
			26423: out = 16'(2221);
			26424: out = 16'(-4572);
			26425: out = 16'(-4095);
			26426: out = 16'(266);
			26427: out = 16'(2010);
			26428: out = 16'(-503);
			26429: out = 16'(359);
			26430: out = 16'(-784);
			26431: out = 16'(-530);
			26432: out = 16'(1131);
			26433: out = 16'(5182);
			26434: out = 16'(-92);
			26435: out = 16'(-4139);
			26436: out = 16'(-3152);
			26437: out = 16'(2376);
			26438: out = 16'(352);
			26439: out = 16'(-295);
			26440: out = 16'(1089);
			26441: out = 16'(3499);
			26442: out = 16'(1574);
			26443: out = 16'(-252);
			26444: out = 16'(-662);
			26445: out = 16'(928);
			26446: out = 16'(1947);
			26447: out = 16'(1501);
			26448: out = 16'(2048);
			26449: out = 16'(3564);
			26450: out = 16'(2943);
			26451: out = 16'(651);
			26452: out = 16'(-2225);
			26453: out = 16'(-3702);
			26454: out = 16'(-3338);
			26455: out = 16'(-2846);
			26456: out = 16'(-1145);
			26457: out = 16'(728);
			26458: out = 16'(2339);
			26459: out = 16'(4785);
			26460: out = 16'(4274);
			26461: out = 16'(853);
			26462: out = 16'(-3290);
			26463: out = 16'(-4155);
			26464: out = 16'(-3283);
			26465: out = 16'(-1777);
			26466: out = 16'(-780);
			26467: out = 16'(-35);
			26468: out = 16'(343);
			26469: out = 16'(1238);
			26470: out = 16'(2534);
			26471: out = 16'(3160);
			26472: out = 16'(3465);
			26473: out = 16'(169);
			26474: out = 16'(-5063);
			26475: out = 16'(-9078);
			26476: out = 16'(-3299);
			26477: out = 16'(252);
			26478: out = 16'(2476);
			26479: out = 16'(3426);
			26480: out = 16'(3519);
			26481: out = 16'(265);
			26482: out = 16'(-1112);
			26483: out = 16'(293);
			26484: out = 16'(195);
			26485: out = 16'(-443);
			26486: out = 16'(-2046);
			26487: out = 16'(-2061);
			26488: out = 16'(96);
			26489: out = 16'(1617);
			26490: out = 16'(2366);
			26491: out = 16'(578);
			26492: out = 16'(-3669);
			26493: out = 16'(-4786);
			26494: out = 16'(-1540);
			26495: out = 16'(3670);
			26496: out = 16'(4352);
			26497: out = 16'(-117);
			26498: out = 16'(-1327);
			26499: out = 16'(2675);
			26500: out = 16'(4030);
			26501: out = 16'(-1230);
			26502: out = 16'(-8784);
			26503: out = 16'(-6159);
			26504: out = 16'(2782);
			26505: out = 16'(4129);
			26506: out = 16'(2506);
			26507: out = 16'(125);
			26508: out = 16'(243);
			26509: out = 16'(388);
			26510: out = 16'(-2722);
			26511: out = 16'(-1817);
			26512: out = 16'(1026);
			26513: out = 16'(1132);
			26514: out = 16'(2327);
			26515: out = 16'(390);
			26516: out = 16'(-673);
			26517: out = 16'(-546);
			26518: out = 16'(4002);
			26519: out = 16'(402);
			26520: out = 16'(-2249);
			26521: out = 16'(-1836);
			26522: out = 16'(2028);
			26523: out = 16'(302);
			26524: out = 16'(-1326);
			26525: out = 16'(-3348);
			26526: out = 16'(-3590);
			26527: out = 16'(43);
			26528: out = 16'(5494);
			26529: out = 16'(5163);
			26530: out = 16'(-804);
			26531: out = 16'(-2343);
			26532: out = 16'(-1709);
			26533: out = 16'(-1419);
			26534: out = 16'(-2513);
			26535: out = 16'(-1056);
			26536: out = 16'(2747);
			26537: out = 16'(2935);
			26538: out = 16'(-1628);
			26539: out = 16'(-5129);
			26540: out = 16'(-770);
			26541: out = 16'(3756);
			26542: out = 16'(2822);
			26543: out = 16'(-67);
			26544: out = 16'(-1261);
			26545: out = 16'(257);
			26546: out = 16'(-431);
			26547: out = 16'(-3484);
			26548: out = 16'(-4862);
			26549: out = 16'(-726);
			26550: out = 16'(4152);
			26551: out = 16'(4341);
			26552: out = 16'(-1778);
			26553: out = 16'(-3073);
			26554: out = 16'(-675);
			26555: out = 16'(1874);
			26556: out = 16'(3372);
			26557: out = 16'(753);
			26558: out = 16'(-460);
			26559: out = 16'(425);
			26560: out = 16'(1839);
			26561: out = 16'(-1597);
			26562: out = 16'(-3439);
			26563: out = 16'(-2757);
			26564: out = 16'(-1650);
			26565: out = 16'(-218);
			26566: out = 16'(656);
			26567: out = 16'(2940);
			26568: out = 16'(5512);
			26569: out = 16'(6861);
			26570: out = 16'(853);
			26571: out = 16'(-6035);
			26572: out = 16'(-7383);
			26573: out = 16'(-412);
			26574: out = 16'(330);
			26575: out = 16'(-388);
			26576: out = 16'(717);
			26577: out = 16'(3258);
			26578: out = 16'(3675);
			26579: out = 16'(594);
			26580: out = 16'(-2198);
			26581: out = 16'(-854);
			26582: out = 16'(-3260);
			26583: out = 16'(-2063);
			26584: out = 16'(206);
			26585: out = 16'(2102);
			26586: out = 16'(32);
			26587: out = 16'(787);
			26588: out = 16'(1803);
			26589: out = 16'(1496);
			26590: out = 16'(-2369);
			26591: out = 16'(-958);
			26592: out = 16'(330);
			26593: out = 16'(-1079);
			26594: out = 16'(-4686);
			26595: out = 16'(-2162);
			26596: out = 16'(1732);
			26597: out = 16'(3697);
			26598: out = 16'(3250);
			26599: out = 16'(1674);
			26600: out = 16'(-383);
			26601: out = 16'(-3310);
			26602: out = 16'(-5544);
			26603: out = 16'(-2177);
			26604: out = 16'(-242);
			26605: out = 16'(37);
			26606: out = 16'(681);
			26607: out = 16'(3786);
			26608: out = 16'(3237);
			26609: out = 16'(-745);
			26610: out = 16'(-3926);
			26611: out = 16'(-800);
			26612: out = 16'(0);
			26613: out = 16'(-311);
			26614: out = 16'(-407);
			26615: out = 16'(1731);
			26616: out = 16'(3679);
			26617: out = 16'(3366);
			26618: out = 16'(644);
			26619: out = 16'(-2653);
			26620: out = 16'(-3079);
			26621: out = 16'(-2963);
			26622: out = 16'(-701);
			26623: out = 16'(2283);
			26624: out = 16'(177);
			26625: out = 16'(-100);
			26626: out = 16'(933);
			26627: out = 16'(2027);
			26628: out = 16'(-4);
			26629: out = 16'(-162);
			26630: out = 16'(-136);
			26631: out = 16'(-636);
			26632: out = 16'(-2306);
			26633: out = 16'(-730);
			26634: out = 16'(3010);
			26635: out = 16'(5287);
			26636: out = 16'(2714);
			26637: out = 16'(-1452);
			26638: out = 16'(-2859);
			26639: out = 16'(-149);
			26640: out = 16'(1847);
			26641: out = 16'(2294);
			26642: out = 16'(-2071);
			26643: out = 16'(-4794);
			26644: out = 16'(-3110);
			26645: out = 16'(1753);
			26646: out = 16'(322);
			26647: out = 16'(-1800);
			26648: out = 16'(-843);
			26649: out = 16'(1251);
			26650: out = 16'(3308);
			26651: out = 16'(1866);
			26652: out = 16'(-1241);
			26653: out = 16'(-3857);
			26654: out = 16'(-795);
			26655: out = 16'(1633);
			26656: out = 16'(919);
			26657: out = 16'(-3419);
			26658: out = 16'(1304);
			26659: out = 16'(499);
			26660: out = 16'(-652);
			26661: out = 16'(-1551);
			26662: out = 16'(2310);
			26663: out = 16'(1255);
			26664: out = 16'(2827);
			26665: out = 16'(3227);
			26666: out = 16'(345);
			26667: out = 16'(-6196);
			26668: out = 16'(-4469);
			26669: out = 16'(1570);
			26670: out = 16'(3894);
			26671: out = 16'(-2042);
			26672: out = 16'(-920);
			26673: out = 16'(2707);
			26674: out = 16'(678);
			26675: out = 16'(-4579);
			26676: out = 16'(-3035);
			26677: out = 16'(2235);
			26678: out = 16'(3725);
			26679: out = 16'(1699);
			26680: out = 16'(1734);
			26681: out = 16'(681);
			26682: out = 16'(-3769);
			26683: out = 16'(-7720);
			26684: out = 16'(-2901);
			26685: out = 16'(3536);
			26686: out = 16'(4616);
			26687: out = 16'(1414);
			26688: out = 16'(-1105);
			26689: out = 16'(-3118);
			26690: out = 16'(-4003);
			26691: out = 16'(-2027);
			26692: out = 16'(1371);
			26693: out = 16'(1559);
			26694: out = 16'(-1482);
			26695: out = 16'(-2357);
			26696: out = 16'(3067);
			26697: out = 16'(5866);
			26698: out = 16'(1545);
			26699: out = 16'(-5644);
			26700: out = 16'(-4660);
			26701: out = 16'(-2762);
			26702: out = 16'(-400);
			26703: out = 16'(118);
			26704: out = 16'(266);
			26705: out = 16'(26);
			26706: out = 16'(1209);
			26707: out = 16'(2533);
			26708: out = 16'(1995);
			26709: out = 16'(1042);
			26710: out = 16'(308);
			26711: out = 16'(744);
			26712: out = 16'(-428);
			26713: out = 16'(398);
			26714: out = 16'(-4072);
			26715: out = 16'(-3983);
			26716: out = 16'(1680);
			26717: out = 16'(3828);
			26718: out = 16'(545);
			26719: out = 16'(-3402);
			26720: out = 16'(-3181);
			26721: out = 16'(-58);
			26722: out = 16'(355);
			26723: out = 16'(-67);
			26724: out = 16'(1239);
			26725: out = 16'(5419);
			26726: out = 16'(862);
			26727: out = 16'(-707);
			26728: out = 16'(-1180);
			26729: out = 16'(-1519);
			26730: out = 16'(-529);
			26731: out = 16'(720);
			26732: out = 16'(-787);
			26733: out = 16'(-2942);
			26734: out = 16'(-454);
			26735: out = 16'(6259);
			26736: out = 16'(8590);
			26737: out = 16'(3017);
			26738: out = 16'(-9537);
			26739: out = 16'(-5920);
			26740: out = 16'(-49);
			26741: out = 16'(1075);
			26742: out = 16'(-674);
			26743: out = 16'(945);
			26744: out = 16'(1187);
			26745: out = 16'(-1500);
			26746: out = 16'(-4518);
			26747: out = 16'(-63);
			26748: out = 16'(2923);
			26749: out = 16'(2851);
			26750: out = 16'(246);
			26751: out = 16'(-1956);
			26752: out = 16'(-1780);
			26753: out = 16'(761);
			26754: out = 16'(2044);
			26755: out = 16'(1029);
			26756: out = 16'(-57);
			26757: out = 16'(902);
			26758: out = 16'(1200);
			26759: out = 16'(895);
			26760: out = 16'(-5339);
			26761: out = 16'(-4039);
			26762: out = 16'(278);
			26763: out = 16'(-79);
			26764: out = 16'(314);
			26765: out = 16'(2017);
			26766: out = 16'(4096);
			26767: out = 16'(2922);
			26768: out = 16'(512);
			26769: out = 16'(-342);
			26770: out = 16'(-722);
			26771: out = 16'(-2898);
			26772: out = 16'(-2001);
			26773: out = 16'(-3361);
			26774: out = 16'(-998);
			26775: out = 16'(2330);
			26776: out = 16'(3438);
			26777: out = 16'(2604);
			26778: out = 16'(1021);
			26779: out = 16'(-260);
			26780: out = 16'(-147);
			26781: out = 16'(-2870);
			26782: out = 16'(-2896);
			26783: out = 16'(-1647);
			26784: out = 16'(559);
			26785: out = 16'(1720);
			26786: out = 16'(4605);
			26787: out = 16'(4174);
			26788: out = 16'(385);
			26789: out = 16'(-4478);
			26790: out = 16'(-3465);
			26791: out = 16'(-1047);
			26792: out = 16'(257);
			26793: out = 16'(-67);
			26794: out = 16'(-296);
			26795: out = 16'(-2214);
			26796: out = 16'(-2406);
			26797: out = 16'(374);
			26798: out = 16'(6301);
			26799: out = 16'(4192);
			26800: out = 16'(-1903);
			26801: out = 16'(-5139);
			26802: out = 16'(-192);
			26803: out = 16'(1983);
			26804: out = 16'(2840);
			26805: out = 16'(4044);
			26806: out = 16'(1522);
			26807: out = 16'(326);
			26808: out = 16'(-62);
			26809: out = 16'(-630);
			26810: out = 16'(-3867);
			26811: out = 16'(-6089);
			26812: out = 16'(-4143);
			26813: out = 16'(585);
			26814: out = 16'(2095);
			26815: out = 16'(3533);
			26816: out = 16'(3889);
			26817: out = 16'(3466);
			26818: out = 16'(128);
			26819: out = 16'(135);
			26820: out = 16'(-912);
			26821: out = 16'(-1003);
			26822: out = 16'(-1803);
			26823: out = 16'(715);
			26824: out = 16'(714);
			26825: out = 16'(3519);
			26826: out = 16'(5050);
			26827: out = 16'(284);
			26828: out = 16'(-5309);
			26829: out = 16'(-4035);
			26830: out = 16'(1961);
			26831: out = 16'(1445);
			26832: out = 16'(1427);
			26833: out = 16'(-698);
			26834: out = 16'(-200);
			26835: out = 16'(1964);
			26836: out = 16'(3086);
			26837: out = 16'(1295);
			26838: out = 16'(-1658);
			26839: out = 16'(-3192);
			26840: out = 16'(-2045);
			26841: out = 16'(-1105);
			26842: out = 16'(-875);
			26843: out = 16'(214);
			26844: out = 16'(1576);
			26845: out = 16'(934);
			26846: out = 16'(-1741);
			26847: out = 16'(-1018);
			26848: out = 16'(4482);
			26849: out = 16'(5652);
			26850: out = 16'(-163);
			26851: out = 16'(-5420);
			26852: out = 16'(-2821);
			26853: out = 16'(2669);
			26854: out = 16'(1718);
			26855: out = 16'(-2332);
			26856: out = 16'(-1969);
			26857: out = 16'(-231);
			26858: out = 16'(-401);
			26859: out = 16'(-2813);
			26860: out = 16'(-2602);
			26861: out = 16'(-670);
			26862: out = 16'(3681);
			26863: out = 16'(5401);
			26864: out = 16'(3836);
			26865: out = 16'(-1662);
			26866: out = 16'(-1455);
			26867: out = 16'(-496);
			26868: out = 16'(-305);
			26869: out = 16'(-1076);
			26870: out = 16'(-2331);
			26871: out = 16'(-1046);
			26872: out = 16'(1258);
			26873: out = 16'(802);
			26874: out = 16'(-373);
			26875: out = 16'(-2449);
			26876: out = 16'(-1154);
			26877: out = 16'(1284);
			26878: out = 16'(1471);
			26879: out = 16'(-2442);
			26880: out = 16'(-3151);
			26881: out = 16'(1019);
			26882: out = 16'(2711);
			26883: out = 16'(1271);
			26884: out = 16'(-2127);
			26885: out = 16'(-2619);
			26886: out = 16'(-178);
			26887: out = 16'(1226);
			26888: out = 16'(528);
			26889: out = 16'(-550);
			26890: out = 16'(-904);
			26891: out = 16'(-135);
			26892: out = 16'(1004);
			26893: out = 16'(2894);
			26894: out = 16'(3479);
			26895: out = 16'(1675);
			26896: out = 16'(-1505);
			26897: out = 16'(-2226);
			26898: out = 16'(-835);
			26899: out = 16'(-295);
			26900: out = 16'(-3532);
			26901: out = 16'(-4089);
			26902: out = 16'(-14);
			26903: out = 16'(3581);
			26904: out = 16'(5185);
			26905: out = 16'(2110);
			26906: out = 16'(-2588);
			26907: out = 16'(-4532);
			26908: out = 16'(-3865);
			26909: out = 16'(-639);
			26910: out = 16'(789);
			26911: out = 16'(602);
			26912: out = 16'(287);
			26913: out = 16'(3505);
			26914: out = 16'(5347);
			26915: out = 16'(4279);
			26916: out = 16'(-94);
			26917: out = 16'(-165);
			26918: out = 16'(-1835);
			26919: out = 16'(-4728);
			26920: out = 16'(-6337);
			26921: out = 16'(-1004);
			26922: out = 16'(853);
			26923: out = 16'(-683);
			26924: out = 16'(-594);
			26925: out = 16'(4020);
			26926: out = 16'(3318);
			26927: out = 16'(-1785);
			26928: out = 16'(-5261);
			26929: out = 16'(-3073);
			26930: out = 16'(-159);
			26931: out = 16'(676);
			26932: out = 16'(161);
			26933: out = 16'(3278);
			26934: out = 16'(2393);
			26935: out = 16'(1293);
			26936: out = 16'(-1123);
			26937: out = 16'(-4253);
			26938: out = 16'(-7751);
			26939: out = 16'(-4419);
			26940: out = 16'(1923);
			26941: out = 16'(5066);
			26942: out = 16'(1022);
			26943: out = 16'(1472);
			26944: out = 16'(3623);
			26945: out = 16'(1166);
			26946: out = 16'(-6319);
			26947: out = 16'(-6778);
			26948: out = 16'(86);
			26949: out = 16'(4828);
			26950: out = 16'(-68);
			26951: out = 16'(-1363);
			26952: out = 16'(1082);
			26953: out = 16'(3336);
			26954: out = 16'(1417);
			26955: out = 16'(-236);
			26956: out = 16'(-1166);
			26957: out = 16'(-453);
			26958: out = 16'(546);
			26959: out = 16'(-2097);
			26960: out = 16'(-3064);
			26961: out = 16'(624);
			26962: out = 16'(4970);
			26963: out = 16'(6154);
			26964: out = 16'(-376);
			26965: out = 16'(-6277);
			26966: out = 16'(-5444);
			26967: out = 16'(-685);
			26968: out = 16'(-389);
			26969: out = 16'(-1778);
			26970: out = 16'(139);
			26971: out = 16'(1717);
			26972: out = 16'(3968);
			26973: out = 16'(2920);
			26974: out = 16'(602);
			26975: out = 16'(-3075);
			26976: out = 16'(954);
			26977: out = 16'(2495);
			26978: out = 16'(1279);
			26979: out = 16'(-908);
			26980: out = 16'(488);
			26981: out = 16'(-54);
			26982: out = 16'(-1333);
			26983: out = 16'(-1553);
			26984: out = 16'(-1637);
			26985: out = 16'(209);
			26986: out = 16'(2524);
			26987: out = 16'(2875);
			26988: out = 16'(382);
			26989: out = 16'(-500);
			26990: out = 16'(1621);
			26991: out = 16'(2816);
			26992: out = 16'(2);
			26993: out = 16'(-3832);
			26994: out = 16'(-4296);
			26995: out = 16'(-2843);
			26996: out = 16'(-3069);
			26997: out = 16'(-3751);
			26998: out = 16'(-1007);
			26999: out = 16'(3204);
			27000: out = 16'(5001);
			27001: out = 16'(2525);
			27002: out = 16'(672);
			27003: out = 16'(-933);
			27004: out = 16'(-1310);
			27005: out = 16'(-332);
			27006: out = 16'(1869);
			27007: out = 16'(67);
			27008: out = 16'(-3151);
			27009: out = 16'(-786);
			27010: out = 16'(2981);
			27011: out = 16'(2640);
			27012: out = 16'(-1055);
			27013: out = 16'(-1937);
			27014: out = 16'(1005);
			27015: out = 16'(2604);
			27016: out = 16'(1349);
			27017: out = 16'(745);
			27018: out = 16'(-76);
			27019: out = 16'(-503);
			27020: out = 16'(-754);
			27021: out = 16'(903);
			27022: out = 16'(1687);
			27023: out = 16'(21);
			27024: out = 16'(-3552);
			27025: out = 16'(-3934);
			27026: out = 16'(-464);
			27027: out = 16'(652);
			27028: out = 16'(-2061);
			27029: out = 16'(-3175);
			27030: out = 16'(-97);
			27031: out = 16'(33);
			27032: out = 16'(-4332);
			27033: out = 16'(-5419);
			27034: out = 16'(2220);
			27035: out = 16'(2148);
			27036: out = 16'(1187);
			27037: out = 16'(544);
			27038: out = 16'(2408);
			27039: out = 16'(891);
			27040: out = 16'(-603);
			27041: out = 16'(-1196);
			27042: out = 16'(659);
			27043: out = 16'(1268);
			27044: out = 16'(696);
			27045: out = 16'(-690);
			27046: out = 16'(-383);
			27047: out = 16'(615);
			27048: out = 16'(4341);
			27049: out = 16'(4703);
			27050: out = 16'(2103);
			27051: out = 16'(-72);
			27052: out = 16'(-1089);
			27053: out = 16'(198);
			27054: out = 16'(-445);
			27055: out = 16'(-3278);
			27056: out = 16'(-4530);
			27057: out = 16'(-846);
			27058: out = 16'(2902);
			27059: out = 16'(2906);
			27060: out = 16'(278);
			27061: out = 16'(1143);
			27062: out = 16'(3007);
			27063: out = 16'(2438);
			27064: out = 16'(-1440);
			27065: out = 16'(-158);
			27066: out = 16'(1639);
			27067: out = 16'(1204);
			27068: out = 16'(-1647);
			27069: out = 16'(-496);
			27070: out = 16'(1726);
			27071: out = 16'(4142);
			27072: out = 16'(5155);
			27073: out = 16'(2387);
			27074: out = 16'(-682);
			27075: out = 16'(-1988);
			27076: out = 16'(-873);
			27077: out = 16'(-424);
			27078: out = 16'(-587);
			27079: out = 16'(-1923);
			27080: out = 16'(-1934);
			27081: out = 16'(1719);
			27082: out = 16'(1970);
			27083: out = 16'(1417);
			27084: out = 16'(1100);
			27085: out = 16'(1025);
			27086: out = 16'(1716);
			27087: out = 16'(26);
			27088: out = 16'(-3273);
			27089: out = 16'(-5313);
			27090: out = 16'(-763);
			27091: out = 16'(678);
			27092: out = 16'(-2265);
			27093: out = 16'(-5274);
			27094: out = 16'(-2897);
			27095: out = 16'(403);
			27096: out = 16'(1279);
			27097: out = 16'(362);
			27098: out = 16'(-877);
			27099: out = 16'(2580);
			27100: out = 16'(4081);
			27101: out = 16'(2431);
			27102: out = 16'(-47);
			27103: out = 16'(-178);
			27104: out = 16'(-557);
			27105: out = 16'(-908);
			27106: out = 16'(-118);
			27107: out = 16'(-1370);
			27108: out = 16'(-2036);
			27109: out = 16'(-193);
			27110: out = 16'(3387);
			27111: out = 16'(3211);
			27112: out = 16'(988);
			27113: out = 16'(-697);
			27114: out = 16'(-11);
			27115: out = 16'(-308);
			27116: out = 16'(-2157);
			27117: out = 16'(-3515);
			27118: out = 16'(-1410);
			27119: out = 16'(1571);
			27120: out = 16'(770);
			27121: out = 16'(-1860);
			27122: out = 16'(-1386);
			27123: out = 16'(1730);
			27124: out = 16'(1217);
			27125: out = 16'(-3037);
			27126: out = 16'(-4825);
			27127: out = 16'(-187);
			27128: out = 16'(3172);
			27129: out = 16'(3273);
			27130: out = 16'(645);
			27131: out = 16'(-889);
			27132: out = 16'(-1156);
			27133: out = 16'(2178);
			27134: out = 16'(4738);
			27135: out = 16'(3977);
			27136: out = 16'(12);
			27137: out = 16'(-1802);
			27138: out = 16'(-1521);
			27139: out = 16'(-1743);
			27140: out = 16'(-3923);
			27141: out = 16'(-1455);
			27142: out = 16'(3749);
			27143: out = 16'(6646);
			27144: out = 16'(4045);
			27145: out = 16'(-3994);
			27146: out = 16'(-6376);
			27147: out = 16'(-3081);
			27148: out = 16'(-184);
			27149: out = 16'(523);
			27150: out = 16'(-234);
			27151: out = 16'(990);
			27152: out = 16'(3362);
			27153: out = 16'(2891);
			27154: out = 16'(857);
			27155: out = 16'(-2596);
			27156: out = 16'(-3640);
			27157: out = 16'(257);
			27158: out = 16'(1592);
			27159: out = 16'(892);
			27160: out = 16'(-732);
			27161: out = 16'(-1023);
			27162: out = 16'(-482);
			27163: out = 16'(-123);
			27164: out = 16'(-588);
			27165: out = 16'(-794);
			27166: out = 16'(3161);
			27167: out = 16'(2512);
			27168: out = 16'(-977);
			27169: out = 16'(-2672);
			27170: out = 16'(4254);
			27171: out = 16'(4414);
			27172: out = 16'(1064);
			27173: out = 16'(-2588);
			27174: out = 16'(-2580);
			27175: out = 16'(-733);
			27176: out = 16'(626);
			27177: out = 16'(-557);
			27178: out = 16'(-1637);
			27179: out = 16'(-1023);
			27180: out = 16'(2239);
			27181: out = 16'(2796);
			27182: out = 16'(-776);
			27183: out = 16'(-2393);
			27184: out = 16'(-1447);
			27185: out = 16'(59);
			27186: out = 16'(-721);
			27187: out = 16'(-2305);
			27188: out = 16'(-1510);
			27189: out = 16'(909);
			27190: out = 16'(1310);
			27191: out = 16'(-959);
			27192: out = 16'(-3028);
			27193: out = 16'(-2445);
			27194: out = 16'(-586);
			27195: out = 16'(-290);
			27196: out = 16'(-1286);
			27197: out = 16'(-1407);
			27198: out = 16'(1397);
			27199: out = 16'(4919);
			27200: out = 16'(4009);
			27201: out = 16'(848);
			27202: out = 16'(-2819);
			27203: out = 16'(-4763);
			27204: out = 16'(-1380);
			27205: out = 16'(-945);
			27206: out = 16'(-718);
			27207: out = 16'(30);
			27208: out = 16'(-190);
			27209: out = 16'(-1142);
			27210: out = 16'(-1974);
			27211: out = 16'(-1168);
			27212: out = 16'(-141);
			27213: out = 16'(183);
			27214: out = 16'(-575);
			27215: out = 16'(-706);
			27216: out = 16'(-189);
			27217: out = 16'(169);
			27218: out = 16'(-648);
			27219: out = 16'(-458);
			27220: out = 16'(647);
			27221: out = 16'(1417);
			27222: out = 16'(757);
			27223: out = 16'(380);
			27224: out = 16'(-260);
			27225: out = 16'(262);
			27226: out = 16'(-2662);
			27227: out = 16'(-588);
			27228: out = 16'(4356);
			27229: out = 16'(4585);
			27230: out = 16'(2340);
			27231: out = 16'(-680);
			27232: out = 16'(-2087);
			27233: out = 16'(-2477);
			27234: out = 16'(-1295);
			27235: out = 16'(-454);
			27236: out = 16'(-282);
			27237: out = 16'(247);
			27238: out = 16'(1469);
			27239: out = 16'(4281);
			27240: out = 16'(3302);
			27241: out = 16'(-623);
			27242: out = 16'(552);
			27243: out = 16'(950);
			27244: out = 16'(56);
			27245: out = 16'(-2039);
			27246: out = 16'(-142);
			27247: out = 16'(-367);
			27248: out = 16'(-39);
			27249: out = 16'(-312);
			27250: out = 16'(-25);
			27251: out = 16'(156);
			27252: out = 16'(330);
			27253: out = 16'(-982);
			27254: out = 16'(-2321);
			27255: out = 16'(-765);
			27256: out = 16'(2483);
			27257: out = 16'(3356);
			27258: out = 16'(413);
			27259: out = 16'(-1299);
			27260: out = 16'(-2333);
			27261: out = 16'(-35);
			27262: out = 16'(1688);
			27263: out = 16'(-111);
			27264: out = 16'(-2647);
			27265: out = 16'(-2170);
			27266: out = 16'(967);
			27267: out = 16'(2981);
			27268: out = 16'(2214);
			27269: out = 16'(1308);
			27270: out = 16'(702);
			27271: out = 16'(-1523);
			27272: out = 16'(-2802);
			27273: out = 16'(-4617);
			27274: out = 16'(-3911);
			27275: out = 16'(-1382);
			27276: out = 16'(-274);
			27277: out = 16'(-229);
			27278: out = 16'(602);
			27279: out = 16'(2466);
			27280: out = 16'(3654);
			27281: out = 16'(-335);
			27282: out = 16'(-4922);
			27283: out = 16'(-5632);
			27284: out = 16'(-2337);
			27285: out = 16'(813);
			27286: out = 16'(1653);
			27287: out = 16'(1068);
			27288: out = 16'(-250);
			27289: out = 16'(-611);
			27290: out = 16'(-1442);
			27291: out = 16'(-1029);
			27292: out = 16'(111);
			27293: out = 16'(228);
			27294: out = 16'(-1925);
			27295: out = 16'(-2623);
			27296: out = 16'(183);
			27297: out = 16'(3073);
			27298: out = 16'(3697);
			27299: out = 16'(2716);
			27300: out = 16'(1413);
			27301: out = 16'(-2395);
			27302: out = 16'(-508);
			27303: out = 16'(563);
			27304: out = 16'(64);
			27305: out = 16'(-3211);
			27306: out = 16'(-1024);
			27307: out = 16'(-341);
			27308: out = 16'(693);
			27309: out = 16'(1424);
			27310: out = 16'(3456);
			27311: out = 16'(1187);
			27312: out = 16'(-214);
			27313: out = 16'(258);
			27314: out = 16'(3895);
			27315: out = 16'(462);
			27316: out = 16'(-495);
			27317: out = 16'(1683);
			27318: out = 16'(1741);
			27319: out = 16'(319);
			27320: out = 16'(-220);
			27321: out = 16'(-1066);
			27322: out = 16'(-4812);
			27323: out = 16'(-4619);
			27324: out = 16'(14);
			27325: out = 16'(3657);
			27326: out = 16'(1493);
			27327: out = 16'(255);
			27328: out = 16'(869);
			27329: out = 16'(1732);
			27330: out = 16'(-1048);
			27331: out = 16'(-4842);
			27332: out = 16'(-5127);
			27333: out = 16'(-2124);
			27334: out = 16'(230);
			27335: out = 16'(2138);
			27336: out = 16'(2913);
			27337: out = 16'(3059);
			27338: out = 16'(1187);
			27339: out = 16'(181);
			27340: out = 16'(-3516);
			27341: out = 16'(-2150);
			27342: out = 16'(775);
			27343: out = 16'(1150);
			27344: out = 16'(153);
			27345: out = 16'(-258);
			27346: out = 16'(116);
			27347: out = 16'(-240);
			27348: out = 16'(-1381);
			27349: out = 16'(-934);
			27350: out = 16'(918);
			27351: out = 16'(2185);
			27352: out = 16'(3311);
			27353: out = 16'(-645);
			27354: out = 16'(-3406);
			27355: out = 16'(-2120);
			27356: out = 16'(1178);
			27357: out = 16'(3253);
			27358: out = 16'(972);
			27359: out = 16'(-2456);
			27360: out = 16'(-1855);
			27361: out = 16'(2055);
			27362: out = 16'(4024);
			27363: out = 16'(1584);
			27364: out = 16'(-789);
			27365: out = 16'(-634);
			27366: out = 16'(1675);
			27367: out = 16'(-136);
			27368: out = 16'(-4275);
			27369: out = 16'(-3307);
			27370: out = 16'(91);
			27371: out = 16'(1145);
			27372: out = 16'(-885);
			27373: out = 16'(-2992);
			27374: out = 16'(1706);
			27375: out = 16'(3132);
			27376: out = 16'(-419);
			27377: out = 16'(-4425);
			27378: out = 16'(-1139);
			27379: out = 16'(2224);
			27380: out = 16'(3459);
			27381: out = 16'(2799);
			27382: out = 16'(-1557);
			27383: out = 16'(-4418);
			27384: out = 16'(-3357);
			27385: out = 16'(217);
			27386: out = 16'(-19);
			27387: out = 16'(340);
			27388: out = 16'(1285);
			27389: out = 16'(2068);
			27390: out = 16'(2088);
			27391: out = 16'(-1383);
			27392: out = 16'(-1673);
			27393: out = 16'(643);
			27394: out = 16'(1047);
			27395: out = 16'(-3896);
			27396: out = 16'(-4062);
			27397: out = 16'(1941);
			27398: out = 16'(5080);
			27399: out = 16'(4379);
			27400: out = 16'(-2427);
			27401: out = 16'(-5171);
			27402: out = 16'(-1815);
			27403: out = 16'(-1014);
			27404: out = 16'(-2219);
			27405: out = 16'(-1809);
			27406: out = 16'(2766);
			27407: out = 16'(4539);
			27408: out = 16'(6922);
			27409: out = 16'(3735);
			27410: out = 16'(-1962);
			27411: out = 16'(-6937);
			27412: out = 16'(-1987);
			27413: out = 16'(2443);
			27414: out = 16'(2282);
			27415: out = 16'(-998);
			27416: out = 16'(-287);
			27417: out = 16'(858);
			27418: out = 16'(780);
			27419: out = 16'(-1144);
			27420: out = 16'(-9);
			27421: out = 16'(-191);
			27422: out = 16'(36);
			27423: out = 16'(-304);
			27424: out = 16'(-768);
			27425: out = 16'(-592);
			27426: out = 16'(1124);
			27427: out = 16'(1440);
			27428: out = 16'(-836);
			27429: out = 16'(-4198);
			27430: out = 16'(-2711);
			27431: out = 16'(834);
			27432: out = 16'(290);
			27433: out = 16'(-1474);
			27434: out = 16'(-3283);
			27435: out = 16'(-1485);
			27436: out = 16'(2589);
			27437: out = 16'(4806);
			27438: out = 16'(2813);
			27439: out = 16'(-1771);
			27440: out = 16'(-4604);
			27441: out = 16'(-4136);
			27442: out = 16'(93);
			27443: out = 16'(1340);
			27444: out = 16'(-250);
			27445: out = 16'(-644);
			27446: out = 16'(278);
			27447: out = 16'(743);
			27448: out = 16'(912);
			27449: out = 16'(2085);
			27450: out = 16'(452);
			27451: out = 16'(-1897);
			27452: out = 16'(-3025);
			27453: out = 16'(-1959);
			27454: out = 16'(481);
			27455: out = 16'(1730);
			27456: out = 16'(2227);
			27457: out = 16'(903);
			27458: out = 16'(-224);
			27459: out = 16'(-4381);
			27460: out = 16'(-3389);
			27461: out = 16'(686);
			27462: out = 16'(155);
			27463: out = 16'(-89);
			27464: out = 16'(2428);
			27465: out = 16'(5732);
			27466: out = 16'(4715);
			27467: out = 16'(-1347);
			27468: out = 16'(-3222);
			27469: out = 16'(-266);
			27470: out = 16'(1178);
			27471: out = 16'(1659);
			27472: out = 16'(372);
			27473: out = 16'(-83);
			27474: out = 16'(142);
			27475: out = 16'(1813);
			27476: out = 16'(2903);
			27477: out = 16'(2860);
			27478: out = 16'(1418);
			27479: out = 16'(-58);
			27480: out = 16'(-1357);
			27481: out = 16'(-2295);
			27482: out = 16'(-2001);
			27483: out = 16'(445);
			27484: out = 16'(1763);
			27485: out = 16'(1035);
			27486: out = 16'(-614);
			27487: out = 16'(-781);
			27488: out = 16'(-354);
			27489: out = 16'(-224);
			27490: out = 16'(-2480);
			27491: out = 16'(-5197);
			27492: out = 16'(-758);
			27493: out = 16'(3469);
			27494: out = 16'(5236);
			27495: out = 16'(2903);
			27496: out = 16'(393);
			27497: out = 16'(-3271);
			27498: out = 16'(-3514);
			27499: out = 16'(-2303);
			27500: out = 16'(-2185);
			27501: out = 16'(-1376);
			27502: out = 16'(1534);
			27503: out = 16'(3400);
			27504: out = 16'(1901);
			27505: out = 16'(287);
			27506: out = 16'(975);
			27507: out = 16'(1647);
			27508: out = 16'(-568);
			27509: out = 16'(-649);
			27510: out = 16'(-521);
			27511: out = 16'(189);
			27512: out = 16'(-238);
			27513: out = 16'(23);
			27514: out = 16'(-1313);
			27515: out = 16'(-974);
			27516: out = 16'(77);
			27517: out = 16'(-909);
			27518: out = 16'(-120);
			27519: out = 16'(31);
			27520: out = 16'(50);
			27521: out = 16'(-49);
			27522: out = 16'(615);
			27523: out = 16'(-895);
			27524: out = 16'(-2193);
			27525: out = 16'(-388);
			27526: out = 16'(142);
			27527: out = 16'(1770);
			27528: out = 16'(1349);
			27529: out = 16'(-95);
			27530: out = 16'(-787);
			27531: out = 16'(83);
			27532: out = 16'(466);
			27533: out = 16'(4);
			27534: out = 16'(539);
			27535: out = 16'(1538);
			27536: out = 16'(1804);
			27537: out = 16'(723);
			27538: out = 16'(-784);
			27539: out = 16'(-497);
			27540: out = 16'(637);
			27541: out = 16'(1346);
			27542: out = 16'(1090);
			27543: out = 16'(186);
			27544: out = 16'(-1385);
			27545: out = 16'(-2726);
			27546: out = 16'(-2712);
			27547: out = 16'(-314);
			27548: out = 16'(219);
			27549: out = 16'(-132);
			27550: out = 16'(330);
			27551: out = 16'(1701);
			27552: out = 16'(1201);
			27553: out = 16'(-699);
			27554: out = 16'(-1110);
			27555: out = 16'(1123);
			27556: out = 16'(1993);
			27557: out = 16'(195);
			27558: out = 16'(-1828);
			27559: out = 16'(-709);
			27560: out = 16'(111);
			27561: out = 16'(-28);
			27562: out = 16'(-1566);
			27563: out = 16'(-1840);
			27564: out = 16'(1224);
			27565: out = 16'(3459);
			27566: out = 16'(2269);
			27567: out = 16'(-1527);
			27568: out = 16'(-2715);
			27569: out = 16'(-2848);
			27570: out = 16'(-1141);
			27571: out = 16'(33);
			27572: out = 16'(3);
			27573: out = 16'(730);
			27574: out = 16'(2457);
			27575: out = 16'(2600);
			27576: out = 16'(523);
			27577: out = 16'(-358);
			27578: out = 16'(937);
			27579: out = 16'(1749);
			27580: out = 16'(921);
			27581: out = 16'(-5179);
			27582: out = 16'(-3283);
			27583: out = 16'(1421);
			27584: out = 16'(998);
			27585: out = 16'(-3545);
			27586: out = 16'(-5374);
			27587: out = 16'(-1818);
			27588: out = 16'(2481);
			27589: out = 16'(3087);
			27590: out = 16'(1358);
			27591: out = 16'(-465);
			27592: out = 16'(-550);
			27593: out = 16'(1200);
			27594: out = 16'(329);
			27595: out = 16'(-1592);
			27596: out = 16'(-3408);
			27597: out = 16'(-2522);
			27598: out = 16'(941);
			27599: out = 16'(3666);
			27600: out = 16'(2301);
			27601: out = 16'(-923);
			27602: out = 16'(318);
			27603: out = 16'(510);
			27604: out = 16'(-2299);
			27605: out = 16'(-4614);
			27606: out = 16'(1546);
			27607: out = 16'(3714);
			27608: out = 16'(1336);
			27609: out = 16'(-3001);
			27610: out = 16'(-2731);
			27611: out = 16'(-808);
			27612: out = 16'(60);
			27613: out = 16'(-1169);
			27614: out = 16'(-402);
			27615: out = 16'(1241);
			27616: out = 16'(3193);
			27617: out = 16'(1783);
			27618: out = 16'(-1849);
			27619: out = 16'(-3614);
			27620: out = 16'(-1155);
			27621: out = 16'(1767);
			27622: out = 16'(1469);
			27623: out = 16'(-365);
			27624: out = 16'(-1283);
			27625: out = 16'(618);
			27626: out = 16'(1707);
			27627: out = 16'(145);
			27628: out = 16'(-1467);
			27629: out = 16'(118);
			27630: out = 16'(1989);
			27631: out = 16'(207);
			27632: out = 16'(-3572);
			27633: out = 16'(-2743);
			27634: out = 16'(2347);
			27635: out = 16'(5001);
			27636: out = 16'(2743);
			27637: out = 16'(-1446);
			27638: out = 16'(-3307);
			27639: out = 16'(-2656);
			27640: out = 16'(364);
			27641: out = 16'(-317);
			27642: out = 16'(-636);
			27643: out = 16'(462);
			27644: out = 16'(1894);
			27645: out = 16'(1989);
			27646: out = 16'(1713);
			27647: out = 16'(520);
			27648: out = 16'(-2268);
			27649: out = 16'(-2432);
			27650: out = 16'(-784);
			27651: out = 16'(740);
			27652: out = 16'(-176);
			27653: out = 16'(168);
			27654: out = 16'(-562);
			27655: out = 16'(-663);
			27656: out = 16'(88);
			27657: out = 16'(1825);
			27658: out = 16'(-70);
			27659: out = 16'(-2934);
			27660: out = 16'(-2825);
			27661: out = 16'(1662);
			27662: out = 16'(1932);
			27663: out = 16'(59);
			27664: out = 16'(-263);
			27665: out = 16'(1755);
			27666: out = 16'(759);
			27667: out = 16'(-2053);
			27668: out = 16'(-1427);
			27669: out = 16'(3774);
			27670: out = 16'(741);
			27671: out = 16'(-2692);
			27672: out = 16'(-1777);
			27673: out = 16'(4527);
			27674: out = 16'(4982);
			27675: out = 16'(2171);
			27676: out = 16'(-1812);
			27677: out = 16'(-1805);
			27678: out = 16'(-754);
			27679: out = 16'(2968);
			27680: out = 16'(2193);
			27681: out = 16'(-997);
			27682: out = 16'(-2161);
			27683: out = 16'(209);
			27684: out = 16'(1101);
			27685: out = 16'(-1206);
			27686: out = 16'(-1719);
			27687: out = 16'(21);
			27688: out = 16'(3668);
			27689: out = 16'(40);
			27690: out = 16'(-8870);
			27691: out = 16'(-8087);
			27692: out = 16'(445);
			27693: out = 16'(5976);
			27694: out = 16'(2480);
			27695: out = 16'(-699);
			27696: out = 16'(-1092);
			27697: out = 16'(1512);
			27698: out = 16'(687);
			27699: out = 16'(-4740);
			27700: out = 16'(-5159);
			27701: out = 16'(-1012);
			27702: out = 16'(2691);
			27703: out = 16'(1810);
			27704: out = 16'(1696);
			27705: out = 16'(1182);
			27706: out = 16'(1403);
			27707: out = 16'(19);
			27708: out = 16'(-2106);
			27709: out = 16'(-5302);
			27710: out = 16'(-3952);
			27711: out = 16'(1080);
			27712: out = 16'(5298);
			27713: out = 16'(649);
			27714: out = 16'(-2649);
			27715: out = 16'(837);
			27716: out = 16'(4276);
			27717: out = 16'(2549);
			27718: out = 16'(-2154);
			27719: out = 16'(-2776);
			27720: out = 16'(-190);
			27721: out = 16'(2246);
			27722: out = 16'(-1106);
			27723: out = 16'(-3165);
			27724: out = 16'(539);
			27725: out = 16'(1793);
			27726: out = 16'(636);
			27727: out = 16'(-1338);
			27728: out = 16'(-1204);
			27729: out = 16'(-195);
			27730: out = 16'(-461);
			27731: out = 16'(-90);
			27732: out = 16'(1961);
			27733: out = 16'(2999);
			27734: out = 16'(2545);
			27735: out = 16'(639);
			27736: out = 16'(-1331);
			27737: out = 16'(-2033);
			27738: out = 16'(-1302);
			27739: out = 16'(223);
			27740: out = 16'(17);
			27741: out = 16'(-1169);
			27742: out = 16'(608);
			27743: out = 16'(4810);
			27744: out = 16'(5535);
			27745: out = 16'(1193);
			27746: out = 16'(-1174);
			27747: out = 16'(-1373);
			27748: out = 16'(-1236);
			27749: out = 16'(-2189);
			27750: out = 16'(611);
			27751: out = 16'(1169);
			27752: out = 16'(240);
			27753: out = 16'(-2162);
			27754: out = 16'(-2749);
			27755: out = 16'(-1505);
			27756: out = 16'(-73);
			27757: out = 16'(289);
			27758: out = 16'(2233);
			27759: out = 16'(1172);
			27760: out = 16'(1901);
			27761: out = 16'(766);
			27762: out = 16'(-2450);
			27763: out = 16'(-2323);
			27764: out = 16'(-111);
			27765: out = 16'(1980);
			27766: out = 16'(1396);
			27767: out = 16'(-1127);
			27768: out = 16'(-2377);
			27769: out = 16'(-1240);
			27770: out = 16'(175);
			27771: out = 16'(47);
			27772: out = 16'(1331);
			27773: out = 16'(3062);
			27774: out = 16'(3032);
			27775: out = 16'(-382);
			27776: out = 16'(-4174);
			27777: out = 16'(-5543);
			27778: out = 16'(-2477);
			27779: out = 16'(2271);
			27780: out = 16'(3121);
			27781: out = 16'(3197);
			27782: out = 16'(2877);
			27783: out = 16'(927);
			27784: out = 16'(-5897);
			27785: out = 16'(-8110);
			27786: out = 16'(-4348);
			27787: out = 16'(1805);
			27788: out = 16'(2999);
			27789: out = 16'(3581);
			27790: out = 16'(2546);
			27791: out = 16'(1986);
			27792: out = 16'(1791);
			27793: out = 16'(452);
			27794: out = 16'(-1924);
			27795: out = 16'(-2501);
			27796: out = 16'(271);
			27797: out = 16'(-136);
			27798: out = 16'(489);
			27799: out = 16'(829);
			27800: out = 16'(1622);
			27801: out = 16'(3379);
			27802: out = 16'(3563);
			27803: out = 16'(1663);
			27804: out = 16'(-343);
			27805: out = 16'(-349);
			27806: out = 16'(-129);
			27807: out = 16'(-362);
			27808: out = 16'(127);
			27809: out = 16'(1643);
			27810: out = 16'(3381);
			27811: out = 16'(1691);
			27812: out = 16'(-889);
			27813: out = 16'(-994);
			27814: out = 16'(-600);
			27815: out = 16'(-1155);
			27816: out = 16'(-1431);
			27817: out = 16'(846);
			27818: out = 16'(744);
			27819: out = 16'(1738);
			27820: out = 16'(911);
			27821: out = 16'(-773);
			27822: out = 16'(-2435);
			27823: out = 16'(-1571);
			27824: out = 16'(-1120);
			27825: out = 16'(-2148);
			27826: out = 16'(-2829);
			27827: out = 16'(273);
			27828: out = 16'(5130);
			27829: out = 16'(6670);
			27830: out = 16'(2296);
			27831: out = 16'(-3743);
			27832: out = 16'(-7598);
			27833: out = 16'(-6533);
			27834: out = 16'(-2586);
			27835: out = 16'(827);
			27836: out = 16'(1910);
			27837: out = 16'(1709);
			27838: out = 16'(1084);
			27839: out = 16'(44);
			27840: out = 16'(-1097);
			27841: out = 16'(-2062);
			27842: out = 16'(-1934);
			27843: out = 16'(-18);
			27844: out = 16'(1470);
			27845: out = 16'(1934);
			27846: out = 16'(526);
			27847: out = 16'(-1444);
			27848: out = 16'(-1813);
			27849: out = 16'(118);
			27850: out = 16'(1242);
			27851: out = 16'(-370);
			27852: out = 16'(-685);
			27853: out = 16'(-460);
			27854: out = 16'(369);
			27855: out = 16'(342);
			27856: out = 16'(-36);
			27857: out = 16'(-795);
			27858: out = 16'(-353);
			27859: out = 16'(604);
			27860: out = 16'(416);
			27861: out = 16'(-437);
			27862: out = 16'(-1108);
			27863: out = 16'(-222);
			27864: out = 16'(1916);
			27865: out = 16'(1443);
			27866: out = 16'(1354);
			27867: out = 16'(2322);
			27868: out = 16'(2680);
			27869: out = 16'(562);
			27870: out = 16'(-3158);
			27871: out = 16'(-4017);
			27872: out = 16'(-145);
			27873: out = 16'(3059);
			27874: out = 16'(2871);
			27875: out = 16'(495);
			27876: out = 16'(-206);
			27877: out = 16'(-695);
			27878: out = 16'(616);
			27879: out = 16'(-1282);
			27880: out = 16'(-2904);
			27881: out = 16'(-315);
			27882: out = 16'(1512);
			27883: out = 16'(879);
			27884: out = 16'(-525);
			27885: out = 16'(170);
			27886: out = 16'(4394);
			27887: out = 16'(3484);
			27888: out = 16'(-1441);
			27889: out = 16'(-5231);
			27890: out = 16'(-2912);
			27891: out = 16'(143);
			27892: out = 16'(1057);
			27893: out = 16'(-426);
			27894: out = 16'(126);
			27895: out = 16'(857);
			27896: out = 16'(3088);
			27897: out = 16'(2564);
			27898: out = 16'(-718);
			27899: out = 16'(-4962);
			27900: out = 16'(-2106);
			27901: out = 16'(2814);
			27902: out = 16'(2521);
			27903: out = 16'(-3222);
			27904: out = 16'(-3109);
			27905: out = 16'(2155);
			27906: out = 16'(3973);
			27907: out = 16'(-585);
			27908: out = 16'(-3850);
			27909: out = 16'(-2473);
			27910: out = 16'(-262);
			27911: out = 16'(-2761);
			27912: out = 16'(-1480);
			27913: out = 16'(2625);
			27914: out = 16'(4956);
			27915: out = 16'(1146);
			27916: out = 16'(-2637);
			27917: out = 16'(-3788);
			27918: out = 16'(-1361);
			27919: out = 16'(-416);
			27920: out = 16'(470);
			27921: out = 16'(-2701);
			27922: out = 16'(-3732);
			27923: out = 16'(509);
			27924: out = 16'(4260);
			27925: out = 16'(2475);
			27926: out = 16'(-1809);
			27927: out = 16'(-2361);
			27928: out = 16'(-642);
			27929: out = 16'(2673);
			27930: out = 16'(1946);
			27931: out = 16'(-230);
			27932: out = 16'(-121);
			27933: out = 16'(1093);
			27934: out = 16'(9);
			27935: out = 16'(-1753);
			27936: out = 16'(-850);
			27937: out = 16'(-54);
			27938: out = 16'(-1806);
			27939: out = 16'(-3912);
			27940: out = 16'(-1603);
			27941: out = 16'(1158);
			27942: out = 16'(3261);
			27943: out = 16'(2266);
			27944: out = 16'(462);
			27945: out = 16'(-84);
			27946: out = 16'(-270);
			27947: out = 16'(-2812);
			27948: out = 16'(-5934);
			27949: out = 16'(-2070);
			27950: out = 16'(741);
			27951: out = 16'(3521);
			27952: out = 16'(2794);
			27953: out = 16'(-1250);
			27954: out = 16'(-2418);
			27955: out = 16'(25);
			27956: out = 16'(2631);
			27957: out = 16'(3120);
			27958: out = 16'(988);
			27959: out = 16'(1365);
			27960: out = 16'(1384);
			27961: out = 16'(-1332);
			27962: out = 16'(-4002);
			27963: out = 16'(-1955);
			27964: out = 16'(1478);
			27965: out = 16'(1513);
			27966: out = 16'(318);
			27967: out = 16'(-405);
			27968: out = 16'(1153);
			27969: out = 16'(1637);
			27970: out = 16'(738);
			27971: out = 16'(-1943);
			27972: out = 16'(-297);
			27973: out = 16'(2270);
			27974: out = 16'(947);
			27975: out = 16'(-2107);
			27976: out = 16'(-1976);
			27977: out = 16'(1677);
			27978: out = 16'(3200);
			27979: out = 16'(855);
			27980: out = 16'(-2087);
			27981: out = 16'(-250);
			27982: out = 16'(3816);
			27983: out = 16'(2008);
			27984: out = 16'(-2403);
			27985: out = 16'(-4830);
			27986: out = 16'(-1521);
			27987: out = 16'(2502);
			27988: out = 16'(2976);
			27989: out = 16'(-871);
			27990: out = 16'(-1918);
			27991: out = 16'(3682);
			27992: out = 16'(3924);
			27993: out = 16'(569);
			27994: out = 16'(-3072);
			27995: out = 16'(-1758);
			27996: out = 16'(2014);
			27997: out = 16'(3013);
			27998: out = 16'(-191);
			27999: out = 16'(-2847);
			28000: out = 16'(-683);
			28001: out = 16'(1182);
			28002: out = 16'(-418);
			28003: out = 16'(-3394);
			28004: out = 16'(-3762);
			28005: out = 16'(-607);
			28006: out = 16'(1025);
			28007: out = 16'(232);
			28008: out = 16'(191);
			28009: out = 16'(3569);
			28010: out = 16'(4077);
			28011: out = 16'(-280);
			28012: out = 16'(-4090);
			28013: out = 16'(-2765);
			28014: out = 16'(2028);
			28015: out = 16'(2621);
			28016: out = 16'(-1436);
			28017: out = 16'(-5514);
			28018: out = 16'(-2702);
			28019: out = 16'(2053);
			28020: out = 16'(3315);
			28021: out = 16'(792);
			28022: out = 16'(-686);
			28023: out = 16'(-665);
			28024: out = 16'(-542);
			28025: out = 16'(-3813);
			28026: out = 16'(-1469);
			28027: out = 16'(-352);
			28028: out = 16'(901);
			28029: out = 16'(3560);
			28030: out = 16'(1042);
			28031: out = 16'(-2448);
			28032: out = 16'(-3041);
			28033: out = 16'(-924);
			28034: out = 16'(-2203);
			28035: out = 16'(-4749);
			28036: out = 16'(-2174);
			28037: out = 16'(4552);
			28038: out = 16'(5503);
			28039: out = 16'(-1217);
			28040: out = 16'(-6111);
			28041: out = 16'(-2735);
			28042: out = 16'(1416);
			28043: out = 16'(1333);
			28044: out = 16'(-1166);
			28045: out = 16'(-270);
			28046: out = 16'(3036);
			28047: out = 16'(2732);
			28048: out = 16'(-361);
			28049: out = 16'(-2299);
			28050: out = 16'(-1258);
			28051: out = 16'(-169);
			28052: out = 16'(1264);
			28053: out = 16'(2732);
			28054: out = 16'(3834);
			28055: out = 16'(3740);
			28056: out = 16'(2167);
			28057: out = 16'(369);
			28058: out = 16'(-236);
			28059: out = 16'(-271);
			28060: out = 16'(88);
			28061: out = 16'(-1978);
			28062: out = 16'(-5223);
			28063: out = 16'(-4823);
			28064: out = 16'(-1581);
			28065: out = 16'(3387);
			28066: out = 16'(5279);
			28067: out = 16'(3437);
			28068: out = 16'(-783);
			28069: out = 16'(-1669);
			28070: out = 16'(-403);
			28071: out = 16'(-163);
			28072: out = 16'(12);
			28073: out = 16'(-119);
			28074: out = 16'(9);
			28075: out = 16'(-72);
			28076: out = 16'(-53);
			28077: out = 16'(890);
			28078: out = 16'(677);
			28079: out = 16'(-1637);
			28080: out = 16'(-2652);
			28081: out = 16'(-3376);
			28082: out = 16'(-707);
			28083: out = 16'(1951);
			28084: out = 16'(2511);
			28085: out = 16'(441);
			28086: out = 16'(-473);
			28087: out = 16'(-1484);
			28088: out = 16'(-3043);
			28089: out = 16'(-4379);
			28090: out = 16'(-1712);
			28091: out = 16'(1347);
			28092: out = 16'(1851);
			28093: out = 16'(185);
			28094: out = 16'(298);
			28095: out = 16'(845);
			28096: out = 16'(600);
			28097: out = 16'(-43);
			28098: out = 16'(396);
			28099: out = 16'(365);
			28100: out = 16'(-609);
			28101: out = 16'(-2126);
			28102: out = 16'(-1110);
			28103: out = 16'(1599);
			28104: out = 16'(5230);
			28105: out = 16'(5801);
			28106: out = 16'(2449);
			28107: out = 16'(-3058);
			28108: out = 16'(-2798);
			28109: out = 16'(2295);
			28110: out = 16'(1915);
			28111: out = 16'(-2465);
			28112: out = 16'(-3697);
			28113: out = 16'(1374);
			28114: out = 16'(3040);
			28115: out = 16'(2957);
			28116: out = 16'(9);
			28117: out = 16'(-664);
			28118: out = 16'(-421);
			28119: out = 16'(818);
			28120: out = 16'(-1562);
			28121: out = 16'(-2563);
			28122: out = 16'(801);
			28123: out = 16'(3192);
			28124: out = 16'(1843);
			28125: out = 16'(-2069);
			28126: out = 16'(-4449);
			28127: out = 16'(-2720);
			28128: out = 16'(-156);
			28129: out = 16'(583);
			28130: out = 16'(-173);
			28131: out = 16'(51);
			28132: out = 16'(-646);
			28133: out = 16'(-1199);
			28134: out = 16'(-1634);
			28135: out = 16'(-1413);
			28136: out = 16'(-381);
			28137: out = 16'(622);
			28138: out = 16'(303);
			28139: out = 16'(-703);
			28140: out = 16'(-1017);
			28141: out = 16'(1656);
			28142: out = 16'(3119);
			28143: out = 16'(880);
			28144: out = 16'(210);
			28145: out = 16'(-296);
			28146: out = 16'(244);
			28147: out = 16'(-242);
			28148: out = 16'(157);
			28149: out = 16'(-1901);
			28150: out = 16'(-1109);
			28151: out = 16'(781);
			28152: out = 16'(26);
			28153: out = 16'(1499);
			28154: out = 16'(2288);
			28155: out = 16'(897);
			28156: out = 16'(-2297);
			28157: out = 16'(-4827);
			28158: out = 16'(-3320);
			28159: out = 16'(-490);
			28160: out = 16'(227);
			28161: out = 16'(3051);
			28162: out = 16'(2368);
			28163: out = 16'(-33);
			28164: out = 16'(-2048);
			28165: out = 16'(-82);
			28166: out = 16'(2707);
			28167: out = 16'(3499);
			28168: out = 16'(1166);
			28169: out = 16'(269);
			28170: out = 16'(-3059);
			28171: out = 16'(-3338);
			28172: out = 16'(-1213);
			28173: out = 16'(2029);
			28174: out = 16'(373);
			28175: out = 16'(218);
			28176: out = 16'(513);
			28177: out = 16'(-68);
			28178: out = 16'(59);
			28179: out = 16'(-92);
			28180: out = 16'(-99);
			28181: out = 16'(182);
			28182: out = 16'(1657);
			28183: out = 16'(1607);
			28184: out = 16'(361);
			28185: out = 16'(-1215);
			28186: out = 16'(-2783);
			28187: out = 16'(-1884);
			28188: out = 16'(-680);
			28189: out = 16'(331);
			28190: out = 16'(588);
			28191: out = 16'(1804);
			28192: out = 16'(1201);
			28193: out = 16'(815);
			28194: out = 16'(1877);
			28195: out = 16'(3367);
			28196: out = 16'(171);
			28197: out = 16'(-5302);
			28198: out = 16'(-7281);
			28199: out = 16'(-396);
			28200: out = 16'(3292);
			28201: out = 16'(2344);
			28202: out = 16'(-30);
			28203: out = 16'(1882);
			28204: out = 16'(1833);
			28205: out = 16'(1161);
			28206: out = 16'(-995);
			28207: out = 16'(-4038);
			28208: out = 16'(-2965);
			28209: out = 16'(249);
			28210: out = 16'(1871);
			28211: out = 16'(412);
			28212: out = 16'(-571);
			28213: out = 16'(-351);
			28214: out = 16'(158);
			28215: out = 16'(-59);
			28216: out = 16'(-1266);
			28217: out = 16'(-608);
			28218: out = 16'(-476);
			28219: out = 16'(-2616);
			28220: out = 16'(-4398);
			28221: out = 16'(-2373);
			28222: out = 16'(1715);
			28223: out = 16'(2679);
			28224: out = 16'(446);
			28225: out = 16'(-3762);
			28226: out = 16'(-3470);
			28227: out = 16'(-82);
			28228: out = 16'(1334);
			28229: out = 16'(653);
			28230: out = 16'(39);
			28231: out = 16'(434);
			28232: out = 16'(-129);
			28233: out = 16'(-3259);
			28234: out = 16'(-4165);
			28235: out = 16'(-586);
			28236: out = 16'(4430);
			28237: out = 16'(4764);
			28238: out = 16'(2748);
			28239: out = 16'(501);
			28240: out = 16'(342);
			28241: out = 16'(-102);
			28242: out = 16'(-85);
			28243: out = 16'(-1918);
			28244: out = 16'(-1761);
			28245: out = 16'(2046);
			28246: out = 16'(3679);
			28247: out = 16'(1873);
			28248: out = 16'(-281);
			28249: out = 16'(287);
			28250: out = 16'(1149);
			28251: out = 16'(260);
			28252: out = 16'(-845);
			28253: out = 16'(511);
			28254: out = 16'(1539);
			28255: out = 16'(1469);
			28256: out = 16'(-687);
			28257: out = 16'(-1966);
			28258: out = 16'(-901);
			28259: out = 16'(26);
			28260: out = 16'(-62);
			28261: out = 16'(138);
			28262: out = 16'(426);
			28263: out = 16'(2763);
			28264: out = 16'(1652);
			28265: out = 16'(-535);
			28266: out = 16'(-568);
			28267: out = 16'(1343);
			28268: out = 16'(1136);
			28269: out = 16'(-1400);
			28270: out = 16'(-3566);
			28271: out = 16'(-3636);
			28272: out = 16'(-1314);
			28273: out = 16'(1656);
			28274: out = 16'(3914);
			28275: out = 16'(4506);
			28276: out = 16'(2373);
			28277: out = 16'(-561);
			28278: out = 16'(-2609);
			28279: out = 16'(-3561);
			28280: out = 16'(-2553);
			28281: out = 16'(-1358);
			28282: out = 16'(-461);
			28283: out = 16'(113);
			28284: out = 16'(51);
			28285: out = 16'(1085);
			28286: out = 16'(2049);
			28287: out = 16'(830);
			28288: out = 16'(-1427);
			28289: out = 16'(-2973);
			28290: out = 16'(-1612);
			28291: out = 16'(294);
			28292: out = 16'(2045);
			28293: out = 16'(490);
			28294: out = 16'(783);
			28295: out = 16'(1949);
			28296: out = 16'(1925);
			28297: out = 16'(-1803);
			28298: out = 16'(-1870);
			28299: out = 16'(489);
			28300: out = 16'(-202);
			28301: out = 16'(4);
			28302: out = 16'(823);
			28303: out = 16'(2170);
			28304: out = 16'(1462);
			28305: out = 16'(-343);
			28306: out = 16'(-1186);
			28307: out = 16'(-383);
			28308: out = 16'(-189);
			28309: out = 16'(-636);
			28310: out = 16'(-1018);
			28311: out = 16'(-160);
			28312: out = 16'(813);
			28313: out = 16'(1785);
			28314: out = 16'(-1038);
			28315: out = 16'(-2692);
			28316: out = 16'(-1471);
			28317: out = 16'(-186);
			28318: out = 16'(260);
			28319: out = 16'(-1421);
			28320: out = 16'(-1487);
			28321: out = 16'(839);
			28322: out = 16'(5628);
			28323: out = 16'(3015);
			28324: out = 16'(-2017);
			28325: out = 16'(-3048);
			28326: out = 16'(-636);
			28327: out = 16'(74);
			28328: out = 16'(-2524);
			28329: out = 16'(-3661);
			28330: out = 16'(-260);
			28331: out = 16'(4837);
			28332: out = 16'(5367);
			28333: out = 16'(1556);
			28334: out = 16'(-1911);
			28335: out = 16'(-2006);
			28336: out = 16'(-933);
			28337: out = 16'(-977);
			28338: out = 16'(-543);
			28339: out = 16'(155);
			28340: out = 16'(2311);
			28341: out = 16'(2237);
			28342: out = 16'(-346);
			28343: out = 16'(-1323);
			28344: out = 16'(-785);
			28345: out = 16'(45);
			28346: out = 16'(-573);
			28347: out = 16'(-2607);
			28348: out = 16'(-1651);
			28349: out = 16'(660);
			28350: out = 16'(1766);
			28351: out = 16'(0);
			28352: out = 16'(950);
			28353: out = 16'(1074);
			28354: out = 16'(-232);
			28355: out = 16'(-2157);
			28356: out = 16'(-2230);
			28357: out = 16'(-690);
			28358: out = 16'(1799);
			28359: out = 16'(3502);
			28360: out = 16'(3152);
			28361: out = 16'(2042);
			28362: out = 16'(1745);
			28363: out = 16'(1216);
			28364: out = 16'(-1271);
			28365: out = 16'(-5254);
			28366: out = 16'(-5817);
			28367: out = 16'(-1100);
			28368: out = 16'(4146);
			28369: out = 16'(5036);
			28370: out = 16'(2226);
			28371: out = 16'(-1046);
			28372: out = 16'(-2851);
			28373: out = 16'(-1397);
			28374: out = 16'(-605);
			28375: out = 16'(-1644);
			28376: out = 16'(-3445);
			28377: out = 16'(-484);
			28378: out = 16'(1304);
			28379: out = 16'(2339);
			28380: out = 16'(2917);
			28381: out = 16'(1205);
			28382: out = 16'(454);
			28383: out = 16'(-1329);
			28384: out = 16'(-2711);
			28385: out = 16'(-77);
			28386: out = 16'(-955);
			28387: out = 16'(-2339);
			28388: out = 16'(-2024);
			28389: out = 16'(1973);
			28390: out = 16'(1913);
			28391: out = 16'(966);
			28392: out = 16'(-315);
			28393: out = 16'(134);
			28394: out = 16'(-921);
			28395: out = 16'(-199);
			28396: out = 16'(-267);
			28397: out = 16'(-723);
			28398: out = 16'(-1014);
			28399: out = 16'(2127);
			28400: out = 16'(3775);
			28401: out = 16'(2317);
			28402: out = 16'(102);
			28403: out = 16'(545);
			28404: out = 16'(1085);
			28405: out = 16'(-510);
			28406: out = 16'(-2681);
			28407: out = 16'(-1049);
			28408: out = 16'(1860);
			28409: out = 16'(2184);
			28410: out = 16'(-1096);
			28411: out = 16'(-1452);
			28412: out = 16'(-1269);
			28413: out = 16'(-752);
			28414: out = 16'(-849);
			28415: out = 16'(-58);
			28416: out = 16'(1003);
			28417: out = 16'(2148);
			28418: out = 16'(1195);
			28419: out = 16'(-420);
			28420: out = 16'(-1478);
			28421: out = 16'(1799);
			28422: out = 16'(5008);
			28423: out = 16'(2695);
			28424: out = 16'(-2132);
			28425: out = 16'(-3795);
			28426: out = 16'(-1217);
			28427: out = 16'(251);
			28428: out = 16'(1248);
			28429: out = 16'(573);
			28430: out = 16'(830);
			28431: out = 16'(1616);
			28432: out = 16'(1728);
			28433: out = 16'(449);
			28434: out = 16'(-261);
			28435: out = 16'(265);
			28436: out = 16'(-1049);
			28437: out = 16'(-1853);
			28438: out = 16'(-2111);
			28439: out = 16'(-445);
			28440: out = 16'(-511);
			28441: out = 16'(1217);
			28442: out = 16'(-590);
			28443: out = 16'(-1946);
			28444: out = 16'(325);
			28445: out = 16'(3910);
			28446: out = 16'(2271);
			28447: out = 16'(-878);
			28448: out = 16'(-93);
			28449: out = 16'(750);
			28450: out = 16'(-993);
			28451: out = 16'(-4142);
			28452: out = 16'(-3630);
			28453: out = 16'(834);
			28454: out = 16'(4015);
			28455: out = 16'(3475);
			28456: out = 16'(1102);
			28457: out = 16'(-851);
			28458: out = 16'(-2522);
			28459: out = 16'(-3201);
			28460: out = 16'(-2740);
			28461: out = 16'(-2263);
			28462: out = 16'(-1134);
			28463: out = 16'(-346);
			28464: out = 16'(76);
			28465: out = 16'(-43);
			28466: out = 16'(517);
			28467: out = 16'(595);
			28468: out = 16'(119);
			28469: out = 16'(-1055);
			28470: out = 16'(-2524);
			28471: out = 16'(-1945);
			28472: out = 16'(937);
			28473: out = 16'(2777);
			28474: out = 16'(310);
			28475: out = 16'(-1192);
			28476: out = 16'(-1422);
			28477: out = 16'(-1499);
			28478: out = 16'(-524);
			28479: out = 16'(-1546);
			28480: out = 16'(61);
			28481: out = 16'(1287);
			28482: out = 16'(787);
			28483: out = 16'(-1830);
			28484: out = 16'(582);
			28485: out = 16'(3627);
			28486: out = 16'(2511);
			28487: out = 16'(-1948);
			28488: out = 16'(-2444);
			28489: out = 16'(-657);
			28490: out = 16'(254);
			28491: out = 16'(2711);
			28492: out = 16'(3584);
			28493: out = 16'(2333);
			28494: out = 16'(213);
			28495: out = 16'(-370);
			28496: out = 16'(-134);
			28497: out = 16'(-1675);
			28498: out = 16'(-2317);
			28499: out = 16'(1821);
			28500: out = 16'(4066);
			28501: out = 16'(3180);
			28502: out = 16'(881);
			28503: out = 16'(-307);
			28504: out = 16'(331);
			28505: out = 16'(-1862);
			28506: out = 16'(-2418);
			28507: out = 16'(1063);
			28508: out = 16'(3955);
			28509: out = 16'(1915);
			28510: out = 16'(-623);
			28511: out = 16'(133);
			28512: out = 16'(1236);
			28513: out = 16'(332);
			28514: out = 16'(-750);
			28515: out = 16'(-423);
			28516: out = 16'(-1312);
			28517: out = 16'(993);
			28518: out = 16'(1723);
			28519: out = 16'(562);
			28520: out = 16'(-2616);
			28521: out = 16'(-1384);
			28522: out = 16'(-391);
			28523: out = 16'(331);
			28524: out = 16'(270);
			28525: out = 16'(206);
			28526: out = 16'(-227);
			28527: out = 16'(-801);
			28528: out = 16'(-878);
			28529: out = 16'(805);
			28530: out = 16'(2712);
			28531: out = 16'(2117);
			28532: out = 16'(-1602);
			28533: out = 16'(-4150);
			28534: out = 16'(-4555);
			28535: out = 16'(-1640);
			28536: out = 16'(-380);
			28537: out = 16'(-1510);
			28538: out = 16'(-2472);
			28539: out = 16'(994);
			28540: out = 16'(4044);
			28541: out = 16'(2926);
			28542: out = 16'(138);
			28543: out = 16'(-278);
			28544: out = 16'(311);
			28545: out = 16'(-390);
			28546: out = 16'(356);
			28547: out = 16'(975);
			28548: out = 16'(2534);
			28549: out = 16'(2779);
			28550: out = 16'(-503);
			28551: out = 16'(-2016);
			28552: out = 16'(-2487);
			28553: out = 16'(-1112);
			28554: out = 16'(-56);
			28555: out = 16'(281);
			28556: out = 16'(-2862);
			28557: out = 16'(-3577);
			28558: out = 16'(1033);
			28559: out = 16'(3925);
			28560: out = 16'(1629);
			28561: out = 16'(-3008);
			28562: out = 16'(-3996);
			28563: out = 16'(-2170);
			28564: out = 16'(-237);
			28565: out = 16'(-1210);
			28566: out = 16'(-1672);
			28567: out = 16'(1638);
			28568: out = 16'(2478);
			28569: out = 16'(831);
			28570: out = 16'(-793);
			28571: out = 16'(1920);
			28572: out = 16'(18);
			28573: out = 16'(-1355);
			28574: out = 16'(-2301);
			28575: out = 16'(-565);
			28576: out = 16'(-1878);
			28577: out = 16'(1299);
			28578: out = 16'(3410);
			28579: out = 16'(3096);
			28580: out = 16'(-791);
			28581: out = 16'(710);
			28582: out = 16'(1318);
			28583: out = 16'(-1328);
			28584: out = 16'(-7083);
			28585: out = 16'(-2624);
			28586: out = 16'(2056);
			28587: out = 16'(2685);
			28588: out = 16'(1858);
			28589: out = 16'(1659);
			28590: out = 16'(934);
			28591: out = 16'(-1049);
			28592: out = 16'(-2886);
			28593: out = 16'(-3618);
			28594: out = 16'(-1744);
			28595: out = 16'(957);
			28596: out = 16'(1662);
			28597: out = 16'(2131);
			28598: out = 16'(-952);
			28599: out = 16'(-1733);
			28600: out = 16'(461);
			28601: out = 16'(1627);
			28602: out = 16'(525);
			28603: out = 16'(-13);
			28604: out = 16'(422);
			28605: out = 16'(-1590);
			28606: out = 16'(-426);
			28607: out = 16'(926);
			28608: out = 16'(1649);
			28609: out = 16'(144);
			28610: out = 16'(-1793);
			28611: out = 16'(-1419);
			28612: out = 16'(890);
			28613: out = 16'(1399);
			28614: out = 16'(386);
			28615: out = 16'(-669);
			28616: out = 16'(1873);
			28617: out = 16'(4826);
			28618: out = 16'(1856);
			28619: out = 16'(-407);
			28620: out = 16'(-979);
			28621: out = 16'(-321);
			28622: out = 16'(-210);
			28623: out = 16'(-2418);
			28624: out = 16'(-2396);
			28625: out = 16'(-360);
			28626: out = 16'(171);
			28627: out = 16'(-82);
			28628: out = 16'(271);
			28629: out = 16'(1423);
			28630: out = 16'(695);
			28631: out = 16'(310);
			28632: out = 16'(-3640);
			28633: out = 16'(-6692);
			28634: out = 16'(-5350);
			28635: out = 16'(2714);
			28636: out = 16'(4857);
			28637: out = 16'(3311);
			28638: out = 16'(1696);
			28639: out = 16'(2185);
			28640: out = 16'(683);
			28641: out = 16'(-2021);
			28642: out = 16'(-3766);
			28643: out = 16'(-2838);
			28644: out = 16'(-575);
			28645: out = 16'(-513);
			28646: out = 16'(-1627);
			28647: out = 16'(-466);
			28648: out = 16'(122);
			28649: out = 16'(-216);
			28650: out = 16'(-2566);
			28651: out = 16'(-2859);
			28652: out = 16'(-649);
			28653: out = 16'(4080);
			28654: out = 16'(3599);
			28655: out = 16'(-1205);
			28656: out = 16'(-5261);
			28657: out = 16'(-559);
			28658: out = 16'(3425);
			28659: out = 16'(2059);
			28660: out = 16'(-464);
			28661: out = 16'(-3166);
			28662: out = 16'(-2857);
			28663: out = 16'(-1285);
			28664: out = 16'(1036);
			28665: out = 16'(3104);
			28666: out = 16'(4530);
			28667: out = 16'(3848);
			28668: out = 16'(1116);
			28669: out = 16'(-4788);
			28670: out = 16'(-5906);
			28671: out = 16'(-2756);
			28672: out = 16'(968);
			28673: out = 16'(1915);
			28674: out = 16'(1807);
			28675: out = 16'(2995);
			28676: out = 16'(4704);
			28677: out = 16'(3203);
			28678: out = 16'(-578);
			28679: out = 16'(-4647);
			28680: out = 16'(-5156);
			28681: out = 16'(-2065);
			28682: out = 16'(745);
			28683: out = 16'(2577);
			28684: out = 16'(4163);
			28685: out = 16'(4031);
			28686: out = 16'(801);
			28687: out = 16'(-3586);
			28688: out = 16'(-4422);
			28689: out = 16'(-1977);
			28690: out = 16'(-2714);
			28691: out = 16'(-2602);
			28692: out = 16'(679);
			28693: out = 16'(5196);
			28694: out = 16'(3290);
			28695: out = 16'(91);
			28696: out = 16'(-2095);
			28697: out = 16'(596);
			28698: out = 16'(3031);
			28699: out = 16'(4144);
			28700: out = 16'(-559);
			28701: out = 16'(-3912);
			28702: out = 16'(-1746);
			28703: out = 16'(2721);
			28704: out = 16'(1843);
			28705: out = 16'(-1402);
			28706: out = 16'(-1898);
			28707: out = 16'(-1247);
			28708: out = 16'(-74);
			28709: out = 16'(-256);
			28710: out = 16'(481);
			28711: out = 16'(2589);
			28712: out = 16'(2517);
			28713: out = 16'(-1197);
			28714: out = 16'(-4257);
			28715: out = 16'(74);
			28716: out = 16'(2112);
			28717: out = 16'(2304);
			28718: out = 16'(-1696);
			28719: out = 16'(-5373);
			28720: out = 16'(-3953);
			28721: out = 16'(1488);
			28722: out = 16'(2888);
			28723: out = 16'(-242);
			28724: out = 16'(-138);
			28725: out = 16'(1416);
			28726: out = 16'(97);
			28727: out = 16'(-3924);
			28728: out = 16'(-2035);
			28729: out = 16'(1829);
			28730: out = 16'(4118);
			28731: out = 16'(1785);
			28732: out = 16'(-1148);
			28733: out = 16'(-3506);
			28734: out = 16'(-1881);
			28735: out = 16'(792);
			28736: out = 16'(1723);
			28737: out = 16'(864);
			28738: out = 16'(6);
			28739: out = 16'(111);
			28740: out = 16'(-317);
			28741: out = 16'(-1662);
			28742: out = 16'(-1872);
			28743: out = 16'(1235);
			28744: out = 16'(3271);
			28745: out = 16'(2320);
			28746: out = 16'(-3326);
			28747: out = 16'(-3452);
			28748: out = 16'(628);
			28749: out = 16'(-155);
			28750: out = 16'(-2059);
			28751: out = 16'(-1765);
			28752: out = 16'(589);
			28753: out = 16'(-149);
			28754: out = 16'(184);
			28755: out = 16'(928);
			28756: out = 16'(2092);
			28757: out = 16'(934);
			28758: out = 16'(-336);
			28759: out = 16'(-1176);
			28760: out = 16'(707);
			28761: out = 16'(3836);
			28762: out = 16'(2761);
			28763: out = 16'(1191);
			28764: out = 16'(-1786);
			28765: out = 16'(-2617);
			28766: out = 16'(-2610);
			28767: out = 16'(3696);
			28768: out = 16'(3414);
			28769: out = 16'(-999);
			28770: out = 16'(-4303);
			28771: out = 16'(-371);
			28772: out = 16'(-1335);
			28773: out = 16'(-3968);
			28774: out = 16'(-2252);
			28775: out = 16'(2773);
			28776: out = 16'(1999);
			28777: out = 16'(-846);
			28778: out = 16'(-386);
			28779: out = 16'(-221);
			28780: out = 16'(933);
			28781: out = 16'(1637);
			28782: out = 16'(1305);
			28783: out = 16'(-1818);
			28784: out = 16'(-3546);
			28785: out = 16'(-1112);
			28786: out = 16'(2115);
			28787: out = 16'(-127);
			28788: out = 16'(-1097);
			28789: out = 16'(89);
			28790: out = 16'(2162);
			28791: out = 16'(214);
			28792: out = 16'(-832);
			28793: out = 16'(-1116);
			28794: out = 16'(1530);
			28795: out = 16'(3368);
			28796: out = 16'(2160);
			28797: out = 16'(309);
			28798: out = 16'(-76);
			28799: out = 16'(-245);
			28800: out = 16'(82);
			28801: out = 16'(-2740);
			28802: out = 16'(-2863);
			28803: out = 16'(311);
			28804: out = 16'(3334);
			28805: out = 16'(2398);
			28806: out = 16'(649);
			28807: out = 16'(-189);
			28808: out = 16'(-86);
			28809: out = 16'(922);
			28810: out = 16'(639);
			28811: out = 16'(-786);
			28812: out = 16'(-1545);
			28813: out = 16'(-3609);
			28814: out = 16'(-1130);
			28815: out = 16'(1338);
			28816: out = 16'(1694);
			28817: out = 16'(518);
			28818: out = 16'(197);
			28819: out = 16'(-735);
			28820: out = 16'(-1338);
			28821: out = 16'(-95);
			28822: out = 16'(1520);
			28823: out = 16'(916);
			28824: out = 16'(-62);
			28825: out = 16'(1949);
			28826: out = 16'(3996);
			28827: out = 16'(2398);
			28828: out = 16'(-2071);
			28829: out = 16'(-3989);
			28830: out = 16'(-1045);
			28831: out = 16'(553);
			28832: out = 16'(-2038);
			28833: out = 16'(-4610);
			28834: out = 16'(-584);
			28835: out = 16'(1699);
			28836: out = 16'(728);
			28837: out = 16'(-757);
			28838: out = 16'(-126);
			28839: out = 16'(2890);
			28840: out = 16'(1610);
			28841: out = 16'(-2728);
			28842: out = 16'(-3892);
			28843: out = 16'(-1193);
			28844: out = 16'(1601);
			28845: out = 16'(1154);
			28846: out = 16'(-856);
			28847: out = 16'(-2461);
			28848: out = 16'(-2025);
			28849: out = 16'(-352);
			28850: out = 16'(1376);
			28851: out = 16'(74);
			28852: out = 16'(1546);
			28853: out = 16'(2475);
			28854: out = 16'(1295);
			28855: out = 16'(725);
			28856: out = 16'(-289);
			28857: out = 16'(1317);
			28858: out = 16'(2681);
			28859: out = 16'(1540);
			28860: out = 16'(-3463);
			28861: out = 16'(-4790);
			28862: out = 16'(-2281);
			28863: out = 16'(-303);
			28864: out = 16'(-1554);
			28865: out = 16'(-925);
			28866: out = 16'(1960);
			28867: out = 16'(3163);
			28868: out = 16'(2226);
			28869: out = 16'(-1643);
			28870: out = 16'(-3599);
			28871: out = 16'(-1678);
			28872: out = 16'(3064);
			28873: out = 16'(3711);
			28874: out = 16'(2566);
			28875: out = 16'(1501);
			28876: out = 16'(1065);
			28877: out = 16'(207);
			28878: out = 16'(-1325);
			28879: out = 16'(-3900);
			28880: out = 16'(-6735);
			28881: out = 16'(-3596);
			28882: out = 16'(233);
			28883: out = 16'(2215);
			28884: out = 16'(1799);
			28885: out = 16'(2876);
			28886: out = 16'(1962);
			28887: out = 16'(187);
			28888: out = 16'(-1477);
			28889: out = 16'(-767);
			28890: out = 16'(-222);
			28891: out = 16'(115);
			28892: out = 16'(-49);
			28893: out = 16'(102);
			28894: out = 16'(1162);
			28895: out = 16'(2560);
			28896: out = 16'(2094);
			28897: out = 16'(-968);
			28898: out = 16'(-5120);
			28899: out = 16'(-5975);
			28900: out = 16'(-2890);
			28901: out = 16'(978);
			28902: out = 16'(4136);
			28903: out = 16'(4029);
			28904: out = 16'(2754);
			28905: out = 16'(1367);
			28906: out = 16'(-1105);
			28907: out = 16'(-2909);
			28908: out = 16'(-2827);
			28909: out = 16'(-1093);
			28910: out = 16'(-2105);
			28911: out = 16'(941);
			28912: out = 16'(2114);
			28913: out = 16'(1657);
			28914: out = 16'(1807);
			28915: out = 16'(346);
			28916: out = 16'(-1031);
			28917: out = 16'(-2555);
			28918: out = 16'(-3196);
			28919: out = 16'(-3410);
			28920: out = 16'(-785);
			28921: out = 16'(3343);
			28922: out = 16'(6144);
			28923: out = 16'(1700);
			28924: out = 16'(-224);
			28925: out = 16'(-1274);
			28926: out = 16'(-2494);
			28927: out = 16'(-5776);
			28928: out = 16'(-3543);
			28929: out = 16'(912);
			28930: out = 16'(3656);
			28931: out = 16'(1767);
			28932: out = 16'(1955);
			28933: out = 16'(1502);
			28934: out = 16'(1110);
			28935: out = 16'(597);
			28936: out = 16'(2125);
			28937: out = 16'(1167);
			28938: out = 16'(-861);
			28939: out = 16'(-1932);
			28940: out = 16'(-997);
			28941: out = 16'(171);
			28942: out = 16'(530);
			28943: out = 16'(-16);
			28944: out = 16'(1804);
			28945: out = 16'(-42);
			28946: out = 16'(-550);
			28947: out = 16'(729);
			28948: out = 16'(1014);
			28949: out = 16'(610);
			28950: out = 16'(736);
			28951: out = 16'(2446);
			28952: out = 16'(4469);
			28953: out = 16'(1865);
			28954: out = 16'(-1724);
			28955: out = 16'(-4343);
			28956: out = 16'(-4716);
			28957: out = 16'(-4449);
			28958: out = 16'(-1659);
			28959: out = 16'(960);
			28960: out = 16'(1568);
			28961: out = 16'(169);
			28962: out = 16'(-90);
			28963: out = 16'(-210);
			28964: out = 16'(-872);
			28965: out = 16'(-54);
			28966: out = 16'(196);
			28967: out = 16'(387);
			28968: out = 16'(-363);
			28969: out = 16'(237);
			28970: out = 16'(-2387);
			28971: out = 16'(-1459);
			28972: out = 16'(589);
			28973: out = 16'(1827);
			28974: out = 16'(174);
			28975: out = 16'(-520);
			28976: out = 16'(-3057);
			28977: out = 16'(-5720);
			28978: out = 16'(-1333);
			28979: out = 16'(2666);
			28980: out = 16'(2461);
			28981: out = 16'(-262);
			28982: out = 16'(76);
			28983: out = 16'(1610);
			28984: out = 16'(-178);
			28985: out = 16'(-3573);
			28986: out = 16'(-915);
			28987: out = 16'(1045);
			28988: out = 16'(2101);
			28989: out = 16'(442);
			28990: out = 16'(-1166);
			28991: out = 16'(-1419);
			28992: out = 16'(-838);
			28993: out = 16'(-78);
			28994: out = 16'(1602);
			28995: out = 16'(1706);
			28996: out = 16'(2010);
			28997: out = 16'(1518);
			28998: out = 16'(1201);
			28999: out = 16'(571);
			29000: out = 16'(176);
			29001: out = 16'(-559);
			29002: out = 16'(-543);
			29003: out = 16'(-39);
			29004: out = 16'(1444);
			29005: out = 16'(1809);
			29006: out = 16'(1738);
			29007: out = 16'(1579);
			29008: out = 16'(854);
			29009: out = 16'(-1069);
			29010: out = 16'(-2187);
			29011: out = 16'(-1358);
			29012: out = 16'(-1467);
			29013: out = 16'(-1133);
			29014: out = 16'(143);
			29015: out = 16'(2054);
			29016: out = 16'(2656);
			29017: out = 16'(2824);
			29018: out = 16'(2302);
			29019: out = 16'(1100);
			29020: out = 16'(-240);
			29021: out = 16'(-2976);
			29022: out = 16'(-2647);
			29023: out = 16'(-292);
			29024: out = 16'(-255);
			29025: out = 16'(1485);
			29026: out = 16'(1626);
			29027: out = 16'(1346);
			29028: out = 16'(171);
			29029: out = 16'(1599);
			29030: out = 16'(44);
			29031: out = 16'(-1449);
			29032: out = 16'(-1269);
			29033: out = 16'(1358);
			29034: out = 16'(555);
			29035: out = 16'(-1042);
			29036: out = 16'(-1017);
			29037: out = 16'(2566);
			29038: out = 16'(2739);
			29039: out = 16'(1093);
			29040: out = 16'(-1961);
			29041: out = 16'(-2568);
			29042: out = 16'(-3412);
			29043: out = 16'(-185);
			29044: out = 16'(1413);
			29045: out = 16'(-272);
			29046: out = 16'(-2093);
			29047: out = 16'(64);
			29048: out = 16'(1648);
			29049: out = 16'(-343);
			29050: out = 16'(-5037);
			29051: out = 16'(-2012);
			29052: out = 16'(2471);
			29053: out = 16'(2502);
			29054: out = 16'(-1786);
			29055: out = 16'(-2337);
			29056: out = 16'(-1987);
			29057: out = 16'(-1670);
			29058: out = 16'(726);
			29059: out = 16'(586);
			29060: out = 16'(303);
			29061: out = 16'(-218);
			29062: out = 16'(27);
			29063: out = 16'(-1198);
			29064: out = 16'(-1177);
			29065: out = 16'(-7);
			29066: out = 16'(1155);
			29067: out = 16'(214);
			29068: out = 16'(-1361);
			29069: out = 16'(-1720);
			29070: out = 16'(-648);
			29071: out = 16'(-1947);
			29072: out = 16'(-2862);
			29073: out = 16'(-2156);
			29074: out = 16'(1565);
			29075: out = 16'(4557);
			29076: out = 16'(3114);
			29077: out = 16'(-973);
			29078: out = 16'(-2019);
			29079: out = 16'(722);
			29080: out = 16'(4064);
			29081: out = 16'(1469);
			29082: out = 16'(-2864);
			29083: out = 16'(-3508);
			29084: out = 16'(1016);
			29085: out = 16'(1946);
			29086: out = 16'(120);
			29087: out = 16'(-1328);
			29088: out = 16'(-793);
			29089: out = 16'(-144);
			29090: out = 16'(575);
			29091: out = 16'(1408);
			29092: out = 16'(1766);
			29093: out = 16'(450);
			29094: out = 16'(51);
			29095: out = 16'(536);
			29096: out = 16'(-154);
			29097: out = 16'(-540);
			29098: out = 16'(-965);
			29099: out = 16'(-341);
			29100: out = 16'(564);
			29101: out = 16'(-579);
			29102: out = 16'(200);
			29103: out = 16'(2053);
			29104: out = 16'(2300);
			29105: out = 16'(-1559);
			29106: out = 16'(-2491);
			29107: out = 16'(-988);
			29108: out = 16'(-344);
			29109: out = 16'(-2383);
			29110: out = 16'(-1107);
			29111: out = 16'(2736);
			29112: out = 16'(4494);
			29113: out = 16'(1659);
			29114: out = 16'(-449);
			29115: out = 16'(-475);
			29116: out = 16'(-484);
			29117: out = 16'(-2197);
			29118: out = 16'(-4495);
			29119: out = 16'(-1900);
			29120: out = 16'(1547);
			29121: out = 16'(1720);
			29122: out = 16'(3391);
			29123: out = 16'(3368);
			29124: out = 16'(2236);
			29125: out = 16'(-898);
			29126: out = 16'(-2362);
			29127: out = 16'(-4536);
			29128: out = 16'(-2915);
			29129: out = 16'(1306);
			29130: out = 16'(4027);
			29131: out = 16'(3097);
			29132: out = 16'(606);
			29133: out = 16'(261);
			29134: out = 16'(651);
			29135: out = 16'(-1128);
			29136: out = 16'(-5564);
			29137: out = 16'(-4862);
			29138: out = 16'(2458);
			29139: out = 16'(3131);
			29140: out = 16'(1330);
			29141: out = 16'(-662);
			29142: out = 16'(370);
			29143: out = 16'(1435);
			29144: out = 16'(-656);
			29145: out = 16'(-2988);
			29146: out = 16'(-1948);
			29147: out = 16'(322);
			29148: out = 16'(457);
			29149: out = 16'(-678);
			29150: out = 16'(-120);
			29151: out = 16'(1652);
			29152: out = 16'(2427);
			29153: out = 16'(-84);
			29154: out = 16'(-2619);
			29155: out = 16'(-1724);
			29156: out = 16'(-1160);
			29157: out = 16'(-771);
			29158: out = 16'(-2336);
			29159: out = 16'(-2819);
			29160: out = 16'(-348);
			29161: out = 16'(2841);
			29162: out = 16'(2355);
			29163: out = 16'(-756);
			29164: out = 16'(-3791);
			29165: out = 16'(-1020);
			29166: out = 16'(311);
			29167: out = 16'(-1283);
			29168: out = 16'(-2214);
			29169: out = 16'(891);
			29170: out = 16'(3073);
			29171: out = 16'(2137);
			29172: out = 16'(100);
			29173: out = 16'(-40);
			29174: out = 16'(907);
			29175: out = 16'(799);
			29176: out = 16'(-878);
			29177: out = 16'(50);
			29178: out = 16'(-580);
			29179: out = 16'(-366);
			29180: out = 16'(312);
			29181: out = 16'(1851);
			29182: out = 16'(502);
			29183: out = 16'(130);
			29184: out = 16'(485);
			29185: out = 16'(85);
			29186: out = 16'(355);
			29187: out = 16'(2055);
			29188: out = 16'(3617);
			29189: out = 16'(2998);
			29190: out = 16'(460);
			29191: out = 16'(-1180);
			29192: out = 16'(-1413);
			29193: out = 16'(-853);
			29194: out = 16'(-1537);
			29195: out = 16'(-949);
			29196: out = 16'(-1283);
			29197: out = 16'(-1720);
			29198: out = 16'(1016);
			29199: out = 16'(2940);
			29200: out = 16'(2141);
			29201: out = 16'(-703);
			29202: out = 16'(-580);
			29203: out = 16'(-2044);
			29204: out = 16'(-2025);
			29205: out = 16'(-1940);
			29206: out = 16'(-429);
			29207: out = 16'(623);
			29208: out = 16'(2852);
			29209: out = 16'(2457);
			29210: out = 16'(-399);
			29211: out = 16'(-2473);
			29212: out = 16'(-2422);
			29213: out = 16'(-1563);
			29214: out = 16'(-436);
			29215: out = 16'(-164);
			29216: out = 16'(2663);
			29217: out = 16'(2327);
			29218: out = 16'(-914);
			29219: out = 16'(-3148);
			29220: out = 16'(-1033);
			29221: out = 16'(34);
			29222: out = 16'(-1160);
			29223: out = 16'(-973);
			29224: out = 16'(584);
			29225: out = 16'(2826);
			29226: out = 16'(3197);
			29227: out = 16'(2123);
			29228: out = 16'(227);
			29229: out = 16'(-192);
			29230: out = 16'(9);
			29231: out = 16'(-243);
			29232: out = 16'(-1277);
			29233: out = 16'(-1238);
			29234: out = 16'(325);
			29235: out = 16'(2082);
			29236: out = 16'(3284);
			29237: out = 16'(2046);
			29238: out = 16'(1471);
			29239: out = 16'(1266);
			29240: out = 16'(-382);
			29241: out = 16'(-2844);
			29242: out = 16'(-3586);
			29243: out = 16'(-1885);
			29244: out = 16'(77);
			29245: out = 16'(2458);
			29246: out = 16'(3718);
			29247: out = 16'(3997);
			29248: out = 16'(1871);
			29249: out = 16'(-954);
			29250: out = 16'(-4401);
			29251: out = 16'(-3051);
			29252: out = 16'(870);
			29253: out = 16'(-324);
			29254: out = 16'(-583);
			29255: out = 16'(-741);
			29256: out = 16'(272);
			29257: out = 16'(957);
			29258: out = 16'(1552);
			29259: out = 16'(1576);
			29260: out = 16'(1341);
			29261: out = 16'(137);
			29262: out = 16'(-1149);
			29263: out = 16'(-3014);
			29264: out = 16'(-2587);
			29265: out = 16'(801);
			29266: out = 16'(745);
			29267: out = 16'(916);
			29268: out = 16'(-683);
			29269: out = 16'(-1244);
			29270: out = 16'(-423);
			29271: out = 16'(348);
			29272: out = 16'(-2344);
			29273: out = 16'(-4287);
			29274: out = 16'(-113);
			29275: out = 16'(2839);
			29276: out = 16'(1888);
			29277: out = 16'(-660);
			29278: out = 16'(155);
			29279: out = 16'(-136);
			29280: out = 16'(-1731);
			29281: out = 16'(-3965);
			29282: out = 16'(-2744);
			29283: out = 16'(-586);
			29284: out = 16'(955);
			29285: out = 16'(-44);
			29286: out = 16'(-393);
			29287: out = 16'(-204);
			29288: out = 16'(1741);
			29289: out = 16'(-194);
			29290: out = 16'(-3738);
			29291: out = 16'(-3017);
			29292: out = 16'(-730);
			29293: out = 16'(601);
			29294: out = 16'(-46);
			29295: out = 16'(403);
			29296: out = 16'(-610);
			29297: out = 16'(-26);
			29298: out = 16'(192);
			29299: out = 16'(315);
			29300: out = 16'(16);
			29301: out = 16'(2033);
			29302: out = 16'(2791);
			29303: out = 16'(757);
			29304: out = 16'(-338);
			29305: out = 16'(-2200);
			29306: out = 16'(-2403);
			29307: out = 16'(-1907);
			29308: out = 16'(-2423);
			29309: out = 16'(-739);
			29310: out = 16'(1992);
			29311: out = 16'(3886);
			29312: out = 16'(3344);
			29313: out = 16'(803);
			29314: out = 16'(-770);
			29315: out = 16'(-278);
			29316: out = 16'(-25);
			29317: out = 16'(287);
			29318: out = 16'(-121);
			29319: out = 16'(466);
			29320: out = 16'(240);
			29321: out = 16'(-260);
			29322: out = 16'(45);
			29323: out = 16'(3876);
			29324: out = 16'(5391);
			29325: out = 16'(513);
			29326: out = 16'(-6704);
			29327: out = 16'(-5233);
			29328: out = 16'(2486);
			29329: out = 16'(3874);
			29330: out = 16'(2704);
			29331: out = 16'(1276);
			29332: out = 16'(1669);
			29333: out = 16'(-541);
			29334: out = 16'(-314);
			29335: out = 16'(-2328);
			29336: out = 16'(-1844);
			29337: out = 16'(553);
			29338: out = 16'(40);
			29339: out = 16'(196);
			29340: out = 16'(1675);
			29341: out = 16'(3157);
			29342: out = 16'(-74);
			29343: out = 16'(-1883);
			29344: out = 16'(-2990);
			29345: out = 16'(-1099);
			29346: out = 16'(707);
			29347: out = 16'(1327);
			29348: out = 16'(-1923);
			29349: out = 16'(-1975);
			29350: out = 16'(3410);
			29351: out = 16'(5023);
			29352: out = 16'(-738);
			29353: out = 16'(-7093);
			29354: out = 16'(-5999);
			29355: out = 16'(-485);
			29356: out = 16'(997);
			29357: out = 16'(-438);
			29358: out = 16'(662);
			29359: out = 16'(814);
			29360: out = 16'(2152);
			29361: out = 16'(123);
			29362: out = 16'(-2106);
			29363: out = 16'(-1946);
			29364: out = 16'(1026);
			29365: out = 16'(1632);
			29366: out = 16'(-196);
			29367: out = 16'(-1706);
			29368: out = 16'(1006);
			29369: out = 16'(2590);
			29370: out = 16'(1579);
			29371: out = 16'(1);
			29372: out = 16'(-1882);
			29373: out = 16'(-577);
			29374: out = 16'(1033);
			29375: out = 16'(1037);
			29376: out = 16'(157);
			29377: out = 16'(-855);
			29378: out = 16'(-2232);
			29379: out = 16'(-3023);
			29380: out = 16'(86);
			29381: out = 16'(84);
			29382: out = 16'(137);
			29383: out = 16'(28);
			29384: out = 16'(107);
			29385: out = 16'(-1547);
			29386: out = 16'(-1151);
			29387: out = 16'(1262);
			29388: out = 16'(3249);
			29389: out = 16'(716);
			29390: out = 16'(-2649);
			29391: out = 16'(-3347);
			29392: out = 16'(-94);
			29393: out = 16'(-175);
			29394: out = 16'(1535);
			29395: out = 16'(1715);
			29396: out = 16'(1130);
			29397: out = 16'(-716);
			29398: out = 16'(-535);
			29399: out = 16'(-1125);
			29400: out = 16'(-903);
			29401: out = 16'(-88);
			29402: out = 16'(1878);
			29403: out = 16'(-324);
			29404: out = 16'(-2588);
			29405: out = 16'(-270);
			29406: out = 16'(3722);
			29407: out = 16'(3114);
			29408: out = 16'(289);
			29409: out = 16'(351);
			29410: out = 16'(1375);
			29411: out = 16'(536);
			29412: out = 16'(-1984);
			29413: out = 16'(-2350);
			29414: out = 16'(-1100);
			29415: out = 16'(1279);
			29416: out = 16'(1631);
			29417: out = 16'(975);
			29418: out = 16'(-51);
			29419: out = 16'(1367);
			29420: out = 16'(1100);
			29421: out = 16'(-759);
			29422: out = 16'(-1872);
			29423: out = 16'(-1212);
			29424: out = 16'(767);
			29425: out = 16'(2322);
			29426: out = 16'(3313);
			29427: out = 16'(1246);
			29428: out = 16'(1084);
			29429: out = 16'(438);
			29430: out = 16'(-1230);
			29431: out = 16'(-2726);
			29432: out = 16'(-1052);
			29433: out = 16'(258);
			29434: out = 16'(-300);
			29435: out = 16'(125);
			29436: out = 16'(997);
			29437: out = 16'(2533);
			29438: out = 16'(1932);
			29439: out = 16'(-923);
			29440: out = 16'(-3197);
			29441: out = 16'(-2291);
			29442: out = 16'(-287);
			29443: out = 16'(-154);
			29444: out = 16'(537);
			29445: out = 16'(1134);
			29446: out = 16'(1771);
			29447: out = 16'(593);
			29448: out = 16'(-418);
			29449: out = 16'(-3889);
			29450: out = 16'(-3231);
			29451: out = 16'(1305);
			29452: out = 16'(1293);
			29453: out = 16'(754);
			29454: out = 16'(-1618);
			29455: out = 16'(-1192);
			29456: out = 16'(1452);
			29457: out = 16'(2212);
			29458: out = 16'(-1790);
			29459: out = 16'(-5037);
			29460: out = 16'(-2944);
			29461: out = 16'(-453);
			29462: out = 16'(-77);
			29463: out = 16'(-668);
			29464: out = 16'(492);
			29465: out = 16'(1610);
			29466: out = 16'(919);
			29467: out = 16'(-297);
			29468: out = 16'(563);
			29469: out = 16'(1510);
			29470: out = 16'(3);
			29471: out = 16'(-3343);
			29472: out = 16'(-3754);
			29473: out = 16'(55);
			29474: out = 16'(1849);
			29475: out = 16'(646);
			29476: out = 16'(-647);
			29477: out = 16'(351);
			29478: out = 16'(3084);
			29479: out = 16'(1190);
			29480: out = 16'(-3150);
			29481: out = 16'(-5053);
			29482: out = 16'(-4271);
			29483: out = 16'(-1075);
			29484: out = 16'(1182);
			29485: out = 16'(2100);
			29486: out = 16'(1927);
			29487: out = 16'(2045);
			29488: out = 16'(969);
			29489: out = 16'(-1451);
			29490: out = 16'(-3642);
			29491: out = 16'(-1683);
			29492: out = 16'(1976);
			29493: out = 16'(3133);
			29494: out = 16'(-17);
			29495: out = 16'(58);
			29496: out = 16'(953);
			29497: out = 16'(2255);
			29498: out = 16'(1299);
			29499: out = 16'(-2396);
			29500: out = 16'(-3922);
			29501: out = 16'(-733);
			29502: out = 16'(3185);
			29503: out = 16'(1458);
			29504: out = 16'(-87);
			29505: out = 16'(-383);
			29506: out = 16'(163);
			29507: out = 16'(-586);
			29508: out = 16'(-1625);
			29509: out = 16'(-1050);
			29510: out = 16'(322);
			29511: out = 16'(-40);
			29512: out = 16'(274);
			29513: out = 16'(959);
			29514: out = 16'(2983);
			29515: out = 16'(4780);
			29516: out = 16'(1735);
			29517: out = 16'(-783);
			29518: out = 16'(-2748);
			29519: out = 16'(-3644);
			29520: out = 16'(-2543);
			29521: out = 16'(-1107);
			29522: out = 16'(253);
			29523: out = 16'(1757);
			29524: out = 16'(2621);
			29525: out = 16'(1256);
			29526: out = 16'(-2596);
			29527: out = 16'(-4804);
			29528: out = 16'(-2252);
			29529: out = 16'(-762);
			29530: out = 16'(-156);
			29531: out = 16'(1523);
			29532: out = 16'(4759);
			29533: out = 16'(2471);
			29534: out = 16'(-1607);
			29535: out = 16'(-3481);
			29536: out = 16'(-466);
			29537: out = 16'(1451);
			29538: out = 16'(1102);
			29539: out = 16'(-256);
			29540: out = 16'(812);
			29541: out = 16'(2469);
			29542: out = 16'(3225);
			29543: out = 16'(940);
			29544: out = 16'(-1949);
			29545: out = 16'(-3673);
			29546: out = 16'(-2263);
			29547: out = 16'(-720);
			29548: out = 16'(884);
			29549: out = 16'(2364);
			29550: out = 16'(3355);
			29551: out = 16'(1234);
			29552: out = 16'(-1637);
			29553: out = 16'(-2004);
			29554: out = 16'(1215);
			29555: out = 16'(1555);
			29556: out = 16'(-941);
			29557: out = 16'(-2958);
			29558: out = 16'(-1346);
			29559: out = 16'(1024);
			29560: out = 16'(2235);
			29561: out = 16'(1966);
			29562: out = 16'(72);
			29563: out = 16'(944);
			29564: out = 16'(775);
			29565: out = 16'(-586);
			29566: out = 16'(-2423);
			29567: out = 16'(-53);
			29568: out = 16'(1122);
			29569: out = 16'(913);
			29570: out = 16'(-14);
			29571: out = 16'(649);
			29572: out = 16'(160);
			29573: out = 16'(253);
			29574: out = 16'(19);
			29575: out = 16'(-3326);
			29576: out = 16'(-4291);
			29577: out = 16'(-981);
			29578: out = 16'(3464);
			29579: out = 16'(3116);
			29580: out = 16'(522);
			29581: out = 16'(-1141);
			29582: out = 16'(-253);
			29583: out = 16'(-188);
			29584: out = 16'(-1751);
			29585: out = 16'(-2675);
			29586: out = 16'(-411);
			29587: out = 16'(2202);
			29588: out = 16'(2126);
			29589: out = 16'(-218);
			29590: out = 16'(-1234);
			29591: out = 16'(-431);
			29592: out = 16'(1715);
			29593: out = 16'(-965);
			29594: out = 16'(-2516);
			29595: out = 16'(-487);
			29596: out = 16'(923);
			29597: out = 16'(1111);
			29598: out = 16'(159);
			29599: out = 16'(538);
			29600: out = 16'(1590);
			29601: out = 16'(1978);
			29602: out = 16'(-87);
			29603: out = 16'(-2540);
			29604: out = 16'(-2920);
			29605: out = 16'(-1607);
			29606: out = 16'(-56);
			29607: out = 16'(1177);
			29608: out = 16'(2431);
			29609: out = 16'(1656);
			29610: out = 16'(1848);
			29611: out = 16'(1044);
			29612: out = 16'(-268);
			29613: out = 16'(-1881);
			29614: out = 16'(-1842);
			29615: out = 16'(-2202);
			29616: out = 16'(-1989);
			29617: out = 16'(110);
			29618: out = 16'(2339);
			29619: out = 16'(1785);
			29620: out = 16'(-892);
			29621: out = 16'(-2291);
			29622: out = 16'(-3181);
			29623: out = 16'(-1334);
			29624: out = 16'(1396);
			29625: out = 16'(3427);
			29626: out = 16'(3363);
			29627: out = 16'(1654);
			29628: out = 16'(-640);
			29629: out = 16'(-1720);
			29630: out = 16'(334);
			29631: out = 16'(285);
			29632: out = 16'(-107);
			29633: out = 16'(48);
			29634: out = 16'(444);
			29635: out = 16'(1427);
			29636: out = 16'(1774);
			29637: out = 16'(1283);
			29638: out = 16'(-82);
			29639: out = 16'(423);
			29640: out = 16'(-17);
			29641: out = 16'(-1743);
			29642: out = 16'(-3910);
			29643: out = 16'(-3283);
			29644: out = 16'(-961);
			29645: out = 16'(2004);
			29646: out = 16'(3070);
			29647: out = 16'(1958);
			29648: out = 16'(-52);
			29649: out = 16'(-1663);
			29650: out = 16'(-3791);
			29651: out = 16'(-4644);
			29652: out = 16'(-6040);
			29653: out = 16'(-1919);
			29654: out = 16'(3793);
			29655: out = 16'(5041);
			29656: out = 16'(3492);
			29657: out = 16'(1862);
			29658: out = 16'(405);
			29659: out = 16'(-1973);
			29660: out = 16'(-1872);
			29661: out = 16'(-364);
			29662: out = 16'(1285);
			29663: out = 16'(1764);
			29664: out = 16'(1707);
			29665: out = 16'(1538);
			29666: out = 16'(-238);
			29667: out = 16'(-2796);
			29668: out = 16'(-2424);
			29669: out = 16'(-240);
			29670: out = 16'(766);
			29671: out = 16'(-155);
			29672: out = 16'(336);
			29673: out = 16'(1967);
			29674: out = 16'(3477);
			29675: out = 16'(2131);
			29676: out = 16'(-714);
			29677: out = 16'(181);
			29678: out = 16'(781);
			29679: out = 16'(-851);
			29680: out = 16'(-3074);
			29681: out = 16'(-25);
			29682: out = 16'(2141);
			29683: out = 16'(2435);
			29684: out = 16'(1185);
			29685: out = 16'(-1260);
			29686: out = 16'(201);
			29687: out = 16'(1405);
			29688: out = 16'(51);
			29689: out = 16'(-4414);
			29690: out = 16'(-2686);
			29691: out = 16'(-1057);
			29692: out = 16'(-519);
			29693: out = 16'(357);
			29694: out = 16'(3790);
			29695: out = 16'(4438);
			29696: out = 16'(1189);
			29697: out = 16'(-2956);
			29698: out = 16'(-7598);
			29699: out = 16'(-3624);
			29700: out = 16'(2733);
			29701: out = 16'(4137);
			29702: out = 16'(2262);
			29703: out = 16'(290);
			29704: out = 16'(2453);
			29705: out = 16'(4112);
			29706: out = 16'(1052);
			29707: out = 16'(-4890);
			29708: out = 16'(-6173);
			29709: out = 16'(-2487);
			29710: out = 16'(-375);
			29711: out = 16'(-225);
			29712: out = 16'(-1292);
			29713: out = 16'(-343);
			29714: out = 16'(1899);
			29715: out = 16'(1733);
			29716: out = 16'(848);
			29717: out = 16'(-764);
			29718: out = 16'(-1881);
			29719: out = 16'(-2523);
			29720: out = 16'(-420);
			29721: out = 16'(1249);
			29722: out = 16'(2227);
			29723: out = 16'(4513);
			29724: out = 16'(2707);
			29725: out = 16'(-652);
			29726: out = 16'(-2597);
			29727: out = 16'(-1300);
			29728: out = 16'(194);
			29729: out = 16'(-668);
			29730: out = 16'(-1956);
			29731: out = 16'(-194);
			29732: out = 16'(2549);
			29733: out = 16'(3437);
			29734: out = 16'(882);
			29735: out = 16'(-2764);
			29736: out = 16'(-1374);
			29737: out = 16'(-958);
			29738: out = 16'(-423);
			29739: out = 16'(69);
			29740: out = 16'(1723);
			29741: out = 16'(1209);
			29742: out = 16'(766);
			29743: out = 16'(-853);
			29744: out = 16'(-2949);
			29745: out = 16'(-4087);
			29746: out = 16'(-1712);
			29747: out = 16'(-84);
			29748: out = 16'(-1022);
			29749: out = 16'(137);
			29750: out = 16'(3681);
			29751: out = 16'(4047);
			29752: out = 16'(-530);
			29753: out = 16'(-1090);
			29754: out = 16'(-263);
			29755: out = 16'(-252);
			29756: out = 16'(-3236);
			29757: out = 16'(-4672);
			29758: out = 16'(-1780);
			29759: out = 16'(2100);
			29760: out = 16'(2282);
			29761: out = 16'(401);
			29762: out = 16'(-124);
			29763: out = 16'(675);
			29764: out = 16'(274);
			29765: out = 16'(-402);
			29766: out = 16'(-1398);
			29767: out = 16'(1422);
			29768: out = 16'(3775);
			29769: out = 16'(2734);
			29770: out = 16'(-1178);
			29771: out = 16'(-1639);
			29772: out = 16'(531);
			29773: out = 16'(1315);
			29774: out = 16'(-1528);
			29775: out = 16'(-1829);
			29776: out = 16'(179);
			29777: out = 16'(1706);
			29778: out = 16'(642);
			29779: out = 16'(1263);
			29780: out = 16'(2579);
			29781: out = 16'(2692);
			29782: out = 16'(190);
			29783: out = 16'(-5690);
			29784: out = 16'(-7197);
			29785: out = 16'(-1989);
			29786: out = 16'(4413);
			29787: out = 16'(5664);
			29788: out = 16'(2274);
			29789: out = 16'(-1579);
			29790: out = 16'(-2971);
			29791: out = 16'(-212);
			29792: out = 16'(-365);
			29793: out = 16'(-431);
			29794: out = 16'(774);
			29795: out = 16'(1014);
			29796: out = 16'(415);
			29797: out = 16'(-244);
			29798: out = 16'(339);
			29799: out = 16'(995);
			29800: out = 16'(2511);
			29801: out = 16'(1380);
			29802: out = 16'(-1136);
			29803: out = 16'(-3071);
			29804: out = 16'(-646);
			29805: out = 16'(1216);
			29806: out = 16'(1037);
			29807: out = 16'(-1000);
			29808: out = 16'(-667);
			29809: out = 16'(-396);
			29810: out = 16'(130);
			29811: out = 16'(-51);
			29812: out = 16'(1740);
			29813: out = 16'(250);
			29814: out = 16'(-52);
			29815: out = 16'(-237);
			29816: out = 16'(162);
			29817: out = 16'(353);
			29818: out = 16'(2592);
			29819: out = 16'(1456);
			29820: out = 16'(-3951);
			29821: out = 16'(-6072);
			29822: out = 16'(-1615);
			29823: out = 16'(2007);
			29824: out = 16'(-629);
			29825: out = 16'(-4396);
			29826: out = 16'(-2414);
			29827: out = 16'(1278);
			29828: out = 16'(800);
			29829: out = 16'(461);
			29830: out = 16'(-124);
			29831: out = 16'(314);
			29832: out = 16'(-208);
			29833: out = 16'(-1079);
			29834: out = 16'(-422);
			29835: out = 16'(-31);
			29836: out = 16'(-1014);
			29837: out = 16'(-1561);
			29838: out = 16'(-305);
			29839: out = 16'(468);
			29840: out = 16'(-734);
			29841: out = 16'(-2159);
			29842: out = 16'(-915);
			29843: out = 16'(1475);
			29844: out = 16'(2306);
			29845: out = 16'(976);
			29846: out = 16'(320);
			29847: out = 16'(-866);
			29848: out = 16'(-901);
			29849: out = 16'(562);
			29850: out = 16'(2637);
			29851: out = 16'(2297);
			29852: out = 16'(-6);
			29853: out = 16'(-2091);
			29854: out = 16'(-1117);
			29855: out = 16'(-220);
			29856: out = 16'(-323);
			29857: out = 16'(-1617);
			29858: out = 16'(-723);
			29859: out = 16'(1006);
			29860: out = 16'(4030);
			29861: out = 16'(3780);
			29862: out = 16'(1601);
			29863: out = 16'(1914);
			29864: out = 16'(3073);
			29865: out = 16'(1584);
			29866: out = 16'(-1067);
			29867: out = 16'(-248);
			29868: out = 16'(2328);
			29869: out = 16'(1422);
			29870: out = 16'(-2694);
			29871: out = 16'(-4190);
			29872: out = 16'(1064);
			29873: out = 16'(4796);
			29874: out = 16'(2474);
			29875: out = 16'(-2761);
			29876: out = 16'(-1443);
			29877: out = 16'(-183);
			29878: out = 16'(-1021);
			29879: out = 16'(-2674);
			29880: out = 16'(-1132);
			29881: out = 16'(844);
			29882: out = 16'(1242);
			29883: out = 16'(-886);
			29884: out = 16'(-3506);
			29885: out = 16'(-1769);
			29886: out = 16'(2675);
			29887: out = 16'(3606);
			29888: out = 16'(-1239);
			29889: out = 16'(-4291);
			29890: out = 16'(-1655);
			29891: out = 16'(2147);
			29892: out = 16'(122);
			29893: out = 16'(139);
			29894: out = 16'(1316);
			29895: out = 16'(3861);
			29896: out = 16'(2254);
			29897: out = 16'(1173);
			29898: out = 16'(-3486);
			29899: out = 16'(-3885);
			29900: out = 16'(-1856);
			29901: out = 16'(131);
			29902: out = 16'(-3006);
			29903: out = 16'(-2587);
			29904: out = 16'(558);
			29905: out = 16'(2223);
			29906: out = 16'(-2505);
			29907: out = 16'(-2291);
			29908: out = 16'(2001);
			29909: out = 16'(3393);
			29910: out = 16'(-289);
			29911: out = 16'(-1148);
			29912: out = 16'(148);
			29913: out = 16'(-987);
			29914: out = 16'(178);
			29915: out = 16'(-467);
			29916: out = 16'(-924);
			29917: out = 16'(-1027);
			29918: out = 16'(1511);
			29919: out = 16'(871);
			29920: out = 16'(-1980);
			29921: out = 16'(-4178);
			29922: out = 16'(-613);
			29923: out = 16'(2440);
			29924: out = 16'(2751);
			29925: out = 16'(553);
			29926: out = 16'(770);
			29927: out = 16'(299);
			29928: out = 16'(290);
			29929: out = 16'(-1938);
			29930: out = 16'(-3438);
			29931: out = 16'(-1467);
			29932: out = 16'(2837);
			29933: out = 16'(3709);
			29934: out = 16'(1308);
			29935: out = 16'(-565);
			29936: out = 16'(88);
			29937: out = 16'(-515);
			29938: out = 16'(-3074);
			29939: out = 16'(-4184);
			29940: out = 16'(-29);
			29941: out = 16'(3010);
			29942: out = 16'(2026);
			29943: out = 16'(186);
			29944: out = 16'(1998);
			29945: out = 16'(2725);
			29946: out = 16'(373);
			29947: out = 16'(-1878);
			29948: out = 16'(-5585);
			29949: out = 16'(-2950);
			29950: out = 16'(712);
			29951: out = 16'(1789);
			29952: out = 16'(1782);
			29953: out = 16'(2721);
			29954: out = 16'(2927);
			29955: out = 16'(1029);
			29956: out = 16'(-425);
			29957: out = 16'(-744);
			29958: out = 16'(1487);
			29959: out = 16'(3095);
			29960: out = 16'(1429);
			29961: out = 16'(271);
			29962: out = 16'(-356);
			29963: out = 16'(77);
			29964: out = 16'(157);
			29965: out = 16'(-602);
			29966: out = 16'(-525);
			29967: out = 16'(1392);
			29968: out = 16'(2873);
			29969: out = 16'(1803);
			29970: out = 16'(-357);
			29971: out = 16'(-235);
			29972: out = 16'(1446);
			29973: out = 16'(-220);
			29974: out = 16'(-1241);
			29975: out = 16'(-1125);
			29976: out = 16'(-141);
			29977: out = 16'(-967);
			29978: out = 16'(-435);
			29979: out = 16'(1330);
			29980: out = 16'(3394);
			29981: out = 16'(2571);
			29982: out = 16'(918);
			29983: out = 16'(-1853);
			29984: out = 16'(-2789);
			29985: out = 16'(-2099);
			29986: out = 16'(-1010);
			29987: out = 16'(-573);
			29988: out = 16'(927);
			29989: out = 16'(3449);
			29990: out = 16'(5418);
			29991: out = 16'(3043);
			29992: out = 16'(-1554);
			29993: out = 16'(-4972);
			29994: out = 16'(-2732);
			29995: out = 16'(-2065);
			29996: out = 16'(-660);
			29997: out = 16'(-377);
			29998: out = 16'(-739);
			29999: out = 16'(-582);
			30000: out = 16'(1010);
			30001: out = 16'(711);
			30002: out = 16'(-1453);
			30003: out = 16'(-1256);
			30004: out = 16'(617);
			30005: out = 16'(-683);
			30006: out = 16'(-4758);
			30007: out = 16'(-3464);
			30008: out = 16'(489);
			30009: out = 16'(1896);
			30010: out = 16'(-781);
			30011: out = 16'(-2263);
			30012: out = 16'(-590);
			30013: out = 16'(450);
			30014: out = 16'(-1670);
			30015: out = 16'(-3454);
			30016: out = 16'(-1044);
			30017: out = 16'(1726);
			30018: out = 16'(2056);
			30019: out = 16'(1698);
			30020: out = 16'(-2010);
			30021: out = 16'(-1992);
			30022: out = 16'(-877);
			30023: out = 16'(-667);
			30024: out = 16'(-555);
			30025: out = 16'(-278);
			30026: out = 16'(143);
			30027: out = 16'(307);
			30028: out = 16'(2292);
			30029: out = 16'(1829);
			30030: out = 16'(2166);
			30031: out = 16'(2521);
			30032: out = 16'(937);
			30033: out = 16'(-2581);
			30034: out = 16'(-5109);
			30035: out = 16'(-3878);
			30036: out = 16'(315);
			30037: out = 16'(2812);
			30038: out = 16'(3522);
			30039: out = 16'(2731);
			30040: out = 16'(1472);
			30041: out = 16'(115);
			30042: out = 16'(-903);
			30043: out = 16'(-1730);
			30044: out = 16'(-1740);
			30045: out = 16'(-148);
			30046: out = 16'(104);
			30047: out = 16'(-138);
			30048: out = 16'(551);
			30049: out = 16'(3070);
			30050: out = 16'(2931);
			30051: out = 16'(1273);
			30052: out = 16'(-540);
			30053: out = 16'(-652);
			30054: out = 16'(947);
			30055: out = 16'(2649);
			30056: out = 16'(2284);
			30057: out = 16'(-459);
			30058: out = 16'(363);
			30059: out = 16'(-1253);
			30060: out = 16'(-2380);
			30061: out = 16'(-1867);
			30062: out = 16'(-1018);
			30063: out = 16'(797);
			30064: out = 16'(2348);
			30065: out = 16'(2925);
			30066: out = 16'(1934);
			30067: out = 16'(380);
			30068: out = 16'(-1308);
			30069: out = 16'(-2092);
			30070: out = 16'(-852);
			30071: out = 16'(-414);
			30072: out = 16'(-46);
			30073: out = 16'(-354);
			30074: out = 16'(-73);
			30075: out = 16'(-1040);
			30076: out = 16'(611);
			30077: out = 16'(1473);
			30078: out = 16'(612);
			30079: out = 16'(-1958);
			30080: out = 16'(101);
			30081: out = 16'(1914);
			30082: out = 16'(915);
			30083: out = 16'(-698);
			30084: out = 16'(-683);
			30085: out = 16'(678);
			30086: out = 16'(1217);
			30087: out = 16'(-342);
			30088: out = 16'(-255);
			30089: out = 16'(-1310);
			30090: out = 16'(-2352);
			30091: out = 16'(-2049);
			30092: out = 16'(-1590);
			30093: out = 16'(-1092);
			30094: out = 16'(-542);
			30095: out = 16'(-95);
			30096: out = 16'(-67);
			30097: out = 16'(141);
			30098: out = 16'(384);
			30099: out = 16'(-614);
			30100: out = 16'(-2207);
			30101: out = 16'(-3192);
			30102: out = 16'(802);
			30103: out = 16'(5594);
			30104: out = 16'(4126);
			30105: out = 16'(-1269);
			30106: out = 16'(-4885);
			30107: out = 16'(-3401);
			30108: out = 16'(-958);
			30109: out = 16'(-427);
			30110: out = 16'(-1615);
			30111: out = 16'(-1328);
			30112: out = 16'(316);
			30113: out = 16'(3035);
			30114: out = 16'(1754);
			30115: out = 16'(-11);
			30116: out = 16'(354);
			30117: out = 16'(1869);
			30118: out = 16'(986);
			30119: out = 16'(-1986);
			30120: out = 16'(-3557);
			30121: out = 16'(-172);
			30122: out = 16'(1686);
			30123: out = 16'(2142);
			30124: out = 16'(1215);
			30125: out = 16'(547);
			30126: out = 16'(-110);
			30127: out = 16'(4);
			30128: out = 16'(-625);
			30129: out = 16'(-2020);
			30130: out = 16'(-1538);
			30131: out = 16'(506);
			30132: out = 16'(1496);
			30133: out = 16'(-490);
			30134: out = 16'(272);
			30135: out = 16'(-68);
			30136: out = 16'(1343);
			30137: out = 16'(803);
			30138: out = 16'(-1539);
			30139: out = 16'(-5449);
			30140: out = 16'(-3336);
			30141: out = 16'(904);
			30142: out = 16'(1616);
			30143: out = 16'(-775);
			30144: out = 16'(151);
			30145: out = 16'(1743);
			30146: out = 16'(-367);
			30147: out = 16'(-2616);
			30148: out = 16'(-1351);
			30149: out = 16'(2135);
			30150: out = 16'(2673);
			30151: out = 16'(-1863);
			30152: out = 16'(-2567);
			30153: out = 16'(-660);
			30154: out = 16'(154);
			30155: out = 16'(-2942);
			30156: out = 16'(-1057);
			30157: out = 16'(999);
			30158: out = 16'(901);
			30159: out = 16'(-492);
			30160: out = 16'(212);
			30161: out = 16'(1089);
			30162: out = 16'(1337);
			30163: out = 16'(1754);
			30164: out = 16'(271);
			30165: out = 16'(-347);
			30166: out = 16'(-1084);
			30167: out = 16'(-1782);
			30168: out = 16'(-741);
			30169: out = 16'(1226);
			30170: out = 16'(3021);
			30171: out = 16'(2813);
			30172: out = 16'(870);
			30173: out = 16'(-626);
			30174: out = 16'(307);
			30175: out = 16'(1591);
			30176: out = 16'(-136);
			30177: out = 16'(-1956);
			30178: out = 16'(-1840);
			30179: out = 16'(1235);
			30180: out = 16'(3407);
			30181: out = 16'(2272);
			30182: out = 16'(-702);
			30183: out = 16'(-2191);
			30184: out = 16'(-2068);
			30185: out = 16'(-2383);
			30186: out = 16'(-2805);
			30187: out = 16'(-715);
			30188: out = 16'(2321);
			30189: out = 16'(1132);
			30190: out = 16'(-856);
			30191: out = 16'(-1901);
			30192: out = 16'(-676);
			30193: out = 16'(466);
			30194: out = 16'(1144);
			30195: out = 16'(608);
			30196: out = 16'(-103);
			30197: out = 16'(120);
			30198: out = 16'(-103);
			30199: out = 16'(236);
			30200: out = 16'(-1260);
			30201: out = 16'(-4206);
			30202: out = 16'(-3731);
			30203: out = 16'(-230);
			30204: out = 16'(2236);
			30205: out = 16'(725);
			30206: out = 16'(-82);
			30207: out = 16'(-437);
			30208: out = 16'(1315);
			30209: out = 16'(1895);
			30210: out = 16'(341);
			30211: out = 16'(-577);
			30212: out = 16'(-50);
			30213: out = 16'(-265);
			30214: out = 16'(-1497);
			30215: out = 16'(-2445);
			30216: out = 16'(465);
			30217: out = 16'(3013);
			30218: out = 16'(1290);
			30219: out = 16'(-1064);
			30220: out = 16'(-1017);
			30221: out = 16'(1085);
			30222: out = 16'(1279);
			30223: out = 16'(-625);
			30224: out = 16'(-1187);
			30225: out = 16'(645);
			30226: out = 16'(1445);
			30227: out = 16'(913);
			30228: out = 16'(-2632);
			30229: out = 16'(-2153);
			30230: out = 16'(1597);
			30231: out = 16'(2803);
			30232: out = 16'(990);
			30233: out = 16'(-1959);
			30234: out = 16'(-2355);
			30235: out = 16'(82);
			30236: out = 16'(-471);
			30237: out = 16'(-254);
			30238: out = 16'(829);
			30239: out = 16'(2187);
			30240: out = 16'(752);
			30241: out = 16'(250);
			30242: out = 16'(0);
			30243: out = 16'(264);
			30244: out = 16'(991);
			30245: out = 16'(913);
			30246: out = 16'(-991);
			30247: out = 16'(-3455);
			30248: out = 16'(-4503);
			30249: out = 16'(-1643);
			30250: out = 16'(1109);
			30251: out = 16'(1499);
			30252: out = 16'(273);
			30253: out = 16'(1401);
			30254: out = 16'(2209);
			30255: out = 16'(1480);
			30256: out = 16'(-803);
			30257: out = 16'(-1479);
			30258: out = 16'(-1251);
			30259: out = 16'(478);
			30260: out = 16'(1583);
			30261: out = 16'(764);
			30262: out = 16'(-898);
			30263: out = 16'(430);
			30264: out = 16'(3470);
			30265: out = 16'(1835);
			30266: out = 16'(1514);
			30267: out = 16'(476);
			30268: out = 16'(553);
			30269: out = 16'(259);
			30270: out = 16'(-236);
			30271: out = 16'(-1683);
			30272: out = 16'(-1021);
			30273: out = 16'(1043);
			30274: out = 16'(1642);
			30275: out = 16'(396);
			30276: out = 16'(-64);
			30277: out = 16'(216);
			30278: out = 16'(67);
			30279: out = 16'(-2712);
			30280: out = 16'(-2666);
			30281: out = 16'(574);
			30282: out = 16'(1903);
			30283: out = 16'(645);
			30284: out = 16'(384);
			30285: out = 16'(1855);
			30286: out = 16'(1281);
			30287: out = 16'(-95);
			30288: out = 16'(-1108);
			30289: out = 16'(-137);
			30290: out = 16'(836);
			30291: out = 16'(-830);
			30292: out = 16'(-788);
			30293: out = 16'(1866);
			30294: out = 16'(3926);
			30295: out = 16'(414);
			30296: out = 16'(-2379);
			30297: out = 16'(-2951);
			30298: out = 16'(-1778);
			30299: out = 16'(-1964);
			30300: out = 16'(-377);
			30301: out = 16'(1646);
			30302: out = 16'(3085);
			30303: out = 16'(2300);
			30304: out = 16'(1356);
			30305: out = 16'(158);
			30306: out = 16'(-399);
			30307: out = 16'(-1563);
			30308: out = 16'(109);
			30309: out = 16'(-9);
			30310: out = 16'(-108);
			30311: out = 16'(-361);
			30312: out = 16'(135);
			30313: out = 16'(-2898);
			30314: out = 16'(-4000);
			30315: out = 16'(-898);
			30316: out = 16'(3860);
			30317: out = 16'(2751);
			30318: out = 16'(-469);
			30319: out = 16'(-2673);
			30320: out = 16'(-1735);
			30321: out = 16'(-730);
			30322: out = 16'(1104);
			30323: out = 16'(649);
			30324: out = 16'(-2330);
			30325: out = 16'(-3291);
			30326: out = 16'(-303);
			30327: out = 16'(1382);
			30328: out = 16'(-886);
			30329: out = 16'(-2845);
			30330: out = 16'(674);
			30331: out = 16'(3252);
			30332: out = 16'(284);
			30333: out = 16'(-718);
			30334: out = 16'(-796);
			30335: out = 16'(462);
			30336: out = 16'(-617);
			30337: out = 16'(-1406);
			30338: out = 16'(-2263);
			30339: out = 16'(59);
			30340: out = 16'(1487);
			30341: out = 16'(14);
			30342: out = 16'(-2450);
			30343: out = 16'(-1999);
			30344: out = 16'(390);
			30345: out = 16'(1553);
			30346: out = 16'(-176);
			30347: out = 16'(-541);
			30348: out = 16'(731);
			30349: out = 16'(1577);
			30350: out = 16'(781);
			30351: out = 16'(1063);
			30352: out = 16'(2406);
			30353: out = 16'(2595);
			30354: out = 16'(132);
			30355: out = 16'(-1953);
			30356: out = 16'(-2117);
			30357: out = 16'(-1000);
			30358: out = 16'(-704);
			30359: out = 16'(191);
			30360: out = 16'(1141);
			30361: out = 16'(1332);
			30362: out = 16'(-253);
			30363: out = 16'(-1960);
			30364: out = 16'(-1762);
			30365: out = 16'(574);
			30366: out = 16'(2029);
			30367: out = 16'(2253);
			30368: out = 16'(819);
			30369: out = 16'(390);
			30370: out = 16'(379);
			30371: out = 16'(594);
			30372: out = 16'(-1778);
			30373: out = 16'(-1944);
			30374: out = 16'(-484);
			30375: out = 16'(-781);
			30376: out = 16'(-1998);
			30377: out = 16'(-1430);
			30378: out = 16'(930);
			30379: out = 16'(1926);
			30380: out = 16'(1872);
			30381: out = 16'(546);
			30382: out = 16'(-113);
			30383: out = 16'(29);
			30384: out = 16'(351);
			30385: out = 16'(190);
			30386: out = 16'(-135);
			30387: out = 16'(204);
			30388: out = 16'(1368);
			30389: out = 16'(1700);
			30390: out = 16'(324);
			30391: out = 16'(-1757);
			30392: out = 16'(-2330);
			30393: out = 16'(71);
			30394: out = 16'(1537);
			30395: out = 16'(-129);
			30396: out = 16'(-3470);
			30397: out = 16'(-1434);
			30398: out = 16'(984);
			30399: out = 16'(1216);
			30400: out = 16'(80);
			30401: out = 16'(1279);
			30402: out = 16'(1844);
			30403: out = 16'(3);
			30404: out = 16'(-3506);
			30405: out = 16'(-4608);
			30406: out = 16'(-1850);
			30407: out = 16'(1403);
			30408: out = 16'(723);
			30409: out = 16'(-3055);
			30410: out = 16'(-3172);
			30411: out = 16'(1044);
			30412: out = 16'(4347);
			30413: out = 16'(2809);
			30414: out = 16'(-2111);
			30415: out = 16'(-3681);
			30416: out = 16'(-726);
			30417: out = 16'(1420);
			30418: out = 16'(766);
			30419: out = 16'(-2360);
			30420: out = 16'(-2553);
			30421: out = 16'(582);
			30422: out = 16'(109);
			30423: out = 16'(1494);
			30424: out = 16'(3509);
			30425: out = 16'(4646);
			30426: out = 16'(1666);
			30427: out = 16'(-1188);
			30428: out = 16'(-2866);
			30429: out = 16'(-1352);
			30430: out = 16'(1521);
			30431: out = 16'(3056);
			30432: out = 16'(1562);
			30433: out = 16'(-375);
			30434: out = 16'(-15);
			30435: out = 16'(-2164);
			30436: out = 16'(-1829);
			30437: out = 16'(-669);
			30438: out = 16'(177);
			30439: out = 16'(540);
			30440: out = 16'(668);
			30441: out = 16'(-171);
			30442: out = 16'(-987);
			30443: out = 16'(1562);
			30444: out = 16'(1317);
			30445: out = 16'(580);
			30446: out = 16'(-73);
			30447: out = 16'(52);
			30448: out = 16'(-974);
			30449: out = 16'(-1068);
			30450: out = 16'(-329);
			30451: out = 16'(-7);
			30452: out = 16'(177);
			30453: out = 16'(-324);
			30454: out = 16'(-765);
			30455: out = 16'(-1184);
			30456: out = 16'(-602);
			30457: out = 16'(722);
			30458: out = 16'(2086);
			30459: out = 16'(1187);
			30460: out = 16'(1041);
			30461: out = 16'(-372);
			30462: out = 16'(2055);
			30463: out = 16'(4039);
			30464: out = 16'(2173);
			30465: out = 16'(-4448);
			30466: out = 16'(-4976);
			30467: out = 16'(-336);
			30468: out = 16'(1768);
			30469: out = 16'(-1356);
			30470: out = 16'(-2235);
			30471: out = 16'(-511);
			30472: out = 16'(-13);
			30473: out = 16'(101);
			30474: out = 16'(1277);
			30475: out = 16'(1781);
			30476: out = 16'(-350);
			30477: out = 16'(241);
			30478: out = 16'(-600);
			30479: out = 16'(-289);
			30480: out = 16'(787);
			30481: out = 16'(2383);
			30482: out = 16'(865);
			30483: out = 16'(-1760);
			30484: out = 16'(-2588);
			30485: out = 16'(458);
			30486: out = 16'(2230);
			30487: out = 16'(1632);
			30488: out = 16'(63);
			30489: out = 16'(26);
			30490: out = 16'(-88);
			30491: out = 16'(-979);
			30492: out = 16'(-2337);
			30493: out = 16'(-1988);
			30494: out = 16'(658);
			30495: out = 16'(1696);
			30496: out = 16'(940);
			30497: out = 16'(-295);
			30498: out = 16'(-1709);
			30499: out = 16'(-2697);
			30500: out = 16'(-2470);
			30501: out = 16'(-333);
			30502: out = 16'(1428);
			30503: out = 16'(2334);
			30504: out = 16'(619);
			30505: out = 16'(-640);
			30506: out = 16'(542);
			30507: out = 16'(1461);
			30508: out = 16'(662);
			30509: out = 16'(-307);
			30510: out = 16'(84);
			30511: out = 16'(-89);
			30512: out = 16'(-66);
			30513: out = 16'(468);
			30514: out = 16'(1458);
			30515: out = 16'(-698);
			30516: out = 16'(-790);
			30517: out = 16'(-278);
			30518: out = 16'(805);
			30519: out = 16'(1386);
			30520: out = 16'(1269);
			30521: out = 16'(-215);
			30522: out = 16'(-1337);
			30523: out = 16'(159);
			30524: out = 16'(979);
			30525: out = 16'(2569);
			30526: out = 16'(2237);
			30527: out = 16'(171);
			30528: out = 16'(-774);
			30529: out = 16'(-395);
			30530: out = 16'(-648);
			30531: out = 16'(-2216);
			30532: out = 16'(-2434);
			30533: out = 16'(-293);
			30534: out = 16'(1699);
			30535: out = 16'(693);
			30536: out = 16'(-2205);
			30537: out = 16'(-3271);
			30538: out = 16'(-1576);
			30539: out = 16'(306);
			30540: out = 16'(479);
			30541: out = 16'(-1399);
			30542: out = 16'(-884);
			30543: out = 16'(803);
			30544: out = 16'(-401);
			30545: out = 16'(-708);
			30546: out = 16'(-2057);
			30547: out = 16'(-473);
			30548: out = 16'(1582);
			30549: out = 16'(1892);
			30550: out = 16'(-1700);
			30551: out = 16'(-2251);
			30552: out = 16'(825);
			30553: out = 16'(2856);
			30554: out = 16'(997);
			30555: out = 16'(-636);
			30556: out = 16'(-430);
			30557: out = 16'(414);
			30558: out = 16'(341);
			30559: out = 16'(1077);
			30560: out = 16'(1253);
			30561: out = 16'(-190);
			30562: out = 16'(-2697);
			30563: out = 16'(-1462);
			30564: out = 16'(284);
			30565: out = 16'(-1069);
			30566: out = 16'(-2069);
			30567: out = 16'(-1570);
			30568: out = 16'(351);
			30569: out = 16'(1456);
			30570: out = 16'(4388);
			30571: out = 16'(3382);
			30572: out = 16'(2336);
			30573: out = 16'(884);
			30574: out = 16'(-753);
			30575: out = 16'(-4086);
			30576: out = 16'(-5003);
			30577: out = 16'(-3054);
			30578: out = 16'(289);
			30579: out = 16'(2606);
			30580: out = 16'(3369);
			30581: out = 16'(2072);
			30582: out = 16'(-249);
			30583: out = 16'(-589);
			30584: out = 16'(-2135);
			30585: out = 16'(-3567);
			30586: out = 16'(-3003);
			30587: out = 16'(143);
			30588: out = 16'(1667);
			30589: out = 16'(1114);
			30590: out = 16'(816);
			30591: out = 16'(1401);
			30592: out = 16'(1536);
			30593: out = 16'(-1377);
			30594: out = 16'(-3426);
			30595: out = 16'(-369);
			30596: out = 16'(1232);
			30597: out = 16'(962);
			30598: out = 16'(-144);
			30599: out = 16'(756);
			30600: out = 16'(-88);
			30601: out = 16'(390);
			30602: out = 16'(-109);
			30603: out = 16'(-1457);
			30604: out = 16'(-1664);
			30605: out = 16'(-1927);
			30606: out = 16'(-930);
			30607: out = 16'(401);
			30608: out = 16'(1704);
			30609: out = 16'(1535);
			30610: out = 16'(2068);
			30611: out = 16'(1054);
			30612: out = 16'(-3001);
			30613: out = 16'(-4178);
			30614: out = 16'(-1188);
			30615: out = 16'(2782);
			30616: out = 16'(2667);
			30617: out = 16'(688);
			30618: out = 16'(180);
			30619: out = 16'(2007);
			30620: out = 16'(2081);
			30621: out = 16'(891);
			30622: out = 16'(-2676);
			30623: out = 16'(-3209);
			30624: out = 16'(-1362);
			30625: out = 16'(587);
			30626: out = 16'(-3319);
			30627: out = 16'(-4131);
			30628: out = 16'(-15);
			30629: out = 16'(3314);
			30630: out = 16'(2872);
			30631: out = 16'(948);
			30632: out = 16'(517);
			30633: out = 16'(-327);
			30634: out = 16'(-1603);
			30635: out = 16'(-4249);
			30636: out = 16'(-3299);
			30637: out = 16'(670);
			30638: out = 16'(3071);
			30639: out = 16'(1252);
			30640: out = 16'(328);
			30641: out = 16'(2184);
			30642: out = 16'(2899);
			30643: out = 16'(1457);
			30644: out = 16'(-286);
			30645: out = 16'(-630);
			30646: out = 16'(-730);
			30647: out = 16'(-1074);
			30648: out = 16'(-703);
			30649: out = 16'(612);
			30650: out = 16'(1478);
			30651: out = 16'(374);
			30652: out = 16'(-542);
			30653: out = 16'(-360);
			30654: out = 16'(587);
			30655: out = 16'(1432);
			30656: out = 16'(1108);
			30657: out = 16'(-864);
			30658: out = 16'(-2920);
			30659: out = 16'(1);
			30660: out = 16'(1117);
			30661: out = 16'(2016);
			30662: out = 16'(1712);
			30663: out = 16'(593);
			30664: out = 16'(-976);
			30665: out = 16'(-593);
			30666: out = 16'(1103);
			30667: out = 16'(1672);
			30668: out = 16'(-2369);
			30669: out = 16'(-5724);
			30670: out = 16'(-4501);
			30671: out = 16'(599);
			30672: out = 16'(1897);
			30673: out = 16'(1118);
			30674: out = 16'(-800);
			30675: out = 16'(-790);
			30676: out = 16'(-185);
			30677: out = 16'(1459);
			30678: out = 16'(988);
			30679: out = 16'(441);
			30680: out = 16'(2926);
			30681: out = 16'(2271);
			30682: out = 16'(-729);
			30683: out = 16'(-2961);
			30684: out = 16'(-476);
			30685: out = 16'(-212);
			30686: out = 16'(-595);
			30687: out = 16'(-940);
			30688: out = 16'(1008);
			30689: out = 16'(2553);
			30690: out = 16'(2650);
			30691: out = 16'(-32);
			30692: out = 16'(-2260);
			30693: out = 16'(-1569);
			30694: out = 16'(2130);
			30695: out = 16'(3226);
			30696: out = 16'(785);
			30697: out = 16'(-954);
			30698: out = 16'(-1615);
			30699: out = 16'(72);
			30700: out = 16'(1757);
			30701: out = 16'(1321);
			30702: out = 16'(-87);
			30703: out = 16'(-1679);
			30704: out = 16'(-1319);
			30705: out = 16'(418);
			30706: out = 16'(1483);
			30707: out = 16'(596);
			30708: out = 16'(-210);
			30709: out = 16'(9);
			30710: out = 16'(919);
			30711: out = 16'(306);
			30712: out = 16'(-197);
			30713: out = 16'(-81);
			30714: out = 16'(489);
			30715: out = 16'(-2080);
			30716: out = 16'(-2547);
			30717: out = 16'(-100);
			30718: out = 16'(-343);
			30719: out = 16'(692);
			30720: out = 16'(-225);
			30721: out = 16'(-468);
			30722: out = 16'(379);
			30723: out = 16'(997);
			30724: out = 16'(1227);
			30725: out = 16'(1670);
			30726: out = 16'(1256);
			30727: out = 16'(1658);
			30728: out = 16'(215);
			30729: out = 16'(48);
			30730: out = 16'(167);
			30731: out = 16'(85);
			30732: out = 16'(-3210);
			30733: out = 16'(-3897);
			30734: out = 16'(-2012);
			30735: out = 16'(-672);
			30736: out = 16'(33);
			30737: out = 16'(2722);
			30738: out = 16'(4686);
			30739: out = 16'(2657);
			30740: out = 16'(-2535);
			30741: out = 16'(-3082);
			30742: out = 16'(-495);
			30743: out = 16'(-295);
			30744: out = 16'(524);
			30745: out = 16'(667);
			30746: out = 16'(911);
			30747: out = 16'(25);
			30748: out = 16'(-1206);
			30749: out = 16'(-1421);
			30750: out = 16'(-1521);
			30751: out = 16'(-1656);
			30752: out = 16'(474);
			30753: out = 16'(593);
			30754: out = 16'(-292);
			30755: out = 16'(-1402);
			30756: out = 16'(-579);
			30757: out = 16'(1031);
			30758: out = 16'(1800);
			30759: out = 16'(1006);
			30760: out = 16'(-326);
			30761: out = 16'(-2115);
			30762: out = 16'(-3322);
			30763: out = 16'(-2911);
			30764: out = 16'(-45);
			30765: out = 16'(1700);
			30766: out = 16'(3093);
			30767: out = 16'(2080);
			30768: out = 16'(15);
			30769: out = 16'(-1188);
			30770: out = 16'(-1668);
			30771: out = 16'(-1947);
			30772: out = 16'(-1049);
			30773: out = 16'(2129);
			30774: out = 16'(2202);
			30775: out = 16'(979);
			30776: out = 16'(40);
			30777: out = 16'(1597);
			30778: out = 16'(-1981);
			30779: out = 16'(-2355);
			30780: out = 16'(-1387);
			30781: out = 16'(-691);
			30782: out = 16'(-1143);
			30783: out = 16'(-480);
			30784: out = 16'(778);
			30785: out = 16'(1736);
			30786: out = 16'(2095);
			30787: out = 16'(1678);
			30788: out = 16'(1496);
			30789: out = 16'(1264);
			30790: out = 16'(-168);
			30791: out = 16'(-551);
			30792: out = 16'(-1683);
			30793: out = 16'(-2546);
			30794: out = 16'(-1512);
			30795: out = 16'(2073);
			30796: out = 16'(3654);
			30797: out = 16'(899);
			30798: out = 16'(-3847);
			30799: out = 16'(-2701);
			30800: out = 16'(151);
			30801: out = 16'(1987);
			30802: out = 16'(1233);
			30803: out = 16'(580);
			30804: out = 16'(175);
			30805: out = 16'(519);
			30806: out = 16'(336);
			30807: out = 16'(451);
			30808: out = 16'(982);
			30809: out = 16'(2638);
			30810: out = 16'(2695);
			30811: out = 16'(-482);
			30812: out = 16'(-4119);
			30813: out = 16'(-4599);
			30814: out = 16'(-1779);
			30815: out = 16'(-320);
			30816: out = 16'(-1314);
			30817: out = 16'(-1310);
			30818: out = 16'(2115);
			30819: out = 16'(3512);
			30820: out = 16'(-1517);
			30821: out = 16'(-5943);
			30822: out = 16'(-2411);
			30823: out = 16'(4729);
			30824: out = 16'(5301);
			30825: out = 16'(639);
			30826: out = 16'(-2327);
			30827: out = 16'(-1355);
			30828: out = 16'(-908);
			30829: out = 16'(-1573);
			30830: out = 16'(-534);
			30831: out = 16'(2038);
			30832: out = 16'(2702);
			30833: out = 16'(431);
			30834: out = 16'(-418);
			30835: out = 16'(-21);
			30836: out = 16'(-128);
			30837: out = 16'(353);
			30838: out = 16'(35);
			30839: out = 16'(-174);
			30840: out = 16'(-139);
			30841: out = 16'(-146);
			30842: out = 16'(-421);
			30843: out = 16'(-1691);
			30844: out = 16'(-1977);
			30845: out = 16'(479);
			30846: out = 16'(1862);
			30847: out = 16'(1107);
			30848: out = 16'(-436);
			30849: out = 16'(-521);
			30850: out = 16'(1222);
			30851: out = 16'(778);
			30852: out = 16'(-353);
			30853: out = 16'(135);
			30854: out = 16'(-208);
			30855: out = 16'(59);
			30856: out = 16'(-191);
			30857: out = 16'(-129);
			30858: out = 16'(-785);
			30859: out = 16'(905);
			30860: out = 16'(1579);
			30861: out = 16'(1093);
			30862: out = 16'(-135);
			30863: out = 16'(-949);
			30864: out = 16'(-1925);
			30865: out = 16'(-2220);
			30866: out = 16'(-1542);
			30867: out = 16'(1400);
			30868: out = 16'(1948);
			30869: out = 16'(849);
			30870: out = 16'(37);
			30871: out = 16'(1212);
			30872: out = 16'(705);
			30873: out = 16'(-1467);
			30874: out = 16'(-3377);
			30875: out = 16'(-735);
			30876: out = 16'(-145);
			30877: out = 16'(-126);
			30878: out = 16'(-866);
			30879: out = 16'(-931);
			30880: out = 16'(589);
			30881: out = 16'(3399);
			30882: out = 16'(3629);
			30883: out = 16'(-336);
			30884: out = 16'(-3341);
			30885: out = 16'(-3775);
			30886: out = 16'(-2015);
			30887: out = 16'(-522);
			30888: out = 16'(443);
			30889: out = 16'(1248);
			30890: out = 16'(983);
			30891: out = 16'(-926);
			30892: out = 16'(-915);
			30893: out = 16'(-557);
			30894: out = 16'(1104);
			30895: out = 16'(1728);
			30896: out = 16'(135);
			30897: out = 16'(-601);
			30898: out = 16'(376);
			30899: out = 16'(1457);
			30900: out = 16'(-205);
			30901: out = 16'(-362);
			30902: out = 16'(-576);
			30903: out = 16'(971);
			30904: out = 16'(2504);
			30905: out = 16'(-829);
			30906: out = 16'(-4258);
			30907: out = 16'(-3986);
			30908: out = 16'(143);
			30909: out = 16'(2542);
			30910: out = 16'(2299);
			30911: out = 16'(452);
			30912: out = 16'(-551);
			30913: out = 16'(351);
			30914: out = 16'(825);
			30915: out = 16'(1242);
			30916: out = 16'(1426);
			30917: out = 16'(1392);
			30918: out = 16'(185);
			30919: out = 16'(-181);
			30920: out = 16'(-92);
			30921: out = 16'(-95);
			30922: out = 16'(-660);
			30923: out = 16'(-338);
			30924: out = 16'(-44);
			30925: out = 16'(-23);
			30926: out = 16'(305);
			30927: out = 16'(289);
			30928: out = 16'(-878);
			30929: out = 16'(-1576);
			30930: out = 16'(-295);
			30931: out = 16'(2507);
			30932: out = 16'(2093);
			30933: out = 16'(-867);
			30934: out = 16'(-1580);
			30935: out = 16'(-321);
			30936: out = 16'(1229);
			30937: out = 16'(859);
			30938: out = 16'(-791);
			30939: out = 16'(-1264);
			30940: out = 16'(-699);
			30941: out = 16'(499);
			30942: out = 16'(1225);
			30943: out = 16'(98);
			30944: out = 16'(-1488);
			30945: out = 16'(-826);
			30946: out = 16'(1686);
			30947: out = 16'(1278);
			30948: out = 16'(-1027);
			30949: out = 16'(-2997);
			30950: out = 16'(-1365);
			30951: out = 16'(1055);
			30952: out = 16'(1940);
			30953: out = 16'(-1074);
			30954: out = 16'(-3411);
			30955: out = 16'(-949);
			30956: out = 16'(980);
			30957: out = 16'(984);
			30958: out = 16'(-663);
			30959: out = 16'(-921);
			30960: out = 16'(-344);
			30961: out = 16'(320);
			30962: out = 16'(-1051);
			30963: out = 16'(-2813);
			30964: out = 16'(-2900);
			30965: out = 16'(517);
			30966: out = 16'(2585);
			30967: out = 16'(1298);
			30968: out = 16'(-1388);
			30969: out = 16'(-1829);
			30970: out = 16'(-1653);
			30971: out = 16'(-2726);
			30972: out = 16'(-4020);
			30973: out = 16'(1292);
			30974: out = 16'(5455);
			30975: out = 16'(4249);
			30976: out = 16'(14);
			30977: out = 16'(-225);
			30978: out = 16'(1498);
			30979: out = 16'(469);
			30980: out = 16'(-3580);
			30981: out = 16'(-739);
			30982: out = 16'(901);
			30983: out = 16'(1266);
			30984: out = 16'(-321);
			30985: out = 16'(-345);
			30986: out = 16'(-378);
			30987: out = 16'(1076);
			30988: out = 16'(1975);
			30989: out = 16'(1432);
			30990: out = 16'(656);
			30991: out = 16'(-770);
			30992: out = 16'(-1794);
			30993: out = 16'(-279);
			30994: out = 16'(1272);
			30995: out = 16'(3522);
			30996: out = 16'(3435);
			30997: out = 16'(1435);
			30998: out = 16'(-2072);
			30999: out = 16'(-1808);
			31000: out = 16'(-1415);
			31001: out = 16'(-2905);
			31002: out = 16'(-6159);
			31003: out = 16'(-1193);
			31004: out = 16'(3963);
			31005: out = 16'(3548);
			31006: out = 16'(380);
			31007: out = 16'(-1704);
			31008: out = 16'(-666);
			31009: out = 16'(-332);
			31010: out = 16'(-1572);
			31011: out = 16'(-2379);
			31012: out = 16'(-437);
			31013: out = 16'(442);
			31014: out = 16'(-491);
			31015: out = 16'(-149);
			31016: out = 16'(3092);
			31017: out = 16'(4039);
			31018: out = 16'(408);
			31019: out = 16'(-3948);
			31020: out = 16'(-4587);
			31021: out = 16'(-2356);
			31022: out = 16'(-74);
			31023: out = 16'(542);
			31024: out = 16'(1542);
			31025: out = 16'(1051);
			31026: out = 16'(1040);
			31027: out = 16'(2779);
			31028: out = 16'(870);
			31029: out = 16'(-3688);
			31030: out = 16'(-6167);
			31031: out = 16'(-1815);
			31032: out = 16'(2069);
			31033: out = 16'(2356);
			31034: out = 16'(-1318);
			31035: out = 16'(-2446);
			31036: out = 16'(2228);
			31037: out = 16'(4616);
			31038: out = 16'(1358);
			31039: out = 16'(-3356);
			31040: out = 16'(-3696);
			31041: out = 16'(-934);
			31042: out = 16'(994);
			31043: out = 16'(1231);
			31044: out = 16'(1666);
			31045: out = 16'(1730);
			31046: out = 16'(31);
			31047: out = 16'(-2021);
			31048: out = 16'(-1169);
			31049: out = 16'(1025);
			31050: out = 16'(1798);
			31051: out = 16'(6);
			31052: out = 16'(-1512);
			31053: out = 16'(-1266);
			31054: out = 16'(-9);
			31055: out = 16'(-618);
			31056: out = 16'(-2447);
			31057: out = 16'(-3603);
			31058: out = 16'(351);
			31059: out = 16'(4021);
			31060: out = 16'(3930);
			31061: out = 16'(617);
			31062: out = 16'(828);
			31063: out = 16'(1348);
			31064: out = 16'(9);
			31065: out = 16'(-3391);
			31066: out = 16'(-1933);
			31067: out = 16'(-325);
			31068: out = 16'(1178);
			31069: out = 16'(2083);
			31070: out = 16'(1613);
			31071: out = 16'(943);
			31072: out = 16'(422);
			31073: out = 16'(595);
			31074: out = 16'(-103);
			31075: out = 16'(-143);
			31076: out = 16'(-2172);
			31077: out = 16'(-3585);
			31078: out = 16'(-366);
			31079: out = 16'(2176);
			31080: out = 16'(3345);
			31081: out = 16'(2131);
			31082: out = 16'(39);
			31083: out = 16'(-33);
			31084: out = 16'(-481);
			31085: out = 16'(-1704);
			31086: out = 16'(-1917);
			31087: out = 16'(92);
			31088: out = 16'(2584);
			31089: out = 16'(2927);
			31090: out = 16'(966);
			31091: out = 16'(-417);
			31092: out = 16'(-1926);
			31093: out = 16'(-2348);
			31094: out = 16'(-2219);
			31095: out = 16'(-2185);
			31096: out = 16'(-1779);
			31097: out = 16'(-666);
			31098: out = 16'(1284);
			31099: out = 16'(2864);
			31100: out = 16'(3102);
			31101: out = 16'(1314);
			31102: out = 16'(-709);
			31103: out = 16'(-1756);
			31104: out = 16'(-2695);
			31105: out = 16'(-2618);
			31106: out = 16'(-894);
			31107: out = 16'(2311);
			31108: out = 16'(5381);
			31109: out = 16'(4937);
			31110: out = 16'(2425);
			31111: out = 16'(-138);
			31112: out = 16'(-2279);
			31113: out = 16'(-2780);
			31114: out = 16'(-2937);
			31115: out = 16'(-2402);
			31116: out = 16'(-497);
			31117: out = 16'(1112);
			31118: out = 16'(1762);
			31119: out = 16'(1052);
			31120: out = 16'(161);
			31121: out = 16'(2342);
			31122: out = 16'(2723);
			31123: out = 16'(-82);
			31124: out = 16'(-4191);
			31125: out = 16'(-2926);
			31126: out = 16'(-2004);
			31127: out = 16'(-1723);
			31128: out = 16'(-1737);
			31129: out = 16'(2033);
			31130: out = 16'(2040);
			31131: out = 16'(2103);
			31132: out = 16'(1611);
			31133: out = 16'(33);
			31134: out = 16'(-1726);
			31135: out = 16'(-2445);
			31136: out = 16'(-1556);
			31137: out = 16'(524);
			31138: out = 16'(-883);
			31139: out = 16'(-501);
			31140: out = 16'(464);
			31141: out = 16'(348);
			31142: out = 16'(-1747);
			31143: out = 16'(-1494);
			31144: out = 16'(1075);
			31145: out = 16'(2956);
			31146: out = 16'(2155);
			31147: out = 16'(-896);
			31148: out = 16'(-2452);
			31149: out = 16'(-816);
			31150: out = 16'(1341);
			31151: out = 16'(1808);
			31152: out = 16'(870);
			31153: out = 16'(447);
			31154: out = 16'(-104);
			31155: out = 16'(1862);
			31156: out = 16'(304);
			31157: out = 16'(-1219);
			31158: out = 16'(352);
			31159: out = 16'(1583);
			31160: out = 16'(724);
			31161: out = 16'(-1705);
			31162: out = 16'(-1672);
			31163: out = 16'(977);
			31164: out = 16'(2858);
			31165: out = 16'(1608);
			31166: out = 16'(-181);
			31167: out = 16'(-135);
			31168: out = 16'(1514);
			31169: out = 16'(863);
			31170: out = 16'(-1168);
			31171: out = 16'(-1003);
			31172: out = 16'(1829);
			31173: out = 16'(3242);
			31174: out = 16'(1495);
			31175: out = 16'(-1324);
			31176: out = 16'(-1464);
			31177: out = 16'(-502);
			31178: out = 16'(-374);
			31179: out = 16'(-1316);
			31180: out = 16'(-241);
			31181: out = 16'(169);
			31182: out = 16'(881);
			31183: out = 16'(1153);
			31184: out = 16'(-639);
			31185: out = 16'(-433);
			31186: out = 16'(652);
			31187: out = 16'(1113);
			31188: out = 16'(-822);
			31189: out = 16'(-817);
			31190: out = 16'(-548);
			31191: out = 16'(-221);
			31192: out = 16'(-251);
			31193: out = 16'(1093);
			31194: out = 16'(1432);
			31195: out = 16'(836);
			31196: out = 16'(-230);
			31197: out = 16'(1201);
			31198: out = 16'(-279);
			31199: out = 16'(-2158);
			31200: out = 16'(-2017);
			31201: out = 16'(63);
			31202: out = 16'(1287);
			31203: out = 16'(669);
			31204: out = 16'(-259);
			31205: out = 16'(-208);
			31206: out = 16'(266);
			31207: out = 16'(-752);
			31208: out = 16'(-2321);
			31209: out = 16'(-2807);
			31210: out = 16'(-184);
			31211: out = 16'(742);
			31212: out = 16'(-116);
			31213: out = 16'(-1284);
			31214: out = 16'(-1268);
			31215: out = 16'(303);
			31216: out = 16'(2460);
			31217: out = 16'(2724);
			31218: out = 16'(291);
			31219: out = 16'(-3902);
			31220: out = 16'(-5246);
			31221: out = 16'(-3535);
			31222: out = 16'(-2876);
			31223: out = 16'(-1915);
			31224: out = 16'(152);
			31225: out = 16'(2713);
			31226: out = 16'(2652);
			31227: out = 16'(856);
			31228: out = 16'(-1259);
			31229: out = 16'(-1082);
			31230: out = 16'(439);
			31231: out = 16'(129);
			31232: out = 16'(-1416);
			31233: out = 16'(-1812);
			31234: out = 16'(773);
			31235: out = 16'(3682);
			31236: out = 16'(4671);
			31237: out = 16'(1891);
			31238: out = 16'(-1715);
			31239: out = 16'(-2202);
			31240: out = 16'(-1455);
			31241: out = 16'(-1530);
			31242: out = 16'(-2097);
			31243: out = 16'(-272);
			31244: out = 16'(3123);
			31245: out = 16'(4740);
			31246: out = 16'(2740);
			31247: out = 16'(-145);
			31248: out = 16'(-2246);
			31249: out = 16'(-1034);
			31250: out = 16'(146);
			31251: out = 16'(-270);
			31252: out = 16'(-2145);
			31253: out = 16'(783);
			31254: out = 16'(4470);
			31255: out = 16'(4317);
			31256: out = 16'(175);
			31257: out = 16'(-2592);
			31258: out = 16'(-2250);
			31259: out = 16'(-304);
			31260: out = 16'(259);
			31261: out = 16'(358);
			31262: out = 16'(-4);
			31263: out = 16'(-156);
			31264: out = 16'(-73);
			31265: out = 16'(1070);
			31266: out = 16'(2448);
			31267: out = 16'(2853);
			31268: out = 16'(585);
			31269: out = 16'(-1844);
			31270: out = 16'(-4497);
			31271: out = 16'(-3395);
			31272: out = 16'(-253);
			31273: out = 16'(1324);
			31274: out = 16'(250);
			31275: out = 16'(604);
			31276: out = 16'(1764);
			31277: out = 16'(-264);
			31278: out = 16'(167);
			31279: out = 16'(819);
			31280: out = 16'(1025);
			31281: out = 16'(-972);
			31282: out = 16'(78);
			31283: out = 16'(148);
			31284: out = 16'(-1282);
			31285: out = 16'(-4179);
			31286: out = 16'(-1005);
			31287: out = 16'(621);
			31288: out = 16'(1754);
			31289: out = 16'(700);
			31290: out = 16'(-2431);
			31291: out = 16'(-3486);
			31292: out = 16'(-259);
			31293: out = 16'(3059);
			31294: out = 16'(1277);
			31295: out = 16'(-2181);
			31296: out = 16'(-3523);
			31297: out = 16'(-1193);
			31298: out = 16'(297);
			31299: out = 16'(-107);
			31300: out = 16'(23);
			31301: out = 16'(3210);
			31302: out = 16'(4564);
			31303: out = 16'(1205);
			31304: out = 16'(-6142);
			31305: out = 16'(-8038);
			31306: out = 16'(-2883);
			31307: out = 16'(-183);
			31308: out = 16'(-82);
			31309: out = 16'(373);
			31310: out = 16'(2857);
			31311: out = 16'(4425);
			31312: out = 16'(2869);
			31313: out = 16'(626);
			31314: out = 16'(-1418);
			31315: out = 16'(-3816);
			31316: out = 16'(-4078);
			31317: out = 16'(-1707);
			31318: out = 16'(911);
			31319: out = 16'(1607);
			31320: out = 16'(1148);
			31321: out = 16'(2248);
			31322: out = 16'(2693);
			31323: out = 16'(1116);
			31324: out = 16'(-1432);
			31325: out = 16'(-433);
			31326: out = 16'(342);
			31327: out = 16'(-929);
			31328: out = 16'(-943);
			31329: out = 16'(1892);
			31330: out = 16'(4448);
			31331: out = 16'(3472);
			31332: out = 16'(-44);
			31333: out = 16'(-1567);
			31334: out = 16'(-2153);
			31335: out = 16'(-2292);
			31336: out = 16'(-1552);
			31337: out = 16'(-373);
			31338: out = 16'(1973);
			31339: out = 16'(3968);
			31340: out = 16'(4102);
			31341: out = 16'(2188);
			31342: out = 16'(-83);
			31343: out = 16'(-985);
			31344: out = 16'(-857);
			31345: out = 16'(-773);
			31346: out = 16'(-1653);
			31347: out = 16'(-1119);
			31348: out = 16'(897);
			31349: out = 16'(2597);
			31350: out = 16'(1668);
			31351: out = 16'(1315);
			31352: out = 16'(1776);
			31353: out = 16'(764);
			31354: out = 16'(-5021);
			31355: out = 16'(-8356);
			31356: out = 16'(-5441);
			31357: out = 16'(1157);
			31358: out = 16'(5155);
			31359: out = 16'(4914);
			31360: out = 16'(2856);
			31361: out = 16'(886);
			31362: out = 16'(-1165);
			31363: out = 16'(-3365);
			31364: out = 16'(-4190);
			31365: out = 16'(-3072);
			31366: out = 16'(-1856);
			31367: out = 16'(-4);
			31368: out = 16'(562);
			31369: out = 16'(155);
			31370: out = 16'(-522);
			31371: out = 16'(1438);
			31372: out = 16'(2052);
			31373: out = 16'(318);
			31374: out = 16'(-2300);
			31375: out = 16'(-2423);
			31376: out = 16'(-560);
			31377: out = 16'(350);
			31378: out = 16'(-852);
			31379: out = 16'(-997);
			31380: out = 16'(-432);
			31381: out = 16'(315);
			31382: out = 16'(-402);
			31383: out = 16'(-1927);
			31384: out = 16'(-1337);
			31385: out = 16'(1392);
			31386: out = 16'(2629);
			31387: out = 16'(-32);
			31388: out = 16'(-875);
			31389: out = 16'(-634);
			31390: out = 16'(322);
			31391: out = 16'(-127);
			31392: out = 16'(-755);
			31393: out = 16'(-751);
			31394: out = 16'(1313);
			31395: out = 16'(2746);
			31396: out = 16'(2329);
			31397: out = 16'(-969);
			31398: out = 16'(-2372);
			31399: out = 16'(-1391);
			31400: out = 16'(-57);
			31401: out = 16'(-565);
			31402: out = 16'(919);
			31403: out = 16'(3162);
			31404: out = 16'(1754);
			31405: out = 16'(9);
			31406: out = 16'(-430);
			31407: out = 16'(973);
			31408: out = 16'(701);
			31409: out = 16'(1201);
			31410: out = 16'(174);
			31411: out = 16'(-7);
			31412: out = 16'(-257);
			31413: out = 16'(-452);
			31414: out = 16'(-1597);
			31415: out = 16'(-1138);
			31416: out = 16'(179);
			31417: out = 16'(1457);
			31418: out = 16'(359);
			31419: out = 16'(-92);
			31420: out = 16'(-420);
			31421: out = 16'(-2112);
			31422: out = 16'(-97);
			31423: out = 16'(3023);
			31424: out = 16'(3194);
			31425: out = 16'(-172);
			31426: out = 16'(-3155);
			31427: out = 16'(-1485);
			31428: out = 16'(831);
			31429: out = 16'(-280);
			31430: out = 16'(45);
			31431: out = 16'(-386);
			31432: out = 16'(-1513);
			31433: out = 16'(-2531);
			31434: out = 16'(1202);
			31435: out = 16'(2684);
			31436: out = 16'(1704);
			31437: out = 16'(-242);
			31438: out = 16'(324);
			31439: out = 16'(98);
			31440: out = 16'(-2030);
			31441: out = 16'(-3979);
			31442: out = 16'(-1350);
			31443: out = 16'(1959);
			31444: out = 16'(2646);
			31445: out = 16'(487);
			31446: out = 16'(-482);
			31447: out = 16'(-931);
			31448: out = 16'(-58);
			31449: out = 16'(-284);
			31450: out = 16'(-838);
			31451: out = 16'(-4435);
			31452: out = 16'(-1348);
			31453: out = 16'(1510);
			31454: out = 16'(1090);
			31455: out = 16'(-828);
			31456: out = 16'(632);
			31457: out = 16'(2116);
			31458: out = 16'(340);
			31459: out = 16'(-3138);
			31460: out = 16'(-5582);
			31461: out = 16'(-3148);
			31462: out = 16'(700);
			31463: out = 16'(1581);
			31464: out = 16'(1752);
			31465: out = 16'(2386);
			31466: out = 16'(2863);
			31467: out = 16'(975);
			31468: out = 16'(-1099);
			31469: out = 16'(-1796);
			31470: out = 16'(264);
			31471: out = 16'(1286);
			31472: out = 16'(272);
			31473: out = 16'(-1997);
			31474: out = 16'(-535);
			31475: out = 16'(1774);
			31476: out = 16'(988);
			31477: out = 16'(-3309);
			31478: out = 16'(-3639);
			31479: out = 16'(-243);
			31480: out = 16'(1434);
			31481: out = 16'(609);
			31482: out = 16'(-722);
			31483: out = 16'(-866);
			31484: out = 16'(-241);
			31485: out = 16'(1393);
			31486: out = 16'(2717);
			31487: out = 16'(2109);
			31488: out = 16'(-248);
			31489: out = 16'(257);
			31490: out = 16'(-57);
			31491: out = 16'(-9);
			31492: out = 16'(-1005);
			31493: out = 16'(-1945);
			31494: out = 16'(-654);
			31495: out = 16'(1870);
			31496: out = 16'(2663);
			31497: out = 16'(1063);
			31498: out = 16'(1349);
			31499: out = 16'(1713);
			31500: out = 16'(112);
			31501: out = 16'(-3701);
			31502: out = 16'(-3835);
			31503: out = 16'(-1424);
			31504: out = 16'(1950);
			31505: out = 16'(2824);
			31506: out = 16'(3567);
			31507: out = 16'(1803);
			31508: out = 16'(1669);
			31509: out = 16'(1410);
			31510: out = 16'(-622);
			31511: out = 16'(-3887);
			31512: out = 16'(-3679);
			31513: out = 16'(-607);
			31514: out = 16'(1381);
			31515: out = 16'(1646);
			31516: out = 16'(639);
			31517: out = 16'(-329);
			31518: out = 16'(-460);
			31519: out = 16'(1069);
			31520: out = 16'(2084);
			31521: out = 16'(344);
			31522: out = 16'(-3242);
			31523: out = 16'(-2774);
			31524: out = 16'(-1777);
			31525: out = 16'(-891);
			31526: out = 16'(-1088);
			31527: out = 16'(224);
			31528: out = 16'(1008);
			31529: out = 16'(1771);
			31530: out = 16'(968);
			31531: out = 16'(186);
			31532: out = 16'(-1854);
			31533: out = 16'(-1509);
			31534: out = 16'(-1172);
			31535: out = 16'(-1981);
			31536: out = 16'(-2544);
			31537: out = 16'(-122);
			31538: out = 16'(2468);
			31539: out = 16'(2619);
			31540: out = 16'(2120);
			31541: out = 16'(22);
			31542: out = 16'(-2074);
			31543: out = 16'(-3077);
			31544: out = 16'(-2587);
			31545: out = 16'(-445);
			31546: out = 16'(178);
			31547: out = 16'(-477);
			31548: out = 16'(242);
			31549: out = 16'(481);
			31550: out = 16'(1006);
			31551: out = 16'(900);
			31552: out = 16'(62);
			31553: out = 16'(-711);
			31554: out = 16'(-1405);
			31555: out = 16'(-829);
			31556: out = 16'(954);
			31557: out = 16'(2613);
			31558: out = 16'(2150);
			31559: out = 16'(766);
			31560: out = 16'(108);
			31561: out = 16'(479);
			31562: out = 16'(-110);
			31563: out = 16'(-1357);
			31564: out = 16'(-1765);
			31565: out = 16'(239);
			31566: out = 16'(2123);
			31567: out = 16'(2754);
			31568: out = 16'(776);
			31569: out = 16'(-1291);
			31570: out = 16'(-606);
			31571: out = 16'(2215);
			31572: out = 16'(1934);
			31573: out = 16'(-1855);
			31574: out = 16'(-2145);
			31575: out = 16'(881);
			31576: out = 16'(2996);
			31577: out = 16'(1091);
			31578: out = 16'(-1157);
			31579: out = 16'(18);
			31580: out = 16'(2686);
			31581: out = 16'(2183);
			31582: out = 16'(-846);
			31583: out = 16'(-3148);
			31584: out = 16'(-1607);
			31585: out = 16'(924);
			31586: out = 16'(1251);
			31587: out = 16'(263);
			31588: out = 16'(287);
			31589: out = 16'(1218);
			31590: out = 16'(1109);
			31591: out = 16'(-284);
			31592: out = 16'(-935);
			31593: out = 16'(-285);
			31594: out = 16'(-216);
			31595: out = 16'(-421);
			31596: out = 16'(-627);
			31597: out = 16'(1125);
			31598: out = 16'(2661);
			31599: out = 16'(3047);
			31600: out = 16'(-2463);
			31601: out = 16'(-4302);
			31602: out = 16'(-623);
			31603: out = 16'(2600);
			31604: out = 16'(1010);
			31605: out = 16'(-2717);
			31606: out = 16'(-4284);
			31607: out = 16'(-2892);
			31608: out = 16'(1158);
			31609: out = 16'(1276);
			31610: out = 16'(-1585);
			31611: out = 16'(-3890);
			31612: out = 16'(69);
			31613: out = 16'(1537);
			31614: out = 16'(413);
			31615: out = 16'(-1583);
			31616: out = 16'(36);
			31617: out = 16'(-1377);
			31618: out = 16'(-2421);
			31619: out = 16'(-1986);
			31620: out = 16'(246);
			31621: out = 16'(1252);
			31622: out = 16'(2330);
			31623: out = 16'(2748);
			31624: out = 16'(1676);
			31625: out = 16'(-1183);
			31626: out = 16'(-3315);
			31627: out = 16'(-2693);
			31628: out = 16'(-309);
			31629: out = 16'(-1287);
			31630: out = 16'(-599);
			31631: out = 16'(922);
			31632: out = 16'(1384);
			31633: out = 16'(467);
			31634: out = 16'(-1141);
			31635: out = 16'(-76);
			31636: out = 16'(2317);
			31637: out = 16'(1377);
			31638: out = 16'(905);
			31639: out = 16'(-101);
			31640: out = 16'(-569);
			31641: out = 16'(-957);
			31642: out = 16'(-47);
			31643: out = 16'(246);
			31644: out = 16'(-50);
			31645: out = 16'(-301);
			31646: out = 16'(1240);
			31647: out = 16'(995);
			31648: out = 16'(-1349);
			31649: out = 16'(-3363);
			31650: out = 16'(-844);
			31651: out = 16'(2339);
			31652: out = 16'(2365);
			31653: out = 16'(-551);
			31654: out = 16'(-1199);
			31655: out = 16'(775);
			31656: out = 16'(2549);
			31657: out = 16'(988);
			31658: out = 16'(-188);
			31659: out = 16'(-2727);
			31660: out = 16'(272);
			31661: out = 16'(3314);
			31662: out = 16'(2819);
			31663: out = 16'(-999);
			31664: out = 16'(-18);
			31665: out = 16'(3032);
			31666: out = 16'(3203);
			31667: out = 16'(-114);
			31668: out = 16'(-2794);
			31669: out = 16'(-2341);
			31670: out = 16'(764);
			31671: out = 16'(2222);
			31672: out = 16'(4133);
			31673: out = 16'(2348);
			31674: out = 16'(-389);
			31675: out = 16'(-1315);
			31676: out = 16'(-792);
			31677: out = 16'(-1647);
			31678: out = 16'(-1788);
			31679: out = 16'(507);
			31680: out = 16'(1617);
			31681: out = 16'(23);
			31682: out = 16'(-1185);
			31683: out = 16'(636);
			31684: out = 16'(2253);
			31685: out = 16'(981);
			31686: out = 16'(-708);
			31687: out = 16'(124);
			31688: out = 16'(878);
			31689: out = 16'(484);
			31690: out = 16'(-2346);
			31691: out = 16'(-4684);
			31692: out = 16'(-3621);
			31693: out = 16'(-12);
			31694: out = 16'(2888);
			31695: out = 16'(1637);
			31696: out = 16'(-2817);
			31697: out = 16'(-4326);
			31698: out = 16'(-1783);
			31699: out = 16'(993);
			31700: out = 16'(67);
			31701: out = 16'(327);
			31702: out = 16'(-579);
			31703: out = 16'(-148);
			31704: out = 16'(357);
			31705: out = 16'(142);
			31706: out = 16'(-510);
			31707: out = 16'(-114);
			31708: out = 16'(529);
			31709: out = 16'(-41);
			31710: out = 16'(-2650);
			31711: out = 16'(-4369);
			31712: out = 16'(-3403);
			31713: out = 16'(-1387);
			31714: out = 16'(498);
			31715: out = 16'(1150);
			31716: out = 16'(2252);
			31717: out = 16'(3007);
			31718: out = 16'(709);
			31719: out = 16'(-2753);
			31720: out = 16'(-3980);
			31721: out = 16'(-1860);
			31722: out = 16'(308);
			31723: out = 16'(1752);
			31724: out = 16'(2437);
			31725: out = 16'(2749);
			31726: out = 16'(1477);
			31727: out = 16'(822);
			31728: out = 16'(32);
			31729: out = 16'(-927);
			31730: out = 16'(-1937);
			31731: out = 16'(-431);
			31732: out = 16'(1958);
			31733: out = 16'(3142);
			31734: out = 16'(1577);
			31735: out = 16'(771);
			31736: out = 16'(767);
			31737: out = 16'(1822);
			31738: out = 16'(1111);
			31739: out = 16'(-2630);
			31740: out = 16'(-4151);
			31741: out = 16'(-1537);
			31742: out = 16'(1937);
			31743: out = 16'(2654);
			31744: out = 16'(1028);
			31745: out = 16'(677);
			31746: out = 16'(1442);
			31747: out = 16'(770);
			31748: out = 16'(456);
			31749: out = 16'(30);
			31750: out = 16'(201);
			31751: out = 16'(1415);
			31752: out = 16'(-92);
			31753: out = 16'(1051);
			31754: out = 16'(1318);
			31755: out = 16'(-299);
			31756: out = 16'(-118);
			31757: out = 16'(1032);
			31758: out = 16'(1693);
			31759: out = 16'(1057);
			31760: out = 16'(1185);
			31761: out = 16'(-154);
			31762: out = 16'(-1974);
			31763: out = 16'(-2500);
			31764: out = 16'(-142);
			31765: out = 16'(1005);
			31766: out = 16'(794);
			31767: out = 16'(198);
			31768: out = 16'(243);
			31769: out = 16'(-7);
			31770: out = 16'(-1506);
			31771: out = 16'(-2052);
			31772: out = 16'(-634);
			31773: out = 16'(-1165);
			31774: out = 16'(-2536);
			31775: out = 16'(-3338);
			31776: out = 16'(-2283);
			31777: out = 16'(-1225);
			31778: out = 16'(132);
			31779: out = 16'(1080);
			31780: out = 16'(1093);
			31781: out = 16'(-1006);
			31782: out = 16'(-2308);
			31783: out = 16'(-1745);
			31784: out = 16'(-51);
			31785: out = 16'(-231);
			31786: out = 16'(-1865);
			31787: out = 16'(-1891);
			31788: out = 16'(1338);
			31789: out = 16'(3616);
			31790: out = 16'(1386);
			31791: out = 16'(-2763);
			31792: out = 16'(-3269);
			31793: out = 16'(256);
			31794: out = 16'(2540);
			31795: out = 16'(1234);
			31796: out = 16'(-848);
			31797: out = 16'(-1258);
			31798: out = 16'(17);
			31799: out = 16'(106);
			31800: out = 16'(767);
			31801: out = 16'(1641);
			31802: out = 16'(1392);
			31803: out = 16'(-516);
			31804: out = 16'(-786);
			31805: out = 16'(591);
			31806: out = 16'(1342);
			31807: out = 16'(315);
			31808: out = 16'(-455);
			31809: out = 16'(6);
			31810: out = 16'(1702);
			31811: out = 16'(1624);
			31812: out = 16'(1811);
			31813: out = 16'(-116);
			31814: out = 16'(-2351);
			31815: out = 16'(-2673);
			31816: out = 16'(1579);
			31817: out = 16'(3474);
			31818: out = 16'(1841);
			31819: out = 16'(81);
			31820: out = 16'(855);
			31821: out = 16'(1124);
			31822: out = 16'(-603);
			31823: out = 16'(-2642);
			31824: out = 16'(-1608);
			31825: out = 16'(1060);
			31826: out = 16'(3454);
			31827: out = 16'(3742);
			31828: out = 16'(1612);
			31829: out = 16'(-371);
			31830: out = 16'(-620);
			31831: out = 16'(-297);
			31832: out = 16'(-655);
			31833: out = 16'(-1753);
			31834: out = 16'(-371);
			31835: out = 16'(1946);
			31836: out = 16'(1441);
			31837: out = 16'(-1748);
			31838: out = 16'(-3156);
			31839: out = 16'(-1511);
			31840: out = 16'(-227);
			31841: out = 16'(1562);
			31842: out = 16'(990);
			31843: out = 16'(-605);
			31844: out = 16'(-2268);
			31845: out = 16'(-279);
			31846: out = 16'(-918);
			31847: out = 16'(-2330);
			31848: out = 16'(-2073);
			31849: out = 16'(2233);
			31850: out = 16'(3260);
			31851: out = 16'(1659);
			31852: out = 16'(-438);
			31853: out = 16'(-652);
			31854: out = 16'(-1092);
			31855: out = 16'(-1944);
			31856: out = 16'(-2609);
			31857: out = 16'(-917);
			31858: out = 16'(-362);
			31859: out = 16'(916);
			31860: out = 16'(1185);
			31861: out = 16'(381);
			31862: out = 16'(-24);
			31863: out = 16'(231);
			31864: out = 16'(43);
			31865: out = 16'(-1527);
			31866: out = 16'(-2926);
			31867: out = 16'(-3139);
			31868: out = 16'(-1221);
			31869: out = 16'(762);
			31870: out = 16'(441);
			31871: out = 16'(-364);
			31872: out = 16'(788);
			31873: out = 16'(3339);
			31874: out = 16'(2596);
			31875: out = 16'(638);
			31876: out = 16'(-4014);
			31877: out = 16'(-5640);
			31878: out = 16'(-2876);
			31879: out = 16'(-1137);
			31880: out = 16'(-715);
			31881: out = 16'(1077);
			31882: out = 16'(4182);
			31883: out = 16'(2930);
			31884: out = 16'(7);
			31885: out = 16'(-2004);
			31886: out = 16'(-1057);
			31887: out = 16'(-62);
			31888: out = 16'(243);
			31889: out = 16'(554);
			31890: out = 16'(2043);
			31891: out = 16'(2919);
			31892: out = 16'(1676);
			31893: out = 16'(-904);
			31894: out = 16'(-1949);
			31895: out = 16'(-423);
			31896: out = 16'(249);
			31897: out = 16'(-18);
			31898: out = 16'(-608);
			31899: out = 16'(511);
			31900: out = 16'(2204);
			31901: out = 16'(3858);
			31902: out = 16'(2206);
			31903: out = 16'(-1549);
			31904: out = 16'(-5817);
			31905: out = 16'(-2549);
			31906: out = 16'(1141);
			31907: out = 16'(1566);
			31908: out = 16'(627);
			31909: out = 16'(1381);
			31910: out = 16'(2018);
			31911: out = 16'(1494);
			31912: out = 16'(1382);
			31913: out = 16'(-16);
			31914: out = 16'(-340);
			31915: out = 16'(-1436);
			31916: out = 16'(-2613);
			31917: out = 16'(-1027);
			31918: out = 16'(812);
			31919: out = 16'(1109);
			31920: out = 16'(405);
			31921: out = 16'(1226);
			31922: out = 16'(826);
			31923: out = 16'(-612);
			31924: out = 16'(-1726);
			31925: out = 16'(-1199);
			31926: out = 16'(129);
			31927: out = 16'(76);
			31928: out = 16'(-1148);
			31929: out = 16'(-2576);
			31930: out = 16'(1047);
			31931: out = 16'(1928);
			31932: out = 16'(703);
			31933: out = 16'(-621);
			31934: out = 16'(375);
			31935: out = 16'(107);
			31936: out = 16'(76);
			31937: out = 16'(280);
			31938: out = 16'(71);
			31939: out = 16'(-223);
			31940: out = 16'(215);
			31941: out = 16'(-994);
			31942: out = 16'(-4947);
			31943: out = 16'(-6120);
			31944: out = 16'(-1196);
			31945: out = 16'(4058);
			31946: out = 16'(3690);
			31947: out = 16'(-868);
			31948: out = 16'(-1721);
			31949: out = 16'(-240);
			31950: out = 16'(-1319);
			31951: out = 16'(-3707);
			31952: out = 16'(-1768);
			31953: out = 16'(1771);
			31954: out = 16'(1524);
			31955: out = 16'(600);
			31956: out = 16'(-227);
			31957: out = 16'(910);
			31958: out = 16'(1217);
			31959: out = 16'(-318);
			31960: out = 16'(-2088);
			31961: out = 16'(-2274);
			31962: out = 16'(-693);
			31963: out = 16'(1506);
			31964: out = 16'(2043);
			31965: out = 16'(993);
			31966: out = 16'(-163);
			31967: out = 16'(311);
			31968: out = 16'(1185);
			31969: out = 16'(978);
			31970: out = 16'(-1089);
			31971: out = 16'(-3099);
			31972: out = 16'(-3194);
			31973: out = 16'(-126);
			31974: out = 16'(2696);
			31975: out = 16'(2907);
			31976: out = 16'(1700);
			31977: out = 16'(305);
			31978: out = 16'(53);
			31979: out = 16'(-97);
			31980: out = 16'(-452);
			31981: out = 16'(-1484);
			31982: out = 16'(-566);
			31983: out = 16'(972);
			31984: out = 16'(1377);
			31985: out = 16'(659);
			31986: out = 16'(946);
			31987: out = 16'(1225);
			31988: out = 16'(-417);
			31989: out = 16'(-2162);
			31990: out = 16'(-2722);
			31991: out = 16'(-606);
			31992: out = 16'(1570);
			31993: out = 16'(1528);
			31994: out = 16'(269);
			31995: out = 16'(986);
			31996: out = 16'(3871);
			31997: out = 16'(4861);
			31998: out = 16'(1568);
			31999: out = 16'(-2695);
			32000: out = 16'(-3062);
			32001: out = 16'(-170);
			32002: out = 16'(2425);
			32003: out = 16'(303);
			32004: out = 16'(-1999);
			32005: out = 16'(-242);
			32006: out = 16'(2048);
			32007: out = 16'(1397);
			32008: out = 16'(-1830);
			32009: out = 16'(-3518);
			32010: out = 16'(-1034);
			32011: out = 16'(65);
			32012: out = 16'(-410);
			32013: out = 16'(-465);
			32014: out = 16'(-159);
			32015: out = 16'(822);
			32016: out = 16'(424);
			32017: out = 16'(-185);
			32018: out = 16'(-700);
			32019: out = 16'(1447);
			32020: out = 16'(923);
			32021: out = 16'(-443);
			32022: out = 16'(-695);
			32023: out = 16'(-1937);
			32024: out = 16'(-2633);
			32025: out = 16'(-2020);
			32026: out = 16'(-311);
			32027: out = 16'(478);
			32028: out = 16'(225);
			32029: out = 16'(222);
			32030: out = 16'(487);
			32031: out = 16'(107);
			32032: out = 16'(-1158);
			32033: out = 16'(-1566);
			32034: out = 16'(-1786);
			32035: out = 16'(-2963);
			32036: out = 16'(-3240);
			32037: out = 16'(-610);
			32038: out = 16'(2247);
			32039: out = 16'(1693);
			32040: out = 16'(-1594);
			32041: out = 16'(-1485);
			32042: out = 16'(1670);
			32043: out = 16'(2243);
			32044: out = 16'(-1000);
			32045: out = 16'(-4656);
			32046: out = 16'(-3375);
			32047: out = 16'(923);
			32048: out = 16'(1514);
			32049: out = 16'(1094);
			32050: out = 16'(524);
			32051: out = 16'(785);
			32052: out = 16'(159);
			32053: out = 16'(674);
			32054: out = 16'(235);
			32055: out = 16'(-713);
			32056: out = 16'(-1189);
			32057: out = 16'(1370);
			32058: out = 16'(2882);
			32059: out = 16'(2032);
			32060: out = 16'(99);
			32061: out = 16'(30);
			32062: out = 16'(1299);
			32063: out = 16'(1931);
			32064: out = 16'(1217);
			32065: out = 16'(156);
			32066: out = 16'(-701);
			32067: out = 16'(-1245);
			32068: out = 16'(-534);
			32069: out = 16'(1298);
			32070: out = 16'(1670);
			32071: out = 16'(365);
			32072: out = 16'(-470);
			32073: out = 16'(-52);
			32074: out = 16'(274);
			32075: out = 16'(-1537);
			32076: out = 16'(-2045);
			32077: out = 16'(730);
			32078: out = 16'(2460);
			32079: out = 16'(2028);
			32080: out = 16'(1233);
			32081: out = 16'(1297);
			32082: out = 16'(1488);
			32083: out = 16'(-2416);
			32084: out = 16'(-4226);
			32085: out = 16'(-929);
			32086: out = 16'(2235);
			32087: out = 16'(2474);
			32088: out = 16'(592);
			32089: out = 16'(128);
			32090: out = 16'(1258);
			32091: out = 16'(2440);
			32092: out = 16'(1367);
			32093: out = 16'(-1116);
			32094: out = 16'(-2592);
			32095: out = 16'(-1681);
			32096: out = 16'(14);
			32097: out = 16'(-559);
			32098: out = 16'(-2600);
			32099: out = 16'(-348);
			32100: out = 16'(1358);
			32101: out = 16'(1390);
			32102: out = 16'(101);
			32103: out = 16'(-612);
			32104: out = 16'(-120);
			32105: out = 16'(-1085);
			32106: out = 16'(-2974);
			32107: out = 16'(-2487);
			32108: out = 16'(-674);
			32109: out = 16'(781);
			32110: out = 16'(1036);
			32111: out = 16'(1458);
			32112: out = 16'(206);
			32113: out = 16'(-347);
			32114: out = 16'(-747);
			32115: out = 16'(-1244);
			32116: out = 16'(-2356);
			32117: out = 16'(-3404);
			32118: out = 16'(-2821);
			32119: out = 16'(-243);
			32120: out = 16'(2566);
			32121: out = 16'(2249);
			32122: out = 16'(311);
			32123: out = 16'(-926);
			32124: out = 16'(227);
			32125: out = 16'(1456);
			32126: out = 16'(2048);
			32127: out = 16'(636);
			32128: out = 16'(-1423);
			32129: out = 16'(-3508);
			32130: out = 16'(-1689);
			32131: out = 16'(1073);
			32132: out = 16'(1814);
			32133: out = 16'(-165);
			32134: out = 16'(73);
			32135: out = 16'(670);
			32136: out = 16'(-175);
			32137: out = 16'(-1262);
			32138: out = 16'(-601);
			32139: out = 16'(1157);
			32140: out = 16'(1580);
			32141: out = 16'(-867);
			32142: out = 16'(1036);
			32143: out = 16'(2713);
			32144: out = 16'(1884);
			32145: out = 16'(-1060);
			32146: out = 16'(-1668);
			32147: out = 16'(-34);
			32148: out = 16'(1931);
			32149: out = 16'(1526);
			32150: out = 16'(1723);
			32151: out = 16'(-915);
			32152: out = 16'(-2172);
			32153: out = 16'(-717);
			32154: out = 16'(1159);
			32155: out = 16'(1708);
			32156: out = 16'(2274);
			32157: out = 16'(2914);
			32158: out = 16'(1196);
			32159: out = 16'(-823);
			32160: out = 16'(-2391);
			32161: out = 16'(-1670);
			32162: out = 16'(-186);
			32163: out = 16'(1563);
			32164: out = 16'(854);
			32165: out = 16'(-322);
			32166: out = 16'(-20);
			32167: out = 16'(-193);
			32168: out = 16'(222);
			32169: out = 16'(-279);
			32170: out = 16'(-1775);
			32171: out = 16'(285);
			32172: out = 16'(-714);
			32173: out = 16'(-892);
			32174: out = 16'(424);
			32175: out = 16'(2453);
			32176: out = 16'(1763);
			32177: out = 16'(571);
			32178: out = 16'(-611);
			32179: out = 16'(-2217);
			32180: out = 16'(-4514);
			32181: out = 16'(-3145);
			32182: out = 16'(631);
			32183: out = 16'(1084);
			32184: out = 16'(2214);
			32185: out = 16'(386);
			32186: out = 16'(933);
			32187: out = 16'(2934);
			32188: out = 16'(1654);
			32189: out = 16'(-1541);
			32190: out = 16'(-2348);
			32191: out = 16'(-563);
			32192: out = 16'(-2182);
			32193: out = 16'(-2632);
			32194: out = 16'(-1075);
			32195: out = 16'(2185);
			32196: out = 16'(2305);
			32197: out = 16'(955);
			32198: out = 16'(-1724);
			32199: out = 16'(-2247);
			32200: out = 16'(-1126);
			32201: out = 16'(-841);
			32202: out = 16'(-2003);
			32203: out = 16'(-1746);
			32204: out = 16'(1054);
			32205: out = 16'(3733);
			32206: out = 16'(2821);
			32207: out = 16'(-419);
			32208: out = 16'(-2290);
			32209: out = 16'(262);
			32210: out = 16'(-523);
			32211: out = 16'(-2738);
			32212: out = 16'(-2757);
			32213: out = 16'(403);
			32214: out = 16'(1925);
			32215: out = 16'(471);
			32216: out = 16'(-682);
			32217: out = 16'(1631);
			32218: out = 16'(2797);
			32219: out = 16'(1636);
			32220: out = 16'(-823);
			32221: out = 16'(-1410);
			32222: out = 16'(-3436);
			32223: out = 16'(-2324);
			32224: out = 16'(-209);
			32225: out = 16'(2284);
			32226: out = 16'(2406);
			32227: out = 16'(3916);
			32228: out = 16'(2701);
			32229: out = 16'(-1343);
			32230: out = 16'(-6586);
			32231: out = 16'(-4543);
			32232: out = 16'(-355);
			32233: out = 16'(1651);
			32234: out = 16'(1564);
			32235: out = 16'(1315);
			32236: out = 16'(2222);
			32237: out = 16'(2208);
			32238: out = 16'(227);
			32239: out = 16'(-1601);
			32240: out = 16'(-2437);
			32241: out = 16'(-2482);
			32242: out = 16'(-2178);
			32243: out = 16'(244);
			32244: out = 16'(1317);
			32245: out = 16'(1208);
			32246: out = 16'(420);
			32247: out = 16'(155);
			32248: out = 16'(76);
			32249: out = 16'(73);
			32250: out = 16'(316);
			32251: out = 16'(1429);
			32252: out = 16'(676);
			32253: out = 16'(26);
			32254: out = 16'(280);
			32255: out = 16'(1369);
			32256: out = 16'(266);
			32257: out = 16'(-660);
			32258: out = 16'(-957);
			32259: out = 16'(-468);
			32260: out = 16'(-550);
			32261: out = 16'(-111);
			32262: out = 16'(144);
			32263: out = 16'(23);
			32264: out = 16'(149);
			32265: out = 16'(224);
			32266: out = 16'(1517);
			32267: out = 16'(2362);
			32268: out = 16'(-64);
			32269: out = 16'(-430);
			32270: out = 16'(-370);
			32271: out = 16'(25);
			32272: out = 16'(-687);
			32273: out = 16'(-75);
			32274: out = 16'(89);
			32275: out = 16'(875);
			32276: out = 16'(1069);
			32277: out = 16'(-134);
			32278: out = 16'(-2745);
			32279: out = 16'(-2681);
			32280: out = 16'(432);
			32281: out = 16'(726);
			32282: out = 16'(1340);
			32283: out = 16'(1337);
			32284: out = 16'(1102);
			32285: out = 16'(-604);
			32286: out = 16'(-971);
			32287: out = 16'(-1129);
			32288: out = 16'(-1032);
			32289: out = 16'(-971);
			32290: out = 16'(897);
			32291: out = 16'(1601);
			32292: out = 16'(743);
			32293: out = 16'(-546);
			32294: out = 16'(-176);
			32295: out = 16'(164);
			32296: out = 16'(-727);
			32297: out = 16'(-1921);
			32298: out = 16'(-162);
			32299: out = 16'(530);
			32300: out = 16'(-136);
			32301: out = 16'(-1067);
			32302: out = 16'(-1082);
			32303: out = 16'(880);
			32304: out = 16'(601);
			32305: out = 16'(-1869);
			32306: out = 16'(-3852);
			32307: out = 16'(-843);
			32308: out = 16'(636);
			32309: out = 16'(-574);
			32310: out = 16'(-1552);
			32311: out = 16'(1179);
			32312: out = 16'(3448);
			32313: out = 16'(3155);
			32314: out = 16'(920);
			32315: out = 16'(-2599);
			32316: out = 16'(-2136);
			32317: out = 16'(741);
			32318: out = 16'(2627);
			32319: out = 16'(1449);
			32320: out = 16'(-1023);
			32321: out = 16'(-2055);
			32322: out = 16'(200);
			32323: out = 16'(3841);
			32324: out = 16'(1268);
			32325: out = 16'(-2314);
			32326: out = 16'(-2869);
			32327: out = 16'(207);
			32328: out = 16'(1573);
			32329: out = 16'(949);
			32330: out = 16'(-538);
			32331: out = 16'(-783);
			32332: out = 16'(1053);
			32333: out = 16'(1787);
			32334: out = 16'(1276);
			32335: out = 16'(96);
			32336: out = 16'(-500);
			32337: out = 16'(-1711);
			32338: out = 16'(-1810);
			32339: out = 16'(-673);
			32340: out = 16'(-28);
			32341: out = 16'(1088);
			32342: out = 16'(1472);
			32343: out = 16'(1016);
			32344: out = 16'(-42);
			32345: out = 16'(-529);
			32346: out = 16'(-154);
			32347: out = 16'(412);
			32348: out = 16'(-169);
			32349: out = 16'(70);
			32350: out = 16'(-145);
			32351: out = 16'(213);
			32352: out = 16'(230);
			32353: out = 16'(-876);
			32354: out = 16'(-634);
			32355: out = 16'(1292);
			32356: out = 16'(2227);
			32357: out = 16'(38);
			32358: out = 16'(-3263);
			32359: out = 16'(-3013);
			32360: out = 16'(802);
			32361: out = 16'(2637);
			32362: out = 16'(2363);
			32363: out = 16'(101);
			32364: out = 16'(-145);
			32365: out = 16'(1162);
			32366: out = 16'(308);
			32367: out = 16'(-2392);
			32368: out = 16'(-3042);
			32369: out = 16'(-11);
			32370: out = 16'(1004);
			32371: out = 16'(727);
			32372: out = 16'(-1209);
			32373: out = 16'(-1680);
			32374: out = 16'(-169);
			32375: out = 16'(1526);
			32376: out = 16'(814);
			32377: out = 16'(-1012);
			32378: out = 16'(-1392);
			32379: out = 16'(661);
			32380: out = 16'(1677);
			32381: out = 16'(696);
			32382: out = 16'(-506);
			32383: out = 16'(-241);
			32384: out = 16'(408);
			32385: out = 16'(54);
			32386: out = 16'(-526);
			32387: out = 16'(-201);
			32388: out = 16'(1280);
			32389: out = 16'(872);
			32390: out = 16'(-1593);
			32391: out = 16'(-1812);
			32392: out = 16'(-895);
			32393: out = 16'(1491);
			32394: out = 16'(2236);
			32395: out = 16'(459);
			32396: out = 16'(-1308);
			32397: out = 16'(-329);
			32398: out = 16'(1829);
			32399: out = 16'(1314);
			32400: out = 16'(526);
			32401: out = 16'(-1890);
			32402: out = 16'(-2032);
			32403: out = 16'(316);
			32404: out = 16'(2617);
			32405: out = 16'(2040);
			32406: out = 16'(504);
			32407: out = 16'(-98);
			32408: out = 16'(276);
			32409: out = 16'(-1318);
			32410: out = 16'(-2561);
			32411: out = 16'(-1392);
			32412: out = 16'(1103);
			32413: out = 16'(1786);
			32414: out = 16'(809);
			32415: out = 16'(-550);
			32416: out = 16'(-1581);
			32417: out = 16'(-96);
			32418: out = 16'(960);
			32419: out = 16'(993);
			32420: out = 16'(-336);
			32421: out = 16'(-422);
			32422: out = 16'(-1783);
			32423: out = 16'(-1568);
			32424: out = 16'(138);
			32425: out = 16'(1174);
			32426: out = 16'(1299);
			32427: out = 16'(929);
			32428: out = 16'(108);
			32429: out = 16'(24);
			32430: out = 16'(-1783);
			32431: out = 16'(-1958);
			32432: out = 16'(-1451);
			32433: out = 16'(-410);
			32434: out = 16'(-419);
			32435: out = 16'(1875);
			32436: out = 16'(2095);
			32437: out = 16'(-1409);
			32438: out = 16'(-2979);
			32439: out = 16'(-580);
			32440: out = 16'(1913);
			32441: out = 16'(756);
			32442: out = 16'(-1638);
			32443: out = 16'(-1032);
			32444: out = 16'(932);
			32445: out = 16'(917);
			32446: out = 16'(-855);
			32447: out = 16'(-465);
			32448: out = 16'(431);
			32449: out = 16'(-119);
			32450: out = 16'(-1413);
			32451: out = 16'(-420);
			32452: out = 16'(708);
			32453: out = 16'(648);
			32454: out = 16'(76);
			32455: out = 16'(1068);
			32456: out = 16'(1023);
			32457: out = 16'(-528);
			32458: out = 16'(-2174);
			32459: out = 16'(-3106);
			32460: out = 16'(-2065);
			32461: out = 16'(-712);
			32462: out = 16'(1197);
			32463: out = 16'(3437);
			32464: out = 16'(4379);
			32465: out = 16'(1734);
			32466: out = 16'(-1769);
			32467: out = 16'(-2008);
			32468: out = 16'(-2120);
			32469: out = 16'(-2340);
			32470: out = 16'(-2102);
			32471: out = 16'(-318);
			32472: out = 16'(1197);
			32473: out = 16'(781);
			32474: out = 16'(-21);
			32475: out = 16'(722);
			32476: out = 16'(1236);
			32477: out = 16'(679);
			32478: out = 16'(-548);
			32479: out = 16'(-1020);
			32480: out = 16'(-1495);
			32481: out = 16'(-1171);
			32482: out = 16'(147);
			32483: out = 16'(2541);
			32484: out = 16'(3796);
			32485: out = 16'(1309);
			32486: out = 16'(-2051);
			32487: out = 16'(-2434);
			32488: out = 16'(23);
			32489: out = 16'(1335);
			32490: out = 16'(502);
			32491: out = 16'(99);
			32492: out = 16'(1092);
			32493: out = 16'(3782);
			32494: out = 16'(914);
			32495: out = 16'(-3692);
			32496: out = 16'(-5404);
			32497: out = 16'(-1464);
			32498: out = 16'(852);
			32499: out = 16'(1576);
			32500: out = 16'(1017);
			32501: out = 16'(-383);
			32502: out = 16'(-787);
			32503: out = 16'(657);
			32504: out = 16'(1590);
			32505: out = 16'(-213);
			32506: out = 16'(-2525);
			32507: out = 16'(-2294);
			32508: out = 16'(-279);
			32509: out = 16'(365);
			32510: out = 16'(1380);
			32511: out = 16'(2268);
			32512: out = 16'(3174);
			32513: out = 16'(2030);
			32514: out = 16'(389);
			32515: out = 16'(-1656);
			32516: out = 16'(-2069);
			32517: out = 16'(-1995);
			32518: out = 16'(-417);
			32519: out = 16'(-528);
			32520: out = 16'(1941);
			32521: out = 16'(4053);
			32522: out = 16'(2337);
			32523: out = 16'(-1922);
			32524: out = 16'(-3014);
			32525: out = 16'(-468);
			32526: out = 16'(1017);
			32527: out = 16'(-479);
			32528: out = 16'(-1282);
			32529: out = 16'(622);
			32530: out = 16'(2381);
			32531: out = 16'(1629);
			32532: out = 16'(-1681);
			32533: out = 16'(-3092);
			32534: out = 16'(-958);
			32535: out = 16'(72);
			32536: out = 16'(1401);
			32537: out = 16'(127);
			32538: out = 16'(-2060);
			32539: out = 16'(-3437);
			32540: out = 16'(152);
			32541: out = 16'(1940);
			32542: out = 16'(604);
			32543: out = 16'(-886);
			32544: out = 16'(-2104);
			32545: out = 16'(-147);
			32546: out = 16'(2068);
			32547: out = 16'(2336);
			32548: out = 16'(339);
			32549: out = 16'(-268);
			32550: out = 16'(150);
			32551: out = 16'(-377);
			32552: out = 16'(-1704);
			32553: out = 16'(-3354);
			32554: out = 16'(-2259);
			32555: out = 16'(904);
			32556: out = 16'(2791);
			32557: out = 16'(2042);
			32558: out = 16'(175);
			32559: out = 16'(-450);
			32560: out = 16'(328);
			32561: out = 16'(1553);
			32562: out = 16'(1099);
			32563: out = 16'(-279);
			32564: out = 16'(-1217);
			32565: out = 16'(-3301);
			32566: out = 16'(-2933);
			32567: out = 16'(-684);
			32568: out = 16'(1639);
			32569: out = 16'(2545);
			32570: out = 16'(1286);
			32571: out = 16'(-223);
			32572: out = 16'(-445);
			32573: out = 16'(-141);
			32574: out = 16'(1084);
			32575: out = 16'(587);
			32576: out = 16'(-924);
			32577: out = 16'(-407);
			32578: out = 16'(718);
			32579: out = 16'(2452);
			32580: out = 16'(2489);
			32581: out = 16'(1126);
			32582: out = 16'(-562);
			32583: out = 16'(342);
			32584: out = 16'(1071);
			32585: out = 16'(-519);
			32586: out = 16'(-946);
			32587: out = 16'(-1431);
			32588: out = 16'(-658);
			32589: out = 16'(-225);
			32590: out = 16'(-1052);
			32591: out = 16'(-317);
			32592: out = 16'(1001);
			32593: out = 16'(671);
			32594: out = 16'(-1526);
			32595: out = 16'(-1887);
			32596: out = 16'(-32);
			32597: out = 16'(1222);
			32598: out = 16'(-278);
			32599: out = 16'(-1307);
			32600: out = 16'(-1224);
			32601: out = 16'(-258);
			32602: out = 16'(-227);
			32603: out = 16'(127);
			32604: out = 16'(61);
			32605: out = 16'(978);
			32606: out = 16'(1524);
			32607: out = 16'(81);
			32608: out = 16'(-1912);
			32609: out = 16'(-2694);
			32610: out = 16'(-1470);
			32611: out = 16'(360);
			32612: out = 16'(1652);
			32613: out = 16'(740);
			32614: out = 16'(-1034);
			32615: out = 16'(-774);
			32616: out = 16'(732);
			32617: out = 16'(1825);
			32618: out = 16'(115);
			32619: out = 16'(-1749);
			32620: out = 16'(659);
			32621: out = 16'(3347);
			32622: out = 16'(1926);
			32623: out = 16'(-2347);
			32624: out = 16'(-5659);
			32625: out = 16'(-1133);
			32626: out = 16'(2465);
			32627: out = 16'(782);
			32628: out = 16'(-1616);
			32629: out = 16'(-877);
			32630: out = 16'(1342);
			32631: out = 16'(1097);
			32632: out = 16'(-877);
			32633: out = 16'(-429);
			32634: out = 16'(1710);
			32635: out = 16'(2068);
			32636: out = 16'(-404);
			32637: out = 16'(-2648);
			32638: out = 16'(-2514);
			32639: out = 16'(-242);
			32640: out = 16'(1446);
			32641: out = 16'(1834);
			32642: out = 16'(1393);
			32643: out = 16'(1381);
			32644: out = 16'(865);
			32645: out = 16'(-972);
			32646: out = 16'(-3915);
			32647: out = 16'(-3903);
			32648: out = 16'(-767);
			32649: out = 16'(1688);
			32650: out = 16'(2762);
			32651: out = 16'(1226);
			32652: out = 16'(-257);
			32653: out = 16'(192);
			32654: out = 16'(1084);
			32655: out = 16'(806);
			32656: out = 16'(-933);
			32657: out = 16'(-1946);
			32658: out = 16'(-2199);
			32659: out = 16'(650);
			32660: out = 16'(1997);
			32661: out = 16'(902);
			32662: out = 16'(-887);
			32663: out = 16'(-1119);
			32664: out = 16'(-551);
			32665: out = 16'(441);
			32666: out = 16'(1231);
			32667: out = 16'(834);
			32668: out = 16'(-1075);
			32669: out = 16'(-1630);
			32670: out = 16'(100);
			32671: out = 16'(161);
			32672: out = 16'(-672);
			32673: out = 16'(-354);
			32674: out = 16'(1564);
			32675: out = 16'(1784);
			32676: out = 16'(575);
			32677: out = 16'(296);
			32678: out = 16'(1328);
			32679: out = 16'(-27);
			32680: out = 16'(-1165);
			32681: out = 16'(-1104);
			32682: out = 16'(271);
			32683: out = 16'(-166);
			32684: out = 16'(425);
			32685: out = 16'(443);
			32686: out = 16'(182);
			32687: out = 16'(-1124);
			32688: out = 16'(-125);
			32689: out = 16'(23);
			32690: out = 16'(65);
			32691: out = 16'(602);
			32692: out = 16'(1506);
			32693: out = 16'(1199);
			32694: out = 16'(-1156);
			32695: out = 16'(-3643);
			32696: out = 16'(-2640);
			32697: out = 16'(1023);
			32698: out = 16'(3181);
			32699: out = 16'(1814);
			32700: out = 16'(-333);
			32701: out = 16'(-147);
			32702: out = 16'(1166);
			32703: out = 16'(478);
			32704: out = 16'(-2007);
			32705: out = 16'(-1962);
			32706: out = 16'(166);
			32707: out = 16'(1055);
			32708: out = 16'(-933);
			32709: out = 16'(-3622);
			32710: out = 16'(-2663);
			32711: out = 16'(456);
			32712: out = 16'(1679);
			32713: out = 16'(1610);
			32714: out = 16'(308);
			32715: out = 16'(49);
			32716: out = 16'(-105);
			32717: out = 16'(177);
			32718: out = 16'(-2015);
			32719: out = 16'(-1576);
			32720: out = 16'(718);
			32721: out = 16'(1623);
			32722: out = 16'(-295);
			32723: out = 16'(-1164);
			32724: out = 16'(232);
			32725: out = 16'(1245);
			32726: out = 16'(1548);
			32727: out = 16'(594);
			32728: out = 16'(640);
			32729: out = 16'(1258);
			32730: out = 16'(1378);
			32731: out = 16'(-1197);
			32732: out = 16'(-3584);
			32733: out = 16'(-3616);
			32734: out = 16'(-133);
			32735: out = 16'(498);
			32736: out = 16'(514);
			32737: out = 16'(376);
			32738: out = 16'(576);
			32739: out = 16'(-384);
			32740: out = 16'(-246);
			32741: out = 16'(-71);
			32742: out = 16'(-519);
			32743: out = 16'(-1076);
			32744: out = 16'(-71);
			32745: out = 16'(327);
			32746: out = 16'(-543);
			32747: out = 16'(-75);
			32748: out = 16'(1749);
			32749: out = 16'(2436);
			32750: out = 16'(873);
			32751: out = 16'(-865);
			32752: out = 16'(-473);
			32753: out = 16'(-4);
			32754: out = 16'(-1005);
			32755: out = 16'(-1916);
			32756: out = 16'(-1760);
			32757: out = 16'(-969);
			32758: out = 16'(-322);
			32759: out = 16'(122);
			32760: out = 16'(1554);
			32761: out = 16'(1673);
			32762: out = 16'(1359);
			32763: out = 16'(1660);
			32764: out = 16'(-742);
			32765: out = 16'(-1586);
			32766: out = 16'(-633);
			32767: out = 16'(1648);
			32768: out = 16'(1158);
			32769: out = 16'(1476);
			32770: out = 16'(660);
			32771: out = 16'(-41);
			32772: out = 16'(301);
			32773: out = 16'(193);
			32774: out = 16'(-1286);
			32775: out = 16'(-2775);
			32776: out = 16'(-1829);
			32777: out = 16'(-155);
			32778: out = 16'(1470);
			32779: out = 16'(1410);
			32780: out = 16'(235);
			32781: out = 16'(-1406);
			32782: out = 16'(-9);
			32783: out = 16'(2136);
			32784: out = 16'(2071);
			32785: out = 16'(-168);
			32786: out = 16'(-2321);
			32787: out = 16'(-1710);
			32788: out = 16'(206);
			32789: out = 16'(-75);
			32790: out = 16'(1192);
			32791: out = 16'(2483);
			32792: out = 16'(2386);
			32793: out = 16'(-220);
			32794: out = 16'(-2532);
			32795: out = 16'(-3513);
			32796: out = 16'(-2429);
			32797: out = 16'(-368);
			32798: out = 16'(2466);
			32799: out = 16'(3249);
			32800: out = 16'(1964);
			32801: out = 16'(-652);
			32802: out = 16'(-4724);
			32803: out = 16'(-6061);
			32804: out = 16'(-4167);
			32805: out = 16'(91);
			32806: out = 16'(2683);
			32807: out = 16'(3584);
			32808: out = 16'(924);
			32809: out = 16'(-1505);
			32810: out = 16'(138);
			32811: out = 16'(2156);
			32812: out = 16'(1626);
			32813: out = 16'(-1137);
			32814: out = 16'(-2927);
			32815: out = 16'(-2267);
			32816: out = 16'(-1052);
			32817: out = 16'(174);
			32818: out = 16'(1656);
			32819: out = 16'(2514);
			32820: out = 16'(1253);
			32821: out = 16'(-1487);
			32822: out = 16'(-3493);
			32823: out = 16'(-2023);
			32824: out = 16'(-278);
			32825: out = 16'(672);
			32826: out = 16'(-155);
			32827: out = 16'(423);
			32828: out = 16'(37);
			32829: out = 16'(1877);
			32830: out = 16'(2095);
			32831: out = 16'(111);
			32832: out = 16'(-3689);
			32833: out = 16'(-1239);
			32834: out = 16'(2100);
			32835: out = 16'(1035);
			32836: out = 16'(-609);
			32837: out = 16'(-211);
			32838: out = 16'(372);
			32839: out = 16'(-1374);
			32840: out = 16'(-1700);
			32841: out = 16'(-565);
			32842: out = 16'(1753);
			32843: out = 16'(2548);
			32844: out = 16'(1413);
			32845: out = 16'(410);
			32846: out = 16'(-613);
			32847: out = 16'(-815);
			32848: out = 16'(10);
			32849: out = 16'(495);
			32850: out = 16'(-927);
			32851: out = 16'(-1731);
			32852: out = 16'(431);
			32853: out = 16'(2267);
			32854: out = 16'(2129);
			32855: out = 16'(1033);
			32856: out = 16'(1530);
			32857: out = 16'(1113);
			32858: out = 16'(662);
			32859: out = 16'(-1133);
			32860: out = 16'(-1955);
			32861: out = 16'(-1708);
			32862: out = 16'(1075);
			32863: out = 16'(1388);
			32864: out = 16'(70);
			32865: out = 16'(-573);
			32866: out = 16'(-1350);
			32867: out = 16'(-1715);
			32868: out = 16'(-690);
			32869: out = 16'(1388);
			32870: out = 16'(2338);
			32871: out = 16'(1694);
			32872: out = 16'(1210);
			32873: out = 16'(1443);
			32874: out = 16'(9);
			32875: out = 16'(-1545);
			32876: out = 16'(-1274);
			32877: out = 16'(604);
			32878: out = 16'(-192);
			32879: out = 16'(-321);
			32880: out = 16'(-750);
			32881: out = 16'(-395);
			32882: out = 16'(-115);
			32883: out = 16'(16);
			32884: out = 16'(-115);
			32885: out = 16'(-182);
			32886: out = 16'(-695);
			32887: out = 16'(-857);
			32888: out = 16'(-1360);
			32889: out = 16'(-920);
			32890: out = 16'(782);
			32891: out = 16'(2450);
			32892: out = 16'(2741);
			32893: out = 16'(1358);
			32894: out = 16'(-412);
			32895: out = 16'(-1919);
			32896: out = 16'(-706);
			32897: out = 16'(187);
			32898: out = 16'(-347);
			32899: out = 16'(-926);
			32900: out = 16'(-804);
			32901: out = 16'(-172);
			32902: out = 16'(0);
			32903: out = 16'(383);
			32904: out = 16'(-1289);
			32905: out = 16'(-691);
			32906: out = 16'(200);
			32907: out = 16'(-177);
			32908: out = 16'(-2031);
			32909: out = 16'(-1139);
			32910: out = 16'(1298);
			32911: out = 16'(2172);
			32912: out = 16'(271);
			32913: out = 16'(-1114);
			32914: out = 16'(-1463);
			32915: out = 16'(-1310);
			32916: out = 16'(-386);
			32917: out = 16'(118);
			32918: out = 16'(1580);
			32919: out = 16'(2537);
			32920: out = 16'(2279);
			32921: out = 16'(-1538);
			32922: out = 16'(-2061);
			32923: out = 16'(0);
			32924: out = 16'(1027);
			32925: out = 16'(-841);
			32926: out = 16'(-2275);
			32927: out = 16'(-1497);
			32928: out = 16'(472);
			32929: out = 16'(2661);
			32930: out = 16'(1207);
			32931: out = 16'(-1402);
			32932: out = 16'(-2467);
			32933: out = 16'(333);
			32934: out = 16'(-113);
			32935: out = 16'(-819);
			32936: out = 16'(-421);
			32937: out = 16'(1373);
			32938: out = 16'(2302);
			32939: out = 16'(1553);
			32940: out = 16'(-32);
			32941: out = 16'(151);
			32942: out = 16'(-259);
			32943: out = 16'(340);
			32944: out = 16'(-1180);
			32945: out = 16'(-3122);
			32946: out = 16'(-1738);
			32947: out = 16'(1431);
			32948: out = 16'(2290);
			32949: out = 16'(1155);
			32950: out = 16'(1213);
			32951: out = 16'(896);
			32952: out = 16'(-1323);
			32953: out = 16'(-3143);
			32954: out = 16'(-837);
			32955: out = 16'(2614);
			32956: out = 16'(3280);
			32957: out = 16'(1900);
			32958: out = 16'(1094);
			32959: out = 16'(572);
			32960: out = 16'(-2451);
			32961: out = 16'(-4386);
			32962: out = 16'(-1807);
			32963: out = 16'(-421);
			32964: out = 16'(608);
			32965: out = 16'(222);
			32966: out = 16'(100);
			32967: out = 16'(-57);
			32968: out = 16'(-15);
			32969: out = 16'(700);
			32970: out = 16'(1619);
			32971: out = 16'(-126);
			32972: out = 16'(-1611);
			32973: out = 16'(-2977);
			32974: out = 16'(-1812);
			32975: out = 16'(1368);
			32976: out = 16'(1772);
			32977: out = 16'(1021);
			32978: out = 16'(555);
			32979: out = 16'(1321);
			32980: out = 16'(106);
			32981: out = 16'(4);
			32982: out = 16'(125);
			32983: out = 16'(396);
			32984: out = 16'(-918);
			32985: out = 16'(-313);
			32986: out = 16'(417);
			32987: out = 16'(831);
			32988: out = 16'(-62);
			32989: out = 16'(111);
			32990: out = 16'(-319);
			32991: out = 16'(-452);
			32992: out = 16'(-651);
			32993: out = 16'(176);
			32994: out = 16'(-1317);
			32995: out = 16'(-2038);
			32996: out = 16'(-243);
			32997: out = 16'(2502);
			32998: out = 16'(1365);
			32999: out = 16'(-404);
			33000: out = 16'(240);
			33001: out = 16'(1408);
			33002: out = 16'(959);
			33003: out = 16'(0);
			33004: out = 16'(-36);
			33005: out = 16'(-631);
			33006: out = 16'(-950);
			33007: out = 16'(-483);
			33008: out = 16'(598);
			33009: out = 16'(89);
			33010: out = 16'(-1660);
			33011: out = 16'(-3278);
			33012: out = 16'(-2570);
			33013: out = 16'(-289);
			33014: out = 16'(2989);
			33015: out = 16'(2782);
			33016: out = 16'(406);
			33017: out = 16'(-1341);
			33018: out = 16'(145);
			33019: out = 16'(1116);
			33020: out = 16'(758);
			33021: out = 16'(-107);
			33022: out = 16'(267);
			33023: out = 16'(-557);
			33024: out = 16'(-1809);
			33025: out = 16'(-2075);
			33026: out = 16'(77);
			33027: out = 16'(2169);
			33028: out = 16'(2890);
			33029: out = 16'(1617);
			33030: out = 16'(-203);
			33031: out = 16'(-4190);
			33032: out = 16'(-4296);
			33033: out = 16'(-1254);
			33034: out = 16'(1318);
			33035: out = 16'(1459);
			33036: out = 16'(1080);
			33037: out = 16'(1947);
			33038: out = 16'(2432);
			33039: out = 16'(655);
			33040: out = 16'(-2466);
			33041: out = 16'(-2604);
			33042: out = 16'(184);
			33043: out = 16'(1414);
			33044: out = 16'(-539);
			33045: out = 16'(-1318);
			33046: out = 16'(1201);
			33047: out = 16'(3009);
			33048: out = 16'(584);
			33049: out = 16'(-3348);
			33050: out = 16'(-3007);
			33051: out = 16'(1548);
			33052: out = 16'(1291);
			33053: out = 16'(352);
			33054: out = 16'(961);
			33055: out = 16'(3667);
			33056: out = 16'(2134);
			33057: out = 16'(239);
			33058: out = 16'(-2608);
			33059: out = 16'(-2978);
			33060: out = 16'(-1304);
			33061: out = 16'(990);
			33062: out = 16'(344);
			33063: out = 16'(-335);
			33064: out = 16'(1271);
			33065: out = 16'(3076);
			33066: out = 16'(1898);
			33067: out = 16'(-594);
			33068: out = 16'(-1580);
			33069: out = 16'(-2902);
			33070: out = 16'(-2804);
			33071: out = 16'(-1487);
			33072: out = 16'(597);
			33073: out = 16'(-68);
			33074: out = 16'(555);
			33075: out = 16'(1070);
			33076: out = 16'(1017);
			33077: out = 16'(-67);
			33078: out = 16'(-1548);
			33079: out = 16'(-1525);
			33080: out = 16'(-158);
			33081: out = 16'(-138);
			33082: out = 16'(497);
			33083: out = 16'(290);
			33084: out = 16'(714);
			33085: out = 16'(1142);
			33086: out = 16'(1345);
			33087: out = 16'(-162);
			33088: out = 16'(-1523);
			33089: out = 16'(-1869);
			33090: out = 16'(-619);
			33091: out = 16'(-245);
			33092: out = 16'(718);
			33093: out = 16'(1420);
			33094: out = 16'(-455);
			33095: out = 16'(-2034);
			33096: out = 16'(-1513);
			33097: out = 16'(481);
			33098: out = 16'(266);
			33099: out = 16'(1260);
			33100: out = 16'(791);
			33101: out = 16'(-38);
			33102: out = 16'(-1046);
			33103: out = 16'(-536);
			33104: out = 16'(-541);
			33105: out = 16'(-296);
			33106: out = 16'(-28);
			33107: out = 16'(-1177);
			33108: out = 16'(-1519);
			33109: out = 16'(-455);
			33110: out = 16'(1030);
			33111: out = 16'(55);
			33112: out = 16'(81);
			33113: out = 16'(524);
			33114: out = 16'(1503);
			33115: out = 16'(1061);
			33116: out = 16'(-852);
			33117: out = 16'(-3316);
			33118: out = 16'(-2799);
			33119: out = 16'(202);
			33120: out = 16'(3235);
			33121: out = 16'(1776);
			33122: out = 16'(-493);
			33123: out = 16'(-191);
			33124: out = 16'(1392);
			33125: out = 16'(873);
			33126: out = 16'(-456);
			33127: out = 16'(-154);
			33128: out = 16'(1422);
			33129: out = 16'(1548);
			33130: out = 16'(740);
			33131: out = 16'(277);
			33132: out = 16'(-83);
			33133: out = 16'(13);
			33134: out = 16'(-292);
			33135: out = 16'(-607);
			33136: out = 16'(-522);
			33137: out = 16'(-129);
			33138: out = 16'(46);
			33139: out = 16'(-63);
			33140: out = 16'(58);
			33141: out = 16'(-113);
			33142: out = 16'(104);
			33143: out = 16'(-396);
			33144: out = 16'(-900);
			33145: out = 16'(-681);
			33146: out = 16'(1496);
			33147: out = 16'(2723);
			33148: out = 16'(2637);
			33149: out = 16'(2582);
			33150: out = 16'(1887);
			33151: out = 16'(-396);
			33152: out = 16'(-3065);
			33153: out = 16'(-2808);
			33154: out = 16'(-2378);
			33155: out = 16'(-870);
			33156: out = 16'(375);
			33157: out = 16'(1171);
			33158: out = 16'(499);
			33159: out = 16'(26);
			33160: out = 16'(-55);
			33161: out = 16'(-359);
			33162: out = 16'(-2953);
			33163: out = 16'(-3670);
			33164: out = 16'(-1858);
			33165: out = 16'(911);
			33166: out = 16'(1172);
			33167: out = 16'(1394);
			33168: out = 16'(716);
			33169: out = 16'(-136);
			33170: out = 16'(18);
			33171: out = 16'(-580);
			33172: out = 16'(421);
			33173: out = 16'(1168);
			33174: out = 16'(-192);
			33175: out = 16'(-1496);
			33176: out = 16'(-1643);
			33177: out = 16'(29);
			33178: out = 16'(1686);
			33179: out = 16'(1731);
			33180: out = 16'(-209);
			33181: out = 16'(-2298);
			33182: out = 16'(-2433);
			33183: out = 16'(-213);
			33184: out = 16'(1923);
			33185: out = 16'(2132);
			33186: out = 16'(864);
			33187: out = 16'(98);
			33188: out = 16'(-155);
			33189: out = 16'(-285);
			33190: out = 16'(-659);
			33191: out = 16'(-444);
			33192: out = 16'(-202);
			33193: out = 16'(922);
			33194: out = 16'(2042);
			33195: out = 16'(2518);
			33196: out = 16'(-615);
			33197: out = 16'(-1813);
			33198: out = 16'(-1949);
			33199: out = 16'(-2031);
			33200: out = 16'(-2755);
			33201: out = 16'(-2583);
			33202: out = 16'(-1350);
			33203: out = 16'(755);
			33204: out = 16'(2690);
			33205: out = 16'(1318);
			33206: out = 16'(-536);
			33207: out = 16'(-617);
			33208: out = 16'(-79);
			33209: out = 16'(1639);
			33210: out = 16'(686);
			33211: out = 16'(541);
			33212: out = 16'(2458);
			33213: out = 16'(2808);
			33214: out = 16'(215);
			33215: out = 16'(-1998);
			33216: out = 16'(-1062);
			33217: out = 16'(870);
			33218: out = 16'(569);
			33219: out = 16'(-342);
			33220: out = 16'(92);
			33221: out = 16'(-193);
			33222: out = 16'(341);
			33223: out = 16'(156);
			33224: out = 16'(-242);
			33225: out = 16'(-1015);
			33226: out = 16'(695);
			33227: out = 16'(1453);
			33228: out = 16'(411);
			33229: out = 16'(-1540);
			33230: out = 16'(-2045);
			33231: out = 16'(-187);
			33232: out = 16'(1930);
			33233: out = 16'(1958);
			33234: out = 16'(-636);
			33235: out = 16'(-1356);
			33236: out = 16'(-473);
			33237: out = 16'(-465);
			33238: out = 16'(-3082);
			33239: out = 16'(-2643);
			33240: out = 16'(330);
			33241: out = 16'(3303);
			33242: out = 16'(3185);
			33243: out = 16'(1268);
			33244: out = 16'(-1166);
			33245: out = 16'(-1543);
			33246: out = 16'(213);
			33247: out = 16'(-1472);
			33248: out = 16'(-2506);
			33249: out = 16'(-1290);
			33250: out = 16'(1515);
			33251: out = 16'(2284);
			33252: out = 16'(982);
			33253: out = 16'(-417);
			33254: out = 16'(288);
			33255: out = 16'(502);
			33256: out = 16'(2086);
			33257: out = 16'(1539);
			33258: out = 16'(-287);
			33259: out = 16'(-1941);
			33260: out = 16'(-585);
			33261: out = 16'(-93);
			33262: out = 16'(-1109);
			33263: out = 16'(-2255);
			33264: out = 16'(1766);
			33265: out = 16'(2269);
			33266: out = 16'(-844);
			33267: out = 16'(-3003);
			33268: out = 16'(-425);
			33269: out = 16'(2198);
			33270: out = 16'(748);
			33271: out = 16'(-2809);
			33272: out = 16'(-4333);
			33273: out = 16'(102);
			33274: out = 16'(3388);
			33275: out = 16'(1837);
			33276: out = 16'(-598);
			33277: out = 16'(453);
			33278: out = 16'(3037);
			33279: out = 16'(2215);
			33280: out = 16'(-1447);
			33281: out = 16'(-4242);
			33282: out = 16'(-2248);
			33283: out = 16'(788);
			33284: out = 16'(955);
			33285: out = 16'(-952);
			33286: out = 16'(-1953);
			33287: out = 16'(-1435);
			33288: out = 16'(-241);
			33289: out = 16'(1115);
			33290: out = 16'(2153);
			33291: out = 16'(2065);
			33292: out = 16'(712);
			33293: out = 16'(-1345);
			33294: out = 16'(-1917);
			33295: out = 16'(-1571);
			33296: out = 16'(-726);
			33297: out = 16'(-609);
			33298: out = 16'(1051);
			33299: out = 16'(1260);
			33300: out = 16'(1170);
			33301: out = 16'(183);
			33302: out = 16'(1426);
			33303: out = 16'(-1072);
			33304: out = 16'(-2002);
			33305: out = 16'(314);
			33306: out = 16'(1461);
			33307: out = 16'(737);
			33308: out = 16'(536);
			33309: out = 16'(936);
			33310: out = 16'(-1323);
			33311: out = 16'(-3112);
			33312: out = 16'(-1696);
			33313: out = 16'(1565);
			33314: out = 16'(2205);
			33315: out = 16'(-552);
			33316: out = 16'(-1161);
			33317: out = 16'(400);
			33318: out = 16'(-336);
			33319: out = 16'(-1005);
			33320: out = 16'(-973);
			33321: out = 16'(1170);
			33322: out = 16'(2547);
			33323: out = 16'(1589);
			33324: out = 16'(-708);
			33325: out = 16'(-1198);
			33326: out = 16'(312);
			33327: out = 16'(1383);
			33328: out = 16'(-883);
			33329: out = 16'(-4089);
			33330: out = 16'(-3990);
			33331: out = 16'(-185);
			33332: out = 16'(1422);
			33333: out = 16'(-287);
			33334: out = 16'(-1680);
			33335: out = 16'(164);
			33336: out = 16'(3026);
			33337: out = 16'(1918);
			33338: out = 16'(-1025);
			33339: out = 16'(-1493);
			33340: out = 16'(1095);
			33341: out = 16'(1125);
			33342: out = 16'(-1496);
			33343: out = 16'(-3035);
			33344: out = 16'(-1230);
			33345: out = 16'(878);
			33346: out = 16'(944);
			33347: out = 16'(-71);
			33348: out = 16'(154);
			33349: out = 16'(2031);
			33350: out = 16'(3197);
			33351: out = 16'(1667);
			33352: out = 16'(-1899);
			33353: out = 16'(-2127);
			33354: out = 16'(-673);
			33355: out = 16'(488);
			33356: out = 16'(-60);
			33357: out = 16'(453);
			33358: out = 16'(410);
			33359: out = 16'(330);
			33360: out = 16'(-128);
			33361: out = 16'(-832);
			33362: out = 16'(-451);
			33363: out = 16'(691);
			33364: out = 16'(973);
			33365: out = 16'(-847);
			33366: out = 16'(-2444);
			33367: out = 16'(-2341);
			33368: out = 16'(-807);
			33369: out = 16'(64);
			33370: out = 16'(1222);
			33371: out = 16'(988);
			33372: out = 16'(382);
			33373: out = 16'(444);
			33374: out = 16'(-385);
			33375: out = 16'(-454);
			33376: out = 16'(-472);
			33377: out = 16'(-453);
			33378: out = 16'(-1297);
			33379: out = 16'(-128);
			33380: out = 16'(1034);
			33381: out = 16'(1108);
			33382: out = 16'(-778);
			33383: out = 16'(-259);
			33384: out = 16'(849);
			33385: out = 16'(1849);
			33386: out = 16'(1136);
			33387: out = 16'(1802);
			33388: out = 16'(298);
			33389: out = 16'(-1256);
			33390: out = 16'(-1368);
			33391: out = 16'(-163);
			33392: out = 16'(-1047);
			33393: out = 16'(-1484);
			33394: out = 16'(419);
			33395: out = 16'(1493);
			33396: out = 16'(1032);
			33397: out = 16'(668);
			33398: out = 16'(1737);
			33399: out = 16'(-83);
			33400: out = 16'(-233);
			33401: out = 16'(-849);
			33402: out = 16'(-825);
			33403: out = 16'(-596);
			33404: out = 16'(359);
			33405: out = 16'(263);
			33406: out = 16'(87);
			33407: out = 16'(447);
			33408: out = 16'(1136);
			33409: out = 16'(661);
			33410: out = 16'(-332);
			33411: out = 16'(-428);
			33412: out = 16'(-199);
			33413: out = 16'(124);
			33414: out = 16'(-775);
			33415: out = 16'(-1900);
			33416: out = 16'(-1487);
			33417: out = 16'(-358);
			33418: out = 16'(154);
			33419: out = 16'(186);
			33420: out = 16'(1245);
			33421: out = 16'(1342);
			33422: out = 16'(318);
			33423: out = 16'(-1525);
			33424: out = 16'(-2151);
			33425: out = 16'(-656);
			33426: out = 16'(1634);
			33427: out = 16'(1970);
			33428: out = 16'(-194);
			33429: out = 16'(-750);
			33430: out = 16'(-1057);
			33431: out = 16'(-743);
			33432: out = 16'(-307);
			33433: out = 16'(1585);
			33434: out = 16'(1682);
			33435: out = 16'(1689);
			33436: out = 16'(1229);
			33437: out = 16'(-1271);
			33438: out = 16'(-3204);
			33439: out = 16'(-3440);
			33440: out = 16'(-1652);
			33441: out = 16'(-538);
			33442: out = 16'(1174);
			33443: out = 16'(1532);
			33444: out = 16'(1780);
			33445: out = 16'(1046);
			33446: out = 16'(901);
			33447: out = 16'(-1656);
			33448: out = 16'(-2312);
			33449: out = 16'(387);
			33450: out = 16'(2502);
			33451: out = 16'(722);
			33452: out = 16'(-2357);
			33453: out = 16'(-2742);
			33454: out = 16'(959);
			33455: out = 16'(1540);
			33456: out = 16'(646);
			33457: out = 16'(-35);
			33458: out = 16'(-15);
			33459: out = 16'(-334);
			33460: out = 16'(-1406);
			33461: out = 16'(-2550);
			33462: out = 16'(-1436);
			33463: out = 16'(1436);
			33464: out = 16'(3945);
			33465: out = 16'(1950);
			33466: out = 16'(-2555);
			33467: out = 16'(-3921);
			33468: out = 16'(-571);
			33469: out = 16'(1498);
			33470: out = 16'(142);
			33471: out = 16'(157);
			33472: out = 16'(1638);
			33473: out = 16'(2431);
			33474: out = 16'(1004);
			33475: out = 16'(-1335);
			33476: out = 16'(-186);
			33477: out = 16'(284);
			33478: out = 16'(-203);
			33479: out = 16'(49);
			33480: out = 16'(1052);
			33481: out = 16'(603);
			33482: out = 16'(87);
			33483: out = 16'(1205);
			33484: out = 16'(-331);
			33485: out = 16'(-1888);
			33486: out = 16'(-1767);
			33487: out = 16'(485);
			33488: out = 16'(-1038);
			33489: out = 16'(-376);
			33490: out = 16'(984);
			33491: out = 16'(2350);
			33492: out = 16'(304);
			33493: out = 16'(-269);
			33494: out = 16'(-548);
			33495: out = 16'(403);
			33496: out = 16'(973);
			33497: out = 16'(-354);
			33498: out = 16'(-2163);
			33499: out = 16'(-1690);
			33500: out = 16'(367);
			33501: out = 16'(1628);
			33502: out = 16'(105);
			33503: out = 16'(-1432);
			33504: out = 16'(-1210);
			33505: out = 16'(287);
			33506: out = 16'(429);
			33507: out = 16'(871);
			33508: out = 16'(1535);
			33509: out = 16'(-22);
			33510: out = 16'(-460);
			33511: out = 16'(-350);
			33512: out = 16'(9);
			33513: out = 16'(-179);
			33514: out = 16'(-1987);
			33515: out = 16'(-1277);
			33516: out = 16'(1396);
			33517: out = 16'(2100);
			33518: out = 16'(1674);
			33519: out = 16'(-206);
			33520: out = 16'(252);
			33521: out = 16'(2346);
			33522: out = 16'(1294);
			33523: out = 16'(-1753);
			33524: out = 16'(-4371);
			33525: out = 16'(-3745);
			33526: out = 16'(-449);
			33527: out = 16'(1185);
			33528: out = 16'(867);
			33529: out = 16'(371);
			33530: out = 16'(-96);
			33531: out = 16'(134);
			33532: out = 16'(-982);
			33533: out = 16'(-2232);
			33534: out = 16'(-2742);
			33535: out = 16'(753);
			33536: out = 16'(1064);
			33537: out = 16'(91);
			33538: out = 16'(252);
			33539: out = 16'(1379);
			33540: out = 16'(744);
			33541: out = 16'(-799);
			33542: out = 16'(-1049);
			33543: out = 16'(-106);
			33544: out = 16'(1254);
			33545: out = 16'(1150);
			33546: out = 16'(131);
			33547: out = 16'(412);
			33548: out = 16'(210);
			33549: out = 16'(314);
			33550: out = 16'(-280);
			33551: out = 16'(-312);
			33552: out = 16'(-304);
			33553: out = 16'(1670);
			33554: out = 16'(2018);
			33555: out = 16'(-271);
			33556: out = 16'(-833);
			33557: out = 16'(244);
			33558: out = 16'(1493);
			33559: out = 16'(1176);
			33560: out = 16'(57);
			33561: out = 16'(-486);
			33562: out = 16'(-921);
			33563: out = 16'(-1367);
			33564: out = 16'(-543);
			33565: out = 16'(-151);
			33566: out = 16'(-42);
			33567: out = 16'(178);
			33568: out = 16'(1118);
			33569: out = 16'(1128);
			33570: out = 16'(272);
			33571: out = 16'(-1291);
			33572: out = 16'(-2669);
			33573: out = 16'(-1154);
			33574: out = 16'(-353);
			33575: out = 16'(764);
			33576: out = 16'(2256);
			33577: out = 16'(1152);
			33578: out = 16'(-733);
			33579: out = 16'(-2538);
			33580: out = 16'(-2175);
			33581: out = 16'(-195);
			33582: out = 16'(1073);
			33583: out = 16'(597);
			33584: out = 16'(33);
			33585: out = 16'(1188);
			33586: out = 16'(239);
			33587: out = 16'(-726);
			33588: out = 16'(-1450);
			33589: out = 16'(-1163);
			33590: out = 16'(-659);
			33591: out = 16'(126);
			33592: out = 16'(317);
			33593: out = 16'(75);
			33594: out = 16'(14);
			33595: out = 16'(803);
			33596: out = 16'(1335);
			33597: out = 16'(954);
			33598: out = 16'(81);
			33599: out = 16'(-1530);
			33600: out = 16'(-2646);
			33601: out = 16'(-2011);
			33602: out = 16'(343);
			33603: out = 16'(1175);
			33604: out = 16'(862);
			33605: out = 16'(544);
			33606: out = 16'(1202);
			33607: out = 16'(289);
			33608: out = 16'(-1242);
			33609: out = 16'(-2183);
			33610: out = 16'(-973);
			33611: out = 16'(-1052);
			33612: out = 16'(172);
			33613: out = 16'(484);
			33614: out = 16'(676);
			33615: out = 16'(1413);
			33616: out = 16'(1776);
			33617: out = 16'(460);
			33618: out = 16'(-1079);
			33619: out = 16'(-1274);
			33620: out = 16'(670);
			33621: out = 16'(821);
			33622: out = 16'(-138);
			33623: out = 16'(462);
			33624: out = 16'(323);
			33625: out = 16'(34);
			33626: out = 16'(-970);
			33627: out = 16'(-1665);
			33628: out = 16'(-1032);
			33629: out = 16'(-71);
			33630: out = 16'(525);
			33631: out = 16'(344);
			33632: out = 16'(-294);
			33633: out = 16'(-270);
			33634: out = 16'(1070);
			33635: out = 16'(2228);
			33636: out = 16'(1160);
			33637: out = 16'(-405);
			33638: out = 16'(-736);
			33639: out = 16'(400);
			33640: out = 16'(1008);
			33641: out = 16'(270);
			33642: out = 16'(305);
			33643: out = 16'(1760);
			33644: out = 16'(2225);
			33645: out = 16'(1489);
			33646: out = 16'(-667);
			33647: out = 16'(-1164);
			33648: out = 16'(50);
			33649: out = 16'(981);
			33650: out = 16'(231);
			33651: out = 16'(-300);
			33652: out = 16'(-94);
			33653: out = 16'(-106);
			33654: out = 16'(-1127);
			33655: out = 16'(-992);
			33656: out = 16'(319);
			33657: out = 16'(945);
			33658: out = 16'(203);
			33659: out = 16'(-478);
			33660: out = 16'(-495);
			33661: out = 16'(-29);
			33662: out = 16'(136);
			33663: out = 16'(1015);
			33664: out = 16'(1028);
			33665: out = 16'(-353);
			33666: out = 16'(-927);
			33667: out = 16'(-1116);
			33668: out = 16'(-1024);
			33669: out = 16'(-888);
			33670: out = 16'(-153);
			33671: out = 16'(1063);
			33672: out = 16'(975);
			33673: out = 16'(-679);
			33674: out = 16'(-2111);
			33675: out = 16'(-1455);
			33676: out = 16'(-233);
			33677: out = 16'(-180);
			33678: out = 16'(-401);
			33679: out = 16'(-1037);
			33680: out = 16'(811);
			33681: out = 16'(2916);
			33682: out = 16'(3133);
			33683: out = 16'(634);
			33684: out = 16'(-1067);
			33685: out = 16'(-1102);
			33686: out = 16'(179);
			33687: out = 16'(841);
			33688: out = 16'(662);
			33689: out = 16'(-702);
			33690: out = 16'(-1183);
			33691: out = 16'(187);
			33692: out = 16'(1044);
			33693: out = 16'(84);
			33694: out = 16'(-1147);
			33695: out = 16'(-560);
			33696: out = 16'(-1939);
			33697: out = 16'(-2492);
			33698: out = 16'(-1254);
			33699: out = 16'(1342);
			33700: out = 16'(2099);
			33701: out = 16'(1768);
			33702: out = 16'(1369);
			33703: out = 16'(1308);
			33704: out = 16'(1126);
			33705: out = 16'(-2109);
			33706: out = 16'(-4107);
			33707: out = 16'(-2138);
			33708: out = 16'(1149);
			33709: out = 16'(2293);
			33710: out = 16'(1553);
			33711: out = 16'(945);
			33712: out = 16'(126);
			33713: out = 16'(125);
			33714: out = 16'(-1367);
			33715: out = 16'(-2467);
			33716: out = 16'(-2123);
			33717: out = 16'(-312);
			33718: out = 16'(68);
			33719: out = 16'(62);
			33720: out = 16'(419);
			33721: out = 16'(347);
			33722: out = 16'(103);
			33723: out = 16'(-375);
			33724: out = 16'(-936);
			33725: out = 16'(360);
			33726: out = 16'(-78);
			33727: out = 16'(721);
			33728: out = 16'(1451);
			33729: out = 16'(1099);
			33730: out = 16'(-1319);
			33731: out = 16'(-1114);
			33732: out = 16'(475);
			33733: out = 16'(1024);
			33734: out = 16'(117);
			33735: out = 16'(-87);
			33736: out = 16'(-764);
			33737: out = 16'(-2179);
			33738: out = 16'(-229);
			33739: out = 16'(1583);
			33740: out = 16'(1466);
			33741: out = 16'(-994);
			33742: out = 16'(-713);
			33743: out = 16'(-492);
			33744: out = 16'(230);
			33745: out = 16'(-352);
			33746: out = 16'(-238);
			33747: out = 16'(682);
			33748: out = 16'(3172);
			33749: out = 16'(3353);
			33750: out = 16'(868);
			33751: out = 16'(-1982);
			33752: out = 16'(-1538);
			33753: out = 16'(-436);
			33754: out = 16'(-733);
			33755: out = 16'(-1809);
			33756: out = 16'(-45);
			33757: out = 16'(1186);
			33758: out = 16'(-168);
			33759: out = 16'(-1570);
			33760: out = 16'(-647);
			33761: out = 16'(996);
			33762: out = 16'(601);
			33763: out = 16'(-815);
			33764: out = 16'(-2486);
			33765: out = 16'(-1990);
			33766: out = 16'(-186);
			33767: out = 16'(1462);
			33768: out = 16'(322);
			33769: out = 16'(-450);
			33770: out = 16'(28);
			33771: out = 16'(1591);
			33772: out = 16'(1123);
			33773: out = 16'(-289);
			33774: out = 16'(-2064);
			33775: out = 16'(-1801);
			33776: out = 16'(-400);
			33777: out = 16'(1679);
			33778: out = 16'(610);
			33779: out = 16'(-1630);
			33780: out = 16'(-1727);
			33781: out = 16'(236);
			33782: out = 16'(437);
			33783: out = 16'(-637);
			33784: out = 16'(93);
			33785: out = 16'(918);
			33786: out = 16'(718);
			33787: out = 16'(-346);
			33788: out = 16'(-452);
			33789: out = 16'(-1653);
			33790: out = 16'(-1763);
			33791: out = 16'(-1192);
			33792: out = 16'(323);
			33793: out = 16'(-47);
			33794: out = 16'(951);
			33795: out = 16'(1300);
			33796: out = 16'(1005);
			33797: out = 16'(-427);
			33798: out = 16'(174);
			33799: out = 16'(414);
			33800: out = 16'(-808);
			33801: out = 16'(-4475);
			33802: out = 16'(-3011);
			33803: out = 16'(-1141);
			33804: out = 16'(1308);
			33805: out = 16'(3661);
			33806: out = 16'(3729);
			33807: out = 16'(1743);
			33808: out = 16'(-384);
			33809: out = 16'(-1464);
			33810: out = 16'(-2872);
			33811: out = 16'(-2407);
			33812: out = 16'(-34);
			33813: out = 16'(2776);
			33814: out = 16'(3409);
			33815: out = 16'(2740);
			33816: out = 16'(1145);
			33817: out = 16'(-448);
			33818: out = 16'(-1256);
			33819: out = 16'(-1800);
			33820: out = 16'(-1269);
			33821: out = 16'(-870);
			33822: out = 16'(-738);
			33823: out = 16'(-199);
			33824: out = 16'(931);
			33825: out = 16'(743);
			33826: out = 16'(-467);
			33827: out = 16'(-952);
			33828: out = 16'(1230);
			33829: out = 16'(2181);
			33830: out = 16'(809);
			33831: out = 16'(-365);
			33832: out = 16'(588);
			33833: out = 16'(1029);
			33834: out = 16'(39);
			33835: out = 16'(-418);
			33836: out = 16'(103);
			33837: out = 16'(72);
			33838: out = 16'(-859);
			33839: out = 16'(-1266);
			33840: out = 16'(-1038);
			33841: out = 16'(-403);
			33842: out = 16'(518);
			33843: out = 16'(1519);
			33844: out = 16'(1568);
			33845: out = 16'(507);
			33846: out = 16'(-57);
			33847: out = 16'(169);
			33848: out = 16'(-1237);
			33849: out = 16'(-1506);
			33850: out = 16'(-353);
			33851: out = 16'(1406);
			33852: out = 16'(1382);
			33853: out = 16'(399);
			33854: out = 16'(-255);
			33855: out = 16'(-122);
			33856: out = 16'(-647);
			33857: out = 16'(-159);
			33858: out = 16'(-103);
			33859: out = 16'(76);
			33860: out = 16'(434);
			33861: out = 16'(1865);
			33862: out = 16'(1769);
			33863: out = 16'(-385);
			33864: out = 16'(-3222);
			33865: out = 16'(-1541);
			33866: out = 16'(506);
			33867: out = 16'(1707);
			33868: out = 16'(664);
			33869: out = 16'(133);
			33870: out = 16'(-1655);
			33871: out = 16'(-865);
			33872: out = 16'(452);
			33873: out = 16'(-95);
			33874: out = 16'(-1104);
			33875: out = 16'(-826);
			33876: out = 16'(504);
			33877: out = 16'(1448);
			33878: out = 16'(1478);
			33879: out = 16'(1264);
			33880: out = 16'(667);
			33881: out = 16'(-214);
			33882: out = 16'(-1738);
			33883: out = 16'(-610);
			33884: out = 16'(273);
			33885: out = 16'(-1099);
			33886: out = 16'(-3221);
			33887: out = 16'(-2161);
			33888: out = 16'(1359);
			33889: out = 16'(3541);
			33890: out = 16'(2445);
			33891: out = 16'(-413);
			33892: out = 16'(-1889);
			33893: out = 16'(-561);
			33894: out = 16'(1260);
			33895: out = 16'(59);
			33896: out = 16'(-2105);
			33897: out = 16'(-1808);
			33898: out = 16'(1429);
			33899: out = 16'(2278);
			33900: out = 16'(1754);
			33901: out = 16'(418);
			33902: out = 16'(-171);
			33903: out = 16'(-641);
			33904: out = 16'(-1178);
			33905: out = 16'(-1439);
			33906: out = 16'(-710);
			33907: out = 16'(-211);
			33908: out = 16'(941);
			33909: out = 16'(568);
			33910: out = 16'(-144);
			33911: out = 16'(292);
			33912: out = 16'(1185);
			33913: out = 16'(958);
			33914: out = 16'(-389);
			33915: out = 16'(-951);
			33916: out = 16'(-1885);
			33917: out = 16'(-1095);
			33918: out = 16'(-2);
			33919: out = 16'(1207);
			33920: out = 16'(-186);
			33921: out = 16'(365);
			33922: out = 16'(-681);
			33923: out = 16'(-1719);
			33924: out = 16'(-703);
			33925: out = 16'(1748);
			33926: out = 16'(617);
			33927: out = 16'(-2407);
			33928: out = 16'(-1996);
			33929: out = 16'(-577);
			33930: out = 16'(292);
			33931: out = 16'(-153);
			33932: out = 16'(73);
			33933: out = 16'(-833);
			33934: out = 16'(-1158);
			33935: out = 16'(-990);
			33936: out = 16'(265);
			33937: out = 16'(294);
			33938: out = 16'(987);
			33939: out = 16'(1543);
			33940: out = 16'(2260);
			33941: out = 16'(1348);
			33942: out = 16'(523);
			33943: out = 16'(-1047);
			33944: out = 16'(-2026);
			33945: out = 16'(-3127);
			33946: out = 16'(1477);
			33947: out = 16'(2491);
			33948: out = 16'(481);
			33949: out = 16'(-1709);
			33950: out = 16'(5);
			33951: out = 16'(506);
			33952: out = 16'(112);
			33953: out = 16'(81);
			33954: out = 16'(1000);
			33955: out = 16'(694);
			33956: out = 16'(110);
			33957: out = 16'(-188);
			33958: out = 16'(-1289);
			33959: out = 16'(-942);
			33960: out = 16'(729);
			33961: out = 16'(2445);
			33962: out = 16'(2367);
			33963: out = 16'(1398);
			33964: out = 16'(550);
			33965: out = 16'(-303);
			33966: out = 16'(-2523);
			33967: out = 16'(-2981);
			33968: out = 16'(-3130);
			33969: out = 16'(-1838);
			33970: out = 16'(381);
			33971: out = 16'(3121);
			33972: out = 16'(3151);
			33973: out = 16'(1401);
			33974: out = 16'(-279);
			33975: out = 16'(-593);
			33976: out = 16'(-1205);
			33977: out = 16'(-1290);
			33978: out = 16'(-92);
			33979: out = 16'(821);
			33980: out = 16'(1145);
			33981: out = 16'(-1544);
			33982: out = 16'(-3556);
			33983: out = 16'(-1067);
			33984: out = 16'(1528);
			33985: out = 16'(1985);
			33986: out = 16'(433);
			33987: out = 16'(183);
			33988: out = 16'(717);
			33989: out = 16'(1411);
			33990: out = 16'(-190);
			33991: out = 16'(-2524);
			33992: out = 16'(-3587);
			33993: out = 16'(-1213);
			33994: out = 16'(838);
			33995: out = 16'(892);
			33996: out = 16'(-398);
			33997: out = 16'(90);
			33998: out = 16'(837);
			33999: out = 16'(1164);
			34000: out = 16'(1057);
			34001: out = 16'(-141);
			34002: out = 16'(-1144);
			34003: out = 16'(-987);
			34004: out = 16'(19);
			34005: out = 16'(46);
			34006: out = 16'(-99);
			34007: out = 16'(529);
			34008: out = 16'(1397);
			34009: out = 16'(152);
			34010: out = 16'(-1058);
			34011: out = 16'(-794);
			34012: out = 16'(554);
			34013: out = 16'(237);
			34014: out = 16'(-590);
			34015: out = 16'(-586);
			34016: out = 16'(566);
			34017: out = 16'(211);
			34018: out = 16'(240);
			34019: out = 16'(-649);
			34020: out = 16'(-705);
			34021: out = 16'(-28);
			34022: out = 16'(57);
			34023: out = 16'(-124);
			34024: out = 16'(468);
			34025: out = 16'(1505);
			34026: out = 16'(1514);
			34027: out = 16'(-523);
			34028: out = 16'(-2823);
			34029: out = 16'(-3334);
			34030: out = 16'(-1852);
			34031: out = 16'(-396);
			34032: out = 16'(650);
			34033: out = 16'(1382);
			34034: out = 16'(1524);
			34035: out = 16'(2326);
			34036: out = 16'(2501);
			34037: out = 16'(1504);
			34038: out = 16'(-765);
			34039: out = 16'(-3446);
			34040: out = 16'(-3949);
			34041: out = 16'(-1816);
			34042: out = 16'(613);
			34043: out = 16'(2517);
			34044: out = 16'(1699);
			34045: out = 16'(1059);
			34046: out = 16'(980);
			34047: out = 16'(92);
			34048: out = 16'(-1927);
			34049: out = 16'(-2438);
			34050: out = 16'(-842);
			34051: out = 16'(-127);
			34052: out = 16'(169);
			34053: out = 16'(-222);
			34054: out = 16'(-675);
			34055: out = 16'(-1704);
			34056: out = 16'(-231);
			34057: out = 16'(732);
			34058: out = 16'(1590);
			34059: out = 16'(2126);
			34060: out = 16'(350);
			34061: out = 16'(-1382);
			34062: out = 16'(-2419);
			34063: out = 16'(-1840);
			34064: out = 16'(-674);
			34065: out = 16'(1531);
			34066: out = 16'(2621);
			34067: out = 16'(2260);
			34068: out = 16'(32);
			34069: out = 16'(841);
			34070: out = 16'(778);
			34071: out = 16'(-518);
			34072: out = 16'(-1671);
			34073: out = 16'(-889);
			34074: out = 16'(459);
			34075: out = 16'(1378);
			34076: out = 16'(1282);
			34077: out = 16'(-801);
			34078: out = 16'(-1780);
			34079: out = 16'(17);
			34080: out = 16'(2443);
			34081: out = 16'(311);
			34082: out = 16'(-1447);
			34083: out = 16'(-703);
			34084: out = 16'(1736);
			34085: out = 16'(975);
			34086: out = 16'(-858);
			34087: out = 16'(-2267);
			34088: out = 16'(-1235);
			34089: out = 16'(-195);
			34090: out = 16'(1356);
			34091: out = 16'(976);
			34092: out = 16'(-65);
			34093: out = 16'(-1431);
			34094: out = 16'(-1245);
			34095: out = 16'(-1687);
			34096: out = 16'(-1131);
			34097: out = 16'(523);
			34098: out = 16'(1156);
			34099: out = 16'(501);
			34100: out = 16'(-109);
			34101: out = 16'(88);
			34102: out = 16'(9);
			34103: out = 16'(-320);
			34104: out = 16'(-211);
			34105: out = 16'(311);
			34106: out = 16'(-941);
			34107: out = 16'(754);
			34108: out = 16'(1369);
			34109: out = 16'(691);
			34110: out = 16'(-884);
			34111: out = 16'(-161);
			34112: out = 16'(126);
			34113: out = 16'(-353);
			34114: out = 16'(-1273);
			34115: out = 16'(-91);
			34116: out = 16'(121);
			34117: out = 16'(-148);
			34118: out = 16'(-393);
			34119: out = 16'(295);
			34120: out = 16'(947);
			34121: out = 16'(1271);
			34122: out = 16'(940);
			34123: out = 16'(42);
			34124: out = 16'(-1317);
			34125: out = 16'(-1948);
			34126: out = 16'(-1225);
			34127: out = 16'(487);
			34128: out = 16'(1079);
			34129: out = 16'(1238);
			34130: out = 16'(882);
			34131: out = 16'(-27);
			34132: out = 16'(1029);
			34133: out = 16'(532);
			34134: out = 16'(-587);
			34135: out = 16'(-1231);
			34136: out = 16'(254);
			34137: out = 16'(903);
			34138: out = 16'(1333);
			34139: out = 16'(1266);
			34140: out = 16'(-12);
			34141: out = 16'(-743);
			34142: out = 16'(-1203);
			34143: out = 16'(-1461);
			34144: out = 16'(-1712);
			34145: out = 16'(-408);
			34146: out = 16'(776);
			34147: out = 16'(1021);
			34148: out = 16'(404);
			34149: out = 16'(1277);
			34150: out = 16'(1616);
			34151: out = 16'(696);
			34152: out = 16'(-1215);
			34153: out = 16'(-1719);
			34154: out = 16'(-821);
			34155: out = 16'(654);
			34156: out = 16'(942);
			34157: out = 16'(480);
			34158: out = 16'(-715);
			34159: out = 16'(-671);
			34160: out = 16'(-117);
			34161: out = 16'(-562);
			34162: out = 16'(-543);
			34163: out = 16'(-244);
			34164: out = 16'(-144);
			34165: out = 16'(-992);
			34166: out = 16'(-1612);
			34167: out = 16'(-893);
			34168: out = 16'(693);
			34169: out = 16'(1040);
			34170: out = 16'(1697);
			34171: out = 16'(-374);
			34172: out = 16'(-1343);
			34173: out = 16'(-115);
			34174: out = 16'(962);
			34175: out = 16'(733);
			34176: out = 16'(32);
			34177: out = 16'(-110);
			34178: out = 16'(-621);
			34179: out = 16'(-409);
			34180: out = 16'(-985);
			34181: out = 16'(-1245);
			34182: out = 16'(-834);
			34183: out = 16'(1169);
			34184: out = 16'(1512);
			34185: out = 16'(758);
			34186: out = 16'(-40);
			34187: out = 16'(280);
			34188: out = 16'(-196);
			34189: out = 16'(-858);
			34190: out = 16'(-1302);
			34191: out = 16'(-485);
			34192: out = 16'(-26);
			34193: out = 16'(847);
			34194: out = 16'(947);
			34195: out = 16'(135);
			34196: out = 16'(-880);
			34197: out = 16'(72);
			34198: out = 16'(1150);
			34199: out = 16'(292);
			34200: out = 16'(-2162);
			34201: out = 16'(-1454);
			34202: out = 16'(1327);
			34203: out = 16'(1949);
			34204: out = 16'(1485);
			34205: out = 16'(-82);
			34206: out = 16'(-499);
			34207: out = 16'(-138);
			34208: out = 16'(-25);
			34209: out = 16'(-837);
			34210: out = 16'(-1459);
			34211: out = 16'(-803);
			34212: out = 16'(1239);
			34213: out = 16'(1258);
			34214: out = 16'(524);
			34215: out = 16'(374);
			34216: out = 16'(930);
			34217: out = 16'(1335);
			34218: out = 16'(320);
			34219: out = 16'(-938);
			34220: out = 16'(-1200);
			34221: out = 16'(956);
			34222: out = 16'(660);
			34223: out = 16'(-624);
			34224: out = 16'(-702);
			34225: out = 16'(729);
			34226: out = 16'(444);
			34227: out = 16'(-771);
			34228: out = 16'(-1235);
			34229: out = 16'(-1027);
			34230: out = 16'(-571);
			34231: out = 16'(-381);
			34232: out = 16'(268);
			34233: out = 16'(879);
			34234: out = 16'(1422);
			34235: out = 16'(551);
			34236: out = 16'(-332);
			34237: out = 16'(-989);
			34238: out = 16'(-452);
			34239: out = 16'(-1292);
			34240: out = 16'(-1248);
			34241: out = 16'(280);
			34242: out = 16'(2954);
			34243: out = 16'(1269);
			34244: out = 16'(-908);
			34245: out = 16'(-1037);
			34246: out = 16'(162);
			34247: out = 16'(-221);
			34248: out = 16'(-451);
			34249: out = 16'(45);
			34250: out = 16'(-126);
			34251: out = 16'(132);
			34252: out = 16'(611);
			34253: out = 16'(763);
			34254: out = 16'(-616);
			34255: out = 16'(124);
			34256: out = 16'(361);
			34257: out = 16'(-479);
			34258: out = 16'(-2568);
			34259: out = 16'(-280);
			34260: out = 16'(471);
			34261: out = 16'(492);
			34262: out = 16'(-193);
			34263: out = 16'(15);
			34264: out = 16'(-135);
			34265: out = 16'(43);
			34266: out = 16'(-267);
			34267: out = 16'(-750);
			34268: out = 16'(-436);
			34269: out = 16'(1124);
			34270: out = 16'(1688);
			34271: out = 16'(-173);
			34272: out = 16'(-1429);
			34273: out = 16'(-924);
			34274: out = 16'(240);
			34275: out = 16'(-221);
			34276: out = 16'(-269);
			34277: out = 16'(-640);
			34278: out = 16'(-193);
			34279: out = 16'(67);
			34280: out = 16'(1990);
			34281: out = 16'(607);
			34282: out = 16'(-725);
			34283: out = 16'(-1178);
			34284: out = 16'(300);
			34285: out = 16'(-152);
			34286: out = 16'(602);
			34287: out = 16'(1194);
			34288: out = 16'(-103);
			34289: out = 16'(-1390);
			34290: out = 16'(-1181);
			34291: out = 16'(-450);
			34292: out = 16'(-1364);
			34293: out = 16'(-1131);
			34294: out = 16'(-841);
			34295: out = 16'(-57);
			34296: out = 16'(604);
			34297: out = 16'(2732);
			34298: out = 16'(2127);
			34299: out = 16'(-66);
			34300: out = 16'(-2162);
			34301: out = 16'(-852);
			34302: out = 16'(-599);
			34303: out = 16'(-131);
			34304: out = 16'(531);
			34305: out = 16'(1389);
			34306: out = 16'(2783);
			34307: out = 16'(2816);
			34308: out = 16'(976);
			34309: out = 16'(-1318);
			34310: out = 16'(-835);
			34311: out = 16'(-170);
			34312: out = 16'(-688);
			34313: out = 16'(-1549);
			34314: out = 16'(625);
			34315: out = 16'(1811);
			34316: out = 16'(1240);
			34317: out = 16'(-309);
			34318: out = 16'(-77);
			34319: out = 16'(-159);
			34320: out = 16'(-281);
			34321: out = 16'(-633);
			34322: out = 16'(-544);
			34323: out = 16'(-318);
			34324: out = 16'(-133);
			34325: out = 16'(-204);
			34326: out = 16'(-4);
			34327: out = 16'(690);
			34328: out = 16'(1244);
			34329: out = 16'(964);
			34330: out = 16'(68);
			34331: out = 16'(-1529);
			34332: out = 16'(-1441);
			34333: out = 16'(-452);
			34334: out = 16'(100);
			34335: out = 16'(-461);
			34336: out = 16'(-110);
			34337: out = 16'(680);
			34338: out = 16'(801);
			34339: out = 16'(342);
			34340: out = 16'(-1015);
			34341: out = 16'(-767);
			34342: out = 16'(838);
			34343: out = 16'(2105);
			34344: out = 16'(1284);
			34345: out = 16'(202);
			34346: out = 16'(-313);
			34347: out = 16'(-688);
			34348: out = 16'(-1272);
			34349: out = 16'(-1047);
			34350: out = 16'(-265);
			34351: out = 16'(-212);
			34352: out = 16'(-10);
			34353: out = 16'(-522);
			34354: out = 16'(-334);
			34355: out = 16'(-209);
			34356: out = 16'(-425);
			34357: out = 16'(-1856);
			34358: out = 16'(-1195);
			34359: out = 16'(872);
			34360: out = 16'(1831);
			34361: out = 16'(445);
			34362: out = 16'(-731);
			34363: out = 16'(-733);
			34364: out = 16'(-31);
			34365: out = 16'(-153);
			34366: out = 16'(28);
			34367: out = 16'(-495);
			34368: out = 16'(-1171);
			34369: out = 16'(-296);
			34370: out = 16'(2146);
			34371: out = 16'(2830);
			34372: out = 16'(591);
			34373: out = 16'(-1448);
			34374: out = 16'(-1449);
			34375: out = 16'(-357);
			34376: out = 16'(-189);
			34377: out = 16'(22);
			34378: out = 16'(-256);
			34379: out = 16'(710);
			34380: out = 16'(992);
			34381: out = 16'(-717);
			34382: out = 16'(-1179);
			34383: out = 16'(-1235);
			34384: out = 16'(-586);
			34385: out = 16'(21);
			34386: out = 16'(1196);
			34387: out = 16'(1332);
			34388: out = 16'(1193);
			34389: out = 16'(737);
			34390: out = 16'(-29);
			34391: out = 16'(-551);
			34392: out = 16'(-379);
			34393: out = 16'(-186);
			34394: out = 16'(-556);
			34395: out = 16'(-1218);
			34396: out = 16'(-803);
			34397: out = 16'(283);
			34398: out = 16'(923);
			34399: out = 16'(986);
			34400: out = 16'(597);
			34401: out = 16'(-514);
			34402: out = 16'(-2198);
			34403: out = 16'(-1041);
			34404: out = 16'(-367);
			34405: out = 16'(341);
			34406: out = 16'(1093);
			34407: out = 16'(908);
			34408: out = 16'(1064);
			34409: out = 16'(341);
			34410: out = 16'(-789);
			34411: out = 16'(-1304);
			34412: out = 16'(-137);
			34413: out = 16'(273);
			34414: out = 16'(-239);
			34415: out = 16'(18);
			34416: out = 16'(-176);
			34417: out = 16'(-194);
			34418: out = 16'(-961);
			34419: out = 16'(-1574);
			34420: out = 16'(-767);
			34421: out = 16'(576);
			34422: out = 16'(895);
			34423: out = 16'(234);
			34424: out = 16'(295);
			34425: out = 16'(-617);
			34426: out = 16'(-2266);
			34427: out = 16'(-2993);
			34428: out = 16'(-534);
			34429: out = 16'(827);
			34430: out = 16'(710);
			34431: out = 16'(-209);
			34432: out = 16'(173);
			34433: out = 16'(1825);
			34434: out = 16'(2039);
			34435: out = 16'(95);
			34436: out = 16'(-1028);
			34437: out = 16'(-1259);
			34438: out = 16'(593);
			34439: out = 16'(244);
			34440: out = 16'(-1653);
			34441: out = 16'(-1032);
			34442: out = 16'(1759);
			34443: out = 16'(2935);
			34444: out = 16'(1503);
			34445: out = 16'(46);
			34446: out = 16'(-1201);
			34447: out = 16'(-2959);
			34448: out = 16'(-3858);
			34449: out = 16'(-625);
			34450: out = 16'(677);
			34451: out = 16'(1319);
			34452: out = 16'(1058);
			34453: out = 16'(1516);
			34454: out = 16'(1838);
			34455: out = 16'(1788);
			34456: out = 16'(458);
			34457: out = 16'(-1445);
			34458: out = 16'(-1587);
			34459: out = 16'(-2022);
			34460: out = 16'(-1413);
			34461: out = 16'(413);
			34462: out = 16'(2164);
			34463: out = 16'(1579);
			34464: out = 16'(363);
			34465: out = 16'(-21);
			34466: out = 16'(-123);
			34467: out = 16'(76);
			34468: out = 16'(-706);
			34469: out = 16'(-1043);
			34470: out = 16'(436);
			34471: out = 16'(1892);
			34472: out = 16'(2537);
			34473: out = 16'(1497);
			34474: out = 16'(-320);
			34475: out = 16'(-1954);
			34476: out = 16'(-1780);
			34477: out = 16'(-768);
			34478: out = 16'(-11);
			34479: out = 16'(-83);
			34480: out = 16'(162);
			34481: out = 16'(552);
			34482: out = 16'(1059);
			34483: out = 16'(821);
			34484: out = 16'(-1140);
			34485: out = 16'(-3370);
			34486: out = 16'(-2949);
			34487: out = 16'(-1);
			34488: out = 16'(2134);
			34489: out = 16'(1096);
			34490: out = 16'(-326);
			34491: out = 16'(338);
			34492: out = 16'(302);
			34493: out = 16'(-401);
			34494: out = 16'(-691);
			34495: out = 16'(322);
			34496: out = 16'(-512);
			34497: out = 16'(-501);
			34498: out = 16'(-168);
			34499: out = 16'(367);
			34500: out = 16'(-49);
			34501: out = 16'(205);
			34502: out = 16'(674);
			34503: out = 16'(926);
			34504: out = 16'(257);
			34505: out = 16'(-352);
			34506: out = 16'(-569);
			34507: out = 16'(-588);
			34508: out = 16'(-904);
			34509: out = 16'(-1213);
			34510: out = 16'(-786);
			34511: out = 16'(-583);
			34512: out = 16'(-1167);
			34513: out = 16'(202);
			34514: out = 16'(1431);
			34515: out = 16'(2266);
			34516: out = 16'(1670);
			34517: out = 16'(454);
			34518: out = 16'(166);
			34519: out = 16'(14);
			34520: out = 16'(-1715);
			34521: out = 16'(-3926);
			34522: out = 16'(-3842);
			34523: out = 16'(-660);
			34524: out = 16'(1969);
			34525: out = 16'(2039);
			34526: out = 16'(1462);
			34527: out = 16'(1809);
			34528: out = 16'(1509);
			34529: out = 16'(-417);
			34530: out = 16'(-3306);
			34531: out = 16'(-3196);
			34532: out = 16'(-1535);
			34533: out = 16'(-93);
			34534: out = 16'(994);
			34535: out = 16'(2530);
			34536: out = 16'(2479);
			34537: out = 16'(972);
			34538: out = 16'(418);
			34539: out = 16'(-57);
			34540: out = 16'(-239);
			34541: out = 16'(-724);
			34542: out = 16'(-1274);
			34543: out = 16'(-1237);
			34544: out = 16'(-694);
			34545: out = 16'(848);
			34546: out = 16'(2279);
			34547: out = 16'(2502);
			34548: out = 16'(211);
			34549: out = 16'(-837);
			34550: out = 16'(453);
			34551: out = 16'(-155);
			34552: out = 16'(-1092);
			34553: out = 16'(-1683);
			34554: out = 16'(-363);
			34555: out = 16'(837);
			34556: out = 16'(1896);
			34557: out = 16'(1538);
			34558: out = 16'(392);
			34559: out = 16'(-1774);
			34560: out = 16'(-1703);
			34561: out = 16'(-1222);
			34562: out = 16'(399);
			34563: out = 16'(2341);
			34564: out = 16'(2322);
			34565: out = 16'(1449);
			34566: out = 16'(503);
			34567: out = 16'(-362);
			34568: out = 16'(-1578);
			34569: out = 16'(-2439);
			34570: out = 16'(-1853);
			34571: out = 16'(-218);
			34572: out = 16'(-141);
			34573: out = 16'(763);
			34574: out = 16'(1092);
			34575: out = 16'(693);
			34576: out = 16'(-541);
			34577: out = 16'(-170);
			34578: out = 16'(-53);
			34579: out = 16'(-132);
			34580: out = 16'(-33);
			34581: out = 16'(188);
			34582: out = 16'(144);
			34583: out = 16'(-337);
			34584: out = 16'(-446);
			34585: out = 16'(-205);
			34586: out = 16'(75);
			34587: out = 16'(-729);
			34588: out = 16'(-1758);
			34589: out = 16'(-2104);
			34590: out = 16'(447);
			34591: out = 16'(1197);
			34592: out = 16'(-865);
			34593: out = 16'(-3014);
			34594: out = 16'(-1881);
			34595: out = 16'(-170);
			34596: out = 16'(-192);
			34597: out = 16'(-542);
			34598: out = 16'(44);
			34599: out = 16'(2306);
			34600: out = 16'(2982);
			34601: out = 16'(1011);
			34602: out = 16'(-833);
			34603: out = 16'(-2361);
			34604: out = 16'(-2930);
			34605: out = 16'(-2335);
			34606: out = 16'(-73);
			34607: out = 16'(1898);
			34608: out = 16'(2264);
			34609: out = 16'(1047);
			34610: out = 16'(100);
			34611: out = 16'(173);
			34612: out = 16'(852);
			34613: out = 16'(853);
			34614: out = 16'(-29);
			34615: out = 16'(261);
			34616: out = 16'(-476);
			34617: out = 16'(-1304);
			34618: out = 16'(-150);
			34619: out = 16'(-284);
			34620: out = 16'(958);
			34621: out = 16'(230);
			34622: out = 16'(-1064);
			34623: out = 16'(816);
			34624: out = 16'(2000);
			34625: out = 16'(835);
			34626: out = 16'(-954);
			34627: out = 16'(243);
			34628: out = 16'(1638);
			34629: out = 16'(1344);
			34630: out = 16'(-30);
			34631: out = 16'(-43);
			34632: out = 16'(-95);
			34633: out = 16'(-739);
			34634: out = 16'(-1146);
			34635: out = 16'(78);
			34636: out = 16'(-116);
			34637: out = 16'(-521);
			34638: out = 16'(-914);
			34639: out = 16'(-358);
			34640: out = 16'(-214);
			34641: out = 16'(653);
			34642: out = 16'(1488);
			34643: out = 16'(1742);
			34644: out = 16'(-43);
			34645: out = 16'(-492);
			34646: out = 16'(-222);
			34647: out = 16'(306);
			34648: out = 16'(-192);
			34649: out = 16'(-998);
			34650: out = 16'(-1147);
			34651: out = 16'(152);
			34652: out = 16'(1194);
			34653: out = 16'(585);
			34654: out = 16'(-988);
			34655: out = 16'(-1905);
			34656: out = 16'(-2069);
			34657: out = 16'(-1973);
			34658: out = 16'(-1401);
			34659: out = 16'(472);
			34660: out = 16'(2261);
			34661: out = 16'(2357);
			34662: out = 16'(631);
			34663: out = 16'(-219);
			34664: out = 16'(-151);
			34665: out = 16'(-1330);
			34666: out = 16'(-2461);
			34667: out = 16'(-2273);
			34668: out = 16'(-326);
			34669: out = 16'(1017);
			34670: out = 16'(1293);
			34671: out = 16'(350);
			34672: out = 16'(376);
			34673: out = 16'(1476);
			34674: out = 16'(1050);
			34675: out = 16'(-53);
			34676: out = 16'(-1747);
			34677: out = 16'(-2990);
			34678: out = 16'(-4062);
			34679: out = 16'(-1858);
			34680: out = 16'(699);
			34681: out = 16'(2073);
			34682: out = 16'(2415);
			34683: out = 16'(2495);
			34684: out = 16'(1355);
			34685: out = 16'(-962);
			34686: out = 16'(-3218);
			34687: out = 16'(-4446);
			34688: out = 16'(-3244);
			34689: out = 16'(-679);
			34690: out = 16'(1390);
			34691: out = 16'(2137);
			34692: out = 16'(2744);
			34693: out = 16'(3030);
			34694: out = 16'(1848);
			34695: out = 16'(-808);
			34696: out = 16'(-2848);
			34697: out = 16'(-2650);
			34698: out = 16'(-1095);
			34699: out = 16'(112);
			34700: out = 16'(964);
			34701: out = 16'(1059);
			34702: out = 16'(-43);
			34703: out = 16'(-855);
			34704: out = 16'(-424);
			34705: out = 16'(2069);
			34706: out = 16'(2373);
			34707: out = 16'(-92);
			34708: out = 16'(-1470);
			34709: out = 16'(250);
			34710: out = 16'(1669);
			34711: out = 16'(898);
			34712: out = 16'(70);
			34713: out = 16'(1678);
			34714: out = 16'(1463);
			34715: out = 16'(-1564);
			34716: out = 16'(-2487);
			34717: out = 16'(-1019);
			34718: out = 16'(1421);
			34719: out = 16'(1721);
			34720: out = 16'(308);
			34721: out = 16'(-370);
			34722: out = 16'(-245);
			34723: out = 16'(164);
			34724: out = 16'(326);
			34725: out = 16'(1042);
			34726: out = 16'(530);
			34727: out = 16'(438);
			34728: out = 16'(957);
			34729: out = 16'(366);
			34730: out = 16'(-1134);
			34731: out = 16'(-1252);
			34732: out = 16'(196);
			34733: out = 16'(-139);
			34734: out = 16'(-275);
			34735: out = 16'(-409);
			34736: out = 16'(279);
			34737: out = 16'(899);
			34738: out = 16'(-1182);
			34739: out = 16'(-2863);
			34740: out = 16'(-1799);
			34741: out = 16'(1201);
			34742: out = 16'(2027);
			34743: out = 16'(989);
			34744: out = 16'(-584);
			34745: out = 16'(-1186);
			34746: out = 16'(-2015);
			34747: out = 16'(-1002);
			34748: out = 16'(-38);
			34749: out = 16'(-26);
			34750: out = 16'(-681);
			34751: out = 16'(-285);
			34752: out = 16'(204);
			34753: out = 16'(-5);
			34754: out = 16'(182);
			34755: out = 16'(-47);
			34756: out = 16'(810);
			34757: out = 16'(1481);
			34758: out = 16'(1018);
			34759: out = 16'(247);
			34760: out = 16'(-792);
			34761: out = 16'(-2301);
			34762: out = 16'(-3493);
			34763: out = 16'(-1874);
			34764: out = 16'(861);
			34765: out = 16'(2819);
			34766: out = 16'(2608);
			34767: out = 16'(-91);
			34768: out = 16'(-1079);
			34769: out = 16'(-891);
			34770: out = 16'(-205);
			34771: out = 16'(23);
			34772: out = 16'(467);
			34773: out = 16'(34);
			34774: out = 16'(-133);
			34775: out = 16'(1203);
			34776: out = 16'(2164);
			34777: out = 16'(1987);
			34778: out = 16'(945);
			34779: out = 16'(352);
			34780: out = 16'(219);
			34781: out = 16'(-763);
			34782: out = 16'(-2395);
			34783: out = 16'(-3102);
			34784: out = 16'(-2184);
			34785: out = 16'(127);
			34786: out = 16'(1875);
			34787: out = 16'(2372);
			34788: out = 16'(2061);
			34789: out = 16'(839);
			34790: out = 16'(-464);
			34791: out = 16'(-1422);
			34792: out = 16'(-1557);
			34793: out = 16'(-410);
			34794: out = 16'(710);
			34795: out = 16'(868);
			34796: out = 16'(-43);
			34797: out = 16'(237);
			34798: out = 16'(252);
			34799: out = 16'(177);
			34800: out = 16'(-29);
			34801: out = 16'(-41);
			34802: out = 16'(184);
			34803: out = 16'(266);
			34804: out = 16'(-109);
			34805: out = 16'(328);
			34806: out = 16'(-1435);
			34807: out = 16'(-1821);
			34808: out = 16'(-418);
			34809: out = 16'(-161);
			34810: out = 16'(1006);
			34811: out = 16'(545);
			34812: out = 16'(-148);
			34813: out = 16'(-477);
			34814: out = 16'(-103);
			34815: out = 16'(-532);
			34816: out = 16'(-667);
			34817: out = 16'(166);
			34818: out = 16'(940);
			34819: out = 16'(1109);
			34820: out = 16'(1112);
			34821: out = 16'(1277);
			34822: out = 16'(321);
			34823: out = 16'(-245);
			34824: out = 16'(-909);
			34825: out = 16'(-1285);
			34826: out = 16'(-858);
			34827: out = 16'(-893);
			34828: out = 16'(-413);
			34829: out = 16'(75);
			34830: out = 16'(-1);
			34831: out = 16'(242);
			34832: out = 16'(203);
			34833: out = 16'(-288);
			34834: out = 16'(-720);
			34835: out = 16'(790);
			34836: out = 16'(1819);
			34837: out = 16'(1517);
			34838: out = 16'(2);
			34839: out = 16'(-1488);
			34840: out = 16'(-561);
			34841: out = 16'(879);
			34842: out = 16'(705);
			34843: out = 16'(-335);
			34844: out = 16'(-1253);
			34845: out = 16'(-964);
			34846: out = 16'(-1246);
			34847: out = 16'(-2717);
			34848: out = 16'(-2320);
			34849: out = 16'(280);
			34850: out = 16'(2794);
			34851: out = 16'(2650);
			34852: out = 16'(189);
			34853: out = 16'(-1251);
			34854: out = 16'(-688);
			34855: out = 16'(-94);
			34856: out = 16'(-948);
			34857: out = 16'(-2173);
			34858: out = 16'(-1513);
			34859: out = 16'(638);
			34860: out = 16'(1974);
			34861: out = 16'(1790);
			34862: out = 16'(747);
			34863: out = 16'(-371);
			34864: out = 16'(-1990);
			34865: out = 16'(-1975);
			34866: out = 16'(-1408);
			34867: out = 16'(-237);
			34868: out = 16'(542);
			34869: out = 16'(2787);
			34870: out = 16'(2078);
			34871: out = 16'(211);
			34872: out = 16'(-1314);
			34873: out = 16'(-1894);
			34874: out = 16'(-1786);
			34875: out = 16'(-852);
			34876: out = 16'(285);
			34877: out = 16'(451);
			34878: out = 16'(239);
			34879: out = 16'(201);
			34880: out = 16'(580);
			34881: out = 16'(1051);
			34882: out = 16'(1048);
			34883: out = 16'(1030);
			34884: out = 16'(830);
			34885: out = 16'(277);
			34886: out = 16'(-893);
			34887: out = 16'(-826);
			34888: out = 16'(-61);
			34889: out = 16'(466);
			34890: out = 16'(1753);
			34891: out = 16'(1948);
			34892: out = 16'(1214);
			34893: out = 16'(-445);
			34894: out = 16'(-1329);
			34895: out = 16'(-1753);
			34896: out = 16'(-519);
			34897: out = 16'(888);
			34898: out = 16'(1244);
			34899: out = 16'(1002);
			34900: out = 16'(952);
			34901: out = 16'(553);
			34902: out = 16'(-857);
			34903: out = 16'(-1437);
			34904: out = 16'(-985);
			34905: out = 16'(-255);
			34906: out = 16'(-467);
			34907: out = 16'(53);
			34908: out = 16'(-40);
			34909: out = 16'(-341);
			34910: out = 16'(-1217);
			34911: out = 16'(-583);
			34912: out = 16'(-377);
			34913: out = 16'(1014);
			34914: out = 16'(1745);
			34915: out = 16'(1043);
			34916: out = 16'(-2073);
			34917: out = 16'(-2976);
			34918: out = 16'(-1467);
			34919: out = 16'(400);
			34920: out = 16'(384);
			34921: out = 16'(942);
			34922: out = 16'(1121);
			34923: out = 16'(-193);
			34924: out = 16'(-1841);
			34925: out = 16'(-1755);
			34926: out = 16'(-132);
			34927: out = 16'(1026);
			34928: out = 16'(156);
			34929: out = 16'(-198);
			34930: out = 16'(-527);
			34931: out = 16'(-467);
			34932: out = 16'(1006);
			34933: out = 16'(1125);
			34934: out = 16'(536);
			34935: out = 16'(188);
			34936: out = 16'(1318);
			34937: out = 16'(536);
			34938: out = 16'(-825);
			34939: out = 16'(-2154);
			34940: out = 16'(-2049);
			34941: out = 16'(-2553);
			34942: out = 16'(-1028);
			34943: out = 16'(1301);
			34944: out = 16'(3103);
			34945: out = 16'(2007);
			34946: out = 16'(1343);
			34947: out = 16'(644);
			34948: out = 16'(229);
			34949: out = 16'(-83);
			34950: out = 16'(229);
			34951: out = 16'(325);
			34952: out = 16'(144);
			34953: out = 16'(-444);
			34954: out = 16'(902);
			34955: out = 16'(1354);
			34956: out = 16'(973);
			34957: out = 16'(187);
			34958: out = 16'(9);
			34959: out = 16'(-380);
			34960: out = 16'(-385);
			34961: out = 16'(-4);
			34962: out = 16'(1133);
			34963: out = 16'(395);
			34964: out = 16'(-162);
			34965: out = 16'(212);
			34966: out = 16'(-116);
			34967: out = 16'(111);
			34968: out = 16'(189);
			34969: out = 16'(-456);
			34970: out = 16'(-1401);
			34971: out = 16'(-1543);
			34972: out = 16'(422);
			34973: out = 16'(1638);
			34974: out = 16'(-224);
			34975: out = 16'(-2231);
			34976: out = 16'(-1198);
			34977: out = 16'(1552);
			34978: out = 16'(1813);
			34979: out = 16'(2076);
			34980: out = 16'(420);
			34981: out = 16'(-282);
			34982: out = 16'(-735);
			34983: out = 16'(-1406);
			34984: out = 16'(-1828);
			34985: out = 16'(-478);
			34986: out = 16'(1053);
			34987: out = 16'(883);
			34988: out = 16'(-440);
			34989: out = 16'(-625);
			34990: out = 16'(-34);
			34991: out = 16'(-968);
			34992: out = 16'(-2177);
			34993: out = 16'(-2209);
			34994: out = 16'(67);
			34995: out = 16'(2132);
			34996: out = 16'(3026);
			34997: out = 16'(1161);
			34998: out = 16'(-895);
			34999: out = 16'(-2054);
			35000: out = 16'(-2502);
			35001: out = 16'(-2066);
			35002: out = 16'(-243);
			35003: out = 16'(1405);
			35004: out = 16'(1013);
			35005: out = 16'(197);
			35006: out = 16'(364);
			35007: out = 16'(893);
			35008: out = 16'(-76);
			35009: out = 16'(-38);
			35010: out = 16'(-3);
			35011: out = 16'(-239);
			35012: out = 16'(-757);
			35013: out = 16'(-595);
			35014: out = 16'(483);
			35015: out = 16'(741);
			35016: out = 16'(-16);
			35017: out = 16'(776);
			35018: out = 16'(1664);
			35019: out = 16'(917);
			35020: out = 16'(-1024);
			35021: out = 16'(-33);
			35022: out = 16'(-59);
			35023: out = 16'(-524);
			35024: out = 16'(-1142);
			35025: out = 16'(51);
			35026: out = 16'(1328);
			35027: out = 16'(1621);
			35028: out = 16'(372);
			35029: out = 16'(59);
			35030: out = 16'(-679);
			35031: out = 16'(394);
			35032: out = 16'(559);
			35033: out = 16'(-630);
			35034: out = 16'(-871);
			35035: out = 16'(-333);
			35036: out = 16'(-279);
			35037: out = 16'(-832);
			35038: out = 16'(153);
			35039: out = 16'(49);
			35040: out = 16'(-156);
			35041: out = 16'(180);
			35042: out = 16'(1067);
			35043: out = 16'(1334);
			35044: out = 16'(-5);
			35045: out = 16'(-1418);
			35046: out = 16'(-747);
			35047: out = 16'(-645);
			35048: out = 16'(-58);
			35049: out = 16'(494);
			35050: out = 16'(789);
			35051: out = 16'(-235);
			35052: out = 16'(-1544);
			35053: out = 16'(-1424);
			35054: out = 16'(185);
			35055: out = 16'(-137);
			35056: out = 16'(26);
			35057: out = 16'(-87);
			35058: out = 16'(-69);
			35059: out = 16'(-829);
			35060: out = 16'(-249);
			35061: out = 16'(-26);
			35062: out = 16'(38);
			35063: out = 16'(293);
			35064: out = 16'(-283);
			35065: out = 16'(-195);
			35066: out = 16'(358);
			35067: out = 16'(-160);
			35068: out = 16'(976);
			35069: out = 16'(229);
			35070: out = 16'(208);
			35071: out = 16'(1004);
			35072: out = 16'(2060);
			35073: out = 16'(-75);
			35074: out = 16'(-1869);
			35075: out = 16'(-1625);
			35076: out = 16'(192);
			35077: out = 16'(263);
			35078: out = 16'(665);
			35079: out = 16'(1222);
			35080: out = 16'(845);
			35081: out = 16'(-248);
			35082: out = 16'(-588);
			35083: out = 16'(-737);
			35084: out = 16'(-1575);
			35085: out = 16'(-1588);
			35086: out = 16'(-588);
			35087: out = 16'(99);
			35088: out = 16'(129);
			35089: out = 16'(1631);
			35090: out = 16'(2710);
			35091: out = 16'(2009);
			35092: out = 16'(-269);
			35093: out = 16'(-1441);
			35094: out = 16'(-1911);
			35095: out = 16'(-2125);
			35096: out = 16'(-1916);
			35097: out = 16'(288);
			35098: out = 16'(1531);
			35099: out = 16'(1574);
			35100: out = 16'(507);
			35101: out = 16'(-54);
			35102: out = 16'(-1076);
			35103: out = 16'(-873);
			35104: out = 16'(-138);
			35105: out = 16'(292);
			35106: out = 16'(891);
			35107: out = 16'(862);
			35108: out = 16'(973);
			35109: out = 16'(541);
			35110: out = 16'(-982);
			35111: out = 16'(-2493);
			35112: out = 16'(-1657);
			35113: out = 16'(295);
			35114: out = 16'(186);
			35115: out = 16'(345);
			35116: out = 16'(563);
			35117: out = 16'(882);
			35118: out = 16'(182);
			35119: out = 16'(28);
			35120: out = 16'(11);
			35121: out = 16'(219);
			35122: out = 16'(-178);
			35123: out = 16'(-674);
			35124: out = 16'(-936);
			35125: out = 16'(-479);
			35126: out = 16'(0);
			35127: out = 16'(-17);
			35128: out = 16'(589);
			35129: out = 16'(1095);
			35130: out = 16'(660);
			35131: out = 16'(60);
			35132: out = 16'(-1296);
			35133: out = 16'(-803);
			35134: out = 16'(673);
			35135: out = 16'(776);
			35136: out = 16'(195);
			35137: out = 16'(-697);
			35138: out = 16'(-592);
			35139: out = 16'(-43);
			35140: out = 16'(283);
			35141: out = 16'(51);
			35142: out = 16'(-63);
			35143: out = 16'(-89);
			35144: out = 16'(1);
			35145: out = 16'(-126);
			35146: out = 16'(137);
			35147: out = 16'(-92);
			35148: out = 16'(-1389);
			35149: out = 16'(-2499);
			35150: out = 16'(-1396);
			35151: out = 16'(1129);
			35152: out = 16'(2557);
			35153: out = 16'(2361);
			35154: out = 16'(1107);
			35155: out = 16'(-266);
			35156: out = 16'(-1231);
			35157: out = 16'(-2532);
			35158: out = 16'(-2063);
			35159: out = 16'(-1041);
			35160: out = 16'(-272);
			35161: out = 16'(-82);
			35162: out = 16'(2497);
			35163: out = 16'(3871);
			35164: out = 16'(2053);
			35165: out = 16'(-827);
			35166: out = 16'(-2070);
			35167: out = 16'(-1183);
			35168: out = 16'(-511);
			35169: out = 16'(-715);
			35170: out = 16'(-912);
			35171: out = 16'(326);
			35172: out = 16'(1384);
			35173: out = 16'(829);
			35174: out = 16'(121);
			35175: out = 16'(416);
			35176: out = 16'(932);
			35177: out = 16'(-49);
			35178: out = 16'(-1195);
			35179: out = 16'(-2022);
			35180: out = 16'(-1259);
			35181: out = 16'(-300);
			35182: out = 16'(402);
			35183: out = 16'(-26);
			35184: out = 16'(837);
			35185: out = 16'(1775);
			35186: out = 16'(251);
			35187: out = 16'(-290);
			35188: out = 16'(-314);
			35189: out = 16'(38);
			35190: out = 16'(-80);
			35191: out = 16'(-659);
			35192: out = 16'(-445);
			35193: out = 16'(133);
			35194: out = 16'(-126);
			35195: out = 16'(38);
			35196: out = 16'(-185);
			35197: out = 16'(667);
			35198: out = 16'(1852);
			35199: out = 16'(915);
			35200: out = 16'(467);
			35201: out = 16'(-101);
			35202: out = 16'(-489);
			35203: out = 16'(-55);
			35204: out = 16'(-111);
			35205: out = 16'(76);
			35206: out = 16'(272);
			35207: out = 16'(217);
			35208: out = 16'(-330);
			35209: out = 16'(-600);
			35210: out = 16'(-282);
			35211: out = 16'(154);
			35212: out = 16'(21);
			35213: out = 16'(-142);
			35214: out = 16'(259);
			35215: out = 16'(861);
			35216: out = 16'(308);
			35217: out = 16'(-292);
			35218: out = 16'(-461);
			35219: out = 16'(-140);
			35220: out = 16'(-550);
			35221: out = 16'(-143);
			35222: out = 16'(-57);
			35223: out = 16'(-84);
			35224: out = 16'(-87);
			35225: out = 16'(-53);
			35226: out = 16'(-97);
			35227: out = 16'(162);
			35228: out = 16'(825);
			35229: out = 16'(-838);
			35230: out = 16'(-1576);
			35231: out = 16'(-1016);
			35232: out = 16'(390);
			35233: out = 16'(1093);
			35234: out = 16'(1280);
			35235: out = 16'(836);
			35236: out = 16'(-180);
			35237: out = 16'(-1815);
			35238: out = 16'(-2030);
			35239: out = 16'(-1421);
			35240: out = 16'(-512);
			35241: out = 16'(292);
			35242: out = 16'(315);
			35243: out = 16'(-91);
			35244: out = 16'(-431);
			35245: out = 16'(148);
			35246: out = 16'(877);
			35247: out = 16'(1952);
			35248: out = 16'(1565);
			35249: out = 16'(-66);
			35250: out = 16'(-2777);
			35251: out = 16'(-1881);
			35252: out = 16'(-82);
			35253: out = 16'(111);
			35254: out = 16'(-954);
			35255: out = 16'(-543);
			35256: out = 16'(901);
			35257: out = 16'(1956);
			35258: out = 16'(1724);
			35259: out = 16'(-262);
			35260: out = 16'(-2645);
			35261: out = 16'(-2676);
			35262: out = 16'(1103);
			35263: out = 16'(1230);
			35264: out = 16'(754);
			35265: out = 16'(78);
			35266: out = 16'(377);
			35267: out = 16'(138);
			35268: out = 16'(101);
			35269: out = 16'(-67);
			35270: out = 16'(380);
			35271: out = 16'(154);
			35272: out = 16'(192);
			35273: out = 16'(-653);
			35274: out = 16'(-1088);
			35275: out = 16'(-943);
			35276: out = 16'(-15);
			35277: out = 16'(-738);
			35278: out = 16'(-1369);
			35279: out = 16'(-373);
			35280: out = 16'(1568);
			35281: out = 16'(861);
			35282: out = 16'(-1022);
			35283: out = 16'(-1252);
			35284: out = 16'(834);
			35285: out = 16'(1499);
			35286: out = 16'(752);
			35287: out = 16'(-115);
			35288: out = 16'(4);
			35289: out = 16'(-169);
			35290: out = 16'(672);
			35291: out = 16'(1821);
			35292: out = 16'(864);
			35293: out = 16'(117);
			35294: out = 16'(-141);
			35295: out = 16'(-434);
			35296: out = 16'(-1912);
			35297: out = 16'(-970);
			35298: out = 16'(1272);
			35299: out = 16'(2497);
			35300: out = 16'(466);
			35301: out = 16'(-2007);
			35302: out = 16'(-3129);
			35303: out = 16'(-1588);
			35304: out = 16'(381);
			35305: out = 16'(368);
			35306: out = 16'(212);
			35307: out = 16'(511);
			35308: out = 16'(1098);
			35309: out = 16'(2039);
			35310: out = 16'(820);
			35311: out = 16'(-805);
			35312: out = 16'(-1505);
			35313: out = 16'(-453);
			35314: out = 16'(-777);
			35315: out = 16'(-846);
			35316: out = 16'(-664);
			35317: out = 16'(75);
			35318: out = 16'(-155);
			35319: out = 16'(1113);
			35320: out = 16'(1527);
			35321: out = 16'(-446);
			35322: out = 16'(-1179);
			35323: out = 16'(-2669);
			35324: out = 16'(-2692);
			35325: out = 16'(-1388);
			35326: out = 16'(925);
			35327: out = 16'(1698);
			35328: out = 16'(2010);
			35329: out = 16'(1547);
			35330: out = 16'(275);
			35331: out = 16'(-1464);
			35332: out = 16'(-1889);
			35333: out = 16'(-1157);
			35334: out = 16'(-397);
			35335: out = 16'(-656);
			35336: out = 16'(-330);
			35337: out = 16'(417);
			35338: out = 16'(920);
			35339: out = 16'(-833);
			35340: out = 16'(-988);
			35341: out = 16'(-334);
			35342: out = 16'(91);
			35343: out = 16'(69);
			35344: out = 16'(28);
			35345: out = 16'(-158);
			35346: out = 16'(-310);
			35347: out = 16'(83);
			35348: out = 16'(283);
			35349: out = 16'(235);
			35350: out = 16'(66);
			35351: out = 16'(431);
			35352: out = 16'(94);
			35353: out = 16'(212);
			35354: out = 16'(365);
			35355: out = 16'(-8);
			35356: out = 16'(59);
			35357: out = 16'(-329);
			35358: out = 16'(90);
			35359: out = 16'(1082);
			35360: out = 16'(362);
			35361: out = 16'(328);
			35362: out = 16'(239);
			35363: out = 16'(261);
			35364: out = 16'(23);
			35365: out = 16'(215);
			35366: out = 16'(14);
			35367: out = 16'(-718);
			35368: out = 16'(-1373);
			35369: out = 16'(-973);
			35370: out = 16'(-25);
			35371: out = 16'(441);
			35372: out = 16'(372);
			35373: out = 16'(-335);
			35374: out = 16'(431);
			35375: out = 16'(1171);
			35376: out = 16'(774);
			35377: out = 16'(-568);
			35378: out = 16'(-413);
			35379: out = 16'(629);
			35380: out = 16'(1142);
			35381: out = 16'(52);
			35382: out = 16'(576);
			35383: out = 16'(1472);
			35384: out = 16'(1562);
			35385: out = 16'(190);
			35386: out = 16'(-1117);
			35387: out = 16'(-1800);
			35388: out = 16'(-770);
			35389: out = 16'(1245);
			35390: out = 16'(1033);
			35391: out = 16'(432);
			35392: out = 16'(362);
			35393: out = 16'(928);
			35394: out = 16'(1165);
			35395: out = 16'(-473);
			35396: out = 16'(-2329);
			35397: out = 16'(-2283);
			35398: out = 16'(-292);
			35399: out = 16'(1047);
			35400: out = 16'(730);
			35401: out = 16'(-75);
			35402: out = 16'(983);
			35403: out = 16'(767);
			35404: out = 16'(1136);
			35405: out = 16'(708);
			35406: out = 16'(-942);
			35407: out = 16'(-1863);
			35408: out = 16'(-1216);
			35409: out = 16'(-364);
			35410: out = 16'(-887);
			35411: out = 16'(291);
			35412: out = 16'(61);
			35413: out = 16'(53);
			35414: out = 16'(386);
			35415: out = 16'(1160);
			35416: out = 16'(401);
			35417: out = 16'(-1104);
			35418: out = 16'(-2422);
			35419: out = 16'(-1737);
			35420: out = 16'(-629);
			35421: out = 16'(1285);
			35422: out = 16'(1978);
			35423: out = 16'(900);
			35424: out = 16'(-523);
			35425: out = 16'(-497);
			35426: out = 16'(99);
			35427: out = 16'(-185);
			35428: out = 16'(-1914);
			35429: out = 16'(-1988);
			35430: out = 16'(-805);
			35431: out = 16'(100);
			35432: out = 16'(322);
			35433: out = 16'(89);
			35434: out = 16'(-189);
			35435: out = 16'(-329);
			35436: out = 16'(38);
			35437: out = 16'(743);
			35438: out = 16'(1111);
			35439: out = 16'(753);
			35440: out = 16'(-8);
			35441: out = 16'(176);
			35442: out = 16'(302);
			35443: out = 16'(224);
			35444: out = 16'(-143);
			35445: out = 16'(-1199);
			35446: out = 16'(-1951);
			35447: out = 16'(-960);
			35448: out = 16'(1177);
			35449: out = 16'(956);
			35450: out = 16'(411);
			35451: out = 16'(-142);
			35452: out = 16'(184);
			35453: out = 16'(851);
			35454: out = 16'(116);
			35455: out = 16'(-837);
			35456: out = 16'(-361);
			35457: out = 16'(853);
			35458: out = 16'(1346);
			35459: out = 16'(670);
			35460: out = 16'(407);
			35461: out = 16'(811);
			35462: out = 16'(210);
			35463: out = 16'(-1061);
			35464: out = 16'(-1241);
			35465: out = 16'(-72);
			35466: out = 16'(18);
			35467: out = 16'(-814);
			35468: out = 16'(-757);
			35469: out = 16'(594);
			35470: out = 16'(1718);
			35471: out = 16'(576);
			35472: out = 16'(-316);
			35473: out = 16'(57);
			35474: out = 16'(-154);
			35475: out = 16'(-29);
			35476: out = 16'(-94);
			35477: out = 16'(-50);
			35478: out = 16'(-58);
			35479: out = 16'(-108);
			35480: out = 16'(140);
			35481: out = 16'(-2);
			35482: out = 16'(-483);
			35483: out = 16'(-895);
			35484: out = 16'(826);
			35485: out = 16'(1894);
			35486: out = 16'(847);
			35487: out = 16'(17);
			35488: out = 16'(-545);
			35489: out = 16'(-446);
			35490: out = 16'(-686);
			35491: out = 16'(-1142);
			35492: out = 16'(-1519);
			35493: out = 16'(-1106);
			35494: out = 16'(-4);
			35495: out = 16'(887);
			35496: out = 16'(1033);
			35497: out = 16'(323);
			35498: out = 16'(113);
			35499: out = 16'(887);
			35500: out = 16'(105);
			35501: out = 16'(-1222);
			35502: out = 16'(-2011);
			35503: out = 16'(-1357);
			35504: out = 16'(-1584);
			35505: out = 16'(150);
			35506: out = 16'(1671);
			35507: out = 16'(1986);
			35508: out = 16'(990);
			35509: out = 16'(-122);
			35510: out = 16'(-772);
			35511: out = 16'(-688);
			35512: out = 16'(-25);
			35513: out = 16'(-368);
			35514: out = 16'(-494);
			35515: out = 16'(-324);
			35516: out = 16'(438);
			35517: out = 16'(714);
			35518: out = 16'(1609);
			35519: out = 16'(1240);
			35520: out = 16'(-235);
			35521: out = 16'(-504);
			35522: out = 16'(21);
			35523: out = 16'(-299);
			35524: out = 16'(-1832);
			35525: out = 16'(-1791);
			35526: out = 16'(-744);
			35527: out = 16'(1049);
			35528: out = 16'(1635);
			35529: out = 16'(239);
			35530: out = 16'(-284);
			35531: out = 16'(-765);
			35532: out = 16'(-552);
			35533: out = 16'(355);
			35534: out = 16'(1081);
			35535: out = 16'(1098);
			35536: out = 16'(752);
			35537: out = 16'(479);
			35538: out = 16'(-392);
			35539: out = 16'(-397);
			35540: out = 16'(479);
			35541: out = 16'(997);
			35542: out = 16'(-373);
			35543: out = 16'(-1690);
			35544: out = 16'(-1150);
			35545: out = 16'(640);
			35546: out = 16'(746);
			35547: out = 16'(225);
			35548: out = 16'(-402);
			35549: out = 16'(257);
			35550: out = 16'(908);
			35551: out = 16'(267);
			35552: out = 16'(-1239);
			35553: out = 16'(-1408);
			35554: out = 16'(96);
			35555: out = 16'(918);
			35556: out = 16'(440);
			35557: out = 16'(-496);
			35558: out = 16'(-761);
			35559: out = 16'(-819);
			35560: out = 16'(-546);
			35561: out = 16'(-283);
			35562: out = 16'(3);
			35563: out = 16'(-100);
			35564: out = 16'(2);
			35565: out = 16'(-369);
			35566: out = 16'(-1045);
			35567: out = 16'(-2007);
			35568: out = 16'(-465);
			35569: out = 16'(582);
			35570: out = 16'(917);
			35571: out = 16'(833);
			35572: out = 16'(348);
			35573: out = 16'(203);
			35574: out = 16'(32);
			35575: out = 16'(-564);
			35576: out = 16'(-1244);
			35577: out = 16'(-1052);
			35578: out = 16'(58);
			35579: out = 16'(1056);
			35580: out = 16'(1676);
			35581: out = 16'(628);
			35582: out = 16'(396);
			35583: out = 16'(819);
			35584: out = 16'(-185);
			35585: out = 16'(2);
			35586: out = 16'(-547);
			35587: out = 16'(-592);
			35588: out = 16'(-13);
			35589: out = 16'(-25);
			35590: out = 16'(56);
			35591: out = 16'(558);
			35592: out = 16'(1004);
			35593: out = 16'(-15);
			35594: out = 16'(-853);
			35595: out = 16'(-828);
			35596: out = 16'(6);
			35597: out = 16'(-129);
			35598: out = 16'(-216);
			35599: out = 16'(-699);
			35600: out = 16'(-384);
			35601: out = 16'(1098);
			35602: out = 16'(1778);
			35603: out = 16'(1400);
			35604: out = 16'(402);
			35605: out = 16'(-97);
			35606: out = 16'(-488);
			35607: out = 16'(-317);
			35608: out = 16'(-165);
			35609: out = 16'(-29);
			35610: out = 16'(644);
			35611: out = 16'(854);
			35612: out = 16'(165);
			35613: out = 16'(-989);
			35614: out = 16'(-1072);
			35615: out = 16'(-971);
			35616: out = 16'(-452);
			35617: out = 16'(204);
			35618: out = 16'(1605);
			35619: out = 16'(531);
			35620: out = 16'(-52);
			35621: out = 16'(-256);
			35622: out = 16'(-469);
			35623: out = 16'(95);
			35624: out = 16'(267);
			35625: out = 16'(-6);
			35626: out = 16'(-503);
			35627: out = 16'(-798);
			35628: out = 16'(-190);
			35629: out = 16'(182);
			35630: out = 16'(-118);
			35631: out = 16'(189);
			35632: out = 16'(497);
			35633: out = 16'(1228);
			35634: out = 16'(1325);
			35635: out = 16'(-125);
			35636: out = 16'(-927);
			35637: out = 16'(-997);
			35638: out = 16'(-50);
			35639: out = 16'(950);
			35640: out = 16'(370);
			35641: out = 16'(-575);
			35642: out = 16'(-443);
			35643: out = 16'(775);
			35644: out = 16'(-27);
			35645: out = 16'(-448);
			35646: out = 16'(-130);
			35647: out = 16'(712);
			35648: out = 16'(-763);
			35649: out = 16'(-1080);
			35650: out = 16'(-804);
			35651: out = 16'(157);
			35652: out = 16'(634);
			35653: out = 16'(272);
			35654: out = 16'(-745);
			35655: out = 16'(-861);
			35656: out = 16'(39);
			35657: out = 16'(141);
			35658: out = 16'(-1077);
			35659: out = 16'(-1450);
			35660: out = 16'(0);
			35661: out = 16'(25);
			35662: out = 16'(-1223);
			35663: out = 16'(-1858);
			35664: out = 16'(14);
			35665: out = 16'(838);
			35666: out = 16'(1220);
			35667: out = 16'(196);
			35668: out = 16'(-301);
			35669: out = 16'(-155);
			35670: out = 16'(913);
			35671: out = 16'(653);
			35672: out = 16'(-491);
			35673: out = 16'(-2351);
			35674: out = 16'(122);
			35675: out = 16'(1235);
			35676: out = 16'(793);
			35677: out = 16'(-116);
			35678: out = 16'(21);
			35679: out = 16'(-1028);
			35680: out = 16'(-1558);
			35681: out = 16'(-146);
			35682: out = 16'(637);
			35683: out = 16'(618);
			35684: out = 16'(4);
			35685: out = 16'(64);
			35686: out = 16'(82);
			35687: out = 16'(277);
			35688: out = 16'(-146);
			35689: out = 16'(-432);
			35690: out = 16'(-436);
			35691: out = 16'(541);
			35692: out = 16'(945);
			35693: out = 16'(404);
			35694: out = 16'(-1072);
			35695: out = 16'(-860);
			35696: out = 16'(190);
			35697: out = 16'(1565);
			35698: out = 16'(1606);
			35699: out = 16'(333);
			35700: out = 16'(-1375);
			35701: out = 16'(-1274);
			35702: out = 16'(98);
			35703: out = 16'(1049);
			35704: out = 16'(208);
			35705: out = 16'(428);
			35706: out = 16'(1657);
			35707: out = 16'(644);
			35708: out = 16'(-341);
			35709: out = 16'(-1334);
			35710: out = 16'(-1407);
			35711: out = 16'(-1098);
			35712: out = 16'(-350);
			35713: out = 16'(984);
			35714: out = 16'(1991);
			35715: out = 16'(1353);
			35716: out = 16'(934);
			35717: out = 16'(-288);
			35718: out = 16'(-1212);
			35719: out = 16'(-1402);
			35720: out = 16'(-258);
			35721: out = 16'(-68);
			35722: out = 16'(-299);
			35723: out = 16'(-452);
			35724: out = 16'(-149);
			35725: out = 16'(127);
			35726: out = 16'(60);
			35727: out = 16'(-92);
			35728: out = 16'(185);
			35729: out = 16'(633);
			35730: out = 16'(372);
			35731: out = 16'(-496);
			35732: out = 16'(-1129);
			35733: out = 16'(-1483);
			35734: out = 16'(-762);
			35735: out = 16'(774);
			35736: out = 16'(2259);
			35737: out = 16'(67);
			35738: out = 16'(-648);
			35739: out = 16'(-874);
			35740: out = 16'(-961);
			35741: out = 16'(-2391);
			35742: out = 16'(-1529);
			35743: out = 16'(-360);
			35744: out = 16'(464);
			35745: out = 16'(800);
			35746: out = 16'(923);
			35747: out = 16'(370);
			35748: out = 16'(-75);
			35749: out = 16'(128);
			35750: out = 16'(-1114);
			35751: out = 16'(-1756);
			35752: out = 16'(-1116);
			35753: out = 16'(435);
			35754: out = 16'(827);
			35755: out = 16'(-218);
			35756: out = 16'(-1415);
			35757: out = 16'(-1041);
			35758: out = 16'(-166);
			35759: out = 16'(802);
			35760: out = 16'(534);
			35761: out = 16'(-40);
			35762: out = 16'(-21);
			35763: out = 16'(52);
			35764: out = 16'(-197);
			35765: out = 16'(-362);
			35766: out = 16'(-381);
			35767: out = 16'(996);
			35768: out = 16'(753);
			35769: out = 16'(104);
			35770: out = 16'(-31);
			35771: out = 16'(8);
			35772: out = 16'(-659);
			35773: out = 16'(-948);
			35774: out = 16'(-214);
			35775: out = 16'(-75);
			35776: out = 16'(623);
			35777: out = 16'(983);
			35778: out = 16'(608);
			35779: out = 16'(-305);
			35780: out = 16'(-1041);
			35781: out = 16'(-120);
			35782: out = 16'(903);
			35783: out = 16'(-171);
			35784: out = 16'(-486);
			35785: out = 16'(-844);
			35786: out = 16'(-438);
			35787: out = 16'(77);
			35788: out = 16'(1017);
			35789: out = 16'(1074);
			35790: out = 16'(517);
			35791: out = 16'(-77);
			35792: out = 16'(-39);
			35793: out = 16'(-453);
			35794: out = 16'(-1098);
			35795: out = 16'(-1068);
			35796: out = 16'(811);
			35797: out = 16'(1154);
			35798: out = 16'(605);
			35799: out = 16'(-176);
			35800: out = 16'(28);
			35801: out = 16'(-90);
			35802: out = 16'(-15);
			35803: out = 16'(-10);
			35804: out = 16'(308);
			35805: out = 16'(691);
			35806: out = 16'(970);
			35807: out = 16'(282);
			35808: out = 16'(-731);
			35809: out = 16'(165);
			35810: out = 16'(1166);
			35811: out = 16'(1612);
			35812: out = 16'(572);
			35813: out = 16'(-1253);
			35814: out = 16'(-2090);
			35815: out = 16'(-1505);
			35816: out = 16'(-492);
			35817: out = 16'(-18);
			35818: out = 16'(640);
			35819: out = 16'(978);
			35820: out = 16'(275);
			35821: out = 16'(-1417);
			35822: out = 16'(-869);
			35823: out = 16'(-265);
			35824: out = 16'(101);
			35825: out = 16'(351);
			35826: out = 16'(743);
			35827: out = 16'(946);
			35828: out = 16'(257);
			35829: out = 16'(-996);
			35830: out = 16'(-1960);
			35831: out = 16'(-1637);
			35832: out = 16'(-647);
			35833: out = 16'(561);
			35834: out = 16'(753);
			35835: out = 16'(428);
			35836: out = 16'(-1174);
			35837: out = 16'(-1785);
			35838: out = 16'(-580);
			35839: out = 16'(1029);
			35840: out = 16'(560);
			35841: out = 16'(232);
			35842: out = 16'(1251);
			35843: out = 16'(1206);
			35844: out = 16'(-793);
			35845: out = 16'(-2208);
			35846: out = 16'(-813);
			35847: out = 16'(625);
			35848: out = 16'(753);
			35849: out = 16'(-166);
			35850: out = 16'(-164);
			35851: out = 16'(-105);
			35852: out = 16'(180);
			35853: out = 16'(-405);
			35854: out = 16'(-361);
			35855: out = 16'(590);
			35856: out = 16'(1197);
			35857: out = 16'(514);
			35858: out = 16'(-20);
			35859: out = 16'(284);
			35860: out = 16'(845);
			35861: out = 16'(140);
			35862: out = 16'(-645);
			35863: out = 16'(-605);
			35864: out = 16'(261);
			35865: out = 16'(-533);
			35866: out = 16'(-1070);
			35867: out = 16'(-459);
			35868: out = 16'(-27);
			35869: out = 16'(257);
			35870: out = 16'(679);
			35871: out = 16'(1227);
			35872: out = 16'(742);
			35873: out = 16'(233);
			35874: out = 16'(-643);
			35875: out = 16'(-1157);
			35876: out = 16'(-1322);
			35877: out = 16'(-489);
			35878: out = 16'(-94);
			35879: out = 16'(61);
			35880: out = 16'(104);
			35881: out = 16'(1107);
			35882: out = 16'(467);
			35883: out = 16'(-476);
			35884: out = 16'(-956);
			35885: out = 16'(-358);
			35886: out = 16'(-352);
			35887: out = 16'(-188);
			35888: out = 16'(323);
			35889: out = 16'(1703);
			35890: out = 16'(356);
			35891: out = 16'(-167);
			35892: out = 16'(215);
			35893: out = 16'(836);
			35894: out = 16'(63);
			35895: out = 16'(67);
			35896: out = 16'(153);
			35897: out = 16'(-78);
			35898: out = 16'(1004);
			35899: out = 16'(1037);
			35900: out = 16'(113);
			35901: out = 16'(-1163);
			35902: out = 16'(-423);
			35903: out = 16'(-151);
			35904: out = 16'(-24);
			35905: out = 16'(58);
			35906: out = 16'(812);
			35907: out = 16'(172);
			35908: out = 16'(-612);
			35909: out = 16'(-1056);
			35910: out = 16'(-380);
			35911: out = 16'(-1576);
			35912: out = 16'(-780);
			35913: out = 16'(967);
			35914: out = 16'(1745);
			35915: out = 16'(295);
			35916: out = 16'(-665);
			35917: out = 16'(-433);
			35918: out = 16'(-58);
			35919: out = 16'(78);
			35920: out = 16'(-1026);
			35921: out = 16'(-905);
			35922: out = 16'(217);
			35923: out = 16'(216);
			35924: out = 16'(-553);
			35925: out = 16'(-1506);
			35926: out = 16'(-1246);
			35927: out = 16'(347);
			35928: out = 16'(87);
			35929: out = 16'(91);
			35930: out = 16'(-52);
			35931: out = 16'(-262);
			35932: out = 16'(148);
			35933: out = 16'(933);
			35934: out = 16'(1127);
			35935: out = 16'(897);
			35936: out = 16'(1073);
			35937: out = 16'(702);
			35938: out = 16'(-746);
			35939: out = 16'(-2113);
			35940: out = 16'(-1703);
			35941: out = 16'(-169);
			35942: out = 16'(264);
			35943: out = 16'(284);
			35944: out = 16'(1720);
			35945: out = 16'(1114);
			35946: out = 16'(-493);
			35947: out = 16'(-1969);
			35948: out = 16'(-1494);
			35949: out = 16'(-874);
			35950: out = 16'(-173);
			35951: out = 16'(398);
			35952: out = 16'(1327);
			35953: out = 16'(1622);
			35954: out = 16'(1237);
			35955: out = 16'(397);
			35956: out = 16'(-96);
			35957: out = 16'(-422);
			35958: out = 16'(-1075);
			35959: out = 16'(-1365);
			35960: out = 16'(-647);
			35961: out = 16'(243);
			35962: out = 16'(422);
			35963: out = 16'(-73);
			35964: out = 16'(-298);
			35965: out = 16'(65);
			35966: out = 16'(1009);
			35967: out = 16'(628);
			35968: out = 16'(-563);
			35969: out = 16'(-1306);
			35970: out = 16'(-1085);
			35971: out = 16'(-262);
			35972: out = 16'(127);
			35973: out = 16'(3);
			35974: out = 16'(10);
			35975: out = 16'(603);
			35976: out = 16'(1081);
			35977: out = 16'(342);
			35978: out = 16'(-1875);
			35979: out = 16'(-947);
			35980: out = 16'(1064);
			35981: out = 16'(1689);
			35982: out = 16'(-93);
			35983: out = 16'(227);
			35984: out = 16'(123);
			35985: out = 16'(-215);
			35986: out = 16'(-706);
			35987: out = 16'(-434);
			35988: out = 16'(-143);
			35989: out = 16'(-42);
			35990: out = 16'(206);
			35991: out = 16'(1564);
			35992: out = 16'(1272);
			35993: out = 16'(-173);
			35994: out = 16'(-1518);
			35995: out = 16'(-1320);
			35996: out = 16'(-149);
			35997: out = 16'(299);
			35998: out = 16'(-88);
			35999: out = 16'(81);
			36000: out = 16'(-62);
			36001: out = 16'(81);
			36002: out = 16'(-132);
			36003: out = 16'(-310);
			36004: out = 16'(-51);
			36005: out = 16'(-264);
			36006: out = 16'(-1257);
			36007: out = 16'(-1781);
			36008: out = 16'(-114);
			36009: out = 16'(987);
			36010: out = 16'(931);
			36011: out = 16'(233);
			36012: out = 16'(370);
			36013: out = 16'(266);
			36014: out = 16'(179);
			36015: out = 16'(-185);
			36016: out = 16'(-1015);
			36017: out = 16'(-1234);
			36018: out = 16'(-893);
			36019: out = 16'(203);
			36020: out = 16'(814);
			36021: out = 16'(339);
			36022: out = 16'(-947);
			36023: out = 16'(-631);
			36024: out = 16'(1153);
			36025: out = 16'(1673);
			36026: out = 16'(787);
			36027: out = 16'(17);
			36028: out = 16'(9);
			36029: out = 16'(30);
			36030: out = 16'(-1268);
			36031: out = 16'(-1032);
			36032: out = 16'(837);
			36033: out = 16'(1537);
			36034: out = 16'(695);
			36035: out = 16'(-455);
			36036: out = 16'(-454);
			36037: out = 16'(334);
			36038: out = 16'(34);
			36039: out = 16'(-9);
			36040: out = 16'(-16);
			36041: out = 16'(93);
			36042: out = 16'(744);
			36043: out = 16'(639);
			36044: out = 16'(-444);
			36045: out = 16'(-1188);
			36046: out = 16'(176);
			36047: out = 16'(1417);
			36048: out = 16'(1148);
			36049: out = 16'(37);
			36050: out = 16'(-7);
			36051: out = 16'(-544);
			36052: out = 16'(-1483);
			36053: out = 16'(-1814);
			36054: out = 16'(-196);
			36055: out = 16'(647);
			36056: out = 16'(669);
			36057: out = 16'(-125);
			36058: out = 16'(-281);
			36059: out = 16'(-126);
			36060: out = 16'(87);
			36061: out = 16'(-232);
			36062: out = 16'(-180);
			36063: out = 16'(993);
			36064: out = 16'(1093);
			36065: out = 16'(90);
			36066: out = 16'(-893);
			36067: out = 16'(-1392);
			36068: out = 16'(-785);
			36069: out = 16'(-734);
			36070: out = 16'(-275);
			36071: out = 16'(924);
			36072: out = 16'(1647);
			36073: out = 16'(783);
			36074: out = 16'(-348);
			36075: out = 16'(-749);
			36076: out = 16'(-1522);
			36077: out = 16'(-1260);
			36078: out = 16'(367);
			36079: out = 16'(1640);
			36080: out = 16'(1083);
			36081: out = 16'(-1454);
			36082: out = 16'(-1817);
			36083: out = 16'(31);
			36084: out = 16'(-77);
			36085: out = 16'(-147);
			36086: out = 16'(-222);
			36087: out = 16'(157);
			36088: out = 16'(46);
			36089: out = 16'(263);
			36090: out = 16'(741);
			36091: out = 16'(425);
			36092: out = 16'(-1403);
			36093: out = 16'(-1589);
			36094: out = 16'(-637);
			36095: out = 16'(379);
			36096: out = 16'(204);
			36097: out = 16'(168);
			36098: out = 16'(22);
			36099: out = 16'(188);
			36100: out = 16'(306);
			36101: out = 16'(31);
			36102: out = 16'(734);
			36103: out = 16'(505);
			36104: out = 16'(-732);
			36105: out = 16'(-1522);
			36106: out = 16'(-938);
			36107: out = 16'(256);
			36108: out = 16'(1340);
			36109: out = 16'(1928);
			36110: out = 16'(1372);
			36111: out = 16'(54);
			36112: out = 16'(-945);
			36113: out = 16'(-900);
			36114: out = 16'(-440);
			36115: out = 16'(-508);
			36116: out = 16'(-490);
			36117: out = 16'(342);
			36118: out = 16'(1564);
			36119: out = 16'(448);
			36120: out = 16'(-1221);
			36121: out = 16'(-1301);
			36122: out = 16'(-38);
			36123: out = 16'(177);
			36124: out = 16'(-266);
			36125: out = 16'(99);
			36126: out = 16'(1143);
			36127: out = 16'(1337);
			36128: out = 16'(-87);
			36129: out = 16'(-1062);
			36130: out = 16'(-556);
			36131: out = 16'(283);
			36132: out = 16'(-303);
			36133: out = 16'(-258);
			36134: out = 16'(1114);
			36135: out = 16'(1083);
			36136: out = 16'(422);
			36137: out = 16'(-190);
			36138: out = 16'(166);
			36139: out = 16'(472);
			36140: out = 16'(-479);
			36141: out = 16'(-1580);
			36142: out = 16'(-1286);
			36143: out = 16'(60);
			36144: out = 16'(764);
			36145: out = 16'(1065);
			36146: out = 16'(1096);
			36147: out = 16'(789);
			36148: out = 16'(333);
			36149: out = 16'(-738);
			36150: out = 16'(-1773);
			36151: out = 16'(-1760);
			36152: out = 16'(-37);
			36153: out = 16'(1373);
			36154: out = 16'(1548);
			36155: out = 16'(971);
			36156: out = 16'(239);
			36157: out = 16'(119);
			36158: out = 16'(-958);
			36159: out = 16'(-2087);
			36160: out = 16'(-865);
			36161: out = 16'(658);
			36162: out = 16'(1322);
			36163: out = 16'(156);
			36164: out = 16'(-1272);
			36165: out = 16'(-659);
			36166: out = 16'(525);
			36167: out = 16'(672);
			36168: out = 16'(-115);
			36169: out = 16'(-661);
			36170: out = 16'(-275);
			36171: out = 16'(181);
			36172: out = 16'(20);
			36173: out = 16'(-1623);
			36174: out = 16'(289);
			36175: out = 16'(1753);
			36176: out = 16'(1053);
			36177: out = 16'(-1300);
			36178: out = 16'(-1752);
			36179: out = 16'(-1139);
			36180: out = 16'(-782);
			36181: out = 16'(-1661);
			36182: out = 16'(-214);
			36183: out = 16'(1159);
			36184: out = 16'(2322);
			36185: out = 16'(1440);
			36186: out = 16'(-944);
			36187: out = 16'(-4278);
			36188: out = 16'(-3576);
			36189: out = 16'(496);
			36190: out = 16'(1834);
			36191: out = 16'(1650);
			36192: out = 16'(774);
			36193: out = 16'(327);
			36194: out = 16'(328);
			36195: out = 16'(-499);
			36196: out = 16'(-293);
			36197: out = 16'(-56);
			36198: out = 16'(-927);
			36199: out = 16'(-488);
			36200: out = 16'(575);
			36201: out = 16'(430);
			36202: out = 16'(-1297);
			36203: out = 16'(-89);
			36204: out = 16'(1271);
			36205: out = 16'(1234);
			36206: out = 16'(-556);
			36207: out = 16'(53);
			36208: out = 16'(4);
			36209: out = 16'(-75);
			36210: out = 16'(-145);
			36211: out = 16'(1204);
			36212: out = 16'(1624);
			36213: out = 16'(842);
			36214: out = 16'(-883);
			36215: out = 16'(-1198);
			36216: out = 16'(-2065);
			36217: out = 16'(-1077);
			36218: out = 16'(168);
			36219: out = 16'(977);
			36220: out = 16'(1458);
			36221: out = 16'(1618);
			36222: out = 16'(1233);
			36223: out = 16'(568);
			36224: out = 16'(-836);
			36225: out = 16'(-811);
			36226: out = 16'(-355);
			36227: out = 16'(71);
			36228: out = 16'(-67);
			36229: out = 16'(830);
			36230: out = 16'(614);
			36231: out = 16'(-320);
			36232: out = 16'(-884);
			36233: out = 16'(-265);
			36234: out = 16'(-142);
			36235: out = 16'(-367);
			36236: out = 16'(-27);
			36237: out = 16'(-339);
			36238: out = 16'(-163);
			36239: out = 16'(553);
			36240: out = 16'(1841);
			36241: out = 16'(935);
			36242: out = 16'(415);
			36243: out = 16'(-833);
			36244: out = 16'(-1398);
			36245: out = 16'(-463);
			36246: out = 16'(791);
			36247: out = 16'(587);
			36248: out = 16'(-209);
			36249: out = 16'(-361);
			36250: out = 16'(-27);
			36251: out = 16'(-635);
			36252: out = 16'(-1217);
			36253: out = 16'(-432);
			36254: out = 16'(1208);
			36255: out = 16'(990);
			36256: out = 16'(-296);
			36257: out = 16'(-453);
			36258: out = 16'(-214);
			36259: out = 16'(671);
			36260: out = 16'(155);
			36261: out = 16'(-1095);
			36262: out = 16'(-1138);
			36263: out = 16'(-381);
			36264: out = 16'(284);
			36265: out = 16'(107);
			36266: out = 16'(-218);
			36267: out = 16'(622);
			36268: out = 16'(1501);
			36269: out = 16'(874);
			36270: out = 16'(-961);
			36271: out = 16'(-1269);
			36272: out = 16'(-636);
			36273: out = 16'(-466);
			36274: out = 16'(-769);
			36275: out = 16'(577);
			36276: out = 16'(1448);
			36277: out = 16'(786);
			36278: out = 16'(-883);
			36279: out = 16'(-1425);
			36280: out = 16'(-540);
			36281: out = 16'(178);
			36282: out = 16'(-62);
			36283: out = 16'(101);
			36284: out = 16'(-55);
			36285: out = 16'(12);
			36286: out = 16'(10);
			36287: out = 16'(5);
			36288: out = 16'(-464);
			36289: out = 16'(-381);
			36290: out = 16'(590);
			36291: out = 16'(1371);
			36292: out = 16'(324);
			36293: out = 16'(-1452);
			36294: out = 16'(-1663);
			36295: out = 16'(19);
			36296: out = 16'(924);
			36297: out = 16'(954);
			36298: out = 16'(741);
			36299: out = 16'(726);
			36300: out = 16'(255);
			36301: out = 16'(-886);
			36302: out = 16'(-706);
			36303: out = 16'(820);
			36304: out = 16'(1541);
			36305: out = 16'(633);
			36306: out = 16'(-806);
			36307: out = 16'(-953);
			36308: out = 16'(80);
			36309: out = 16'(857);
			36310: out = 16'(928);
			36311: out = 16'(428);
			36312: out = 16'(-87);
			36313: out = 16'(154);
			36314: out = 16'(-735);
			36315: out = 16'(-1576);
			36316: out = 16'(-1132);
			36317: out = 16'(602);
			36318: out = 16'(1453);
			36319: out = 16'(1079);
			36320: out = 16'(875);
			36321: out = 16'(1553);
			36322: out = 16'(373);
			36323: out = 16'(-1756);
			36324: out = 16'(-2547);
			36325: out = 16'(-457);
			36326: out = 16'(34);
			36327: out = 16'(344);
			36328: out = 16'(98);
			36329: out = 16'(-20);
			36330: out = 16'(-47);
			36331: out = 16'(103);
			36332: out = 16'(387);
			36333: out = 16'(691);
			36334: out = 16'(-99);
			36335: out = 16'(-316);
			36336: out = 16'(-289);
			36337: out = 16'(56);
			36338: out = 16'(148);
			36339: out = 16'(219);
			36340: out = 16'(-173);
			36341: out = 16'(-487);
			36342: out = 16'(-676);
			36343: out = 16'(52);
			36344: out = 16'(-256);
			36345: out = 16'(-736);
			36346: out = 16'(-217);
			36347: out = 16'(-166);
			36348: out = 16'(592);
			36349: out = 16'(476);
			36350: out = 16'(-78);
			36351: out = 16'(-69);
			36352: out = 16'(542);
			36353: out = 16'(474);
			36354: out = 16'(-163);
			36355: out = 16'(191);
			36356: out = 16'(-293);
			36357: out = 16'(-574);
			36358: out = 16'(-577);
			36359: out = 16'(25);
			36360: out = 16'(556);
			36361: out = 16'(824);
			36362: out = 16'(443);
			36363: out = 16'(-97);
			36364: out = 16'(-86);
			36365: out = 16'(-240);
			36366: out = 16'(-514);
			36367: out = 16'(-304);
			36368: out = 16'(-159);
			36369: out = 16'(715);
			36370: out = 16'(750);
			36371: out = 16'(-221);
			36372: out = 16'(-1503);
			36373: out = 16'(-978);
			36374: out = 16'(-188);
			36375: out = 16'(213);
			36376: out = 16'(232);
			36377: out = 16'(837);
			36378: out = 16'(651);
			36379: out = 16'(-236);
			36380: out = 16'(-599);
			36381: out = 16'(-58);
			36382: out = 16'(735);
			36383: out = 16'(881);
			36384: out = 16'(569);
			36385: out = 16'(-645);
			36386: out = 16'(-572);
			36387: out = 16'(-399);
			36388: out = 16'(-516);
			36389: out = 16'(-1269);
			36390: out = 16'(-176);
			36391: out = 16'(350);
			36392: out = 16'(117);
			36393: out = 16'(-26);
			36394: out = 16'(-52);
			36395: out = 16'(-355);
			36396: out = 16'(-707);
			36397: out = 16'(-257);
			36398: out = 16'(530);
			36399: out = 16'(883);
			36400: out = 16'(248);
			36401: out = 16'(-719);
			36402: out = 16'(-416);
			36403: out = 16'(-41);
			36404: out = 16'(243);
			36405: out = 16'(145);
			36406: out = 16'(-28);
			36407: out = 16'(84);
			36408: out = 16'(181);
			36409: out = 16'(-315);
			36410: out = 16'(-860);
			36411: out = 16'(-689);
			36412: out = 16'(673);
			36413: out = 16'(1401);
			36414: out = 16'(639);
			36415: out = 16'(26);
			36416: out = 16'(-257);
			36417: out = 16'(-816);
			36418: out = 16'(-1531);
			36419: out = 16'(-1124);
			36420: out = 16'(779);
			36421: out = 16'(1946);
			36422: out = 16'(1361);
			36423: out = 16'(20);
			36424: out = 16'(-29);
			36425: out = 16'(48);
			36426: out = 16'(-38);
			36427: out = 16'(649);
			36428: out = 16'(109);
			36429: out = 16'(-779);
			36430: out = 16'(-1273);
			36431: out = 16'(-621);
			36432: out = 16'(1262);
			36433: out = 16'(1335);
			36434: out = 16'(29);
			36435: out = 16'(-1008);
			36436: out = 16'(-535);
			36437: out = 16'(-1073);
			36438: out = 16'(-1710);
			36439: out = 16'(-908);
			36440: out = 16'(478);
			36441: out = 16'(1136);
			36442: out = 16'(215);
			36443: out = 16'(-571);
			36444: out = 16'(695);
			36445: out = 16'(1308);
			36446: out = 16'(815);
			36447: out = 16'(-460);
			36448: out = 16'(-566);
			36449: out = 16'(-384);
			36450: out = 16'(501);
			36451: out = 16'(373);
			36452: out = 16'(-488);
			36453: out = 16'(-1553);
			36454: out = 16'(-696);
			36455: out = 16'(135);
			36456: out = 16'(122);
			36457: out = 16'(-88);
			36458: out = 16'(654);
			36459: out = 16'(657);
			36460: out = 16'(-199);
			36461: out = 16'(216);
			36462: out = 16'(528);
			36463: out = 16'(432);
			36464: out = 16'(-431);
			36465: out = 16'(-890);
			36466: out = 16'(-371);
			36467: out = 16'(437);
			36468: out = 16'(573);
			36469: out = 16'(58);
			36470: out = 16'(-374);
			36471: out = 16'(-332);
			36472: out = 16'(0);
			36473: out = 16'(124);
			36474: out = 16'(-32);
			36475: out = 16'(-217);
			36476: out = 16'(558);
			36477: out = 16'(1574);
			36478: out = 16'(-174);
			36479: out = 16'(-532);
			36480: out = 16'(-998);
			36481: out = 16'(-865);
			36482: out = 16'(-507);
			36483: out = 16'(538);
			36484: out = 16'(472);
			36485: out = 16'(90);
			36486: out = 16'(92);
			36487: out = 16'(-42);
			36488: out = 16'(-362);
			36489: out = 16'(-146);
			36490: out = 16'(745);
			36491: out = 16'(674);
			36492: out = 16'(-55);
			36493: out = 16'(-457);
			36494: out = 16'(361);
			36495: out = 16'(1209);
			36496: out = 16'(1207);
			36497: out = 16'(-70);
			36498: out = 16'(-1144);
			36499: out = 16'(-485);
			36500: out = 16'(-1133);
			36501: out = 16'(-1725);
			36502: out = 16'(-1692);
			36503: out = 16'(-285);
			36504: out = 16'(-216);
			36505: out = 16'(600);
			36506: out = 16'(754);
			36507: out = 16'(-199);
			36508: out = 16'(-335);
			36509: out = 16'(-463);
			36510: out = 16'(-466);
			36511: out = 16'(-734);
			36512: out = 16'(-638);
			36513: out = 16'(-509);
			36514: out = 16'(-77);
			36515: out = 16'(387);
			36516: out = 16'(996);
			36517: out = 16'(229);
			36518: out = 16'(-164);
			36519: out = 16'(169);
			36520: out = 16'(655);
			36521: out = 16'(-90);
			36522: out = 16'(-1297);
			36523: out = 16'(-1692);
			36524: out = 16'(-449);
			36525: out = 16'(-171);
			36526: out = 16'(692);
			36527: out = 16'(1021);
			36528: out = 16'(602);
			36529: out = 16'(-528);
			36530: out = 16'(-720);
			36531: out = 16'(-512);
			36532: out = 16'(-276);
			36533: out = 16'(-9);
			36534: out = 16'(565);
			36535: out = 16'(840);
			36536: out = 16'(606);
			36537: out = 16'(269);
			36538: out = 16'(760);
			36539: out = 16'(1319);
			36540: out = 16'(1068);
			36541: out = 16'(-230);
			36542: out = 16'(-587);
			36543: out = 16'(-823);
			36544: out = 16'(-475);
			36545: out = 16'(9);
			36546: out = 16'(882);
			36547: out = 16'(311);
			36548: out = 16'(-520);
			36549: out = 16'(-1049);
			36550: out = 16'(-1226);
			36551: out = 16'(-477);
			36552: out = 16'(736);
			36553: out = 16'(1395);
			36554: out = 16'(672);
			36555: out = 16'(-183);
			36556: out = 16'(-286);
			36557: out = 16'(376);
			36558: out = 16'(586);
			36559: out = 16'(101);
			36560: out = 16'(-400);
			36561: out = 16'(-298);
			36562: out = 16'(-79);
			36563: out = 16'(656);
			36564: out = 16'(4);
			36565: out = 16'(-569);
			36566: out = 16'(-459);
			36567: out = 16'(-1289);
			36568: out = 16'(-272);
			36569: out = 16'(557);
			36570: out = 16'(521);
			36571: out = 16'(-367);
			36572: out = 16'(-491);
			36573: out = 16'(-182);
			36574: out = 16'(-123);
			36575: out = 16'(-389);
			36576: out = 16'(-462);
			36577: out = 16'(242);
			36578: out = 16'(728);
			36579: out = 16'(89);
			36580: out = 16'(206);
			36581: out = 16'(-20);
			36582: out = 16'(-238);
			36583: out = 16'(-807);
			36584: out = 16'(-866);
			36585: out = 16'(-1052);
			36586: out = 16'(-513);
			36587: out = 16'(99);
			36588: out = 16'(775);
			36589: out = 16'(701);
			36590: out = 16'(807);
			36591: out = 16'(486);
			36592: out = 16'(-30);
			36593: out = 16'(-1380);
			36594: out = 16'(-1012);
			36595: out = 16'(-130);
			36596: out = 16'(200);
			36597: out = 16'(165);
			36598: out = 16'(649);
			36599: out = 16'(158);
			36600: out = 16'(-1329);
			36601: out = 16'(-983);
			36602: out = 16'(343);
			36603: out = 16'(1113);
			36604: out = 16'(625);
			36605: out = 16'(755);
			36606: out = 16'(196);
			36607: out = 16'(-927);
			36608: out = 16'(-1845);
			36609: out = 16'(-570);
			36610: out = 16'(-14);
			36611: out = 16'(14);
			36612: out = 16'(-495);
			36613: out = 16'(-271);
			36614: out = 16'(-413);
			36615: out = 16'(-102);
			36616: out = 16'(73);
			36617: out = 16'(269);
			36618: out = 16'(-64);
			36619: out = 16'(-238);
			36620: out = 16'(-398);
			36621: out = 16'(-256);
			36622: out = 16'(151);
			36623: out = 16'(110);
			36624: out = 16'(20);
			36625: out = 16'(377);
			36626: out = 16'(695);
			36627: out = 16'(1418);
			36628: out = 16'(798);
			36629: out = 16'(-660);
			36630: out = 16'(-2100);
			36631: out = 16'(-205);
			36632: out = 16'(376);
			36633: out = 16'(-78);
			36634: out = 16'(-305);
			36635: out = 16'(-69);
			36636: out = 16'(-155);
			36637: out = 16'(-537);
			36638: out = 16'(-524);
			36639: out = 16'(-61);
			36640: out = 16'(432);
			36641: out = 16'(344);
			36642: out = 16'(-130);
			36643: out = 16'(-299);
			36644: out = 16'(-389);
			36645: out = 16'(-154);
			36646: out = 16'(73);
			36647: out = 16'(303);
			36648: out = 16'(912);
			36649: out = 16'(577);
			36650: out = 16'(-546);
			36651: out = 16'(-977);
			36652: out = 16'(389);
			36653: out = 16'(2037);
			36654: out = 16'(1531);
			36655: out = 16'(-804);
			36656: out = 16'(-1959);
			36657: out = 16'(-1083);
			36658: out = 16'(184);
			36659: out = 16'(106);
			36660: out = 16'(141);
			36661: out = 16'(17);
			36662: out = 16'(980);
			36663: out = 16'(1357);
			36664: out = 16'(673);
			36665: out = 16'(-1170);
			36666: out = 16'(-1570);
			36667: out = 16'(-928);
			36668: out = 16'(-316);
			36669: out = 16'(-52);
			36670: out = 16'(459);
			36671: out = 16'(858);
			36672: out = 16'(668);
			36673: out = 16'(234);
			36674: out = 16'(164);
			36675: out = 16'(166);
			36676: out = 16'(-103);
			36677: out = 16'(262);
			36678: out = 16'(-860);
			36679: out = 16'(-1667);
			36680: out = 16'(-1497);
			36681: out = 16'(368);
			36682: out = 16'(-19);
			36683: out = 16'(446);
			36684: out = 16'(814);
			36685: out = 16'(723);
			36686: out = 16'(-259);
			36687: out = 16'(-190);
			36688: out = 16'(-8);
			36689: out = 16'(-24);
			36690: out = 16'(-76);
			36691: out = 16'(60);
			36692: out = 16'(-613);
			36693: out = 16'(-1627);
			36694: out = 16'(-1481);
			36695: out = 16'(-373);
			36696: out = 16'(270);
			36697: out = 16'(404);
			36698: out = 16'(1075);
			36699: out = 16'(861);
			36700: out = 16'(237);
			36701: out = 16'(-638);
			36702: out = 16'(-1164);
			36703: out = 16'(-937);
			36704: out = 16'(-376);
			36705: out = 16'(625);
			36706: out = 16'(1462);
			36707: out = 16'(227);
			36708: out = 16'(-710);
			36709: out = 16'(-456);
			36710: out = 16'(340);
			36711: out = 16'(70);
			36712: out = 16'(-1077);
			36713: out = 16'(-1125);
			36714: out = 16'(-15);
			36715: out = 16'(-19);
			36716: out = 16'(325);
			36717: out = 16'(424);
			36718: out = 16'(578);
			36719: out = 16'(240);
			36720: out = 16'(114);
			36721: out = 16'(-31);
			36722: out = 16'(56);
			36723: out = 16'(24);
			36724: out = 16'(256);
			36725: out = 16'(605);
			36726: out = 16'(697);
			36727: out = 16'(109);
			36728: out = 16'(41);
			36729: out = 16'(-928);
			36730: out = 16'(-1252);
			36731: out = 16'(-1048);
			36732: out = 16'(-255);
			36733: out = 16'(-91);
			36734: out = 16'(906);
			36735: out = 16'(1897);
			36736: out = 16'(1376);
			36737: out = 16'(964);
			36738: out = 16'(241);
			36739: out = 16'(-226);
			36740: out = 16'(-768);
			36741: out = 16'(-1664);
			36742: out = 16'(-1446);
			36743: out = 16'(-157);
			36744: out = 16'(898);
			36745: out = 16'(1738);
			36746: out = 16'(1055);
			36747: out = 16'(500);
			36748: out = 16'(-110);
			36749: out = 16'(-1154);
			36750: out = 16'(-2697);
			36751: out = 16'(-2713);
			36752: out = 16'(-1071);
			36753: out = 16'(864);
			36754: out = 16'(1987);
			36755: out = 16'(2030);
			36756: out = 16'(835);
			36757: out = 16'(-637);
			36758: out = 16'(-1770);
			36759: out = 16'(-918);
			36760: out = 16'(-241);
			36761: out = 16'(-529);
			36762: out = 16'(232);
			36763: out = 16'(914);
			36764: out = 16'(530);
			36765: out = 16'(-760);
			36766: out = 16'(-506);
			36767: out = 16'(-586);
			36768: out = 16'(-706);
			36769: out = 16'(-558);
			36770: out = 16'(887);
			36771: out = 16'(1450);
			36772: out = 16'(1003);
			36773: out = 16'(-30);
			36774: out = 16'(134);
			36775: out = 16'(-370);
			36776: out = 16'(-78);
			36777: out = 16'(48);
			36778: out = 16'(191);
			36779: out = 16'(-1112);
			36780: out = 16'(-460);
			36781: out = 16'(411);
			36782: out = 16'(853);
			36783: out = 16'(745);
			36784: out = 16'(1010);
			36785: out = 16'(508);
			36786: out = 16'(-888);
			36787: out = 16'(-2655);
			36788: out = 16'(-1714);
			36789: out = 16'(58);
			36790: out = 16'(1355);
			36791: out = 16'(1409);
			36792: out = 16'(815);
			36793: out = 16'(-533);
			36794: out = 16'(-1258);
			36795: out = 16'(-829);
			36796: out = 16'(-907);
			36797: out = 16'(-539);
			36798: out = 16'(217);
			36799: out = 16'(1243);
			36800: out = 16'(1685);
			36801: out = 16'(1180);
			36802: out = 16'(335);
			36803: out = 16'(-185);
			36804: out = 16'(-1201);
			36805: out = 16'(-570);
			36806: out = 16'(-35);
			36807: out = 16'(275);
			36808: out = 16'(250);
			36809: out = 16'(91);
			36810: out = 16'(-221);
			36811: out = 16'(-265);
			36812: out = 16'(58);
			36813: out = 16'(698);
			36814: out = 16'(219);
			36815: out = 16'(-885);
			36816: out = 16'(-1388);
			36817: out = 16'(-458);
			36818: out = 16'(676);
			36819: out = 16'(1165);
			36820: out = 16'(811);
			36821: out = 16'(-292);
			36822: out = 16'(-608);
			36823: out = 16'(-626);
			36824: out = 16'(-627);
			36825: out = 16'(-579);
			36826: out = 16'(-105);
			36827: out = 16'(208);
			36828: out = 16'(386);
			36829: out = 16'(856);
			36830: out = 16'(754);
			36831: out = 16'(808);
			36832: out = 16'(562);
			36833: out = 16'(208);
			36834: out = 16'(-63);
			36835: out = 16'(-14);
			36836: out = 16'(-551);
			36837: out = 16'(-1271);
			36838: out = 16'(-922);
			36839: out = 16'(442);
			36840: out = 16'(1439);
			36841: out = 16'(1181);
			36842: out = 16'(-51);
			36843: out = 16'(114);
			36844: out = 16'(-222);
			36845: out = 16'(-811);
			36846: out = 16'(-536);
			36847: out = 16'(-5);
			36848: out = 16'(1055);
			36849: out = 16'(1355);
			36850: out = 16'(479);
			36851: out = 16'(-747);
			36852: out = 16'(-1330);
			36853: out = 16'(-799);
			36854: out = 16'(153);
			36855: out = 16'(922);
			36856: out = 16'(813);
			36857: out = 16'(493);
			36858: out = 16'(35);
			36859: out = 16'(-371);
			36860: out = 16'(-1128);
			36861: out = 16'(-1057);
			36862: out = 16'(-422);
			36863: out = 16'(213);
			36864: out = 16'(616);
			36865: out = 16'(939);
			36866: out = 16'(735);
			36867: out = 16'(33);
			36868: out = 16'(-1945);
			36869: out = 16'(-1417);
			36870: out = 16'(98);
			36871: out = 16'(1033);
			36872: out = 16'(954);
			36873: out = 16'(845);
			36874: out = 16'(225);
			36875: out = 16'(-545);
			36876: out = 16'(-697);
			36877: out = 16'(-464);
			36878: out = 16'(-535);
			36879: out = 16'(-533);
			36880: out = 16'(168);
			36881: out = 16'(-266);
			36882: out = 16'(-464);
			36883: out = 16'(-7);
			36884: out = 16'(692);
			36885: out = 16'(166);
			36886: out = 16'(-1361);
			36887: out = 16'(-2041);
			36888: out = 16'(-862);
			36889: out = 16'(21);
			36890: out = 16'(1223);
			36891: out = 16'(1863);
			36892: out = 16'(1838);
			36893: out = 16'(198);
			36894: out = 16'(-426);
			36895: out = 16'(-453);
			36896: out = 16'(69);
			36897: out = 16'(-186);
			36898: out = 16'(-542);
			36899: out = 16'(-1456);
			36900: out = 16'(-1171);
			36901: out = 16'(278);
			36902: out = 16'(1425);
			36903: out = 16'(668);
			36904: out = 16'(-244);
			36905: out = 16'(81);
			36906: out = 16'(-130);
			36907: out = 16'(-122);
			36908: out = 16'(-639);
			36909: out = 16'(-704);
			36910: out = 16'(-408);
			36911: out = 16'(642);
			36912: out = 16'(850);
			36913: out = 16'(510);
			36914: out = 16'(-80);
			36915: out = 16'(206);
			36916: out = 16'(-347);
			36917: out = 16'(-848);
			36918: out = 16'(-209);
			36919: out = 16'(1046);
			36920: out = 16'(1074);
			36921: out = 16'(119);
			36922: out = 16'(-674);
			36923: out = 16'(-1336);
			36924: out = 16'(-592);
			36925: out = 16'(601);
			36926: out = 16'(1273);
			36927: out = 16'(875);
			36928: out = 16'(-195);
			36929: out = 16'(-974);
			36930: out = 16'(-1057);
			36931: out = 16'(-830);
			36932: out = 16'(-218);
			36933: out = 16'(398);
			36934: out = 16'(560);
			36935: out = 16'(-80);
			36936: out = 16'(-8);
			36937: out = 16'(70);
			36938: out = 16'(366);
			36939: out = 16'(647);
			36940: out = 16'(849);
			36941: out = 16'(299);
			36942: out = 16'(-367);
			36943: out = 16'(-650);
			36944: out = 16'(-1138);
			36945: out = 16'(-759);
			36946: out = 16'(-285);
			36947: out = 16'(332);
			36948: out = 16'(544);
			36949: out = 16'(263);
			36950: out = 16'(-932);
			36951: out = 16'(-1568);
			36952: out = 16'(-748);
			36953: out = 16'(466);
			36954: out = 16'(410);
			36955: out = 16'(-157);
			36956: out = 16'(127);
			36957: out = 16'(1300);
			36958: out = 16'(1137);
			36959: out = 16'(0);
			36960: out = 16'(-835);
			36961: out = 16'(-174);
			36962: out = 16'(-367);
			36963: out = 16'(-890);
			36964: out = 16'(-891);
			36965: out = 16'(142);
			36966: out = 16'(254);
			36967: out = 16'(104);
			36968: out = 16'(84);
			36969: out = 16'(691);
			36970: out = 16'(69);
			36971: out = 16'(-31);
			36972: out = 16'(-165);
			36973: out = 16'(-603);
			36974: out = 16'(-1272);
			36975: out = 16'(-217);
			36976: out = 16'(1248);
			36977: out = 16'(1267);
			36978: out = 16'(227);
			36979: out = 16'(-1225);
			36980: out = 16'(-1487);
			36981: out = 16'(-898);
			36982: out = 16'(-284);
			36983: out = 16'(-80);
			36984: out = 16'(694);
			36985: out = 16'(1728);
			36986: out = 16'(1368);
			36987: out = 16'(202);
			36988: out = 16'(-1031);
			36989: out = 16'(-462);
			36990: out = 16'(1280);
			36991: out = 16'(840);
			36992: out = 16'(-326);
			36993: out = 16'(-730);
			36994: out = 16'(24);
			36995: out = 16'(-329);
			36996: out = 16'(-376);
			36997: out = 16'(76);
			36998: out = 16'(947);
			36999: out = 16'(587);
			37000: out = 16'(-324);
			37001: out = 16'(-1200);
			37002: out = 16'(-811);
			37003: out = 16'(-121);
			37004: out = 16'(637);
			37005: out = 16'(258);
			37006: out = 16'(116);
			37007: out = 16'(862);
			37008: out = 16'(713);
			37009: out = 16'(43);
			37010: out = 16'(-381);
			37011: out = 16'(-53);
			37012: out = 16'(-791);
			37013: out = 16'(-630);
			37014: out = 16'(93);
			37015: out = 16'(564);
			37016: out = 16'(-255);
			37017: out = 16'(-805);
			37018: out = 16'(-263);
			37019: out = 16'(726);
			37020: out = 16'(-115);
			37021: out = 16'(516);
			37022: out = 16'(406);
			37023: out = 16'(-559);
			37024: out = 16'(-2091);
			37025: out = 16'(-758);
			37026: out = 16'(552);
			37027: out = 16'(525);
			37028: out = 16'(-839);
			37029: out = 16'(32);
			37030: out = 16'(900);
			37031: out = 16'(1238);
			37032: out = 16'(489);
			37033: out = 16'(735);
			37034: out = 16'(-111);
			37035: out = 16'(-557);
			37036: out = 16'(-967);
			37037: out = 16'(-723);
			37038: out = 16'(-992);
			37039: out = 16'(29);
			37040: out = 16'(935);
			37041: out = 16'(644);
			37042: out = 16'(-991);
			37043: out = 16'(-964);
			37044: out = 16'(-130);
			37045: out = 16'(-394);
			37046: out = 16'(-696);
			37047: out = 16'(-279);
			37048: out = 16'(545);
			37049: out = 16'(635);
			37050: out = 16'(912);
			37051: out = 16'(719);
			37052: out = 16'(408);
			37053: out = 16'(-70);
			37054: out = 16'(641);
			37055: out = 16'(-420);
			37056: out = 16'(-1116);
			37057: out = 16'(-877);
			37058: out = 16'(-75);
			37059: out = 16'(43);
			37060: out = 16'(-84);
			37061: out = 16'(170);
			37062: out = 16'(597);
			37063: out = 16'(186);
			37064: out = 16'(-1019);
			37065: out = 16'(-1533);
			37066: out = 16'(-594);
			37067: out = 16'(514);
			37068: out = 16'(793);
			37069: out = 16'(629);
			37070: out = 16'(640);
			37071: out = 16'(-47);
			37072: out = 16'(-214);
			37073: out = 16'(-387);
			37074: out = 16'(-279);
			37075: out = 16'(-367);
			37076: out = 16'(642);
			37077: out = 16'(866);
			37078: out = 16'(386);
			37079: out = 16'(-373);
			37080: out = 16'(-362);
			37081: out = 16'(-209);
			37082: out = 16'(182);
			37083: out = 16'(640);
			37084: out = 16'(652);
			37085: out = 16'(189);
			37086: out = 16'(-80);
			37087: out = 16'(102);
			37088: out = 16'(-1105);
			37089: out = 16'(-424);
			37090: out = 16'(331);
			37091: out = 16'(541);
			37092: out = 16'(-54);
			37093: out = 16'(425);
			37094: out = 16'(805);
			37095: out = 16'(492);
			37096: out = 16'(-905);
			37097: out = 16'(-261);
			37098: out = 16'(433);
			37099: out = 16'(777);
			37100: out = 16'(-81);
			37101: out = 16'(-600);
			37102: out = 16'(-1474);
			37103: out = 16'(-494);
			37104: out = 16'(1403);
			37105: out = 16'(1466);
			37106: out = 16'(-783);
			37107: out = 16'(-2369);
			37108: out = 16'(-1361);
			37109: out = 16'(458);
			37110: out = 16'(962);
			37111: out = 16'(672);
			37112: out = 16'(555);
			37113: out = 16'(-202);
			37114: out = 16'(44);
			37115: out = 16'(-731);
			37116: out = 16'(-1057);
			37117: out = 16'(-548);
			37118: out = 16'(529);
			37119: out = 16'(265);
			37120: out = 16'(-155);
			37121: out = 16'(75);
			37122: out = 16'(1359);
			37123: out = 16'(349);
			37124: out = 16'(-939);
			37125: out = 16'(-879);
			37126: out = 16'(522);
			37127: out = 16'(680);
			37128: out = 16'(359);
			37129: out = 16'(-57);
			37130: out = 16'(-371);
			37131: out = 16'(-430);
			37132: out = 16'(-212);
			37133: out = 16'(-87);
			37134: out = 16'(-32);
			37135: out = 16'(53);
			37136: out = 16'(251);
			37137: out = 16'(-496);
			37138: out = 16'(-1641);
			37139: out = 16'(-510);
			37140: out = 16'(404);
			37141: out = 16'(507);
			37142: out = 16'(203);
			37143: out = 16'(594);
			37144: out = 16'(701);
			37145: out = 16'(12);
			37146: out = 16'(-618);
			37147: out = 16'(-154);
			37148: out = 16'(-246);
			37149: out = 16'(-826);
			37150: out = 16'(-890);
			37151: out = 16'(-37);
			37152: out = 16'(236);
			37153: out = 16'(-671);
			37154: out = 16'(-512);
			37155: out = 16'(1531);
			37156: out = 16'(1738);
			37157: out = 16'(877);
			37158: out = 16'(-426);
			37159: out = 16'(-936);
			37160: out = 16'(-1397);
			37161: out = 16'(-1077);
			37162: out = 16'(62);
			37163: out = 16'(1544);
			37164: out = 16'(1303);
			37165: out = 16'(16);
			37166: out = 16'(-1339);
			37167: out = 16'(-819);
			37168: out = 16'(814);
			37169: out = 16'(935);
			37170: out = 16'(98);
			37171: out = 16'(-457);
			37172: out = 16'(-368);
			37173: out = 16'(-46);
			37174: out = 16'(-319);
			37175: out = 16'(-10);
			37176: out = 16'(995);
			37177: out = 16'(1358);
			37178: out = 16'(1041);
			37179: out = 16'(348);
			37180: out = 16'(-364);
			37181: out = 16'(-1128);
			37182: out = 16'(-1473);
			37183: out = 16'(-821);
			37184: out = 16'(186);
			37185: out = 16'(551);
			37186: out = 16'(252);
			37187: out = 16'(-12);
			37188: out = 16'(-219);
			37189: out = 16'(-672);
			37190: out = 16'(-841);
			37191: out = 16'(-312);
			37192: out = 16'(533);
			37193: out = 16'(737);
			37194: out = 16'(263);
			37195: out = 16'(-560);
			37196: out = 16'(-1048);
			37197: out = 16'(-1021);
			37198: out = 16'(-353);
			37199: out = 16'(-99);
			37200: out = 16'(20);
			37201: out = 16'(-181);
			37202: out = 16'(-781);
			37203: out = 16'(-226);
			37204: out = 16'(423);
			37205: out = 16'(690);
			37206: out = 16'(632);
			37207: out = 16'(23);
			37208: out = 16'(-32);
			37209: out = 16'(-276);
			37210: out = 16'(-911);
			37211: out = 16'(-1058);
			37212: out = 16'(-344);
			37213: out = 16'(596);
			37214: out = 16'(783);
			37215: out = 16'(206);
			37216: out = 16'(-9);
			37217: out = 16'(-135);
			37218: out = 16'(-554);
			37219: out = 16'(-1292);
			37220: out = 16'(-1021);
			37221: out = 16'(-13);
			37222: out = 16'(760);
			37223: out = 16'(97);
			37224: out = 16'(103);
			37225: out = 16'(-588);
			37226: out = 16'(-540);
			37227: out = 16'(323);
			37228: out = 16'(638);
			37229: out = 16'(835);
			37230: out = 16'(722);
			37231: out = 16'(0);
			37232: out = 16'(-168);
			37233: out = 16'(-1376);
			37234: out = 16'(-1166);
			37235: out = 16'(-56);
			37236: out = 16'(690);
			37237: out = 16'(99);
			37238: out = 16'(295);
			37239: out = 16'(616);
			37240: out = 16'(193);
			37241: out = 16'(-520);
			37242: out = 16'(99);
			37243: out = 16'(606);
			37244: out = 16'(-148);
			37245: out = 16'(-750);
			37246: out = 16'(30);
			37247: out = 16'(853);
			37248: out = 16'(438);
			37249: out = 16'(-710);
			37250: out = 16'(-253);
			37251: out = 16'(241);
			37252: out = 16'(-154);
			37253: out = 16'(26);
			37254: out = 16'(-64);
			37255: out = 16'(-26);
			37256: out = 16'(71);
			37257: out = 16'(649);
			37258: out = 16'(314);
			37259: out = 16'(-501);
			37260: out = 16'(-1216);
			37261: out = 16'(-661);
			37262: out = 16'(-13);
			37263: out = 16'(968);
			37264: out = 16'(1231);
			37265: out = 16'(626);
			37266: out = 16'(-910);
			37267: out = 16'(-1117);
			37268: out = 16'(-133);
			37269: out = 16'(1036);
			37270: out = 16'(1201);
			37271: out = 16'(375);
			37272: out = 16'(-678);
			37273: out = 16'(-1034);
			37274: out = 16'(-364);
			37275: out = 16'(-77);
			37276: out = 16'(-49);
			37277: out = 16'(110);
			37278: out = 16'(643);
			37279: out = 16'(33);
			37280: out = 16'(-493);
			37281: out = 16'(-1095);
			37282: out = 16'(-1257);
			37283: out = 16'(-483);
			37284: out = 16'(463);
			37285: out = 16'(482);
			37286: out = 16'(-143);
			37287: out = 16'(-501);
			37288: out = 16'(-424);
			37289: out = 16'(-49);
			37290: out = 16'(370);
			37291: out = 16'(633);
			37292: out = 16'(728);
			37293: out = 16'(295);
			37294: out = 16'(-178);
			37295: out = 16'(-629);
			37296: out = 16'(-312);
			37297: out = 16'(-783);
			37298: out = 16'(-816);
			37299: out = 16'(347);
			37300: out = 16'(775);
			37301: out = 16'(450);
			37302: out = 16'(-533);
			37303: out = 16'(-983);
			37304: out = 16'(-363);
			37305: out = 16'(419);
			37306: out = 16'(867);
			37307: out = 16'(747);
			37308: out = 16'(-23);
			37309: out = 16'(-807);
			37310: out = 16'(-1222);
			37311: out = 16'(-765);
			37312: out = 16'(29);
			37313: out = 16'(609);
			37314: out = 16'(717);
			37315: out = 16'(527);
			37316: out = 16'(-117);
			37317: out = 16'(32);
			37318: out = 16'(-756);
			37319: out = 16'(-922);
			37320: out = 16'(-35);
			37321: out = 16'(1427);
			37322: out = 16'(1018);
			37323: out = 16'(342);
			37324: out = 16'(116);
			37325: out = 16'(-39);
			37326: out = 16'(-265);
			37327: out = 16'(-239);
			37328: out = 16'(136);
			37329: out = 16'(641);
			37330: out = 16'(257);
			37331: out = 16'(40);
			37332: out = 16'(-172);
			37333: out = 16'(-318);
			37334: out = 16'(-439);
			37335: out = 16'(316);
			37336: out = 16'(408);
			37337: out = 16'(-472);
			37338: out = 16'(-555);
			37339: out = 16'(-444);
			37340: out = 16'(-332);
			37341: out = 16'(-90);
			37342: out = 16'(1234);
			37343: out = 16'(1534);
			37344: out = 16'(553);
			37345: out = 16'(-846);
			37346: out = 16'(-234);
			37347: out = 16'(-706);
			37348: out = 16'(-156);
			37349: out = 16'(310);
			37350: out = 16'(635);
			37351: out = 16'(154);
			37352: out = 16'(92);
			37353: out = 16'(41);
			37354: out = 16'(-128);
			37355: out = 16'(-824);
			37356: out = 16'(-577);
			37357: out = 16'(-181);
			37358: out = 16'(-28);
			37359: out = 16'(-83);
			37360: out = 16'(122);
			37361: out = 16'(-85);
			37362: out = 16'(-333);
			37363: out = 16'(-30);
			37364: out = 16'(113);
			37365: out = 16'(-80);
			37366: out = 16'(-473);
			37367: out = 16'(-578);
			37368: out = 16'(-1027);
			37369: out = 16'(-714);
			37370: out = 16'(116);
			37371: out = 16'(641);
			37372: out = 16'(318);
			37373: out = 16'(-349);
			37374: out = 16'(-323);
			37375: out = 16'(194);
			37376: out = 16'(-786);
			37377: out = 16'(-1533);
			37378: out = 16'(-1661);
			37379: out = 16'(-628);
			37380: out = 16'(-48);
			37381: out = 16'(931);
			37382: out = 16'(486);
			37383: out = 16'(149);
			37384: out = 16'(718);
			37385: out = 16'(217);
			37386: out = 16'(-643);
			37387: out = 16'(-815);
			37388: out = 16'(260);
			37389: out = 16'(1382);
			37390: out = 16'(1175);
			37391: out = 16'(124);
			37392: out = 16'(-512);
			37393: out = 16'(-41);
			37394: out = 16'(30);
			37395: out = 16'(33);
			37396: out = 16'(217);
			37397: out = 16'(-44);
			37398: out = 16'(40);
			37399: out = 16'(-173);
			37400: out = 16'(-427);
			37401: out = 16'(-1073);
			37402: out = 16'(16);
			37403: out = 16'(188);
			37404: out = 16'(-142);
			37405: out = 16'(-489);
			37406: out = 16'(799);
			37407: out = 16'(820);
			37408: out = 16'(662);
			37409: out = 16'(652);
			37410: out = 16'(710);
			37411: out = 16'(-61);
			37412: out = 16'(-329);
			37413: out = 16'(-23);
			37414: out = 16'(-24);
			37415: out = 16'(-800);
			37416: out = 16'(-750);
			37417: out = 16'(347);
			37418: out = 16'(1272);
			37419: out = 16'(814);
			37420: out = 16'(586);
			37421: out = 16'(515);
			37422: out = 16'(-250);
			37423: out = 16'(-1342);
			37424: out = 16'(-1728);
			37425: out = 16'(-532);
			37426: out = 16'(959);
			37427: out = 16'(898);
			37428: out = 16'(251);
			37429: out = 16'(-128);
			37430: out = 16'(-40);
			37431: out = 16'(-358);
			37432: out = 16'(-333);
			37433: out = 16'(-447);
			37434: out = 16'(-510);
			37435: out = 16'(10);
			37436: out = 16'(-50);
			37437: out = 16'(39);
			37438: out = 16'(-141);
			37439: out = 16'(-248);
			37440: out = 16'(-123);
			37441: out = 16'(483);
			37442: out = 16'(419);
			37443: out = 16'(-410);
			37444: out = 16'(-781);
			37445: out = 16'(-201);
			37446: out = 16'(328);
			37447: out = 16'(111);
			37448: out = 16'(-516);
			37449: out = 16'(-169);
			37450: out = 16'(-24);
			37451: out = 16'(-465);
			37452: out = 16'(-992);
			37453: out = 16'(-93);
			37454: out = 16'(637);
			37455: out = 16'(540);
			37456: out = 16'(-15);
			37457: out = 16'(-254);
			37458: out = 16'(-151);
			37459: out = 16'(128);
			37460: out = 16'(161);
			37461: out = 16'(-154);
			37462: out = 16'(-861);
			37463: out = 16'(-755);
			37464: out = 16'(100);
			37465: out = 16'(218);
			37466: out = 16'(139);
			37467: out = 16'(-14);
			37468: out = 16'(-50);
			37469: out = 16'(-741);
			37470: out = 16'(-188);
			37471: out = 16'(529);
			37472: out = 16'(834);
			37473: out = 16'(-33);
			37474: out = 16'(210);
			37475: out = 16'(84);
			37476: out = 16'(53);
			37477: out = 16'(243);
			37478: out = 16'(39);
			37479: out = 16'(-28);
			37480: out = 16'(80);
			37481: out = 16'(234);
			37482: out = 16'(-3);
			37483: out = 16'(115);
			37484: out = 16'(155);
			37485: out = 16'(-146);
			37486: out = 16'(-746);
			37487: out = 16'(-303);
			37488: out = 16'(534);
			37489: out = 16'(689);
			37490: out = 16'(-567);
			37491: out = 16'(-26);
			37492: out = 16'(616);
			37493: out = 16'(726);
			37494: out = 16'(-109);
			37495: out = 16'(10);
			37496: out = 16'(-350);
			37497: out = 16'(-735);
			37498: out = 16'(-737);
			37499: out = 16'(-118);
			37500: out = 16'(602);
			37501: out = 16'(893);
			37502: out = 16'(493);
			37503: out = 16'(29);
			37504: out = 16'(-132);
			37505: out = 16'(91);
			37506: out = 16'(-42);
			37507: out = 16'(-541);
			37508: out = 16'(-253);
			37509: out = 16'(389);
			37510: out = 16'(524);
			37511: out = 16'(112);
			37512: out = 16'(-787);
			37513: out = 16'(-327);
			37514: out = 16'(202);
			37515: out = 16'(-100);
			37516: out = 16'(-43);
			37517: out = 16'(404);
			37518: out = 16'(494);
			37519: out = 16'(-128);
			37520: out = 16'(674);
			37521: out = 16'(120);
			37522: out = 16'(-245);
			37523: out = 16'(-244);
			37524: out = 16'(620);
			37525: out = 16'(255);
			37526: out = 16'(19);
			37527: out = 16'(-103);
			37528: out = 16'(-90);
			37529: out = 16'(-352);
			37530: out = 16'(-238);
			37531: out = 16'(38);
			37532: out = 16'(99);
			37533: out = 16'(-287);
			37534: out = 16'(-897);
			37535: out = 16'(-1035);
			37536: out = 16'(-449);
			37537: out = 16'(-134);
			37538: out = 16'(37);
			37539: out = 16'(-198);
			37540: out = 16'(-267);
			37541: out = 16'(-67);
			37542: out = 16'(544);
			37543: out = 16'(366);
			37544: out = 16'(-179);
			37545: out = 16'(-320);
			37546: out = 16'(72);
			37547: out = 16'(-329);
			37548: out = 16'(-934);
			37549: out = 16'(-398);
			37550: out = 16'(-178);
			37551: out = 16'(257);
			37552: out = 16'(-79);
			37553: out = 16'(-195);
			37554: out = 16'(-137);
			37555: out = 16'(1022);
			37556: out = 16'(947);
			37557: out = 16'(-95);
			37558: out = 16'(-804);
			37559: out = 16'(-431);
			37560: out = 16'(-466);
			37561: out = 16'(-643);
			37562: out = 16'(32);
			37563: out = 16'(522);
			37564: out = 16'(393);
			37565: out = 16'(278);
			37566: out = 16'(763);
			37567: out = 16'(638);
			37568: out = 16'(-388);
			37569: out = 16'(-875);
			37570: out = 16'(151);
			37571: out = 16'(39);
			37572: out = 16'(215);
			37573: out = 16'(2);
			37574: out = 16'(-54);
			37575: out = 16'(-553);
			37576: out = 16'(-59);
			37577: out = 16'(347);
			37578: out = 16'(605);
			37579: out = 16'(485);
			37580: out = 16'(105);
			37581: out = 16'(-297);
			37582: out = 16'(-243);
			37583: out = 16'(-53);
			37584: out = 16'(667);
			37585: out = 16'(289);
			37586: out = 16'(-243);
			37587: out = 16'(-296);
			37588: out = 16'(94);
			37589: out = 16'(-252);
			37590: out = 16'(-891);
			37591: out = 16'(-1132);
			37592: out = 16'(-335);
			37593: out = 16'(323);
			37594: out = 16'(771);
			37595: out = 16'(478);
			37596: out = 16'(-502);
			37597: out = 16'(-1323);
			37598: out = 16'(-1025);
			37599: out = 16'(-224);
			37600: out = 16'(177);
			37601: out = 16'(510);
			37602: out = 16'(963);
			37603: out = 16'(913);
			37604: out = 16'(22);
			37605: out = 16'(144);
			37606: out = 16'(4);
			37607: out = 16'(-257);
			37608: out = 16'(-829);
			37609: out = 16'(-668);
			37610: out = 16'(-177);
			37611: out = 16'(782);
			37612: out = 16'(1331);
			37613: out = 16'(1260);
			37614: out = 16'(240);
			37615: out = 16'(-322);
			37616: out = 16'(-221);
			37617: out = 16'(114);
			37618: out = 16'(-444);
			37619: out = 16'(-367);
			37620: out = 16'(231);
			37621: out = 16'(647);
			37622: out = 16'(31);
			37623: out = 16'(-419);
			37624: out = 16'(-590);
			37625: out = 16'(-495);
			37626: out = 16'(-87);
			37627: out = 16'(70);
			37628: out = 16'(47);
			37629: out = 16'(-83);
			37630: out = 16'(-47);
			37631: out = 16'(95);
			37632: out = 16'(96);
			37633: out = 16'(-129);
			37634: out = 16'(-8);
			37635: out = 16'(52);
			37636: out = 16'(417);
			37637: out = 16'(434);
			37638: out = 16'(112);
			37639: out = 16'(-315);
			37640: out = 16'(-52);
			37641: out = 16'(161);
			37642: out = 16'(49);
			37643: out = 16'(-948);
			37644: out = 16'(-575);
			37645: out = 16'(-321);
			37646: out = 16'(-532);
			37647: out = 16'(-78);
			37648: out = 16'(910);
			37649: out = 16'(1369);
			37650: out = 16'(717);
			37651: out = 16'(-316);
			37652: out = 16'(-1110);
			37653: out = 16'(-1285);
			37654: out = 16'(-1009);
			37655: out = 16'(-180);
			37656: out = 16'(1021);
			37657: out = 16'(1447);
			37658: out = 16'(796);
			37659: out = 16'(-257);
			37660: out = 16'(-944);
			37661: out = 16'(-750);
			37662: out = 16'(-416);
			37663: out = 16'(-277);
			37664: out = 16'(-69);
			37665: out = 16'(515);
			37666: out = 16'(750);
			37667: out = 16'(308);
			37668: out = 16'(-288);
			37669: out = 16'(-205);
			37670: out = 16'(289);
			37671: out = 16'(381);
			37672: out = 16'(-389);
			37673: out = 16'(409);
			37674: out = 16'(137);
			37675: out = 16'(-806);
			37676: out = 16'(-1354);
			37677: out = 16'(-77);
			37678: out = 16'(870);
			37679: out = 16'(837);
			37680: out = 16'(-48);
			37681: out = 16'(-436);
			37682: out = 16'(-954);
			37683: out = 16'(-631);
			37684: out = 16'(122);
			37685: out = 16'(503);
			37686: out = 16'(-50);
			37687: out = 16'(-651);
			37688: out = 16'(-655);
			37689: out = 16'(-298);
			37690: out = 16'(449);
			37691: out = 16'(394);
			37692: out = 16'(-197);
			37693: out = 16'(-707);
			37694: out = 16'(41);
			37695: out = 16'(761);
			37696: out = 16'(1222);
			37697: out = 16'(882);
			37698: out = 16'(231);
			37699: out = 16'(-795);
			37700: out = 16'(-717);
			37701: out = 16'(17);
			37702: out = 16'(-122);
			37703: out = 16'(-245);
			37704: out = 16'(-381);
			37705: out = 16'(-263);
			37706: out = 16'(-38);
			37707: out = 16'(375);
			37708: out = 16'(741);
			37709: out = 16'(329);
			37710: out = 16'(-798);
			37711: out = 16'(-268);
			37712: out = 16'(769);
			37713: out = 16'(1166);
			37714: out = 16'(308);
			37715: out = 16'(163);
			37716: out = 16'(-448);
			37717: out = 16'(-618);
			37718: out = 16'(-526);
			37719: out = 16'(-105);
			37720: out = 16'(-99);
			37721: out = 16'(-84);
			37722: out = 16'(-130);
			37723: out = 16'(-339);
			37724: out = 16'(-164);
			37725: out = 16'(216);
			37726: out = 16'(588);
			37727: out = 16'(429);
			37728: out = 16'(567);
			37729: out = 16'(-43);
			37730: out = 16'(-470);
			37731: out = 16'(-296);
			37732: out = 16'(429);
			37733: out = 16'(127);
			37734: out = 16'(-205);
			37735: out = 16'(-15);
			37736: out = 16'(432);
			37737: out = 16'(98);
			37738: out = 16'(-395);
			37739: out = 16'(-516);
			37740: out = 16'(50);
			37741: out = 16'(374);
			37742: out = 16'(557);
			37743: out = 16'(283);
			37744: out = 16'(-106);
			37745: out = 16'(-410);
			37746: out = 16'(-90);
			37747: out = 16'(-33);
			37748: out = 16'(-376);
			37749: out = 16'(-192);
			37750: out = 16'(337);
			37751: out = 16'(148);
			37752: out = 16'(-786);
			37753: out = 16'(-1439);
			37754: out = 16'(-596);
			37755: out = 16'(316);
			37756: out = 16'(512);
			37757: out = 16'(501);
			37758: out = 16'(674);
			37759: out = 16'(238);
			37760: out = 16'(-657);
			37761: out = 16'(-938);
			37762: out = 16'(-173);
			37763: out = 16'(562);
			37764: out = 16'(490);
			37765: out = 16'(-180);
			37766: out = 16'(-523);
			37767: out = 16'(-497);
			37768: out = 16'(-210);
			37769: out = 16'(-85);
			37770: out = 16'(523);
			37771: out = 16'(65);
			37772: out = 16'(-127);
			37773: out = 16'(-156);
			37774: out = 16'(-322);
			37775: out = 16'(-1100);
			37776: out = 16'(-705);
			37777: out = 16'(301);
			37778: out = 16'(58);
			37779: out = 16'(192);
			37780: out = 16'(-15);
			37781: out = 16'(-24);
			37782: out = 16'(65);
			37783: out = 16'(-686);
			37784: out = 16'(-406);
			37785: out = 16'(114);
			37786: out = 16'(82);
			37787: out = 16'(-7);
			37788: out = 16'(-100);
			37789: out = 16'(-34);
			37790: out = 16'(-66);
			37791: out = 16'(125);
			37792: out = 16'(113);
			37793: out = 16'(81);
			37794: out = 16'(-192);
			37795: out = 16'(-480);
			37796: out = 16'(-232);
			37797: out = 16'(442);
			37798: out = 16'(597);
			37799: out = 16'(-212);
			37800: out = 16'(-838);
			37801: out = 16'(-715);
			37802: out = 16'(94);
			37803: out = 16'(577);
			37804: out = 16'(1114);
			37805: out = 16'(460);
			37806: out = 16'(-35);
			37807: out = 16'(-6);
			37808: out = 16'(488);
			37809: out = 16'(254);
			37810: out = 16'(-191);
			37811: out = 16'(-759);
			37812: out = 16'(-1179);
			37813: out = 16'(-635);
			37814: out = 16'(527);
			37815: out = 16'(1055);
			37816: out = 16'(409);
			37817: out = 16'(-744);
			37818: out = 16'(-908);
			37819: out = 16'(-119);
			37820: out = 16'(573);
			37821: out = 16'(1050);
			37822: out = 16'(759);
			37823: out = 16'(256);
			37824: out = 16'(52);
			37825: out = 16'(-137);
			37826: out = 16'(69);
			37827: out = 16'(-193);
			37828: out = 16'(-609);
			37829: out = 16'(-361);
			37830: out = 16'(-126);
			37831: out = 16'(-232);
			37832: out = 16'(-195);
			37833: out = 16'(545);
			37834: out = 16'(518);
			37835: out = 16'(44);
			37836: out = 16'(-540);
			37837: out = 16'(-505);
			37838: out = 16'(-182);
			37839: out = 16'(-31);
			37840: out = 16'(-101);
			37841: out = 16'(178);
			37842: out = 16'(422);
			37843: out = 16'(307);
			37844: out = 16'(-560);
			37845: out = 16'(-1194);
			37846: out = 16'(-366);
			37847: out = 16'(-115);
			37848: out = 16'(-257);
			37849: out = 16'(-650);
			37850: out = 16'(-699);
			37851: out = 16'(-225);
			37852: out = 16'(439);
			37853: out = 16'(751);
			37854: out = 16'(451);
			37855: out = 16'(50);
			37856: out = 16'(-438);
			37857: out = 16'(-382);
			37858: out = 16'(150);
			37859: out = 16'(54);
			37860: out = 16'(-177);
			37861: out = 16'(-398);
			37862: out = 16'(-207);
			37863: out = 16'(51);
			37864: out = 16'(499);
			37865: out = 16'(279);
			37866: out = 16'(-131);
			37867: out = 16'(-17);
			37868: out = 16'(376);
			37869: out = 16'(639);
			37870: out = 16'(115);
			37871: out = 16'(-1035);
			37872: out = 16'(-808);
			37873: out = 16'(-345);
			37874: out = 16'(86);
			37875: out = 16'(96);
			37876: out = 16'(3);
			37877: out = 16'(-5);
			37878: out = 16'(145);
			37879: out = 16'(38);
			37880: out = 16'(162);
			37881: out = 16'(-119);
			37882: out = 16'(323);
			37883: out = 16'(638);
			37884: out = 16'(91);
			37885: out = 16'(-691);
			37886: out = 16'(-339);
			37887: out = 16'(90);
			37888: out = 16'(-604);
			37889: out = 16'(-577);
			37890: out = 16'(154);
			37891: out = 16'(905);
			37892: out = 16'(554);
			37893: out = 16'(59);
			37894: out = 16'(-448);
			37895: out = 16'(-641);
			37896: out = 16'(-712);
			37897: out = 16'(115);
			37898: out = 16'(554);
			37899: out = 16'(723);
			37900: out = 16'(317);
			37901: out = 16'(-274);
			37902: out = 16'(-761);
			37903: out = 16'(-457);
			37904: out = 16'(119);
			37905: out = 16'(503);
			37906: out = 16'(-140);
			37907: out = 16'(-760);
			37908: out = 16'(-928);
			37909: out = 16'(-430);
			37910: out = 16'(-149);
			37911: out = 16'(68);
			37912: out = 16'(-333);
			37913: out = 16'(-626);
			37914: out = 16'(-153);
			37915: out = 16'(987);
			37916: out = 16'(875);
			37917: out = 16'(-353);
			37918: out = 16'(-645);
			37919: out = 16'(-168);
			37920: out = 16'(493);
			37921: out = 16'(415);
			37922: out = 16'(-30);
			37923: out = 16'(-119);
			37924: out = 16'(-197);
			37925: out = 16'(-255);
			37926: out = 16'(260);
			37927: out = 16'(425);
			37928: out = 16'(652);
			37929: out = 16'(210);
			37930: out = 16'(-406);
			37931: out = 16'(-1199);
			37932: out = 16'(-110);
			37933: out = 16'(1029);
			37934: out = 16'(1076);
			37935: out = 16'(-28);
			37936: out = 16'(-443);
			37937: out = 16'(-759);
			37938: out = 16'(-1112);
			37939: out = 16'(-1405);
			37940: out = 16'(-358);
			37941: out = 16'(413);
			37942: out = 16'(447);
			37943: out = 16'(-30);
			37944: out = 16'(483);
			37945: out = 16'(279);
			37946: out = 16'(-341);
			37947: out = 16'(-688);
			37948: out = 16'(-130);
			37949: out = 16'(356);
			37950: out = 16'(681);
			37951: out = 16'(651);
			37952: out = 16'(163);
			37953: out = 16'(-223);
			37954: out = 16'(-384);
			37955: out = 16'(-317);
			37956: out = 16'(-347);
			37957: out = 16'(29);
			37958: out = 16'(107);
			37959: out = 16'(-260);
			37960: out = 16'(-740);
			37961: out = 16'(-451);
			37962: out = 16'(248);
			37963: out = 16'(520);
			37964: out = 16'(116);
			37965: out = 16'(718);
			37966: out = 16'(266);
			37967: out = 16'(-405);
			37968: out = 16'(-719);
			37969: out = 16'(-375);
			37970: out = 16'(56);
			37971: out = 16'(8);
			37972: out = 16'(-466);
			37973: out = 16'(-931);
			37974: out = 16'(-649);
			37975: out = 16'(-255);
			37976: out = 16'(241);
			37977: out = 16'(1163);
			37978: out = 16'(667);
			37979: out = 16'(185);
			37980: out = 16'(-71);
			37981: out = 16'(181);
			37982: out = 16'(-85);
			37983: out = 16'(-287);
			37984: out = 16'(-792);
			37985: out = 16'(-843);
			37986: out = 16'(-150);
			37987: out = 16'(478);
			37988: out = 16'(323);
			37989: out = 16'(-106);
			37990: out = 16'(164);
			37991: out = 16'(626);
			37992: out = 16'(417);
			37993: out = 16'(-144);
			37994: out = 16'(200);
			37995: out = 16'(-68);
			37996: out = 16'(-196);
			37997: out = 16'(-268);
			37998: out = 16'(247);
			37999: out = 16'(422);
			38000: out = 16'(329);
			38001: out = 16'(-859);
			38002: out = 16'(-2165);
			38003: out = 16'(-1043);
			38004: out = 16'(-179);
			38005: out = 16'(407);
			38006: out = 16'(543);
			38007: out = 16'(-12);
			38008: out = 16'(437);
			38009: out = 16'(612);
			38010: out = 16'(554);
			38011: out = 16'(534);
			38012: out = 16'(253);
			38013: out = 16'(-238);
			38014: out = 16'(-606);
			38015: out = 16'(-501);
			38016: out = 16'(-104);
			38017: out = 16'(-34);
			38018: out = 16'(-48);
			38019: out = 16'(-56);
			38020: out = 16'(2);
			38021: out = 16'(-689);
			38022: out = 16'(-888);
			38023: out = 16'(-347);
			38024: out = 16'(-60);
			38025: out = 16'(10);
			38026: out = 16'(220);
			38027: out = 16'(695);
			38028: out = 16'(477);
			38029: out = 16'(-146);
			38030: out = 16'(-1332);
			38031: out = 16'(-1815);
			38032: out = 16'(-958);
			38033: out = 16'(804);
			38034: out = 16'(1534);
			38035: out = 16'(853);
			38036: out = 16'(-78);
			38037: out = 16'(-897);
			38038: out = 16'(-500);
			38039: out = 16'(-228);
			38040: out = 16'(-212);
			38041: out = 16'(-17);
			38042: out = 16'(872);
			38043: out = 16'(1046);
			38044: out = 16'(286);
			38045: out = 16'(-445);
			38046: out = 16'(-378);
			38047: out = 16'(-216);
			38048: out = 16'(-265);
			38049: out = 16'(71);
			38050: out = 16'(-49);
			38051: out = 16'(70);
			38052: out = 16'(-101);
			38053: out = 16'(-197);
			38054: out = 16'(-96);
			38055: out = 16'(895);
			38056: out = 16'(1232);
			38057: out = 16'(313);
			38058: out = 16'(-353);
			38059: out = 16'(-960);
			38060: out = 16'(-542);
			38061: out = 16'(76);
			38062: out = 16'(172);
			38063: out = 16'(-465);
			38064: out = 16'(-782);
			38065: out = 16'(-599);
			38066: out = 16'(-492);
			38067: out = 16'(-773);
			38068: out = 16'(-522);
			38069: out = 16'(705);
			38070: out = 16'(1815);
			38071: out = 16'(1329);
			38072: out = 16'(218);
			38073: out = 16'(-524);
			38074: out = 16'(-665);
			38075: out = 16'(-27);
			38076: out = 16'(348);
			38077: out = 16'(998);
			38078: out = 16'(1073);
			38079: out = 16'(43);
			38080: out = 16'(-1183);
			38081: out = 16'(-1016);
			38082: out = 16'(-58);
			38083: out = 16'(150);
			38084: out = 16'(-177);
			38085: out = 16'(-76);
			38086: out = 16'(243);
			38087: out = 16'(103);
			38088: out = 16'(-243);
			38089: out = 16'(221);
			38090: out = 16'(665);
			38091: out = 16'(479);
			38092: out = 16'(178);
			38093: out = 16'(84);
			38094: out = 16'(-12);
			38095: out = 16'(-506);
			38096: out = 16'(-1608);
			38097: out = 16'(-700);
			38098: out = 16'(2);
			38099: out = 16'(-73);
			38100: out = 16'(-226);
			38101: out = 16'(56);
			38102: out = 16'(1);
			38103: out = 16'(-278);
			38104: out = 16'(138);
			38105: out = 16'(1060);
			38106: out = 16'(1498);
			38107: out = 16'(828);
			38108: out = 16'(-154);
			38109: out = 16'(-885);
			38110: out = 16'(-1138);
			38111: out = 16'(-1080);
			38112: out = 16'(-440);
			38113: out = 16'(650);
			38114: out = 16'(819);
			38115: out = 16'(-128);
			38116: out = 16'(-972);
			38117: out = 16'(-445);
			38118: out = 16'(504);
			38119: out = 16'(812);
			38120: out = 16'(365);
			38121: out = 16'(-4);
			38122: out = 16'(119);
			38123: out = 16'(-19);
			38124: out = 16'(-508);
			38125: out = 16'(-632);
			38126: out = 16'(-1);
			38127: out = 16'(611);
			38128: out = 16'(738);
			38129: out = 16'(417);
			38130: out = 16'(-643);
			38131: out = 16'(-935);
			38132: out = 16'(-812);
			38133: out = 16'(-276);
			38134: out = 16'(562);
			38135: out = 16'(1175);
			38136: out = 16'(1121);
			38137: out = 16'(419);
			38138: out = 16'(-295);
			38139: out = 16'(-562);
			38140: out = 16'(-264);
			38141: out = 16'(-29);
			38142: out = 16'(-49);
			38143: out = 16'(-67);
			38144: out = 16'(-36);
			38145: out = 16'(-156);
			38146: out = 16'(-312);
			38147: out = 16'(-542);
			38148: out = 16'(-157);
			38149: out = 16'(-116);
			38150: out = 16'(-260);
			38151: out = 16'(-34);
			38152: out = 16'(987);
			38153: out = 16'(1098);
			38154: out = 16'(238);
			38155: out = 16'(-261);
			38156: out = 16'(-176);
			38157: out = 16'(-192);
			38158: out = 16'(-933);
			38159: out = 16'(-1588);
			38160: out = 16'(-1134);
			38161: out = 16'(53);
			38162: out = 16'(724);
			38163: out = 16'(562);
			38164: out = 16'(772);
			38165: out = 16'(640);
			38166: out = 16'(323);
			38167: out = 16'(-132);
			38168: out = 16'(-279);
			38169: out = 16'(-359);
			38170: out = 16'(-172);
			38171: out = 16'(78);
			38172: out = 16'(548);
			38173: out = 16'(72);
			38174: out = 16'(-108);
			38175: out = 16'(-76);
			38176: out = 16'(-57);
			38177: out = 16'(97);
			38178: out = 16'(-346);
			38179: out = 16'(-942);
			38180: out = 16'(-830);
			38181: out = 16'(-191);
			38182: out = 16'(474);
			38183: out = 16'(422);
			38184: out = 16'(166);
			38185: out = 16'(115);
			38186: out = 16'(246);
			38187: out = 16'(-384);
			38188: out = 16'(-850);
			38189: out = 16'(142);
			38190: out = 16'(931);
			38191: out = 16'(664);
			38192: out = 16'(-444);
			38193: out = 16'(-882);
			38194: out = 16'(-862);
			38195: out = 16'(-645);
			38196: out = 16'(-740);
			38197: out = 16'(-344);
			38198: out = 16'(-162);
			38199: out = 16'(831);
			38200: out = 16'(1040);
			38201: out = 16'(453);
			38202: out = 16'(-14);
			38203: out = 16'(-59);
			38204: out = 16'(-195);
			38205: out = 16'(-236);
			38206: out = 16'(116);
			38207: out = 16'(59);
			38208: out = 16'(-291);
			38209: out = 16'(-517);
			38210: out = 16'(-506);
			38211: out = 16'(-89);
			38212: out = 16'(-71);
			38213: out = 16'(353);
			38214: out = 16'(1057);
			38215: out = 16'(204);
			38216: out = 16'(-1016);
			38217: out = 16'(-1024);
			38218: out = 16'(466);
			38219: out = 16'(1009);
			38220: out = 16'(450);
			38221: out = 16'(-464);
			38222: out = 16'(-734);
			38223: out = 16'(-990);
			38224: out = 16'(-931);
			38225: out = 16'(-553);
			38226: out = 16'(329);
			38227: out = 16'(734);
			38228: out = 16'(1178);
			38229: out = 16'(547);
			38230: out = 16'(-369);
			38231: out = 16'(-1031);
			38232: out = 16'(-846);
			38233: out = 16'(-572);
			38234: out = 16'(-172);
			38235: out = 16'(299);
			38236: out = 16'(1067);
			38237: out = 16'(472);
			38238: out = 16'(-550);
			38239: out = 16'(-870);
			38240: out = 16'(-29);
			38241: out = 16'(424);
			38242: out = 16'(345);
			38243: out = 16'(-216);
			38244: out = 16'(-739);
			38245: out = 16'(-184);
			38246: out = 16'(354);
			38247: out = 16'(456);
			38248: out = 16'(151);
			38249: out = 16'(0);
			38250: out = 16'(252);
			38251: out = 16'(581);
			38252: out = 16'(373);
			38253: out = 16'(-137);
			38254: out = 16'(-582);
			38255: out = 16'(-485);
			38256: out = 16'(-146);
			38257: out = 16'(495);
			38258: out = 16'(126);
			38259: out = 16'(-152);
			38260: out = 16'(-210);
			38261: out = 16'(215);
			38262: out = 16'(324);
			38263: out = 16'(1097);
			38264: out = 16'(1357);
			38265: out = 16'(488);
			38266: out = 16'(-813);
			38267: out = 16'(-948);
			38268: out = 16'(-469);
			38269: out = 16'(-273);
			38270: out = 16'(-66);
			38271: out = 16'(301);
			38272: out = 16'(278);
			38273: out = 16'(-414);
			38274: out = 16'(-566);
			38275: out = 16'(-282);
			38276: out = 16'(266);
			38277: out = 16'(471);
			38278: out = 16'(470);
			38279: out = 16'(64);
			38280: out = 16'(-426);
			38281: out = 16'(-1003);
			38282: out = 16'(-1129);
			38283: out = 16'(-299);
			38284: out = 16'(659);
			38285: out = 16'(917);
			38286: out = 16'(533);
			38287: out = 16'(-492);
			38288: out = 16'(-805);
			38289: out = 16'(-817);
			38290: out = 16'(-777);
			38291: out = 16'(-801);
			38292: out = 16'(108);
			38293: out = 16'(730);
			38294: out = 16'(493);
			38295: out = 16'(-157);
			38296: out = 16'(-301);
			38297: out = 16'(-61);
			38298: out = 16'(-4);
			38299: out = 16'(0);
			38300: out = 16'(-30);
			38301: out = 16'(36);
			38302: out = 16'(-44);
			38303: out = 16'(55);
			38304: out = 16'(-94);
			38305: out = 16'(375);
			38306: out = 16'(241);
			38307: out = 16'(-490);
			38308: out = 16'(-413);
			38309: out = 16'(-140);
			38310: out = 16'(30);
			38311: out = 16'(6);
			38312: out = 16'(121);
			38313: out = 16'(875);
			38314: out = 16'(963);
			38315: out = 16'(8);
			38316: out = 16'(-1336);
			38317: out = 16'(-557);
			38318: out = 16'(127);
			38319: out = 16'(-22);
			38320: out = 16'(-121);
			38321: out = 16'(324);
			38322: out = 16'(988);
			38323: out = 16'(773);
			38324: out = 16'(-135);
			38325: out = 16'(-396);
			38326: out = 16'(118);
			38327: out = 16'(595);
			38328: out = 16'(318);
			38329: out = 16'(44);
			38330: out = 16'(-46);
			38331: out = 16'(611);
			38332: out = 16'(939);
			38333: out = 16'(35);
			38334: out = 16'(-249);
			38335: out = 16'(-196);
			38336: out = 16'(-162);
			38337: out = 16'(-725);
			38338: out = 16'(-785);
			38339: out = 16'(-580);
			38340: out = 16'(36);
			38341: out = 16'(483);
			38342: out = 16'(919);
			38343: out = 16'(426);
			38344: out = 16'(-170);
			38345: out = 16'(-392);
			38346: out = 16'(393);
			38347: out = 16'(99);
			38348: out = 16'(-219);
			38349: out = 16'(-259);
			38350: out = 16'(-106);
			38351: out = 16'(-112);
			38352: out = 16'(193);
			38353: out = 16'(387);
			38354: out = 16'(-134);
			38355: out = 16'(-539);
			38356: out = 16'(-629);
			38357: out = 16'(-339);
			38358: out = 16'(-296);
			38359: out = 16'(77);
			38360: out = 16'(-6);
			38361: out = 16'(-44);
			38362: out = 16'(-30);
			38363: out = 16'(459);
			38364: out = 16'(430);
			38365: out = 16'(372);
			38366: out = 16'(-148);
			38367: out = 16'(-910);
			38368: out = 16'(-1636);
			38369: out = 16'(-597);
			38370: out = 16'(946);
			38371: out = 16'(967);
			38372: out = 16'(87);
			38373: out = 16'(-430);
			38374: out = 16'(-104);
			38375: out = 16'(-113);
			38376: out = 16'(13);
			38377: out = 16'(-205);
			38378: out = 16'(-251);
			38379: out = 16'(-255);
			38380: out = 16'(142);
			38381: out = 16'(10);
			38382: out = 16'(0);
			38383: out = 16'(177);
			38384: out = 16'(448);
			38385: out = 16'(-19);
			38386: out = 16'(-507);
			38387: out = 16'(-470);
			38388: out = 16'(465);
			38389: out = 16'(225);
			38390: out = 16'(-1);
			38391: out = 16'(50);
			38392: out = 16'(476);
			38393: out = 16'(1);
			38394: out = 16'(-75);
			38395: out = 16'(-118);
			38396: out = 16'(-265);
			38397: out = 16'(-123);
			38398: out = 16'(80);
			38399: out = 16'(57);
			38400: out = 16'(-99);
			38401: out = 16'(-245);
			38402: out = 16'(-133);
			38403: out = 16'(28);
			38404: out = 16'(72);
			38405: out = 16'(-104);
			38406: out = 16'(-33);
			38407: out = 16'(-196);
			38408: out = 16'(-222);
			38409: out = 16'(-81);
			38410: out = 16'(520);
			38411: out = 16'(500);
			38412: out = 16'(587);
			38413: out = 16'(966);
			38414: out = 16'(91);
			38415: out = 16'(-1161);
			38416: out = 16'(-1418);
			38417: out = 16'(-42);
			38418: out = 16'(431);
			38419: out = 16'(617);
			38420: out = 16'(57);
			38421: out = 16'(-341);
			38422: out = 16'(-526);
			38423: out = 16'(-325);
			38424: out = 16'(-330);
			38425: out = 16'(-207);
			38426: out = 16'(-64);
			38427: out = 16'(493);
			38428: out = 16'(398);
			38429: out = 16'(-334);
			38430: out = 16'(-1241);
			38431: out = 16'(-253);
			38432: out = 16'(0);
			38433: out = 16'(-70);
			38434: out = 16'(-8);
			38435: out = 16'(413);
			38436: out = 16'(245);
			38437: out = 16'(-166);
			38438: out = 16'(-510);
			38439: out = 16'(-428);
			38440: out = 16'(-146);
			38441: out = 16'(623);
			38442: out = 16'(973);
			38443: out = 16'(57);
			38444: out = 16'(-368);
			38445: out = 16'(-509);
			38446: out = 16'(-512);
			38447: out = 16'(-615);
			38448: out = 16'(-169);
			38449: out = 16'(596);
			38450: out = 16'(778);
			38451: out = 16'(-110);
			38452: out = 16'(-699);
			38453: out = 16'(-460);
			38454: out = 16'(313);
			38455: out = 16'(286);
			38456: out = 16'(-136);
			38457: out = 16'(-822);
			38458: out = 16'(-247);
			38459: out = 16'(566);
			38460: out = 16'(437);
			38461: out = 16'(-111);
			38462: out = 16'(-155);
			38463: out = 16'(271);
			38464: out = 16'(404);
			38465: out = 16'(-158);
			38466: out = 16'(-532);
			38467: out = 16'(-730);
			38468: out = 16'(-764);
			38469: out = 16'(-133);
			38470: out = 16'(455);
			38471: out = 16'(467);
			38472: out = 16'(-143);
			38473: out = 16'(0);
			38474: out = 16'(-342);
			38475: out = 16'(-567);
			38476: out = 16'(-518);
			38477: out = 16'(-25);
			38478: out = 16'(381);
			38479: out = 16'(284);
			38480: out = 16'(-128);
			38481: out = 16'(25);
			38482: out = 16'(43);
			38483: out = 16'(123);
			38484: out = 16'(-282);
			38485: out = 16'(-588);
			38486: out = 16'(-884);
			38487: out = 16'(43);
			38488: out = 16'(613);
			38489: out = 16'(425);
			38490: out = 16'(123);
			38491: out = 16'(152);
			38492: out = 16'(-211);
			38493: out = 16'(-1002);
			38494: out = 16'(-1326);
			38495: out = 16'(-568);
			38496: out = 16'(285);
			38497: out = 16'(515);
			38498: out = 16'(541);
			38499: out = 16'(610);
			38500: out = 16'(714);
			38501: out = 16'(404);
			38502: out = 16'(-348);
			38503: out = 16'(-897);
			38504: out = 16'(-509);
			38505: out = 16'(533);
			38506: out = 16'(1022);
			38507: out = 16'(275);
			38508: out = 16'(-600);
			38509: out = 16'(-551);
			38510: out = 16'(104);
			38511: out = 16'(123);
			38512: out = 16'(41);
			38513: out = 16'(-34);
			38514: out = 16'(-61);
			38515: out = 16'(-425);
			38516: out = 16'(-102);
			38517: out = 16'(299);
			38518: out = 16'(446);
			38519: out = 16'(74);
			38520: out = 16'(23);
			38521: out = 16'(-156);
			38522: out = 16'(-488);
			38523: out = 16'(-984);
			38524: out = 16'(-257);
			38525: out = 16'(242);
			38526: out = 16'(766);
			38527: out = 16'(886);
			38528: out = 16'(518);
			38529: out = 16'(77);
			38530: out = 16'(-219);
			38531: out = 16'(-601);
			38532: out = 16'(-962);
			38533: out = 16'(-629);
			38534: out = 16'(152);
			38535: out = 16'(421);
			38536: out = 16'(-43);
			38537: out = 16'(-376);
			38538: out = 16'(-111);
			38539: out = 16'(88);
			38540: out = 16'(-267);
			38541: out = 16'(10);
			38542: out = 16'(81);
			38543: out = 16'(24);
			38544: out = 16'(-273);
			38545: out = 16'(-186);
			38546: out = 16'(-94);
			38547: out = 16'(76);
			38548: out = 16'(223);
			38549: out = 16'(657);
			38550: out = 16'(150);
			38551: out = 16'(-400);
			38552: out = 16'(-921);
			38553: out = 16'(-892);
			38554: out = 16'(-201);
			38555: out = 16'(405);
			38556: out = 16'(409);
			38557: out = 16'(-49);
			38558: out = 16'(-518);
			38559: out = 16'(-386);
			38560: out = 16'(-5);
			38561: out = 16'(225);
			38562: out = 16'(497);
			38563: out = 16'(640);
			38564: out = 16'(499);
			38565: out = 16'(66);
			38566: out = 16'(173);
			38567: out = 16'(-490);
			38568: out = 16'(-381);
			38569: out = 16'(274);
			38570: out = 16'(1102);
			38571: out = 16'(737);
			38572: out = 16'(261);
			38573: out = 16'(-227);
			38574: out = 16'(-453);
			38575: out = 16'(-1187);
			38576: out = 16'(-439);
			38577: out = 16'(466);
			38578: out = 16'(588);
			38579: out = 16'(666);
			38580: out = 16'(166);
			38581: out = 16'(-263);
			38582: out = 16'(-419);
			38583: out = 16'(-64);
			38584: out = 16'(449);
			38585: out = 16'(480);
			38586: out = 16'(-176);
			38587: out = 16'(-572);
			38588: out = 16'(-432);
			38589: out = 16'(252);
			38590: out = 16'(653);
			38591: out = 16'(575);
			38592: out = 16'(9);
			38593: out = 16'(-113);
			38594: out = 16'(-40);
			38595: out = 16'(59);
			38596: out = 16'(-811);
			38597: out = 16'(-378);
			38598: out = 16'(213);
			38599: out = 16'(414);
			38600: out = 16'(85);
			38601: out = 16'(143);
			38602: out = 16'(-212);
			38603: out = 16'(-798);
			38604: out = 16'(-1014);
			38605: out = 16'(-577);
			38606: out = 16'(-222);
			38607: out = 16'(129);
			38608: out = 16'(397);
			38609: out = 16'(-340);
			38610: out = 16'(-1452);
			38611: out = 16'(-1377);
			38612: out = 16'(202);
			38613: out = 16'(1008);
			38614: out = 16'(525);
			38615: out = 16'(-326);
			38616: out = 16'(-290);
			38617: out = 16'(25);
			38618: out = 16'(107);
			38619: out = 16'(-95);
			38620: out = 16'(88);
			38621: out = 16'(46);
			38622: out = 16'(192);
			38623: out = 16'(-198);
			38624: out = 16'(-398);
			38625: out = 16'(-215);
			38626: out = 16'(400);
			38627: out = 16'(344);
			38628: out = 16'(96);
			38629: out = 16'(151);
			38630: out = 16'(-212);
			38631: out = 16'(-281);
			38632: out = 16'(-168);
			38633: out = 16'(8);
			38634: out = 16'(141);
			38635: out = 16'(27);
			38636: out = 16'(-52);
			38637: out = 16'(-19);
			38638: out = 16'(-15);
			38639: out = 16'(79);
			38640: out = 16'(314);
			38641: out = 16'(439);
			38642: out = 16'(119);
			38643: out = 16'(118);
			38644: out = 16'(312);
			38645: out = 16'(376);
			38646: out = 16'(-125);
			38647: out = 16'(-207);
			38648: out = 16'(-200);
			38649: out = 16'(221);
			38650: out = 16'(548);
			38651: out = 16'(26);
			38652: out = 16'(-628);
			38653: out = 16'(-700);
			38654: out = 16'(-71);
			38655: out = 16'(566);
			38656: out = 16'(680);
			38657: out = 16'(295);
			38658: out = 16'(-227);
			38659: out = 16'(-442);
			38660: out = 16'(-680);
			38661: out = 16'(-107);
			38662: out = 16'(714);
			38663: out = 16'(797);
			38664: out = 16'(282);
			38665: out = 16'(-541);
			38666: out = 16'(-920);
			38667: out = 16'(-772);
			38668: out = 16'(-125);
			38669: out = 16'(-36);
			38670: out = 16'(-92);
			38671: out = 16'(56);
			38672: out = 16'(579);
			38673: out = 16'(175);
			38674: out = 16'(-393);
			38675: out = 16'(-544);
			38676: out = 16'(140);
			38677: out = 16'(370);
			38678: out = 16'(348);
			38679: out = 16'(-75);
			38680: out = 16'(-248);
			38681: out = 16'(-846);
			38682: out = 16'(-407);
			38683: out = 16'(0);
			38684: out = 16'(105);
			38685: out = 16'(-83);
			38686: out = 16'(354);
			38687: out = 16'(-4);
			38688: out = 16'(-1158);
			38689: out = 16'(-772);
			38690: out = 16'(79);
			38691: out = 16'(529);
			38692: out = 16'(-162);
			38693: out = 16'(-489);
			38694: out = 16'(-603);
			38695: out = 16'(130);
			38696: out = 16'(517);
			38697: out = 16'(494);
			38698: out = 16'(-321);
			38699: out = 16'(-234);
			38700: out = 16'(21);
			38701: out = 16'(-84);
			38702: out = 16'(-1079);
			38703: out = 16'(-690);
			38704: out = 16'(228);
			38705: out = 16'(639);
			38706: out = 16'(17);
			38707: out = 16'(353);
			38708: out = 16'(433);
			38709: out = 16'(-175);
			38710: out = 16'(-1315);
			38711: out = 16'(-998);
			38712: out = 16'(-337);
			38713: out = 16'(194);
			38714: out = 16'(496);
			38715: out = 16'(165);
			38716: out = 16'(-296);
			38717: out = 16'(-111);
			38718: out = 16'(740);
			38719: out = 16'(961);
			38720: out = 16'(403);
			38721: out = 16'(-200);
			38722: out = 16'(-269);
			38723: out = 16'(-1005);
			38724: out = 16'(-509);
			38725: out = 16'(209);
			38726: out = 16'(706);
			38727: out = 16'(486);
			38728: out = 16'(469);
			38729: out = 16'(579);
			38730: out = 16'(421);
			38731: out = 16'(-677);
			38732: out = 16'(-482);
			38733: out = 16'(-185);
			38734: out = 16'(276);
			38735: out = 16'(438);
			38736: out = 16'(670);
			38737: out = 16'(73);
			38738: out = 16'(-369);
			38739: out = 16'(-254);
			38740: out = 16'(-466);
			38741: out = 16'(-334);
			38742: out = 16'(-149);
			38743: out = 16'(-7);
			38744: out = 16'(-46);
			38745: out = 16'(84);
			38746: out = 16'(133);
			38747: out = 16'(155);
			38748: out = 16'(140);
			38749: out = 16'(396);
			38750: out = 16'(365);
			38751: out = 16'(-153);
			38752: out = 16'(-778);
			38753: out = 16'(-221);
			38754: out = 16'(365);
			38755: out = 16'(269);
			38756: out = 16'(-293);
			38757: out = 16'(-299);
			38758: out = 16'(-57);
			38759: out = 16'(-300);
			38760: out = 16'(-825);
			38761: out = 16'(-443);
			38762: out = 16'(384);
			38763: out = 16'(490);
			38764: out = 16'(-200);
			38765: out = 16'(-130);
			38766: out = 16'(-153);
			38767: out = 16'(141);
			38768: out = 16'(59);
			38769: out = 16'(21);
			38770: out = 16'(-433);
			38771: out = 16'(-64);
			38772: out = 16'(79);
			38773: out = 16'(-296);
			38774: out = 16'(-576);
			38775: out = 16'(-239);
			38776: out = 16'(86);
			38777: out = 16'(-5);
			38778: out = 16'(174);
			38779: out = 16'(186);
			38780: out = 16'(106);
			38781: out = 16'(58);
			38782: out = 16'(487);
			38783: out = 16'(125);
			38784: out = 16'(-243);
			38785: out = 16'(-334);
			38786: out = 16'(122);
			38787: out = 16'(-456);
			38788: out = 16'(-779);
			38789: out = 16'(-397);
			38790: out = 16'(802);
			38791: out = 16'(884);
			38792: out = 16'(493);
			38793: out = 16'(-739);
			38794: out = 16'(-1487);
			38795: out = 16'(-918);
			38796: out = 16'(658);
			38797: out = 16'(1106);
			38798: out = 16'(472);
			38799: out = 16'(-189);
			38800: out = 16'(320);
			38801: out = 16'(352);
			38802: out = 16'(-98);
			38803: out = 16'(196);
			38804: out = 16'(-327);
			38805: out = 16'(-655);
			38806: out = 16'(-637);
			38807: out = 16'(80);
			38808: out = 16'(105);
			38809: out = 16'(131);
			38810: out = 16'(-120);
			38811: out = 16'(-173);
			38812: out = 16'(-58);
			38813: out = 16'(363);
			38814: out = 16'(540);
			38815: out = 16'(421);
			38816: out = 16'(1);
			38817: out = 16'(-454);
			38818: out = 16'(-438);
			38819: out = 16'(214);
			38820: out = 16'(376);
			38821: out = 16'(357);
			38822: out = 16'(-756);
			38823: out = 16'(-1164);
			38824: out = 16'(96);
			38825: out = 16'(574);
			38826: out = 16'(333);
			38827: out = 16'(-62);
			38828: out = 16'(195);
			38829: out = 16'(-11);
			38830: out = 16'(-346);
			38831: out = 16'(-676);
			38832: out = 16'(-478);
			38833: out = 16'(-47);
			38834: out = 16'(172);
			38835: out = 16'(115);
			38836: out = 16'(-42);
			38837: out = 16'(-190);
			38838: out = 16'(-129);
			38839: out = 16'(277);
			38840: out = 16'(446);
			38841: out = 16'(-23);
			38842: out = 16'(-28);
			38843: out = 16'(277);
			38844: out = 16'(440);
			38845: out = 16'(-118);
			38846: out = 16'(-147);
			38847: out = 16'(-414);
			38848: out = 16'(-289);
			38849: out = 16'(-54);
			38850: out = 16'(-201);
			38851: out = 16'(-117);
			38852: out = 16'(241);
			38853: out = 16'(451);
			38854: out = 16'(0);
			38855: out = 16'(-191);
			38856: out = 16'(-141);
			38857: out = 16'(5);
			38858: out = 16'(-20);
			38859: out = 16'(3);
			38860: out = 16'(-54);
			38861: out = 16'(120);
			38862: out = 16'(687);
			38863: out = 16'(445);
			38864: out = 16'(522);
			38865: out = 16'(149);
			38866: out = 16'(-554);
			38867: out = 16'(-990);
			38868: out = 16'(-783);
			38869: out = 16'(-578);
			38870: out = 16'(-548);
			38871: out = 16'(-7);
			38872: out = 16'(376);
			38873: out = 16'(536);
			38874: out = 16'(468);
			38875: out = 16'(482);
			38876: out = 16'(482);
			38877: out = 16'(130);
			38878: out = 16'(-499);
			38879: out = 16'(-760);
			38880: out = 16'(-220);
			38881: out = 16'(449);
			38882: out = 16'(527);
			38883: out = 16'(83);
			38884: out = 16'(-35);
			38885: out = 16'(-43);
			38886: out = 16'(-160);
			38887: out = 16'(-545);
			38888: out = 16'(-757);
			38889: out = 16'(-635);
			38890: out = 16'(50);
			38891: out = 16'(554);
			38892: out = 16'(644);
			38893: out = 16'(205);
			38894: out = 16'(-84);
			38895: out = 16'(-481);
			38896: out = 16'(-997);
			38897: out = 16'(-1073);
			38898: out = 16'(-157);
			38899: out = 16'(806);
			38900: out = 16'(762);
			38901: out = 16'(-221);
			38902: out = 16'(-255);
			38903: out = 16'(215);
			38904: out = 16'(320);
			38905: out = 16'(129);
			38906: out = 16'(-302);
			38907: out = 16'(-193);
			38908: out = 16'(153);
			38909: out = 16'(-75);
			38910: out = 16'(106);
			38911: out = 16'(-72);
			38912: out = 16'(-116);
			38913: out = 16'(413);
			38914: out = 16'(484);
			38915: out = 16'(167);
			38916: out = 16'(-572);
			38917: out = 16'(-998);
			38918: out = 16'(-1046);
			38919: out = 16'(-381);
			38920: out = 16'(224);
			38921: out = 16'(407);
			38922: out = 16'(407);
			38923: out = 16'(126);
			38924: out = 16'(-151);
			38925: out = 16'(-132);
			38926: out = 16'(91);
			38927: out = 16'(461);
			38928: out = 16'(220);
			38929: out = 16'(-386);
			38930: out = 16'(-461);
			38931: out = 16'(-142);
			38932: out = 16'(30);
			38933: out = 16'(-209);
			38934: out = 16'(-289);
			38935: out = 16'(-121);
			38936: out = 16'(536);
			38937: out = 16'(709);
			38938: out = 16'(259);
			38939: out = 16'(-308);
			38940: out = 16'(-410);
			38941: out = 16'(-297);
			38942: out = 16'(-237);
			38943: out = 16'(-508);
			38944: out = 16'(-143);
			38945: out = 16'(79);
			38946: out = 16'(38);
			38947: out = 16'(-205);
			38948: out = 16'(-16);
			38949: out = 16'(-121);
			38950: out = 16'(-131);
			38951: out = 16'(133);
			38952: out = 16'(738);
			38953: out = 16'(352);
			38954: out = 16'(-289);
			38955: out = 16'(-407);
			38956: out = 16'(442);
			38957: out = 16'(214);
			38958: out = 16'(-242);
			38959: out = 16'(-306);
			38960: out = 16'(-102);
			38961: out = 16'(-120);
			38962: out = 16'(-358);
			38963: out = 16'(-493);
			38964: out = 16'(-311);
			38965: out = 16'(-82);
			38966: out = 16'(243);
			38967: out = 16'(459);
			38968: out = 16'(379);
			38969: out = 16'(38);
			38970: out = 16'(-43);
			38971: out = 16'(0);
			38972: out = 16'(-27);
			38973: out = 16'(-207);
			38974: out = 16'(-11);
			38975: out = 16'(107);
			38976: out = 16'(-63);
			38977: out = 16'(7);
			38978: out = 16'(-266);
			38979: out = 16'(-365);
			38980: out = 16'(-285);
			38981: out = 16'(5);
			38982: out = 16'(-16);
			38983: out = 16'(69);
			38984: out = 16'(76);
			38985: out = 16'(0);
			38986: out = 16'(-38);
			38987: out = 16'(285);
			38988: out = 16'(686);
			38989: out = 16'(882);
			38990: out = 16'(773);
			38991: out = 16'(257);
			38992: out = 16'(-473);
			38993: out = 16'(-793);
			38994: out = 16'(-301);
			38995: out = 16'(31);
			38996: out = 16'(-13);
			38997: out = 16'(178);
			38998: out = 16'(1171);
			38999: out = 16'(1033);
			39000: out = 16'(-11);
			39001: out = 16'(-1048);
			39002: out = 16'(-778);
			39003: out = 16'(-138);
			39004: out = 16'(109);
			39005: out = 16'(-119);
			39006: out = 16'(123);
			39007: out = 16'(-423);
			39008: out = 16'(-154);
			39009: out = 16'(-245);
			39010: out = 16'(-500);
			39011: out = 16'(-408);
			39012: out = 16'(251);
			39013: out = 16'(575);
			39014: out = 16'(433);
			39015: out = 16'(92);
			39016: out = 16'(301);
			39017: out = 16'(182);
			39018: out = 16'(-161);
			39019: out = 16'(-385);
			39020: out = 16'(-120);
			39021: out = 16'(-190);
			39022: out = 16'(-494);
			39023: out = 16'(-691);
			39024: out = 16'(-682);
			39025: out = 16'(-374);
			39026: out = 16'(406);
			39027: out = 16'(1063);
			39028: out = 16'(240);
			39029: out = 16'(-1013);
			39030: out = 16'(-1404);
			39031: out = 16'(-312);
			39032: out = 16'(384);
			39033: out = 16'(870);
			39034: out = 16'(426);
			39035: out = 16'(57);
			39036: out = 16'(-75);
			39037: out = 16'(25);
			39038: out = 16'(-302);
			39039: out = 16'(-473);
			39040: out = 16'(-186);
			39041: out = 16'(0);
			39042: out = 16'(-256);
			39043: out = 16'(-133);
			39044: out = 16'(417);
			39045: out = 16'(175);
			39046: out = 16'(-234);
			39047: out = 16'(-93);
			39048: out = 16'(609);
			39049: out = 16'(474);
			39050: out = 16'(421);
			39051: out = 16'(343);
			39052: out = 16'(293);
			39053: out = 16'(-74);
			39054: out = 16'(-2);
			39055: out = 16'(220);
			39056: out = 16'(269);
			39057: out = 16'(-109);
			39058: out = 16'(-497);
			39059: out = 16'(-316);
			39060: out = 16'(-1);
			39061: out = 16'(-79);
			39062: out = 16'(46);
			39063: out = 16'(269);
			39064: out = 16'(192);
			39065: out = 16'(-352);
			39066: out = 16'(-509);
			39067: out = 16'(-492);
			39068: out = 16'(-222);
			39069: out = 16'(-19);
			39070: out = 16'(380);
			39071: out = 16'(35);
			39072: out = 16'(-96);
			39073: out = 16'(-35);
			39074: out = 16'(-72);
			39075: out = 16'(-58);
			39076: out = 16'(-277);
			39077: out = 16'(-314);
			39078: out = 16'(0);
			39079: out = 16'(429);
			39080: out = 16'(293);
			39081: out = 16'(-40);
			39082: out = 16'(-32);
			39083: out = 16'(-252);
			39084: out = 16'(-231);
			39085: out = 16'(-259);
			39086: out = 16'(-205);
			39087: out = 16'(-244);
			39088: out = 16'(240);
			39089: out = 16'(287);
			39090: out = 16'(38);
			39091: out = 16'(80);
			39092: out = 16'(-51);
			39093: out = 16'(-62);
			39094: out = 16'(-18);
			39095: out = 16'(90);
			39096: out = 16'(80);
			39097: out = 16'(5);
			39098: out = 16'(-88);
			39099: out = 16'(-30);
			39100: out = 16'(29);
			39101: out = 16'(123);
			39102: out = 16'(-312);
			39103: out = 16'(-864);
			39104: out = 16'(-227);
			39105: out = 16'(-236);
			39106: out = 16'(-142);
			39107: out = 16'(75);
			39108: out = 16'(509);
			39109: out = 16'(537);
			39110: out = 16'(195);
			39111: out = 16'(-40);
			39112: out = 16'(402);
			39113: out = 16'(-37);
			39114: out = 16'(-61);
			39115: out = 16'(-105);
			39116: out = 16'(-79);
			39117: out = 16'(-828);
			39118: out = 16'(-578);
			39119: out = 16'(-286);
			39120: out = 16'(-182);
			39121: out = 16'(-60);
			39122: out = 16'(310);
			39123: out = 16'(146);
			39124: out = 16'(-260);
			39125: out = 16'(-3);
			39126: out = 16'(279);
			39127: out = 16'(217);
			39128: out = 16'(-207);
			39129: out = 16'(-175);
			39130: out = 16'(-28);
			39131: out = 16'(287);
			39132: out = 16'(389);
			39133: out = 16'(479);
			39134: out = 16'(95);
			39135: out = 16'(-200);
			39136: out = 16'(-636);
			39137: out = 16'(-779);
			39138: out = 16'(-128);
			39139: out = 16'(128);
			39140: out = 16'(-179);
			39141: out = 16'(-540);
			39142: out = 16'(-358);
			39143: out = 16'(302);
			39144: out = 16'(707);
			39145: out = 16'(672);
			39146: out = 16'(321);
			39147: out = 16'(-107);
			39148: out = 16'(-559);
			39149: out = 16'(-543);
			39150: out = 16'(115);
			39151: out = 16'(334);
			39152: out = 16'(202);
			39153: out = 16'(-22);
			39154: out = 16'(-61);
			39155: out = 16'(-70);
			39156: out = 16'(-180);
			39157: out = 16'(-202);
			39158: out = 16'(-7);
			39159: out = 16'(31);
			39160: out = 16'(-46);
			39161: out = 16'(-49);
			39162: out = 16'(176);
			39163: out = 16'(313);
			39164: out = 16'(65);
			39165: out = 16'(-455);
			39166: out = 16'(-705);
			39167: out = 16'(-481);
			39168: out = 16'(255);
			39169: out = 16'(285);
			39170: out = 16'(-77);
			39171: out = 16'(-202);
			39172: out = 16'(-82);
			39173: out = 16'(-24);
			39174: out = 16'(-75);
			39175: out = 16'(-29);
			39176: out = 16'(-71);
			39177: out = 16'(64);
			39178: out = 16'(-7);
			39179: out = 16'(28);
			39180: out = 16'(344);
			39181: out = 16'(194);
			39182: out = 16'(-227);
			39183: out = 16'(-275);
			39184: out = 16'(84);
			39185: out = 16'(367);
			39186: out = 16'(-83);
			39187: out = 16'(-364);
			39188: out = 16'(13);
			39189: out = 16'(440);
			39190: out = 16'(148);
			39191: out = 16'(-97);
			39192: out = 16'(1);
			39193: out = 16'(-709);
			39194: out = 16'(-720);
			39195: out = 16'(-455);
			39196: out = 16'(120);
			39197: out = 16'(324);
			39198: out = 16'(518);
			39199: out = 16'(222);
			39200: out = 16'(-190);
			39201: out = 16'(-392);
			39202: out = 16'(-672);
			39203: out = 16'(-606);
			39204: out = 16'(-464);
			39205: out = 16'(-290);
			39206: out = 16'(437);
			39207: out = 16'(814);
			39208: out = 16'(738);
			39209: out = 16'(251);
			39210: out = 16'(-184);
			39211: out = 16'(-587);
			39212: out = 16'(-741);
			39213: out = 16'(-575);
			39214: out = 16'(-28);
			39215: out = 16'(-165);
			39216: out = 16'(-153);
			39217: out = 16'(109);
			39218: out = 16'(354);
			39219: out = 16'(63);
			39220: out = 16'(-109);
			39221: out = 16'(160);
			39222: out = 16'(448);
			39223: out = 16'(-80);
			39224: out = 16'(-597);
			39225: out = 16'(-298);
			39226: out = 16'(618);
			39227: out = 16'(352);
			39228: out = 16'(137);
			39229: out = 16'(-257);
			39230: out = 16'(-649);
			39231: out = 16'(-1290);
			39232: out = 16'(-953);
			39233: out = 16'(-376);
			39234: out = 16'(124);
			39235: out = 16'(139);
			39236: out = 16'(726);
			39237: out = 16'(655);
			39238: out = 16'(257);
			39239: out = 16'(134);
			39240: out = 16'(327);
			39241: out = 16'(441);
			39242: out = 16'(168);
			39243: out = 16'(-209);
			39244: out = 16'(16);
			39245: out = 16'(399);
			39246: out = 16'(404);
			39247: out = 16'(-85);
			39248: out = 16'(-950);
			39249: out = 16'(-366);
			39250: out = 16'(339);
			39251: out = 16'(394);
			39252: out = 16'(-209);
			39253: out = 16'(-463);
			39254: out = 16'(-416);
			39255: out = 16'(1);
			39256: out = 16'(403);
			39257: out = 16'(738);
			39258: out = 16'(418);
			39259: out = 16'(-233);
			39260: out = 16'(-879);
			39261: out = 16'(-664);
			39262: out = 16'(-523);
			39263: out = 16'(15);
			39264: out = 16'(590);
			39265: out = 16'(770);
			39266: out = 16'(84);
			39267: out = 16'(-318);
			39268: out = 16'(-146);
			39269: out = 16'(-51);
			39270: out = 16'(-264);
			39271: out = 16'(-353);
			39272: out = 16'(-36);
			39273: out = 16'(390);
			39274: out = 16'(158);
			39275: out = 16'(99);
			39276: out = 16'(33);
			39277: out = 16'(-239);
			39278: out = 16'(-350);
			39279: out = 16'(-97);
			39280: out = 16'(313);
			39281: out = 16'(462);
			39282: out = 16'(-8);
			39283: out = 16'(-64);
			39284: out = 16'(-192);
			39285: out = 16'(-406);
			39286: out = 16'(-344);
			39287: out = 16'(-12);
			39288: out = 16'(102);
			39289: out = 16'(-144);
			39290: out = 16'(-313);
			39291: out = 16'(-528);
			39292: out = 16'(-222);
			39293: out = 16'(20);
			39294: out = 16'(-35);
			39295: out = 16'(-295);
			39296: out = 16'(-357);
			39297: out = 16'(-275);
			39298: out = 16'(-151);
			39299: out = 16'(77);
			39300: out = 16'(334);
			39301: out = 16'(433);
			39302: out = 16'(354);
			39303: out = 16'(-18);
			39304: out = 16'(-2);
			39305: out = 16'(-158);
			39306: out = 16'(-376);
			39307: out = 16'(-155);
			39308: out = 16'(242);
			39309: out = 16'(645);
			39310: out = 16'(705);
			39311: out = 16'(298);
			39312: out = 16'(44);
			39313: out = 16'(-462);
			39314: out = 16'(-708);
			39315: out = 16'(-426);
			39316: out = 16'(388);
			39317: out = 16'(489);
			39318: out = 16'(177);
			39319: out = 16'(-68);
			39320: out = 16'(-75);
			39321: out = 16'(241);
			39322: out = 16'(291);
			39323: out = 16'(-58);
			39324: out = 16'(-352);
			39325: out = 16'(-727);
			39326: out = 16'(-334);
			39327: out = 16'(128);
			39328: out = 16'(-73);
			39329: out = 16'(70);
			39330: out = 16'(304);
			39331: out = 16'(553);
			39332: out = 16'(434);
			39333: out = 16'(523);
			39334: out = 16'(98);
			39335: out = 16'(-226);
			39336: out = 16'(-492);
			39337: out = 16'(-836);
			39338: out = 16'(-722);
			39339: out = 16'(-125);
			39340: out = 16'(430);
			39341: out = 16'(334);
			39342: out = 16'(-71);
			39343: out = 16'(-453);
			39344: out = 16'(-549);
			39345: out = 16'(-529);
			39346: out = 16'(-290);
			39347: out = 16'(-185);
			39348: out = 16'(-318);
			39349: out = 16'(-470);
			39350: out = 16'(18);
			39351: out = 16'(555);
			39352: out = 16'(837);
			39353: out = 16'(665);
			39354: out = 16'(122);
			39355: out = 16'(-528);
			39356: out = 16'(-1121);
			39357: out = 16'(-964);
			39358: out = 16'(-111);
			39359: out = 16'(427);
			39360: out = 16'(-119);
			39361: out = 16'(-619);
			39362: out = 16'(33);
			39363: out = 16'(763);
			39364: out = 16'(561);
			39365: out = 16'(-235);
			39366: out = 16'(-624);
			39367: out = 16'(-129);
			39368: out = 16'(16);
			39369: out = 16'(0);
			39370: out = 16'(131);
			39371: out = 16'(-26);
			39372: out = 16'(-242);
			39373: out = 16'(-288);
			39374: out = 16'(100);
			39375: out = 16'(335);
			39376: out = 16'(221);
			39377: out = 16'(-233);
			39378: out = 16'(-617);
			39379: out = 16'(-802);
			39380: out = 16'(-218);
			39381: out = 16'(261);
			39382: out = 16'(330);
			39383: out = 16'(-56);
			39384: out = 16'(-417);
			39385: out = 16'(-547);
			39386: out = 16'(-384);
			39387: out = 16'(-160);
			39388: out = 16'(-169);
			39389: out = 16'(20);
			39390: out = 16'(294);
			39391: out = 16'(385);
			39392: out = 16'(161);
			39393: out = 16'(21);
			39394: out = 16'(32);
			39395: out = 16'(193);
			39396: out = 16'(401);
			39397: out = 16'(65);
			39398: out = 16'(-53);
			39399: out = 16'(-19);
			39400: out = 16'(-251);
			39401: out = 16'(-173);
			39402: out = 16'(-308);
			39403: out = 16'(-210);
			39404: out = 16'(216);
			39405: out = 16'(468);
			39406: out = 16'(332);
			39407: out = 16'(-112);
			39408: out = 16'(-358);
			39409: out = 16'(-364);
			39410: out = 16'(-12);
			39411: out = 16'(92);
			39412: out = 16'(-18);
			39413: out = 16'(156);
			39414: out = 16'(-16);
			39415: out = 16'(190);
			39416: out = 16'(390);
			39417: out = 16'(65);
			39418: out = 16'(406);
			39419: out = 16'(-99);
			39420: out = 16'(-763);
			39421: out = 16'(-864);
			39422: out = 16'(355);
			39423: out = 16'(860);
			39424: out = 16'(726);
			39425: out = 16'(289);
			39426: out = 16'(-1);
			39427: out = 16'(-3);
			39428: out = 16'(229);
			39429: out = 16'(296);
			39430: out = 16'(-48);
			39431: out = 16'(-784);
			39432: out = 16'(-1001);
			39433: out = 16'(-379);
			39434: out = 16'(386);
			39435: out = 16'(422);
			39436: out = 16'(133);
			39437: out = 16'(-197);
			39438: out = 16'(-350);
			39439: out = 16'(-77);
			39440: out = 16'(-13);
			39441: out = 16'(-96);
			39442: out = 16'(-221);
			39443: out = 16'(-211);
			39444: out = 16'(169);
			39445: out = 16'(660);
			39446: out = 16'(794);
			39447: out = 16'(80);
			39448: out = 16'(-19);
			39449: out = 16'(-448);
			39450: out = 16'(-924);
			39451: out = 16'(-599);
			39452: out = 16'(-228);
			39453: out = 16'(376);
			39454: out = 16'(306);
			39455: out = 16'(-412);
			39456: out = 16'(-939);
			39457: out = 16'(-479);
			39458: out = 16'(362);
			39459: out = 16'(733);
			39460: out = 16'(50);
			39461: out = 16'(-78);
			39462: out = 16'(0);
			39463: out = 16'(-77);
			39464: out = 16'(-203);
			39465: out = 16'(219);
			39466: out = 16'(475);
			39467: out = 16'(261);
			39468: out = 16'(-217);
			39469: out = 16'(-339);
			39470: out = 16'(-360);
			39471: out = 16'(-431);
			39472: out = 16'(-663);
			39473: out = 16'(-363);
			39474: out = 16'(-159);
			39475: out = 16'(217);
			39476: out = 16'(529);
			39477: out = 16'(460);
			39478: out = 16'(-388);
			39479: out = 16'(-851);
			39480: out = 16'(-266);
			39481: out = 16'(435);
			39482: out = 16'(646);
			39483: out = 16'(140);
			39484: out = 16'(-472);
			39485: out = 16'(-593);
			39486: out = 16'(103);
			39487: out = 16'(896);
			39488: out = 16'(951);
			39489: out = 16'(55);
			39490: out = 16'(101);
			39491: out = 16'(20);
			39492: out = 16'(-111);
			39493: out = 16'(-215);
			39494: out = 16'(-74);
			39495: out = 16'(-29);
			39496: out = 16'(-122);
			39497: out = 16'(-223);
			39498: out = 16'(-248);
			39499: out = 16'(22);
			39500: out = 16'(70);
			39501: out = 16'(-113);
			39502: out = 16'(-341);
			39503: out = 16'(-115);
			39504: out = 16'(2);
			39505: out = 16'(-50);
			39506: out = 16'(9);
			39507: out = 16'(397);
			39508: out = 16'(585);
			39509: out = 16'(369);
			39510: out = 16'(76);
			39511: out = 16'(-68);
			39512: out = 16'(-195);
			39513: out = 16'(-680);
			39514: out = 16'(-1149);
			39515: out = 16'(-708);
			39516: out = 16'(71);
			39517: out = 16'(661);
			39518: out = 16'(720);
			39519: out = 16'(398);
			39520: out = 16'(-166);
			39521: out = 16'(-592);
			39522: out = 16'(-556);
			39523: out = 16'(-10);
			39524: out = 16'(314);
			39525: out = 16'(349);
			39526: out = 16'(156);
			39527: out = 16'(-53);
			39528: out = 16'(-195);
			39529: out = 16'(-152);
			39530: out = 16'(137);
			39531: out = 16'(317);
			39532: out = 16'(-269);
			39533: out = 16'(-648);
			39534: out = 16'(-413);
			39535: out = 16'(202);
			39536: out = 16'(85);
			39537: out = 16'(22);
			39538: out = 16'(-93);
			39539: out = 16'(58);
			39540: out = 16'(373);
			39541: out = 16'(68);
			39542: out = 16'(-89);
			39543: out = 16'(-15);
			39544: out = 16'(-97);
			39545: out = 16'(114);
			39546: out = 16'(0);
			39547: out = 16'(-7);
			39548: out = 16'(108);
			39549: out = 16'(383);
			39550: out = 16'(-23);
			39551: out = 16'(-251);
			39552: out = 16'(79);
			39553: out = 16'(422);
			39554: out = 16'(185);
			39555: out = 16'(-500);
			39556: out = 16'(-777);
			39557: out = 16'(-222);
			39558: out = 16'(-64);
			39559: out = 16'(30);
			39560: out = 16'(220);
			39561: out = 16'(485);
			39562: out = 16'(427);
			39563: out = 16'(10);
			39564: out = 16'(-316);
			39565: out = 16'(-377);
			39566: out = 16'(38);
			39567: out = 16'(-395);
			39568: out = 16'(-645);
			39569: out = 16'(29);
			39570: out = 16'(923);
			39571: out = 16'(805);
			39572: out = 16'(150);
			39573: out = 16'(-442);
			39574: out = 16'(-702);
			39575: out = 16'(-604);
			39576: out = 16'(-422);
			39577: out = 16'(-224);
			39578: out = 16'(-23);
			39579: out = 16'(-50);
			39580: out = 16'(134);
			39581: out = 16'(358);
			39582: out = 16'(346);
			39583: out = 16'(-12);
			39584: out = 16'(-193);
			39585: out = 16'(-135);
			39586: out = 16'(-32);
			39587: out = 16'(-66);
			39588: out = 16'(-49);
			39589: out = 16'(-6);
			39590: out = 16'(73);
			39591: out = 16'(-68);
			39592: out = 16'(39);
			39593: out = 16'(10);
			39594: out = 16'(-56);
			39595: out = 16'(-74);
			39596: out = 16'(-441);
			39597: out = 16'(-620);
			39598: out = 16'(-301);
			39599: out = 16'(328);
			39600: out = 16'(309);
			39601: out = 16'(-61);
			39602: out = 16'(-296);
			39603: out = 16'(68);
			39604: out = 16'(221);
			39605: out = 16'(408);
			39606: out = 16'(205);
			39607: out = 16'(-79);
			39608: out = 16'(-87);
			39609: out = 16'(-47);
			39610: out = 16'(-113);
			39611: out = 16'(-202);
			39612: out = 16'(-185);
			39613: out = 16'(277);
			39614: out = 16'(369);
			39615: out = 16'(173);
			39616: out = 16'(58);
			39617: out = 16'(-50);
			39618: out = 16'(-74);
			39619: out = 16'(-143);
			39620: out = 16'(-193);
			39621: out = 16'(-54);
			39622: out = 16'(2);
			39623: out = 16'(144);
			39624: out = 16'(267);
			39625: out = 16'(261);
			39626: out = 16'(79);
			39627: out = 16'(-145);
			39628: out = 16'(-405);
			39629: out = 16'(-548);
			39630: out = 16'(-521);
			39631: out = 16'(-131);
			39632: out = 16'(58);
			39633: out = 16'(-33);
			39634: out = 16'(-5);
			39635: out = 16'(360);
			39636: out = 16'(520);
			39637: out = 16'(58);
			39638: out = 16'(-244);
			39639: out = 16'(-459);
			39640: out = 16'(-296);
			39641: out = 16'(-5);
			39642: out = 16'(159);
			39643: out = 16'(307);
			39644: out = 16'(313);
			39645: out = 16'(38);
			39646: out = 16'(-304);
			39647: out = 16'(-374);
			39648: out = 16'(-164);
			39649: out = 16'(-33);
			39650: out = 16'(50);
			39651: out = 16'(-92);
			39652: out = 16'(156);
			39653: out = 16'(130);
			39654: out = 16'(-363);
			39655: out = 16'(-181);
			39656: out = 16'(-129);
			39657: out = 16'(-43);
			39658: out = 16'(-88);
			39659: out = 16'(-32);
			39660: out = 16'(-73);
			39661: out = 16'(-46);
			39662: out = 16'(-72);
			39663: out = 16'(-193);
			39664: out = 16'(-32);
			39665: out = 16'(171);
			39666: out = 16'(282);
			39667: out = 16'(249);
			39668: out = 16'(-198);
			39669: out = 16'(-578);
			39670: out = 16'(-590);
			39671: out = 16'(-113);
			39672: out = 16'(216);
			39673: out = 16'(326);
			39674: out = 16'(150);
			39675: out = 16'(-44);
			39676: out = 16'(44);
			39677: out = 16'(81);
			39678: out = 16'(-1);
			39679: out = 16'(-41);
			39680: out = 16'(71);
			39681: out = 16'(-41);
			39682: out = 16'(-9);
			39683: out = 16'(67);
			39684: out = 16'(-77);
			39685: out = 16'(-139);
			39686: out = 16'(-354);
			39687: out = 16'(-322);
			39688: out = 16'(-12);
			39689: out = 16'(252);
			39690: out = 16'(-21);
			39691: out = 16'(-459);
			39692: out = 16'(-462);
			39693: out = 16'(-100);
			39694: out = 16'(171);
			39695: out = 16'(98);
			39696: out = 16'(-9);
			39697: out = 16'(280);
			39698: out = 16'(228);
			39699: out = 16'(66);
			39700: out = 16'(-80);
			39701: out = 16'(-27);
			39702: out = 16'(-56);
			39703: out = 16'(11);
			39704: out = 16'(23);
			39705: out = 16'(46);
			39706: out = 16'(-38);
			39707: out = 16'(-47);
			39708: out = 16'(-124);
			39709: out = 16'(-300);
			39710: out = 16'(-211);
			39711: out = 16'(120);
			39712: out = 16'(285);
			39713: out = 16'(113);
			39714: out = 16'(-30);
			39715: out = 16'(-101);
			39716: out = 16'(51);
			39717: out = 16'(149);
			39718: out = 16'(-58);
			39719: out = 16'(-60);
			39720: out = 16'(-59);
			39721: out = 16'(-180);
			39722: out = 16'(-550);
			39723: out = 16'(-147);
			39724: out = 16'(32);
			39725: out = 16'(45);
			39726: out = 16'(-63);
			39727: out = 16'(-15);
			39728: out = 16'(-68);
			39729: out = 16'(76);
			39730: out = 16'(287);
			39731: out = 16'(289);
			39732: out = 16'(44);
			39733: out = 16'(-82);
			39734: out = 16'(-63);
			39735: out = 16'(63);
			39736: out = 16'(-37);
			39737: out = 16'(83);
			39738: out = 16'(256);
			39739: out = 16'(149);
			39740: out = 16'(-334);
			39741: out = 16'(-291);
			39742: out = 16'(68);
			39743: out = 16'(112);
			39744: out = 16'(100);
			39745: out = 16'(-123);
			39746: out = 16'(-212);
			39747: out = 16'(-190);
			39748: out = 16'(-74);
			39749: out = 16'(14);
			39750: out = 16'(60);
			39751: out = 16'(50);
			39752: out = 16'(6);
			39753: out = 16'(-13);
			39754: out = 16'(-138);
			39755: out = 16'(-204);
			39756: out = 16'(-204);
			39757: out = 16'(-86);
			39758: out = 16'(-75);
			39759: out = 16'(42);
			39760: out = 16'(356);
			39761: out = 16'(394);
			39762: out = 16'(-32);
			39763: out = 16'(-462);
			39764: out = 16'(-400);
			39765: out = 16'(-163);
			39766: out = 16'(28);
			39767: out = 16'(30);
			39768: out = 16'(17);
			39769: out = 16'(-61);
			39770: out = 16'(151);
			39771: out = 16'(305);
			39772: out = 16'(164);
			39773: out = 16'(-50);
			39774: out = 16'(-474);
			39775: out = 16'(-565);
			39776: out = 16'(-329);
			39777: out = 16'(-49);
			39778: out = 16'(26);
			39779: out = 16'(152);
			39780: out = 16'(309);
			39781: out = 16'(223);
			39782: out = 16'(-36);
			39783: out = 16'(-266);
			39784: out = 16'(-402);
			39785: out = 16'(-599);
			39786: out = 16'(-655);
			39787: out = 16'(-541);
			39788: out = 16'(-88);
			39789: out = 16'(0);
			default: out = 0;
		endcase
	end
endmodule
