module kick_lookup(index, out);
	input logic unsigned [12:0] index;
	output logic signed [15:0] out;
	always_comb begin
		case(index)
			0: out = 16'(0);
			1: out = 16'(1259);
			2: out = 16'(1690);
			3: out = 16'(3209);
			4: out = 16'(3182);
			5: out = 16'(3069);
			6: out = 16'(4561);
			7: out = 16'(6078);
			8: out = 16'(6316);
			9: out = 16'(6881);
			10: out = 16'(6789);
			11: out = 16'(5283);
			12: out = 16'(5057);
			13: out = 16'(5497);
			14: out = 16'(7415);
			15: out = 16'(9756);
			16: out = 16'(14459);
			17: out = 16'(19484);
			18: out = 16'(24088);
			19: out = 16'(32312);
			20: out = 16'(32112);
			21: out = 16'(32061);
			22: out = 16'(31955);
			23: out = 16'(31859);
			24: out = 16'(31768);
			25: out = 16'(31670);
			26: out = 16'(31578);
			27: out = 16'(31474);
			28: out = 16'(31120);
			29: out = 16'(24857);
			30: out = 16'(22038);
			31: out = 16'(18218);
			32: out = 16'(11622);
			33: out = 16'(6324);
			34: out = 16'(696);
			35: out = 16'(-6732);
			36: out = 16'(-12712);
			37: out = 16'(-16357);
			38: out = 16'(-20442);
			39: out = 16'(-24487);
			40: out = 16'(-28912);
			41: out = 16'(-32561);
			42: out = 16'(-32521);
			43: out = 16'(-32432);
			44: out = 16'(-32354);
			45: out = 16'(-32262);
			46: out = 16'(-32161);
			47: out = 16'(-32061);
			48: out = 16'(-31963);
			49: out = 16'(-31859);
			50: out = 16'(-31750);
			51: out = 16'(-31614);
			52: out = 16'(-31410);
			53: out = 16'(-28673);
			54: out = 16'(-26871);
			55: out = 16'(-25403);
			56: out = 16'(-23297);
			57: out = 16'(-19508);
			58: out = 16'(-14095);
			59: out = 16'(-9140);
			60: out = 16'(-3197);
			61: out = 16'(2533);
			62: out = 16'(6175);
			63: out = 16'(10067);
			64: out = 16'(15980);
			65: out = 16'(20281);
			66: out = 16'(23240);
			67: out = 16'(24488);
			68: out = 16'(27362);
			69: out = 16'(31668);
			70: out = 16'(32481);
			71: out = 16'(32396);
			72: out = 16'(32294);
			73: out = 16'(32196);
			74: out = 16'(32101);
			75: out = 16'(31999);
			76: out = 16'(29814);
			77: out = 16'(26983);
			78: out = 16'(25692);
			79: out = 16'(24339);
			80: out = 16'(22692);
			81: out = 16'(19372);
			82: out = 16'(18178);
			83: out = 16'(16173);
			84: out = 16'(11296);
			85: out = 16'(8592);
			86: out = 16'(5284);
			87: out = 16'(1232);
			88: out = 16'(-4886);
			89: out = 16'(-9846);
			90: out = 16'(-14380);
			91: out = 16'(-18116);
			92: out = 16'(-20700);
			93: out = 16'(-24121);
			94: out = 16'(-26445);
			95: out = 16'(-29308);
			96: out = 16'(-32199);
			97: out = 16'(-32122);
			98: out = 16'(-32035);
			99: out = 16'(-31955);
			100: out = 16'(-31885);
			101: out = 16'(-31797);
			102: out = 16'(-31661);
			103: out = 16'(-31564);
			104: out = 16'(-31398);
			105: out = 16'(-31144);
			106: out = 16'(-28786);
			107: out = 16'(-27072);
			108: out = 16'(-26226);
			109: out = 16'(-26579);
			110: out = 16'(-23476);
			111: out = 16'(-20624);
			112: out = 16'(-17889);
			113: out = 16'(-16220);
			114: out = 16'(-13886);
			115: out = 16'(-11318);
			116: out = 16'(-8723);
			117: out = 16'(-5202);
			118: out = 16'(-1557);
			119: out = 16'(2459);
			120: out = 16'(5527);
			121: out = 16'(7832);
			122: out = 16'(11282);
			123: out = 16'(14702);
			124: out = 16'(17850);
			125: out = 16'(20041);
			126: out = 16'(24693);
			127: out = 16'(26560);
			128: out = 16'(29029);
			129: out = 16'(30251);
			130: out = 16'(32429);
			131: out = 16'(32679);
			132: out = 16'(32582);
			133: out = 16'(32479);
			134: out = 16'(32383);
			135: out = 16'(32289);
			136: out = 16'(32189);
			137: out = 16'(32098);
			138: out = 16'(31343);
			139: out = 16'(28658);
			140: out = 16'(26841);
			141: out = 16'(25576);
			142: out = 16'(24311);
			143: out = 16'(22031);
			144: out = 16'(19618);
			145: out = 16'(18304);
			146: out = 16'(15896);
			147: out = 16'(12664);
			148: out = 16'(11362);
			149: out = 16'(9401);
			150: out = 16'(6280);
			151: out = 16'(4229);
			152: out = 16'(1229);
			153: out = 16'(-1329);
			154: out = 16'(-4862);
			155: out = 16'(-8205);
			156: out = 16'(-12193);
			157: out = 16'(-15226);
			158: out = 16'(-18221);
			159: out = 16'(-20249);
			160: out = 16'(-22653);
			161: out = 16'(-25328);
			162: out = 16'(-26945);
			163: out = 16'(-28369);
			164: out = 16'(-29324);
			165: out = 16'(-30874);
			166: out = 16'(-29739);
			167: out = 16'(-30481);
			168: out = 16'(-31698);
			169: out = 16'(-31655);
			170: out = 16'(-31388);
			171: out = 16'(-31363);
			172: out = 16'(-30607);
			173: out = 16'(-28871);
			174: out = 16'(-27226);
			175: out = 16'(-26401);
			176: out = 16'(-25104);
			177: out = 16'(-24681);
			178: out = 16'(-23898);
			179: out = 16'(-23277);
			180: out = 16'(-21378);
			181: out = 16'(-18943);
			182: out = 16'(-16700);
			183: out = 16'(-15422);
			184: out = 16'(-14646);
			185: out = 16'(-12879);
			186: out = 16'(-10507);
			187: out = 16'(-9526);
			188: out = 16'(-7139);
			189: out = 16'(-5638);
			190: out = 16'(-4659);
			191: out = 16'(-1993);
			192: out = 16'(823);
			193: out = 16'(2450);
			194: out = 16'(4885);
			195: out = 16'(7214);
			196: out = 16'(9390);
			197: out = 16'(11307);
			198: out = 16'(13037);
			199: out = 16'(14326);
			200: out = 16'(15761);
			201: out = 16'(18576);
			202: out = 16'(20391);
			203: out = 16'(22512);
			204: out = 16'(24664);
			205: out = 16'(25025);
			206: out = 16'(26348);
			207: out = 16'(27576);
			208: out = 16'(28649);
			209: out = 16'(30042);
			210: out = 16'(31368);
			211: out = 16'(31613);
			212: out = 16'(31104);
			213: out = 16'(30282);
			214: out = 16'(29682);
			215: out = 16'(29331);
			216: out = 16'(28403);
			217: out = 16'(27032);
			218: out = 16'(25982);
			219: out = 16'(24680);
			220: out = 16'(23742);
			221: out = 16'(21842);
			222: out = 16'(20849);
			223: out = 16'(19003);
			224: out = 16'(17571);
			225: out = 16'(15591);
			226: out = 16'(14335);
			227: out = 16'(13101);
			228: out = 16'(11828);
			229: out = 16'(10187);
			230: out = 16'(9865);
			231: out = 16'(8369);
			232: out = 16'(7566);
			233: out = 16'(6482);
			234: out = 16'(4651);
			235: out = 16'(2968);
			236: out = 16'(1087);
			237: out = 16'(-1187);
			238: out = 16'(-3633);
			239: out = 16'(-5880);
			240: out = 16'(-8893);
			241: out = 16'(-11778);
			242: out = 16'(-13863);
			243: out = 16'(-15936);
			244: out = 16'(-17568);
			245: out = 16'(-19162);
			246: out = 16'(-20687);
			247: out = 16'(-21615);
			248: out = 16'(-22504);
			249: out = 16'(-23498);
			250: out = 16'(-24208);
			251: out = 16'(-25423);
			252: out = 16'(-26753);
			253: out = 16'(-27244);
			254: out = 16'(-27397);
			255: out = 16'(-28007);
			256: out = 16'(-27981);
			257: out = 16'(-28311);
			258: out = 16'(-28484);
			259: out = 16'(-28803);
			260: out = 16'(-28503);
			261: out = 16'(-27687);
			262: out = 16'(-27119);
			263: out = 16'(-26085);
			264: out = 16'(-25220);
			265: out = 16'(-24537);
			266: out = 16'(-23428);
			267: out = 16'(-22071);
			268: out = 16'(-20494);
			269: out = 16'(-19640);
			270: out = 16'(-18451);
			271: out = 16'(-18045);
			272: out = 16'(-17257);
			273: out = 16'(-16254);
			274: out = 16'(-15511);
			275: out = 16'(-14245);
			276: out = 16'(-12607);
			277: out = 16'(-11144);
			278: out = 16'(-10027);
			279: out = 16'(-8818);
			280: out = 16'(-7969);
			281: out = 16'(-6882);
			282: out = 16'(-5890);
			283: out = 16'(-5379);
			284: out = 16'(-4481);
			285: out = 16'(-3386);
			286: out = 16'(-2151);
			287: out = 16'(-756);
			288: out = 16'(798);
			289: out = 16'(1939);
			290: out = 16'(3190);
			291: out = 16'(5202);
			292: out = 16'(6834);
			293: out = 16'(8468);
			294: out = 16'(10126);
			295: out = 16'(11344);
			296: out = 16'(12446);
			297: out = 16'(13878);
			298: out = 16'(15129);
			299: out = 16'(16275);
			300: out = 16'(17468);
			301: out = 16'(18380);
			302: out = 16'(19446);
			303: out = 16'(20357);
			304: out = 16'(21237);
			305: out = 16'(22175);
			306: out = 16'(23211);
			307: out = 16'(24050);
			308: out = 16'(24948);
			309: out = 16'(25549);
			310: out = 16'(26295);
			311: out = 16'(26758);
			312: out = 16'(27155);
			313: out = 16'(27872);
			314: out = 16'(27872);
			315: out = 16'(27597);
			316: out = 16'(27329);
			317: out = 16'(26517);
			318: out = 16'(25912);
			319: out = 16'(25244);
			320: out = 16'(24352);
			321: out = 16'(23808);
			322: out = 16'(22833);
			323: out = 16'(21735);
			324: out = 16'(20700);
			325: out = 16'(19807);
			326: out = 16'(18822);
			327: out = 16'(17716);
			328: out = 16'(17008);
			329: out = 16'(16102);
			330: out = 16'(15304);
			331: out = 16'(14353);
			332: out = 16'(13357);
			333: out = 16'(12489);
			334: out = 16'(11267);
			335: out = 16'(10087);
			336: out = 16'(9014);
			337: out = 16'(8121);
			338: out = 16'(7304);
			339: out = 16'(6392);
			340: out = 16'(5519);
			341: out = 16'(4613);
			342: out = 16'(3607);
			343: out = 16'(2885);
			344: out = 16'(1863);
			345: out = 16'(990);
			346: out = 16'(73);
			347: out = 16'(-984);
			348: out = 16'(-1946);
			349: out = 16'(-3217);
			350: out = 16'(-4602);
			351: out = 16'(-5868);
			352: out = 16'(-7205);
			353: out = 16'(-8906);
			354: out = 16'(-10492);
			355: out = 16'(-12017);
			356: out = 16'(-13184);
			357: out = 16'(-14464);
			358: out = 16'(-15818);
			359: out = 16'(-16855);
			360: out = 16'(-17874);
			361: out = 16'(-18870);
			362: out = 16'(-19598);
			363: out = 16'(-20312);
			364: out = 16'(-21078);
			365: out = 16'(-21737);
			366: out = 16'(-22297);
			367: out = 16'(-22824);
			368: out = 16'(-23162);
			369: out = 16'(-23468);
			370: out = 16'(-23589);
			371: out = 16'(-23866);
			372: out = 16'(-24034);
			373: out = 16'(-24191);
			374: out = 16'(-24289);
			375: out = 16'(-24291);
			376: out = 16'(-24499);
			377: out = 16'(-24464);
			378: out = 16'(-24609);
			379: out = 16'(-24375);
			380: out = 16'(-24087);
			381: out = 16'(-23621);
			382: out = 16'(-23045);
			383: out = 16'(-22545);
			384: out = 16'(-21847);
			385: out = 16'(-21100);
			386: out = 16'(-20299);
			387: out = 16'(-19313);
			388: out = 16'(-18485);
			389: out = 16'(-17507);
			390: out = 16'(-16648);
			391: out = 16'(-15843);
			392: out = 16'(-15127);
			393: out = 16'(-14376);
			394: out = 16'(-13567);
			395: out = 16'(-12911);
			396: out = 16'(-12230);
			397: out = 16'(-11609);
			398: out = 16'(-10994);
			399: out = 16'(-10296);
			400: out = 16'(-9520);
			401: out = 16'(-8619);
			402: out = 16'(-7772);
			403: out = 16'(-6936);
			404: out = 16'(-6187);
			405: out = 16'(-5521);
			406: out = 16'(-4821);
			407: out = 16'(-4140);
			408: out = 16'(-3472);
			409: out = 16'(-2807);
			410: out = 16'(-2043);
			411: out = 16'(-1399);
			412: out = 16'(-760);
			413: out = 16'(-93);
			414: out = 16'(575);
			415: out = 16'(1268);
			416: out = 16'(1960);
			417: out = 16'(2838);
			418: out = 16'(3704);
			419: out = 16'(4681);
			420: out = 16'(5665);
			421: out = 16'(6749);
			422: out = 16'(7802);
			423: out = 16'(8725);
			424: out = 16'(9704);
			425: out = 16'(10601);
			426: out = 16'(11528);
			427: out = 16'(12322);
			428: out = 16'(13094);
			429: out = 16'(13899);
			430: out = 16'(14695);
			431: out = 16'(15412);
			432: out = 16'(16103);
			433: out = 16'(16734);
			434: out = 16'(17292);
			435: out = 16'(17852);
			436: out = 16'(18367);
			437: out = 16'(18887);
			438: out = 16'(19365);
			439: out = 16'(19878);
			440: out = 16'(20370);
			441: out = 16'(20766);
			442: out = 16'(21191);
			443: out = 16'(21569);
			444: out = 16'(21901);
			445: out = 16'(22242);
			446: out = 16'(22569);
			447: out = 16'(22868);
			448: out = 16'(23119);
			449: out = 16'(23271);
			450: out = 16'(23334);
			451: out = 16'(23278);
			452: out = 16'(23041);
			453: out = 16'(22678);
			454: out = 16'(22205);
			455: out = 16'(21656);
			456: out = 16'(21056);
			457: out = 16'(20422);
			458: out = 16'(19752);
			459: out = 16'(19035);
			460: out = 16'(18323);
			461: out = 16'(17607);
			462: out = 16'(16909);
			463: out = 16'(16165);
			464: out = 16'(15447);
			465: out = 16'(14779);
			466: out = 16'(14118);
			467: out = 16'(13474);
			468: out = 16'(12797);
			469: out = 16'(12194);
			470: out = 16'(11575);
			471: out = 16'(11038);
			472: out = 16'(10495);
			473: out = 16'(9979);
			474: out = 16'(9491);
			475: out = 16'(9014);
			476: out = 16'(8528);
			477: out = 16'(8069);
			478: out = 16'(7666);
			479: out = 16'(7036);
			480: out = 16'(6198);
			481: out = 16'(5412);
			482: out = 16'(4664);
			483: out = 16'(3988);
			484: out = 16'(3346);
			485: out = 16'(2711);
			486: out = 16'(2110);
			487: out = 16'(1531);
			488: out = 16'(949);
			489: out = 16'(412);
			490: out = 16'(-176);
			491: out = 16'(-736);
			492: out = 16'(-1271);
			493: out = 16'(-1808);
			494: out = 16'(-2346);
			495: out = 16'(-2950);
			496: out = 16'(-3552);
			497: out = 16'(-4173);
			498: out = 16'(-4857);
			499: out = 16'(-5582);
			500: out = 16'(-6363);
			501: out = 16'(-7226);
			502: out = 16'(-8125);
			503: out = 16'(-9056);
			504: out = 16'(-10012);
			505: out = 16'(-10989);
			506: out = 16'(-11952);
			507: out = 16'(-12872);
			508: out = 16'(-13759);
			509: out = 16'(-14561);
			510: out = 16'(-15320);
			511: out = 16'(-16040);
			512: out = 16'(-16689);
			513: out = 16'(-17277);
			514: out = 16'(-17839);
			515: out = 16'(-18278);
			516: out = 16'(-18718);
			517: out = 16'(-19061);
			518: out = 16'(-19407);
			519: out = 16'(-19716);
			520: out = 16'(-19959);
			521: out = 16'(-20155);
			522: out = 16'(-20363);
			523: out = 16'(-20494);
			524: out = 16'(-20620);
			525: out = 16'(-20712);
			526: out = 16'(-20774);
			527: out = 16'(-20801);
			528: out = 16'(-20841);
			529: out = 16'(-20852);
			530: out = 16'(-20830);
			531: out = 16'(-20783);
			532: out = 16'(-20746);
			533: out = 16'(-20668);
			534: out = 16'(-20546);
			535: out = 16'(-20376);
			536: out = 16'(-20214);
			537: out = 16'(-20016);
			538: out = 16'(-19755);
			539: out = 16'(-19419);
			540: out = 16'(-19056);
			541: out = 16'(-18611);
			542: out = 16'(-18108);
			543: out = 16'(-17533);
			544: out = 16'(-16918);
			545: out = 16'(-16254);
			546: out = 16'(-15623);
			547: out = 16'(-14929);
			548: out = 16'(-14245);
			549: out = 16'(-13594);
			550: out = 16'(-12921);
			551: out = 16'(-12308);
			552: out = 16'(-11686);
			553: out = 16'(-11087);
			554: out = 16'(-10527);
			555: out = 16'(-9971);
			556: out = 16'(-9435);
			557: out = 16'(-8915);
			558: out = 16'(-8431);
			559: out = 16'(-7953);
			560: out = 16'(-7504);
			561: out = 16'(-7074);
			562: out = 16'(-6675);
			563: out = 16'(-6102);
			564: out = 16'(-5464);
			565: out = 16'(-4873);
			566: out = 16'(-4300);
			567: out = 16'(-3741);
			568: out = 16'(-3251);
			569: out = 16'(-2759);
			570: out = 16'(-2301);
			571: out = 16'(-1863);
			572: out = 16'(-1411);
			573: out = 16'(-999);
			574: out = 16'(-563);
			575: out = 16'(-138);
			576: out = 16'(268);
			577: out = 16'(684);
			578: out = 16'(1138);
			579: out = 16'(1530);
			580: out = 16'(1957);
			581: out = 16'(2446);
			582: out = 16'(2965);
			583: out = 16'(3494);
			584: out = 16'(4085);
			585: out = 16'(4705);
			586: out = 16'(5369);
			587: out = 16'(6071);
			588: out = 16'(6790);
			589: out = 16'(7524);
			590: out = 16'(8220);
			591: out = 16'(8917);
			592: out = 16'(9588);
			593: out = 16'(10264);
			594: out = 16'(10876);
			595: out = 16'(11473);
			596: out = 16'(12048);
			597: out = 16'(12563);
			598: out = 16'(13086);
			599: out = 16'(13614);
			600: out = 16'(14067);
			601: out = 16'(14548);
			602: out = 16'(14940);
			603: out = 16'(15340);
			604: out = 16'(15723);
			605: out = 16'(16101);
			606: out = 16'(16447);
			607: out = 16'(16777);
			608: out = 16'(17091);
			609: out = 16'(17393);
			610: out = 16'(17700);
			611: out = 16'(17969);
			612: out = 16'(18244);
			613: out = 16'(18532);
			614: out = 16'(18774);
			615: out = 16'(19012);
			616: out = 16'(19234);
			617: out = 16'(19283);
			618: out = 16'(19389);
			619: out = 16'(19258);
			620: out = 16'(19194);
			621: out = 16'(19156);
			622: out = 16'(19085);
			623: out = 16'(19045);
			624: out = 16'(18858);
			625: out = 16'(18788);
			626: out = 16'(18533);
			627: out = 16'(18392);
			628: out = 16'(18181);
			629: out = 16'(17937);
			630: out = 16'(17613);
			631: out = 16'(17247);
			632: out = 16'(16825);
			633: out = 16'(16399);
			634: out = 16'(15898);
			635: out = 16'(15428);
			636: out = 16'(14925);
			637: out = 16'(14348);
			638: out = 16'(13858);
			639: out = 16'(13314);
			640: out = 16'(12829);
			641: out = 16'(12238);
			642: out = 16'(11775);
			643: out = 16'(11273);
			644: out = 16'(10751);
			645: out = 16'(10281);
			646: out = 16'(9828);
			647: out = 16'(9389);
			648: out = 16'(8943);
			649: out = 16'(8523);
			650: out = 16'(8107);
			651: out = 16'(7729);
			652: out = 16'(7344);
			653: out = 16'(6992);
			654: out = 16'(6635);
			655: out = 16'(6314);
			656: out = 16'(5989);
			657: out = 16'(5662);
			658: out = 16'(5385);
			659: out = 16'(5087);
			660: out = 16'(4807);
			661: out = 16'(4467);
			662: out = 16'(3853);
			663: out = 16'(3251);
			664: out = 16'(2699);
			665: out = 16'(2192);
			666: out = 16'(1712);
			667: out = 16'(1248);
			668: out = 16'(775);
			669: out = 16'(342);
			670: out = 16'(-83);
			671: out = 16'(-489);
			672: out = 16'(-894);
			673: out = 16'(-1288);
			674: out = 16'(-1631);
			675: out = 16'(-2060);
			676: out = 16'(-2474);
			677: out = 16'(-2859);
			678: out = 16'(-3274);
			679: out = 16'(-3691);
			680: out = 16'(-4083);
			681: out = 16'(-4521);
			682: out = 16'(-4982);
			683: out = 16'(-5466);
			684: out = 16'(-5980);
			685: out = 16'(-6529);
			686: out = 16'(-7115);
			687: out = 16'(-7753);
			688: out = 16'(-8409);
			689: out = 16'(-9129);
			690: out = 16'(-9830);
			691: out = 16'(-10563);
			692: out = 16'(-11343);
			693: out = 16'(-12003);
			694: out = 16'(-12688);
			695: out = 16'(-13321);
			696: out = 16'(-13901);
			697: out = 16'(-14458);
			698: out = 16'(-14979);
			699: out = 16'(-15441);
			700: out = 16'(-15863);
			701: out = 16'(-16251);
			702: out = 16'(-16600);
			703: out = 16'(-16907);
			704: out = 16'(-17159);
			705: out = 16'(-17403);
			706: out = 16'(-17642);
			707: out = 16'(-17807);
			708: out = 16'(-17919);
			709: out = 16'(-18062);
			710: out = 16'(-18170);
			711: out = 16'(-18218);
			712: out = 16'(-18266);
			713: out = 16'(-18274);
			714: out = 16'(-18326);
			715: out = 16'(-18320);
			716: out = 16'(-18305);
			717: out = 16'(-18297);
			718: out = 16'(-18244);
			719: out = 16'(-18192);
			720: out = 16'(-18129);
			721: out = 16'(-18026);
			722: out = 16'(-17911);
			723: out = 16'(-17807);
			724: out = 16'(-17647);
			725: out = 16'(-17531);
			726: out = 16'(-17393);
			727: out = 16'(-17214);
			728: out = 16'(-17003);
			729: out = 16'(-16789);
			730: out = 16'(-16523);
			731: out = 16'(-16207);
			732: out = 16'(-15878);
			733: out = 16'(-15482);
			734: out = 16'(-15042);
			735: out = 16'(-14576);
			736: out = 16'(-14089);
			737: out = 16'(-13551);
			738: out = 16'(-13033);
			739: out = 16'(-12449);
			740: out = 16'(-11887);
			741: out = 16'(-11347);
			742: out = 16'(-10806);
			743: out = 16'(-10266);
			744: out = 16'(-9763);
			745: out = 16'(-9260);
			746: out = 16'(-8789);
			747: out = 16'(-8305);
			748: out = 16'(-7853);
			749: out = 16'(-7403);
			750: out = 16'(-6974);
			751: out = 16'(-6570);
			752: out = 16'(-6198);
			753: out = 16'(-5834);
			754: out = 16'(-5495);
			755: out = 16'(-5153);
			756: out = 16'(-4826);
			757: out = 16'(-4510);
			758: out = 16'(-4114);
			759: out = 16'(-3620);
			760: out = 16'(-3133);
			761: out = 16'(-2719);
			762: out = 16'(-2293);
			763: out = 16'(-1914);
			764: out = 16'(-1531);
			765: out = 16'(-1169);
			766: out = 16'(-829);
			767: out = 16'(-495);
			768: out = 16'(-175);
			769: out = 16'(140);
			770: out = 16'(463);
			771: out = 16'(719);
			772: out = 16'(1031);
			773: out = 16'(1298);
			774: out = 16'(1582);
			775: out = 16'(1861);
			776: out = 16'(2191);
			777: out = 16'(2514);
			778: out = 16'(2848);
			779: out = 16'(3210);
			780: out = 16'(3575);
			781: out = 16'(3977);
			782: out = 16'(4379);
			783: out = 16'(4840);
			784: out = 16'(5338);
			785: out = 16'(5830);
			786: out = 16'(6364);
			787: out = 16'(6882);
			788: out = 16'(7412);
			789: out = 16'(7934);
			790: out = 16'(8421);
			791: out = 16'(8900);
			792: out = 16'(9382);
			793: out = 16'(9812);
			794: out = 16'(10244);
			795: out = 16'(10652);
			796: out = 16'(11060);
			797: out = 16'(11405);
			798: out = 16'(11741);
			799: out = 16'(12085);
			800: out = 16'(12383);
			801: out = 16'(12676);
			802: out = 16'(12978);
			803: out = 16'(13246);
			804: out = 16'(13518);
			805: out = 16'(13746);
			806: out = 16'(13935);
			807: out = 16'(14172);
			808: out = 16'(14387);
			809: out = 16'(14575);
			810: out = 16'(14772);
			811: out = 16'(14952);
			812: out = 16'(15120);
			813: out = 16'(15284);
			814: out = 16'(15425);
			815: out = 16'(15484);
			816: out = 16'(15437);
			817: out = 16'(15405);
			818: out = 16'(15309);
			819: out = 16'(15267);
			820: out = 16'(15240);
			821: out = 16'(15145);
			822: out = 16'(15114);
			823: out = 16'(15021);
			824: out = 16'(15046);
			825: out = 16'(14895);
			826: out = 16'(14891);
			827: out = 16'(14845);
			828: out = 16'(14743);
			829: out = 16'(14565);
			830: out = 16'(14477);
			831: out = 16'(14282);
			832: out = 16'(14111);
			833: out = 16'(13873);
			834: out = 16'(13614);
			835: out = 16'(13333);
			836: out = 16'(13037);
			837: out = 16'(12598);
			838: out = 16'(12257);
			839: out = 16'(11896);
			840: out = 16'(11476);
			841: out = 16'(11058);
			842: out = 16'(10668);
			843: out = 16'(10269);
			844: out = 16'(9850);
			845: out = 16'(9437);
			846: out = 16'(9058);
			847: out = 16'(8642);
			848: out = 16'(8267);
			849: out = 16'(7880);
			850: out = 16'(7538);
			851: out = 16'(7183);
			852: out = 16'(6845);
			853: out = 16'(6481);
			854: out = 16'(6194);
			855: out = 16'(5866);
			856: out = 16'(5559);
			857: out = 16'(5288);
			858: out = 16'(5040);
			859: out = 16'(4766);
			860: out = 16'(4529);
			861: out = 16'(4272);
			862: out = 16'(4050);
			863: out = 16'(3819);
			864: out = 16'(3594);
			865: out = 16'(3386);
			866: out = 16'(3200);
			867: out = 16'(2997);
			868: out = 16'(2827);
			869: out = 16'(2404);
			870: out = 16'(1963);
			871: out = 16'(1567);
			872: out = 16'(1169);
			873: out = 16'(786);
			874: out = 16'(434);
			875: out = 16'(67);
			876: out = 16'(-274);
			877: out = 16'(-597);
			878: out = 16'(-884);
			879: out = 16'(-1152);
			880: out = 16'(-1450);
			881: out = 16'(-1724);
			882: out = 16'(-2010);
			883: out = 16'(-2280);
			884: out = 16'(-2570);
			885: out = 16'(-2819);
			886: out = 16'(-3110);
			887: out = 16'(-3393);
			888: out = 16'(-3661);
			889: out = 16'(-3950);
			890: out = 16'(-4250);
			891: out = 16'(-4589);
			892: out = 16'(-4926);
			893: out = 16'(-5323);
			894: out = 16'(-5714);
			895: out = 16'(-6132);
			896: out = 16'(-6593);
			897: out = 16'(-7084);
			898: out = 16'(-7571);
			899: out = 16'(-8118);
			900: out = 16'(-8654);
			901: out = 16'(-9201);
			902: out = 16'(-9717);
			903: out = 16'(-10248);
			904: out = 16'(-10720);
			905: out = 16'(-11197);
			906: out = 16'(-11615);
			907: out = 16'(-12030);
			908: out = 16'(-12410);
			909: out = 16'(-12738);
			910: out = 16'(-13045);
			911: out = 16'(-13333);
			912: out = 16'(-13563);
			913: out = 16'(-13766);
			914: out = 16'(-13976);
			915: out = 16'(-14109);
			916: out = 16'(-14264);
			917: out = 16'(-14403);
			918: out = 16'(-14521);
			919: out = 16'(-14595);
			920: out = 16'(-14633);
			921: out = 16'(-14692);
			922: out = 16'(-14717);
			923: out = 16'(-14714);
			924: out = 16'(-14719);
			925: out = 16'(-14705);
			926: out = 16'(-14675);
			927: out = 16'(-14644);
			928: out = 16'(-14591);
			929: out = 16'(-14563);
			930: out = 16'(-14502);
			931: out = 16'(-14421);
			932: out = 16'(-14336);
			933: out = 16'(-14226);
			934: out = 16'(-14135);
			935: out = 16'(-14035);
			936: out = 16'(-13929);
			937: out = 16'(-13799);
			938: out = 16'(-13663);
			939: out = 16'(-13519);
			940: out = 16'(-13332);
			941: out = 16'(-13153);
			942: out = 16'(-12929);
			943: out = 16'(-12698);
			944: out = 16'(-12426);
			945: out = 16'(-12132);
			946: out = 16'(-11804);
			947: out = 16'(-11448);
			948: out = 16'(-11068);
			949: out = 16'(-10666);
			950: out = 16'(-10251);
			951: out = 16'(-9829);
			952: out = 16'(-9414);
			953: out = 16'(-8978);
			954: out = 16'(-8535);
			955: out = 16'(-8120);
			956: out = 16'(-7724);
			957: out = 16'(-7334);
			958: out = 16'(-6944);
			959: out = 16'(-6561);
			960: out = 16'(-6220);
			961: out = 16'(-5866);
			962: out = 16'(-5522);
			963: out = 16'(-5203);
			964: out = 16'(-4901);
			965: out = 16'(-4616);
			966: out = 16'(-4333);
			967: out = 16'(-4052);
			968: out = 16'(-3812);
			969: out = 16'(-3558);
			970: out = 16'(-3323);
			971: out = 16'(-3098);
			972: out = 16'(-2813);
			973: out = 16'(-2441);
			974: out = 16'(-2080);
			975: out = 16'(-1756);
			976: out = 16'(-1427);
			977: out = 16'(-1146);
			978: out = 16'(-854);
			979: out = 16'(-590);
			980: out = 16'(-330);
			981: out = 16'(-86);
			982: out = 16'(136);
			983: out = 16'(391);
			984: out = 16'(600);
			985: out = 16'(820);
			986: out = 16'(1057);
			987: out = 16'(1247);
			988: out = 16'(1459);
			989: out = 16'(1674);
			990: out = 16'(1888);
			991: out = 16'(2112);
			992: out = 16'(2339);
			993: out = 16'(2600);
			994: out = 16'(2850);
			995: out = 16'(3117);
			996: out = 16'(3430);
			997: out = 16'(3753);
			998: out = 16'(4116);
			999: out = 16'(4479);
			1000: out = 16'(4855);
			1001: out = 16'(5246);
			1002: out = 16'(5639);
			1003: out = 16'(6025);
			1004: out = 16'(6444);
			1005: out = 16'(6826);
			1006: out = 16'(7179);
			1007: out = 16'(7580);
			1008: out = 16'(7913);
			1009: out = 16'(8249);
			1010: out = 16'(8561);
			1011: out = 16'(8874);
			1012: out = 16'(9162);
			1013: out = 16'(9433);
			1014: out = 16'(9693);
			1015: out = 16'(9937);
			1016: out = 16'(10192);
			1017: out = 16'(10421);
			1018: out = 16'(10636);
			1019: out = 16'(10828);
			1020: out = 16'(11019);
			1021: out = 16'(11201);
			1022: out = 16'(11363);
			1023: out = 16'(11547);
			1024: out = 16'(11708);
			1025: out = 16'(11856);
			1026: out = 16'(12013);
			1027: out = 16'(12163);
			1028: out = 16'(12307);
			1029: out = 16'(12415);
			1030: out = 16'(12489);
			1031: out = 16'(12452);
			1032: out = 16'(12421);
			1033: out = 16'(12380);
			1034: out = 16'(12344);
			1035: out = 16'(12246);
			1036: out = 16'(12248);
			1037: out = 16'(12169);
			1038: out = 16'(12108);
			1039: out = 16'(12144);
			1040: out = 16'(12012);
			1041: out = 16'(12020);
			1042: out = 16'(11965);
			1043: out = 16'(11953);
			1044: out = 16'(11927);
			1045: out = 16'(11835);
			1046: out = 16'(11711);
			1047: out = 16'(11692);
			1048: out = 16'(11517);
			1049: out = 16'(11439);
			1050: out = 16'(11213);
			1051: out = 16'(11026);
			1052: out = 16'(10864);
			1053: out = 16'(10601);
			1054: out = 16'(10345);
			1055: out = 16'(10108);
			1056: out = 16'(9789);
			1057: out = 16'(9476);
			1058: out = 16'(9187);
			1059: out = 16'(8870);
			1060: out = 16'(8547);
			1061: out = 16'(8234);
			1062: out = 16'(7909);
			1063: out = 16'(7586);
			1064: out = 16'(7282);
			1065: out = 16'(6974);
			1066: out = 16'(6660);
			1067: out = 16'(6356);
			1068: out = 16'(6081);
			1069: out = 16'(5808);
			1070: out = 16'(5528);
			1071: out = 16'(5253);
			1072: out = 16'(5000);
			1073: out = 16'(4769);
			1074: out = 16'(4507);
			1075: out = 16'(4280);
			1076: out = 16'(4065);
			1077: out = 16'(3833);
			1078: out = 16'(3643);
			1079: out = 16'(3459);
			1080: out = 16'(3286);
			1081: out = 16'(3103);
			1082: out = 16'(2933);
			1083: out = 16'(2737);
			1084: out = 16'(2607);
			1085: out = 16'(2446);
			1086: out = 16'(2294);
			1087: out = 16'(2134);
			1088: out = 16'(1772);
			1089: out = 16'(1417);
			1090: out = 16'(1058);
			1091: out = 16'(749);
			1092: out = 16'(448);
			1093: out = 16'(154);
			1094: out = 16'(-95);
			1095: out = 16'(-358);
			1096: out = 16'(-619);
			1097: out = 16'(-859);
			1098: out = 16'(-1056);
			1099: out = 16'(-1321);
			1100: out = 16'(-1546);
			1101: out = 16'(-1759);
			1102: out = 16'(-1969);
			1103: out = 16'(-2194);
			1104: out = 16'(-2406);
			1105: out = 16'(-2607);
			1106: out = 16'(-2812);
			1107: out = 16'(-3034);
			1108: out = 16'(-3256);
			1109: out = 16'(-3509);
			1110: out = 16'(-3787);
			1111: out = 16'(-4060);
			1112: out = 16'(-4369);
			1113: out = 16'(-4684);
			1114: out = 16'(-4994);
			1115: out = 16'(-5346);
			1116: out = 16'(-5722);
			1117: out = 16'(-6128);
			1118: out = 16'(-6525);
			1119: out = 16'(-6935);
			1120: out = 16'(-7381);
			1121: out = 16'(-7835);
			1122: out = 16'(-8254);
			1123: out = 16'(-8663);
			1124: out = 16'(-9043);
			1125: out = 16'(-9402);
			1126: out = 16'(-9706);
			1127: out = 16'(-10032);
			1128: out = 16'(-10309);
			1129: out = 16'(-10577);
			1130: out = 16'(-10818);
			1131: out = 16'(-11039);
			1132: out = 16'(-11225);
			1133: out = 16'(-11401);
			1134: out = 16'(-11539);
			1135: out = 16'(-11649);
			1136: out = 16'(-11772);
			1137: out = 16'(-11864);
			1138: out = 16'(-11915);
			1139: out = 16'(-11970);
			1140: out = 16'(-12014);
			1141: out = 16'(-12036);
			1142: out = 16'(-12051);
			1143: out = 16'(-12073);
			1144: out = 16'(-12043);
			1145: out = 16'(-12039);
			1146: out = 16'(-12012);
			1147: out = 16'(-11971);
			1148: out = 16'(-11936);
			1149: out = 16'(-11887);
			1150: out = 16'(-11825);
			1151: out = 16'(-11756);
			1152: out = 16'(-11684);
			1153: out = 16'(-11613);
			1154: out = 16'(-11511);
			1155: out = 16'(-11420);
			1156: out = 16'(-11330);
			1157: out = 16'(-11216);
			1158: out = 16'(-11112);
			1159: out = 16'(-10982);
			1160: out = 16'(-10837);
			1161: out = 16'(-10702);
			1162: out = 16'(-10537);
			1163: out = 16'(-10340);
			1164: out = 16'(-10142);
			1165: out = 16'(-9919);
			1166: out = 16'(-9653);
			1167: out = 16'(-9371);
			1168: out = 16'(-9079);
			1169: out = 16'(-8762);
			1170: out = 16'(-8404);
			1171: out = 16'(-8084);
			1172: out = 16'(-7740);
			1173: out = 16'(-7380);
			1174: out = 16'(-7045);
			1175: out = 16'(-6718);
			1176: out = 16'(-6398);
			1177: out = 16'(-6048);
			1178: out = 16'(-5748);
			1179: out = 16'(-5427);
			1180: out = 16'(-5129);
			1181: out = 16'(-4831);
			1182: out = 16'(-4574);
			1183: out = 16'(-4293);
			1184: out = 16'(-4045);
			1185: out = 16'(-3805);
			1186: out = 16'(-3571);
			1187: out = 16'(-3343);
			1188: out = 16'(-3144);
			1189: out = 16'(-2950);
			1190: out = 16'(-2738);
			1191: out = 16'(-2561);
			1192: out = 16'(-2382);
			1193: out = 16'(-2134);
			1194: out = 16'(-1823);
			1195: out = 16'(-1552);
			1196: out = 16'(-1279);
			1197: out = 16'(-1036);
			1198: out = 16'(-802);
			1199: out = 16'(-577);
			1200: out = 16'(-348);
			1201: out = 16'(-147);
			1202: out = 16'(27);
			1203: out = 16'(227);
			1204: out = 16'(401);
			1205: out = 16'(574);
			1206: out = 16'(756);
			1207: out = 16'(920);
			1208: out = 16'(1092);
			1209: out = 16'(1276);
			1210: out = 16'(1436);
			1211: out = 16'(1607);
			1212: out = 16'(1774);
			1213: out = 16'(1953);
			1214: out = 16'(2152);
			1215: out = 16'(2338);
			1216: out = 16'(2564);
			1217: out = 16'(2805);
			1218: out = 16'(3069);
			1219: out = 16'(3340);
			1220: out = 16'(3618);
			1221: out = 16'(3926);
			1222: out = 16'(4234);
			1223: out = 16'(4560);
			1224: out = 16'(4884);
			1225: out = 16'(5201);
			1226: out = 16'(5522);
			1227: out = 16'(5832);
			1228: out = 16'(6125);
			1229: out = 16'(6423);
			1230: out = 16'(6692);
			1231: out = 16'(6940);
			1232: out = 16'(7188);
			1233: out = 16'(7432);
			1234: out = 16'(7669);
			1235: out = 16'(7894);
			1236: out = 16'(8115);
			1237: out = 16'(8333);
			1238: out = 16'(8497);
			1239: out = 16'(8661);
			1240: out = 16'(8843);
			1241: out = 16'(8990);
			1242: out = 16'(9150);
			1243: out = 16'(9308);
			1244: out = 16'(9459);
			1245: out = 16'(9597);
			1246: out = 16'(9730);
			1247: out = 16'(9850);
			1248: out = 16'(9977);
			1249: out = 16'(10085);
			1250: out = 16'(10182);
			1251: out = 16'(10267);
			1252: out = 16'(10280);
			1253: out = 16'(10246);
			1254: out = 16'(10148);
			1255: out = 16'(10157);
			1256: out = 16'(10143);
			1257: out = 16'(10094);
			1258: out = 16'(10102);
			1259: out = 16'(10065);
			1260: out = 16'(10031);
			1261: out = 16'(10004);
			1262: out = 16'(10002);
			1263: out = 16'(9952);
			1264: out = 16'(9976);
			1265: out = 16'(9915);
			1266: out = 16'(9831);
			1267: out = 16'(9747);
			1268: out = 16'(9730);
			1269: out = 16'(9594);
			1270: out = 16'(9529);
			1271: out = 16'(9439);
			1272: out = 16'(9294);
			1273: out = 16'(9125);
			1274: out = 16'(8914);
			1275: out = 16'(8716);
			1276: out = 16'(8548);
			1277: out = 16'(8296);
			1278: out = 16'(8074);
			1279: out = 16'(7775);
			1280: out = 16'(7519);
			1281: out = 16'(7285);
			1282: out = 16'(6987);
			1283: out = 16'(6744);
			1284: out = 16'(6483);
			1285: out = 16'(6240);
			1286: out = 16'(5965);
			1287: out = 16'(5722);
			1288: out = 16'(5477);
			1289: out = 16'(5231);
			1290: out = 16'(4988);
			1291: out = 16'(4769);
			1292: out = 16'(4527);
			1293: out = 16'(4326);
			1294: out = 16'(4107);
			1295: out = 16'(3910);
			1296: out = 16'(3726);
			1297: out = 16'(3543);
			1298: out = 16'(3343);
			1299: out = 16'(3190);
			1300: out = 16'(3038);
			1301: out = 16'(2834);
			1302: out = 16'(2694);
			1303: out = 16'(2561);
			1304: out = 16'(2429);
			1305: out = 16'(2266);
			1306: out = 16'(2147);
			1307: out = 16'(2037);
			1308: out = 16'(1878);
			1309: out = 16'(1796);
			1310: out = 16'(1493);
			1311: out = 16'(1204);
			1312: out = 16'(925);
			1313: out = 16'(654);
			1314: out = 16'(416);
			1315: out = 16'(202);
			1316: out = 16'(-32);
			1317: out = 16'(-257);
			1318: out = 16'(-469);
			1319: out = 16'(-680);
			1320: out = 16'(-886);
			1321: out = 16'(-1081);
			1322: out = 16'(-1269);
			1323: out = 16'(-1429);
			1324: out = 16'(-1617);
			1325: out = 16'(-1800);
			1326: out = 16'(-1956);
			1327: out = 16'(-2149);
			1328: out = 16'(-2309);
			1329: out = 16'(-2498);
			1330: out = 16'(-2705);
			1331: out = 16'(-2903);
			1332: out = 16'(-3111);
			1333: out = 16'(-3350);
			1334: out = 16'(-3572);
			1335: out = 16'(-3820);
			1336: out = 16'(-4090);
			1337: out = 16'(-4381);
			1338: out = 16'(-4682);
			1339: out = 16'(-5003);
			1340: out = 16'(-5342);
			1341: out = 16'(-5711);
			1342: out = 16'(-6071);
			1343: out = 16'(-6411);
			1344: out = 16'(-6758);
			1345: out = 16'(-7128);
			1346: out = 16'(-7449);
			1347: out = 16'(-7740);
			1348: out = 16'(-8022);
			1349: out = 16'(-8292);
			1350: out = 16'(-8515);
			1351: out = 16'(-8746);
			1352: out = 16'(-8940);
			1353: out = 16'(-9118);
			1354: out = 16'(-9280);
			1355: out = 16'(-9400);
			1356: out = 16'(-9538);
			1357: out = 16'(-9643);
			1358: out = 16'(-9726);
			1359: out = 16'(-9796);
			1360: out = 16'(-9860);
			1361: out = 16'(-9895);
			1362: out = 16'(-9936);
			1363: out = 16'(-9977);
			1364: out = 16'(-9959);
			1365: out = 16'(-9961);
			1366: out = 16'(-9962);
			1367: out = 16'(-9968);
			1368: out = 16'(-9911);
			1369: out = 16'(-9885);
			1370: out = 16'(-9847);
			1371: out = 16'(-9806);
			1372: out = 16'(-9749);
			1373: out = 16'(-9686);
			1374: out = 16'(-9625);
			1375: out = 16'(-9566);
			1376: out = 16'(-9492);
			1377: out = 16'(-9401);
			1378: out = 16'(-9333);
			1379: out = 16'(-9235);
			1380: out = 16'(-9143);
			1381: out = 16'(-9053);
			1382: out = 16'(-8943);
			1383: out = 16'(-8799);
			1384: out = 16'(-8656);
			1385: out = 16'(-8521);
			1386: out = 16'(-8338);
			1387: out = 16'(-8158);
			1388: out = 16'(-7956);
			1389: out = 16'(-7731);
			1390: out = 16'(-7497);
			1391: out = 16'(-7244);
			1392: out = 16'(-6967);
			1393: out = 16'(-6690);
			1394: out = 16'(-6398);
			1395: out = 16'(-6121);
			1396: out = 16'(-5842);
			1397: out = 16'(-5558);
			1398: out = 16'(-5294);
			1399: out = 16'(-5039);
			1400: out = 16'(-4766);
			1401: out = 16'(-4505);
			1402: out = 16'(-4269);
			1403: out = 16'(-4027);
			1404: out = 16'(-3790);
			1405: out = 16'(-3577);
			1406: out = 16'(-3356);
			1407: out = 16'(-3148);
			1408: out = 16'(-2953);
			1409: out = 16'(-2781);
			1410: out = 16'(-2596);
			1411: out = 16'(-2436);
			1412: out = 16'(-2266);
			1413: out = 16'(-2126);
			1414: out = 16'(-1970);
			1415: out = 16'(-1813);
			1416: out = 16'(-1566);
			1417: out = 16'(-1314);
			1418: out = 16'(-1095);
			1419: out = 16'(-900);
			1420: out = 16'(-680);
			1421: out = 16'(-499);
			1422: out = 16'(-329);
			1423: out = 16'(-152);
			1424: out = 16'(3);
			1425: out = 16'(163);
			1426: out = 16'(317);
			1427: out = 16'(462);
			1428: out = 16'(596);
			1429: out = 16'(760);
			1430: out = 16'(880);
			1431: out = 16'(1006);
			1432: out = 16'(1143);
			1433: out = 16'(1299);
			1434: out = 16'(1427);
			1435: out = 16'(1590);
			1436: out = 16'(1723);
			1437: out = 16'(1885);
			1438: out = 16'(2068);
			1439: out = 16'(2266);
			1440: out = 16'(2467);
			1441: out = 16'(2665);
			1442: out = 16'(2903);
			1443: out = 16'(3139);
			1444: out = 16'(3390);
			1445: out = 16'(3651);
			1446: out = 16'(3909);
			1447: out = 16'(4186);
			1448: out = 16'(4441);
			1449: out = 16'(4693);
			1450: out = 16'(4944);
			1451: out = 16'(5173);
			1452: out = 16'(5397);
			1453: out = 16'(5617);
			1454: out = 16'(5828);
			1455: out = 16'(6017);
			1456: out = 16'(6218);
			1457: out = 16'(6406);
			1458: out = 16'(6571);
			1459: out = 16'(6746);
			1460: out = 16'(6891);
			1461: out = 16'(7048);
			1462: out = 16'(7195);
			1463: out = 16'(7339);
			1464: out = 16'(7468);
			1465: out = 16'(7575);
			1466: out = 16'(7706);
			1467: out = 16'(7823);
			1468: out = 16'(7934);
			1469: out = 16'(8062);
			1470: out = 16'(8149);
			1471: out = 16'(8246);
			1472: out = 16'(8346);
			1473: out = 16'(8427);
			1474: out = 16'(8467);
			1475: out = 16'(8405);
			1476: out = 16'(8444);
			1477: out = 16'(8368);
			1478: out = 16'(8372);
			1479: out = 16'(8304);
			1480: out = 16'(8332);
			1481: out = 16'(8292);
			1482: out = 16'(8269);
			1483: out = 16'(8281);
			1484: out = 16'(8218);
			1485: out = 16'(8238);
			1486: out = 16'(8248);
			1487: out = 16'(8159);
			1488: out = 16'(8102);
			1489: out = 16'(8113);
			1490: out = 16'(8080);
			1491: out = 16'(7998);
			1492: out = 16'(7914);
			1493: out = 16'(7849);
			1494: out = 16'(7737);
			1495: out = 16'(7637);
			1496: out = 16'(7504);
			1497: out = 16'(7332);
			1498: out = 16'(7146);
			1499: out = 16'(6960);
			1500: out = 16'(6826);
			1501: out = 16'(6602);
			1502: out = 16'(6376);
			1503: out = 16'(6182);
			1504: out = 16'(5954);
			1505: out = 16'(5748);
			1506: out = 16'(5520);
			1507: out = 16'(5287);
			1508: out = 16'(5072);
			1509: out = 16'(4867);
			1510: out = 16'(4656);
			1511: out = 16'(4442);
			1512: out = 16'(4264);
			1513: out = 16'(4071);
			1514: out = 16'(3896);
			1515: out = 16'(3713);
			1516: out = 16'(3532);
			1517: out = 16'(3329);
			1518: out = 16'(3182);
			1519: out = 16'(3034);
			1520: out = 16'(2889);
			1521: out = 16'(2741);
			1522: out = 16'(2601);
			1523: out = 16'(2453);
			1524: out = 16'(2330);
			1525: out = 16'(2192);
			1526: out = 16'(2077);
			1527: out = 16'(1963);
			1528: out = 16'(1868);
			1529: out = 16'(1761);
			1530: out = 16'(1660);
			1531: out = 16'(1551);
			1532: out = 16'(1376);
			1533: out = 16'(1108);
			1534: out = 16'(872);
			1535: out = 16'(670);
			1536: out = 16'(469);
			1537: out = 16'(243);
			1538: out = 16'(51);
			1539: out = 16'(-123);
			1540: out = 16'(-326);
			1541: out = 16'(-478);
			1542: out = 16'(-647);
			1543: out = 16'(-817);
			1544: out = 16'(-989);
			1545: out = 16'(-1107);
			1546: out = 16'(-1286);
			1547: out = 16'(-1404);
			1548: out = 16'(-1566);
			1549: out = 16'(-1713);
			1550: out = 16'(-1844);
			1551: out = 16'(-1992);
			1552: out = 16'(-2171);
			1553: out = 16'(-2332);
			1554: out = 16'(-2501);
			1555: out = 16'(-2678);
			1556: out = 16'(-2877);
			1557: out = 16'(-3086);
			1558: out = 16'(-3286);
			1559: out = 16'(-3515);
			1560: out = 16'(-3772);
			1561: out = 16'(-4046);
			1562: out = 16'(-4314);
			1563: out = 16'(-4602);
			1564: out = 16'(-4896);
			1565: out = 16'(-5187);
			1566: out = 16'(-5473);
			1567: out = 16'(-5777);
			1568: out = 16'(-6044);
			1569: out = 16'(-6312);
			1570: out = 16'(-6554);
			1571: out = 16'(-6777);
			1572: out = 16'(-6985);
			1573: out = 16'(-7160);
			1574: out = 16'(-7339);
			1575: out = 16'(-7486);
			1576: out = 16'(-7630);
			1577: out = 16'(-7745);
			1578: out = 16'(-7864);
			1579: out = 16'(-7943);
			1580: out = 16'(-8027);
			1581: out = 16'(-8091);
			1582: out = 16'(-8140);
			1583: out = 16'(-8178);
			1584: out = 16'(-8199);
			1585: out = 16'(-8220);
			1586: out = 16'(-8227);
			1587: out = 16'(-8223);
			1588: out = 16'(-8226);
			1589: out = 16'(-8206);
			1590: out = 16'(-8207);
			1591: out = 16'(-8184);
			1592: out = 16'(-8133);
			1593: out = 16'(-8096);
			1594: out = 16'(-8049);
			1595: out = 16'(-8005);
			1596: out = 16'(-7947);
			1597: out = 16'(-7887);
			1598: out = 16'(-7823);
			1599: out = 16'(-7758);
			1600: out = 16'(-7702);
			1601: out = 16'(-7624);
			1602: out = 16'(-7548);
			1603: out = 16'(-7457);
			1604: out = 16'(-7351);
			1605: out = 16'(-7256);
			1606: out = 16'(-7150);
			1607: out = 16'(-7039);
			1608: out = 16'(-6895);
			1609: out = 16'(-6760);
			1610: out = 16'(-6578);
			1611: out = 16'(-6416);
			1612: out = 16'(-6204);
			1613: out = 16'(-6012);
			1614: out = 16'(-5802);
			1615: out = 16'(-5578);
			1616: out = 16'(-5342);
			1617: out = 16'(-5099);
			1618: out = 16'(-4868);
			1619: out = 16'(-4640);
			1620: out = 16'(-4416);
			1621: out = 16'(-4194);
			1622: out = 16'(-3983);
			1623: out = 16'(-3756);
			1624: out = 16'(-3546);
			1625: out = 16'(-3345);
			1626: out = 16'(-3169);
			1627: out = 16'(-2986);
			1628: out = 16'(-2805);
			1629: out = 16'(-2635);
			1630: out = 16'(-2459);
			1631: out = 16'(-2317);
			1632: out = 16'(-2175);
			1633: out = 16'(-2016);
			1634: out = 16'(-1891);
			1635: out = 16'(-1778);
			1636: out = 16'(-1652);
			1637: out = 16'(-1535);
			1638: out = 16'(-1375);
			1639: out = 16'(-1166);
			1640: out = 16'(-978);
			1641: out = 16'(-795);
			1642: out = 16'(-636);
			1643: out = 16'(-483);
			1644: out = 16'(-346);
			1645: out = 16'(-203);
			1646: out = 16'(-56);
			1647: out = 16'(60);
			1648: out = 16'(183);
			1649: out = 16'(312);
			1650: out = 16'(423);
			1651: out = 16'(545);
			1652: out = 16'(647);
			1653: out = 16'(759);
			1654: out = 16'(856);
			1655: out = 16'(975);
			1656: out = 16'(1098);
			1657: out = 16'(1219);
			1658: out = 16'(1344);
			1659: out = 16'(1480);
			1660: out = 16'(1608);
			1661: out = 16'(1753);
			1662: out = 16'(1908);
			1663: out = 16'(2063);
			1664: out = 16'(2253);
			1665: out = 16'(2440);
			1666: out = 16'(2658);
			1667: out = 16'(2855);
			1668: out = 16'(3075);
			1669: out = 16'(3296);
			1670: out = 16'(3499);
			1671: out = 16'(3701);
			1672: out = 16'(3914);
			1673: out = 16'(4127);
			1674: out = 16'(4292);
			1675: out = 16'(4489);
			1676: out = 16'(4669);
			1677: out = 16'(4845);
			1678: out = 16'(5000);
			1679: out = 16'(5174);
			1680: out = 16'(5312);
			1681: out = 16'(5442);
			1682: out = 16'(5565);
			1683: out = 16'(5714);
			1684: out = 16'(5841);
			1685: out = 16'(5942);
			1686: out = 16'(6067);
			1687: out = 16'(6169);
			1688: out = 16'(6270);
			1689: out = 16'(6379);
			1690: out = 16'(6468);
			1691: out = 16'(6557);
			1692: out = 16'(6657);
			1693: out = 16'(6739);
			1694: out = 16'(6810);
			1695: out = 16'(6896);
			1696: out = 16'(6959);
			1697: out = 16'(6970);
			1698: out = 16'(6940);
			1699: out = 16'(6929);
			1700: out = 16'(6889);
			1701: out = 16'(6861);
			1702: out = 16'(6881);
			1703: out = 16'(6870);
			1704: out = 16'(6836);
			1705: out = 16'(6833);
			1706: out = 16'(6783);
			1707: out = 16'(6794);
			1708: out = 16'(6783);
			1709: out = 16'(6781);
			1710: out = 16'(6741);
			1711: out = 16'(6705);
			1712: out = 16'(6687);
			1713: out = 16'(6616);
			1714: out = 16'(6557);
			1715: out = 16'(6505);
			1716: out = 16'(6445);
			1717: out = 16'(6344);
			1718: out = 16'(6254);
			1719: out = 16'(6166);
			1720: out = 16'(6012);
			1721: out = 16'(5861);
			1722: out = 16'(5710);
			1723: out = 16'(5548);
			1724: out = 16'(5389);
			1725: out = 16'(5214);
			1726: out = 16'(5025);
			1727: out = 16'(4858);
			1728: out = 16'(4683);
			1729: out = 16'(4491);
			1730: out = 16'(4332);
			1731: out = 16'(4159);
			1732: out = 16'(3958);
			1733: out = 16'(3795);
			1734: out = 16'(3633);
			1735: out = 16'(3466);
			1736: out = 16'(3310);
			1737: out = 16'(3160);
			1738: out = 16'(3020);
			1739: out = 16'(2881);
			1740: out = 16'(2737);
			1741: out = 16'(2607);
			1742: out = 16'(2491);
			1743: out = 16'(2361);
			1744: out = 16'(2238);
			1745: out = 16'(2123);
			1746: out = 16'(2020);
			1747: out = 16'(1890);
			1748: out = 16'(1808);
			1749: out = 16'(1700);
			1750: out = 16'(1607);
			1751: out = 16'(1510);
			1752: out = 16'(1425);
			1753: out = 16'(1359);
			1754: out = 16'(1258);
			1755: out = 16'(1087);
			1756: out = 16'(867);
			1757: out = 16'(666);
			1758: out = 16'(486);
			1759: out = 16'(310);
			1760: out = 16'(135);
			1761: out = 16'(-10);
			1762: out = 16'(-173);
			1763: out = 16'(-325);
			1764: out = 16'(-460);
			1765: out = 16'(-576);
			1766: out = 16'(-725);
			1767: out = 16'(-849);
			1768: out = 16'(-967);
			1769: out = 16'(-1101);
			1770: out = 16'(-1222);
			1771: out = 16'(-1341);
			1772: out = 16'(-1469);
			1773: out = 16'(-1566);
			1774: out = 16'(-1716);
			1775: out = 16'(-1860);
			1776: out = 16'(-1990);
			1777: out = 16'(-2133);
			1778: out = 16'(-2282);
			1779: out = 16'(-2444);
			1780: out = 16'(-2614);
			1781: out = 16'(-2783);
			1782: out = 16'(-2987);
			1783: out = 16'(-3180);
			1784: out = 16'(-3415);
			1785: out = 16'(-3640);
			1786: out = 16'(-3880);
			1787: out = 16'(-4142);
			1788: out = 16'(-4374);
			1789: out = 16'(-4604);
			1790: out = 16'(-4836);
			1791: out = 16'(-5055);
			1792: out = 16'(-5261);
			1793: out = 16'(-5458);
			1794: out = 16'(-5639);
			1795: out = 16'(-5814);
			1796: out = 16'(-5974);
			1797: out = 16'(-6101);
			1798: out = 16'(-6230);
			1799: out = 16'(-6331);
			1800: out = 16'(-6427);
			1801: out = 16'(-6513);
			1802: out = 16'(-6569);
			1803: out = 16'(-6627);
			1804: out = 16'(-6666);
			1805: out = 16'(-6705);
			1806: out = 16'(-6748);
			1807: out = 16'(-6759);
			1808: out = 16'(-6775);
			1809: out = 16'(-6785);
			1810: out = 16'(-6782);
			1811: out = 16'(-6772);
			1812: out = 16'(-6744);
			1813: out = 16'(-6729);
			1814: out = 16'(-6700);
			1815: out = 16'(-6681);
			1816: out = 16'(-6639);
			1817: out = 16'(-6606);
			1818: out = 16'(-6572);
			1819: out = 16'(-6513);
			1820: out = 16'(-6474);
			1821: out = 16'(-6415);
			1822: out = 16'(-6374);
			1823: out = 16'(-6296);
			1824: out = 16'(-6234);
			1825: out = 16'(-6176);
			1826: out = 16'(-6096);
			1827: out = 16'(-6024);
			1828: out = 16'(-5941);
			1829: out = 16'(-5856);
			1830: out = 16'(-5745);
			1831: out = 16'(-5629);
			1832: out = 16'(-5511);
			1833: out = 16'(-5363);
			1834: out = 16'(-5212);
			1835: out = 16'(-5046);
			1836: out = 16'(-4889);
			1837: out = 16'(-4694);
			1838: out = 16'(-4512);
			1839: out = 16'(-4312);
			1840: out = 16'(-4131);
			1841: out = 16'(-3934);
			1842: out = 16'(-3754);
			1843: out = 16'(-3549);
			1844: out = 16'(-3388);
			1845: out = 16'(-3197);
			1846: out = 16'(-3035);
			1847: out = 16'(-2872);
			1848: out = 16'(-2707);
			1849: out = 16'(-2555);
			1850: out = 16'(-2398);
			1851: out = 16'(-2258);
			1852: out = 16'(-2129);
			1853: out = 16'(-1992);
			1854: out = 16'(-1862);
			1855: out = 16'(-1750);
			1856: out = 16'(-1627);
			1857: out = 16'(-1515);
			1858: out = 16'(-1426);
			1859: out = 16'(-1316);
			1860: out = 16'(-1219);
			1861: out = 16'(-1073);
			1862: out = 16'(-895);
			1863: out = 16'(-761);
			1864: out = 16'(-623);
			1865: out = 16'(-482);
			1866: out = 16'(-352);
			1867: out = 16'(-231);
			1868: out = 16'(-128);
			1869: out = 16'(-15);
			1870: out = 16'(79);
			1871: out = 16'(182);
			1872: out = 16'(288);
			1873: out = 16'(379);
			1874: out = 16'(470);
			1875: out = 16'(559);
			1876: out = 16'(644);
			1877: out = 16'(742);
			1878: out = 16'(834);
			1879: out = 16'(932);
			1880: out = 16'(1035);
			1881: out = 16'(1121);
			1882: out = 16'(1226);
			1883: out = 16'(1341);
			1884: out = 16'(1468);
			1885: out = 16'(1600);
			1886: out = 16'(1749);
			1887: out = 16'(1865);
			1888: out = 16'(2032);
			1889: out = 16'(2193);
			1890: out = 16'(2370);
			1891: out = 16'(2548);
			1892: out = 16'(2722);
			1893: out = 16'(2898);
			1894: out = 16'(3066);
			1895: out = 16'(3245);
			1896: out = 16'(3397);
			1897: out = 16'(3555);
			1898: out = 16'(3706);
			1899: out = 16'(3838);
			1900: out = 16'(3988);
			1901: out = 16'(4115);
			1902: out = 16'(4247);
			1903: out = 16'(4364);
			1904: out = 16'(4472);
			1905: out = 16'(4577);
			1906: out = 16'(4687);
			1907: out = 16'(4786);
			1908: out = 16'(4873);
			1909: out = 16'(4976);
			1910: out = 16'(5066);
			1911: out = 16'(5149);
			1912: out = 16'(5223);
			1913: out = 16'(5314);
			1914: out = 16'(5397);
			1915: out = 16'(5456);
			1916: out = 16'(5523);
			1917: out = 16'(5603);
			1918: out = 16'(5669);
			1919: out = 16'(5674);
			1920: out = 16'(5694);
			1921: out = 16'(5694);
			1922: out = 16'(5708);
			1923: out = 16'(5681);
			1924: out = 16'(5648);
			1925: out = 16'(5633);
			1926: out = 16'(5610);
			1927: out = 16'(5622);
			1928: out = 16'(5594);
			1929: out = 16'(5594);
			1930: out = 16'(5592);
			1931: out = 16'(5602);
			1932: out = 16'(5580);
			1933: out = 16'(5537);
			1934: out = 16'(5506);
			1935: out = 16'(5504);
			1936: out = 16'(5476);
			1937: out = 16'(5423);
			1938: out = 16'(5361);
			1939: out = 16'(5294);
			1940: out = 16'(5240);
			1941: out = 16'(5114);
			1942: out = 16'(5042);
			1943: out = 16'(4930);
			1944: out = 16'(4789);
			1945: out = 16'(4684);
			1946: out = 16'(4527);
			1947: out = 16'(4409);
			1948: out = 16'(4252);
			1949: out = 16'(4097);
			1950: out = 16'(3945);
			1951: out = 16'(3833);
			1952: out = 16'(3654);
			1953: out = 16'(3511);
			1954: out = 16'(3380);
			1955: out = 16'(3244);
			1956: out = 16'(3082);
			1957: out = 16'(2963);
			1958: out = 16'(2836);
			1959: out = 16'(2680);
			1960: out = 16'(2584);
			1961: out = 16'(2444);
			1962: out = 16'(2347);
			1963: out = 16'(2215);
			1964: out = 16'(2128);
			1965: out = 16'(2021);
			1966: out = 16'(1913);
			1967: out = 16'(1815);
			1968: out = 16'(1720);
			1969: out = 16'(1629);
			1970: out = 16'(1536);
			1971: out = 16'(1465);
			1972: out = 16'(1383);
			1973: out = 16'(1321);
			1974: out = 16'(1233);
			1975: out = 16'(1175);
			1976: out = 16'(1114);
			1977: out = 16'(1028);
			1978: out = 16'(843);
			1979: out = 16'(677);
			1980: out = 16'(529);
			1981: out = 16'(389);
			1982: out = 16'(225);
			1983: out = 16'(108);
			1984: out = 16'(-36);
			1985: out = 16'(-151);
			1986: out = 16'(-281);
			1987: out = 16'(-387);
			1988: out = 16'(-493);
			1989: out = 16'(-618);
			1990: out = 16'(-709);
			1991: out = 16'(-813);
			1992: out = 16'(-928);
			1993: out = 16'(-1016);
			1994: out = 16'(-1121);
			1995: out = 16'(-1226);
			1996: out = 16'(-1328);
			1997: out = 16'(-1438);
			1998: out = 16'(-1536);
			1999: out = 16'(-1659);
			2000: out = 16'(-1765);
			2001: out = 16'(-1900);
			2002: out = 16'(-2034);
			2003: out = 16'(-2196);
			2004: out = 16'(-2346);
			2005: out = 16'(-2501);
			2006: out = 16'(-2669);
			2007: out = 16'(-2860);
			2008: out = 16'(-3045);
			2009: out = 16'(-3255);
			2010: out = 16'(-3470);
			2011: out = 16'(-3666);
			2012: out = 16'(-3862);
			2013: out = 16'(-4062);
			2014: out = 16'(-4234);
			2015: out = 16'(-4393);
			2016: out = 16'(-4553);
			2017: out = 16'(-4713);
			2018: out = 16'(-4829);
			2019: out = 16'(-4956);
			2020: out = 16'(-5067);
			2021: out = 16'(-5160);
			2022: out = 16'(-5253);
			2023: out = 16'(-5328);
			2024: out = 16'(-5389);
			2025: out = 16'(-5425);
			2026: out = 16'(-5484);
			2027: out = 16'(-5500);
			2028: out = 16'(-5548);
			2029: out = 16'(-5562);
			2030: out = 16'(-5581);
			2031: out = 16'(-5577);
			2032: out = 16'(-5591);
			2033: out = 16'(-5580);
			2034: out = 16'(-5569);
			2035: out = 16'(-5563);
			2036: out = 16'(-5534);
			2037: out = 16'(-5517);
			2038: out = 16'(-5505);
			2039: out = 16'(-5453);
			2040: out = 16'(-5421);
			2041: out = 16'(-5398);
			2042: out = 16'(-5354);
			2043: out = 16'(-5314);
			2044: out = 16'(-5259);
			2045: out = 16'(-5204);
			2046: out = 16'(-5149);
			2047: out = 16'(-5090);
			2048: out = 16'(-5044);
			2049: out = 16'(-4982);
			2050: out = 16'(-4907);
			2051: out = 16'(-4842);
			2052: out = 16'(-4756);
			2053: out = 16'(-4673);
			2054: out = 16'(-4589);
			2055: out = 16'(-4487);
			2056: out = 16'(-4359);
			2057: out = 16'(-4250);
			2058: out = 16'(-4104);
			2059: out = 16'(-3954);
			2060: out = 16'(-3813);
			2061: out = 16'(-3652);
			2062: out = 16'(-3510);
			2063: out = 16'(-3335);
			2064: out = 16'(-3186);
			2065: out = 16'(-3027);
			2066: out = 16'(-2878);
			2067: out = 16'(-2722);
			2068: out = 16'(-2593);
			2069: out = 16'(-2446);
			2070: out = 16'(-2302);
			2071: out = 16'(-2188);
			2072: out = 16'(-2048);
			2073: out = 16'(-1931);
			2074: out = 16'(-1816);
			2075: out = 16'(-1703);
			2076: out = 16'(-1592);
			2077: out = 16'(-1495);
			2078: out = 16'(-1410);
			2079: out = 16'(-1300);
			2080: out = 16'(-1221);
			2081: out = 16'(-1131);
			2082: out = 16'(-1052);
			2083: out = 16'(-972);
			2084: out = 16'(-848);
			2085: out = 16'(-704);
			2086: out = 16'(-595);
			2087: out = 16'(-488);
			2088: out = 16'(-393);
			2089: out = 16'(-286);
			2090: out = 16'(-176);
			2091: out = 16'(-81);
			2092: out = 16'(-14);
			2093: out = 16'(75);
			2094: out = 16'(162);
			2095: out = 16'(231);
			2096: out = 16'(301);
			2097: out = 16'(395);
			2098: out = 16'(462);
			2099: out = 16'(538);
			2100: out = 16'(614);
			2101: out = 16'(685);
			2102: out = 16'(762);
			2103: out = 16'(836);
			2104: out = 16'(921);
			2105: out = 16'(1011);
			2106: out = 16'(1108);
			2107: out = 16'(1205);
			2108: out = 16'(1305);
			2109: out = 16'(1414);
			2110: out = 16'(1552);
			2111: out = 16'(1674);
			2112: out = 16'(1806);
			2113: out = 16'(1950);
			2114: out = 16'(2098);
			2115: out = 16'(2240);
			2116: out = 16'(2384);
			2117: out = 16'(2512);
			2118: out = 16'(2654);
			2119: out = 16'(2782);
			2120: out = 16'(2906);
			2121: out = 16'(3035);
			2122: out = 16'(3152);
			2123: out = 16'(3264);
			2124: out = 16'(3363);
			2125: out = 16'(3458);
			2126: out = 16'(3575);
			2127: out = 16'(3645);
			2128: out = 16'(3736);
			2129: out = 16'(3830);
			2130: out = 16'(3917);
			2131: out = 16'(3996);
			2132: out = 16'(4072);
			2133: out = 16'(4120);
			2134: out = 16'(4203);
			2135: out = 16'(4255);
			2136: out = 16'(4340);
			2137: out = 16'(4404);
			2138: out = 16'(4447);
			2139: out = 16'(4524);
			2140: out = 16'(4584);
			2141: out = 16'(4635);
			2142: out = 16'(4661);
			2143: out = 16'(4651);
			2144: out = 16'(4630);
			2145: out = 16'(4642);
			2146: out = 16'(4634);
			2147: out = 16'(4616);
			2148: out = 16'(4620);
			2149: out = 16'(4598);
			2150: out = 16'(4587);
			2151: out = 16'(4593);
			2152: out = 16'(4573);
			2153: out = 16'(4568);
			2154: out = 16'(4565);
			2155: out = 16'(4554);
			2156: out = 16'(4533);
			2157: out = 16'(4535);
			2158: out = 16'(4510);
			2159: out = 16'(4481);
			2160: out = 16'(4445);
			2161: out = 16'(4414);
			2162: out = 16'(4383);
			2163: out = 16'(4301);
			2164: out = 16'(4209);
			2165: out = 16'(4140);
			2166: out = 16'(4052);
			2167: out = 16'(3936);
			2168: out = 16'(3844);
			2169: out = 16'(3726);
			2170: out = 16'(3601);
			2171: out = 16'(3499);
			2172: out = 16'(3378);
			2173: out = 16'(3250);
			2174: out = 16'(3130);
			2175: out = 16'(3013);
			2176: out = 16'(2889);
			2177: out = 16'(2752);
			2178: out = 16'(2642);
			2179: out = 16'(2540);
			2180: out = 16'(2435);
			2181: out = 16'(2317);
			2182: out = 16'(2219);
			2183: out = 16'(2115);
			2184: out = 16'(2002);
			2185: out = 16'(1923);
			2186: out = 16'(1823);
			2187: out = 16'(1725);
			2188: out = 16'(1648);
			2189: out = 16'(1574);
			2190: out = 16'(1483);
			2191: out = 16'(1415);
			2192: out = 16'(1334);
			2193: out = 16'(1259);
			2194: out = 16'(1177);
			2195: out = 16'(1125);
			2196: out = 16'(1057);
			2197: out = 16'(1003);
			2198: out = 16'(948);
			2199: out = 16'(893);
			2200: out = 16'(811);
			2201: out = 16'(663);
			2202: out = 16'(535);
			2203: out = 16'(382);
			2204: out = 16'(270);
			2205: out = 16'(154);
			2206: out = 16'(37);
			2207: out = 16'(-70);
			2208: out = 16'(-156);
			2209: out = 16'(-257);
			2210: out = 16'(-356);
			2211: out = 16'(-439);
			2212: out = 16'(-529);
			2213: out = 16'(-621);
			2214: out = 16'(-707);
			2215: out = 16'(-798);
			2216: out = 16'(-872);
			2217: out = 16'(-959);
			2218: out = 16'(-1036);
			2219: out = 16'(-1116);
			2220: out = 16'(-1221);
			2221: out = 16'(-1306);
			2222: out = 16'(-1394);
			2223: out = 16'(-1505);
			2224: out = 16'(-1600);
			2225: out = 16'(-1717);
			2226: out = 16'(-1840);
			2227: out = 16'(-1969);
			2228: out = 16'(-2089);
			2229: out = 16'(-2230);
			2230: out = 16'(-2384);
			2231: out = 16'(-2557);
			2232: out = 16'(-2723);
			2233: out = 16'(-2885);
			2234: out = 16'(-3048);
			2235: out = 16'(-3214);
			2236: out = 16'(-3362);
			2237: out = 16'(-3499);
			2238: out = 16'(-3640);
			2239: out = 16'(-3779);
			2240: out = 16'(-3890);
			2241: out = 16'(-4010);
			2242: out = 16'(-4096);
			2243: out = 16'(-4178);
			2244: out = 16'(-4265);
			2245: out = 16'(-4343);
			2246: out = 16'(-4381);
			2247: out = 16'(-4434);
			2248: out = 16'(-4475);
			2249: out = 16'(-4513);
			2250: out = 16'(-4523);
			2251: out = 16'(-4559);
			2252: out = 16'(-4562);
			2253: out = 16'(-4575);
			2254: out = 16'(-4571);
			2255: out = 16'(-4590);
			2256: out = 16'(-4574);
			2257: out = 16'(-4554);
			2258: out = 16'(-4558);
			2259: out = 16'(-4531);
			2260: out = 16'(-4507);
			2261: out = 16'(-4491);
			2262: out = 16'(-4460);
			2263: out = 16'(-4435);
			2264: out = 16'(-4405);
			2265: out = 16'(-4370);
			2266: out = 16'(-4345);
			2267: out = 16'(-4289);
			2268: out = 16'(-4254);
			2269: out = 16'(-4205);
			2270: out = 16'(-4172);
			2271: out = 16'(-4117);
			2272: out = 16'(-4064);
			2273: out = 16'(-4010);
			2274: out = 16'(-3953);
			2275: out = 16'(-3886);
			2276: out = 16'(-3804);
			2277: out = 16'(-3731);
			2278: out = 16'(-3647);
			2279: out = 16'(-3549);
			2280: out = 16'(-3442);
			2281: out = 16'(-3324);
			2282: out = 16'(-3212);
			2283: out = 16'(-3094);
			2284: out = 16'(-2960);
			2285: out = 16'(-2836);
			2286: out = 16'(-2700);
			2287: out = 16'(-2571);
			2288: out = 16'(-2441);
			2289: out = 16'(-2333);
			2290: out = 16'(-2211);
			2291: out = 16'(-2091);
			2292: out = 16'(-1980);
			2293: out = 16'(-1862);
			2294: out = 16'(-1765);
			2295: out = 16'(-1650);
			2296: out = 16'(-1553);
			2297: out = 16'(-1466);
			2298: out = 16'(-1369);
			2299: out = 16'(-1298);
			2300: out = 16'(-1205);
			2301: out = 16'(-1131);
			2302: out = 16'(-1046);
			2303: out = 16'(-979);
			2304: out = 16'(-920);
			2305: out = 16'(-854);
			2306: out = 16'(-776);
			2307: out = 16'(-661);
			2308: out = 16'(-570);
			2309: out = 16'(-457);
			2310: out = 16'(-372);
			2311: out = 16'(-289);
			2312: out = 16'(-218);
			2313: out = 16'(-148);
			2314: out = 16'(-70);
			2315: out = 16'(5);
			2316: out = 16'(74);
			2317: out = 16'(134);
			2318: out = 16'(204);
			2319: out = 16'(252);
			2320: out = 16'(316);
			2321: out = 16'(372);
			2322: out = 16'(434);
			2323: out = 16'(502);
			2324: out = 16'(566);
			2325: out = 16'(622);
			2326: out = 16'(693);
			2327: out = 16'(755);
			2328: out = 16'(821);
			2329: out = 16'(901);
			2330: out = 16'(980);
			2331: out = 16'(1066);
			2332: out = 16'(1165);
			2333: out = 16'(1259);
			2334: out = 16'(1363);
			2335: out = 16'(1475);
			2336: out = 16'(1598);
			2337: out = 16'(1710);
			2338: out = 16'(1835);
			2339: out = 16'(1946);
			2340: out = 16'(2067);
			2341: out = 16'(2168);
			2342: out = 16'(2275);
			2343: out = 16'(2381);
			2344: out = 16'(2481);
			2345: out = 16'(2574);
			2346: out = 16'(2670);
			2347: out = 16'(2752);
			2348: out = 16'(2831);
			2349: out = 16'(2916);
			2350: out = 16'(2984);
			2351: out = 16'(3063);
			2352: out = 16'(3134);
			2353: out = 16'(3211);
			2354: out = 16'(3262);
			2355: out = 16'(3326);
			2356: out = 16'(3376);
			2357: out = 16'(3433);
			2358: out = 16'(3483);
			2359: out = 16'(3552);
			2360: out = 16'(3600);
			2361: out = 16'(3646);
			2362: out = 16'(3693);
			2363: out = 16'(3735);
			2364: out = 16'(3780);
			2365: out = 16'(3813);
			2366: out = 16'(3792);
			2367: out = 16'(3791);
			2368: out = 16'(3773);
			2369: out = 16'(3765);
			2370: out = 16'(3775);
			2371: out = 16'(3777);
			2372: out = 16'(3757);
			2373: out = 16'(3756);
			2374: out = 16'(3745);
			2375: out = 16'(3728);
			2376: out = 16'(3745);
			2377: out = 16'(3736);
			2378: out = 16'(3729);
			2379: out = 16'(3708);
			2380: out = 16'(3686);
			2381: out = 16'(3665);
			2382: out = 16'(3675);
			2383: out = 16'(3607);
			2384: out = 16'(3569);
			2385: out = 16'(3529);
			2386: out = 16'(3495);
			2387: out = 16'(3442);
			2388: out = 16'(3347);
			2389: out = 16'(3274);
			2390: out = 16'(3201);
			2391: out = 16'(3117);
			2392: out = 16'(3032);
			2393: out = 16'(2929);
			2394: out = 16'(2823);
			2395: out = 16'(2751);
			2396: out = 16'(2649);
			2397: out = 16'(2539);
			2398: out = 16'(2446);
			2399: out = 16'(2350);
			2400: out = 16'(2262);
			2401: out = 16'(2137);
			2402: out = 16'(2051);
			2403: out = 16'(1967);
			2404: out = 16'(1879);
			2405: out = 16'(1792);
			2406: out = 16'(1697);
			2407: out = 16'(1607);
			2408: out = 16'(1549);
			2409: out = 16'(1465);
			2410: out = 16'(1402);
			2411: out = 16'(1312);
			2412: out = 16'(1256);
			2413: out = 16'(1210);
			2414: out = 16'(1135);
			2415: out = 16'(1086);
			2416: out = 16'(1035);
			2417: out = 16'(974);
			2418: out = 16'(916);
			2419: out = 16'(862);
			2420: out = 16'(817);
			2421: out = 16'(778);
			2422: out = 16'(715);
			2423: out = 16'(646);
			2424: out = 16'(519);
			2425: out = 16'(409);
			2426: out = 16'(318);
			2427: out = 16'(222);
			2428: out = 16'(121);
			2429: out = 16'(16);
			2430: out = 16'(-62);
			2431: out = 16'(-137);
			2432: out = 16'(-237);
			2433: out = 16'(-301);
			2434: out = 16'(-384);
			2435: out = 16'(-456);
			2436: out = 16'(-522);
			2437: out = 16'(-592);
			2438: out = 16'(-664);
			2439: out = 16'(-722);
			2440: out = 16'(-793);
			2441: out = 16'(-859);
			2442: out = 16'(-938);
			2443: out = 16'(-1018);
			2444: out = 16'(-1085);
			2445: out = 16'(-1166);
			2446: out = 16'(-1234);
			2447: out = 16'(-1338);
			2448: out = 16'(-1425);
			2449: out = 16'(-1525);
			2450: out = 16'(-1637);
			2451: out = 16'(-1748);
			2452: out = 16'(-1872);
			2453: out = 16'(-1992);
			2454: out = 16'(-2110);
			2455: out = 16'(-2258);
			2456: out = 16'(-2400);
			2457: out = 16'(-2541);
			2458: out = 16'(-2658);
			2459: out = 16'(-2790);
			2460: out = 16'(-2907);
			2461: out = 16'(-3016);
			2462: out = 16'(-3123);
			2463: out = 16'(-3213);
			2464: out = 16'(-3298);
			2465: out = 16'(-3371);
			2466: out = 16'(-3448);
			2467: out = 16'(-3495);
			2468: out = 16'(-3559);
			2469: out = 16'(-3611);
			2470: out = 16'(-3640);
			2471: out = 16'(-3681);
			2472: out = 16'(-3698);
			2473: out = 16'(-3719);
			2474: out = 16'(-3734);
			2475: out = 16'(-3736);
			2476: out = 16'(-3747);
			2477: out = 16'(-3746);
			2478: out = 16'(-3741);
			2479: out = 16'(-3746);
			2480: out = 16'(-3731);
			2481: out = 16'(-3720);
			2482: out = 16'(-3707);
			2483: out = 16'(-3697);
			2484: out = 16'(-3666);
			2485: out = 16'(-3652);
			2486: out = 16'(-3636);
			2487: out = 16'(-3588);
			2488: out = 16'(-3568);
			2489: out = 16'(-3544);
			2490: out = 16'(-3501);
			2491: out = 16'(-3477);
			2492: out = 16'(-3435);
			2493: out = 16'(-3397);
			2494: out = 16'(-3352);
			2495: out = 16'(-3308);
			2496: out = 16'(-3278);
			2497: out = 16'(-3223);
			2498: out = 16'(-3160);
			2499: out = 16'(-3096);
			2500: out = 16'(-3030);
			2501: out = 16'(-2969);
			2502: out = 16'(-2882);
			2503: out = 16'(-2795);
			2504: out = 16'(-2710);
			2505: out = 16'(-2606);
			2506: out = 16'(-2507);
			2507: out = 16'(-2386);
			2508: out = 16'(-2294);
			2509: out = 16'(-2193);
			2510: out = 16'(-2085);
			2511: out = 16'(-1986);
			2512: out = 16'(-1874);
			2513: out = 16'(-1789);
			2514: out = 16'(-1690);
			2515: out = 16'(-1604);
			2516: out = 16'(-1505);
			2517: out = 16'(-1416);
			2518: out = 16'(-1344);
			2519: out = 16'(-1270);
			2520: out = 16'(-1188);
			2521: out = 16'(-1107);
			2522: out = 16'(-1038);
			2523: out = 16'(-968);
			2524: out = 16'(-917);
			2525: out = 16'(-854);
			2526: out = 16'(-789);
			2527: out = 16'(-735);
			2528: out = 16'(-682);
			2529: out = 16'(-608);
			2530: out = 16'(-531);
			2531: out = 16'(-457);
			2532: out = 16'(-373);
			2533: out = 16'(-303);
			2534: out = 16'(-233);
			2535: out = 16'(-166);
			2536: out = 16'(-104);
			2537: out = 16'(-57);
			2538: out = 16'(18);
			2539: out = 16'(72);
			2540: out = 16'(124);
			2541: out = 16'(168);
			2542: out = 16'(217);
			2543: out = 16'(267);
			2544: out = 16'(321);
			2545: out = 16'(371);
			2546: out = 16'(416);
			2547: out = 16'(470);
			2548: out = 16'(531);
			2549: out = 16'(577);
			2550: out = 16'(640);
			2551: out = 16'(692);
			2552: out = 16'(747);
			2553: out = 16'(824);
			2554: out = 16'(904);
			2555: out = 16'(986);
			2556: out = 16'(1057);
			2557: out = 16'(1132);
			2558: out = 16'(1241);
			2559: out = 16'(1327);
			2560: out = 16'(1426);
			2561: out = 16'(1503);
			2562: out = 16'(1608);
			2563: out = 16'(1696);
			2564: out = 16'(1794);
			2565: out = 16'(1871);
			2566: out = 16'(1954);
			2567: out = 16'(2030);
			2568: out = 16'(2102);
			2569: out = 16'(2175);
			2570: out = 16'(2257);
			2571: out = 16'(2315);
			2572: out = 16'(2386);
			2573: out = 16'(2446);
			2574: out = 16'(2502);
			2575: out = 16'(2554);
			2576: out = 16'(2614);
			2577: out = 16'(2646);
			2578: out = 16'(2710);
			2579: out = 16'(2750);
			2580: out = 16'(2815);
			2581: out = 16'(2846);
			2582: out = 16'(2892);
			2583: out = 16'(2936);
			2584: out = 16'(2983);
			2585: out = 16'(3009);
			2586: out = 16'(3047);
			2587: out = 16'(3075);
			2588: out = 16'(3095);
			2589: out = 16'(3069);
			2590: out = 16'(3079);
			2591: out = 16'(3054);
			2592: out = 16'(3052);
			2593: out = 16'(3047);
			2594: out = 16'(3038);
			2595: out = 16'(3050);
			2596: out = 16'(3054);
			2597: out = 16'(3044);
			2598: out = 16'(3052);
			2599: out = 16'(3052);
			2600: out = 16'(3013);
			2601: out = 16'(3038);
			2602: out = 16'(3004);
			2603: out = 16'(3026);
			2604: out = 16'(2972);
			2605: out = 16'(2951);
			2606: out = 16'(2938);
			2607: out = 16'(2923);
			2608: out = 16'(2867);
			2609: out = 16'(2823);
			2610: out = 16'(2763);
			2611: out = 16'(2715);
			2612: out = 16'(2660);
			2613: out = 16'(2581);
			2614: out = 16'(2516);
			2615: out = 16'(2430);
			2616: out = 16'(2350);
			2617: out = 16'(2264);
			2618: out = 16'(2198);
			2619: out = 16'(2119);
			2620: out = 16'(2034);
			2621: out = 16'(1960);
			2622: out = 16'(1883);
			2623: out = 16'(1802);
			2624: out = 16'(1722);
			2625: out = 16'(1639);
			2626: out = 16'(1577);
			2627: out = 16'(1493);
			2628: out = 16'(1433);
			2629: out = 16'(1361);
			2630: out = 16'(1294);
			2631: out = 16'(1250);
			2632: out = 16'(1158);
			2633: out = 16'(1115);
			2634: out = 16'(1058);
			2635: out = 16'(1010);
			2636: out = 16'(955);
			2637: out = 16'(904);
			2638: out = 16'(868);
			2639: out = 16'(820);
			2640: out = 16'(771);
			2641: out = 16'(736);
			2642: out = 16'(689);
			2643: out = 16'(642);
			2644: out = 16'(600);
			2645: out = 16'(567);
			2646: out = 16'(480);
			2647: out = 16'(385);
			2648: out = 16'(290);
			2649: out = 16'(220);
			2650: out = 16'(128);
			2651: out = 16'(42);
			2652: out = 16'(-43);
			2653: out = 16'(-100);
			2654: out = 16'(-161);
			2655: out = 16'(-227);
			2656: out = 16'(-280);
			2657: out = 16'(-339);
			2658: out = 16'(-399);
			2659: out = 16'(-448);
			2660: out = 16'(-519);
			2661: out = 16'(-578);
			2662: out = 16'(-626);
			2663: out = 16'(-692);
			2664: out = 16'(-741);
			2665: out = 16'(-797);
			2666: out = 16'(-872);
			2667: out = 16'(-927);
			2668: out = 16'(-988);
			2669: out = 16'(-1051);
			2670: out = 16'(-1134);
			2671: out = 16'(-1197);
			2672: out = 16'(-1279);
			2673: out = 16'(-1374);
			2674: out = 16'(-1466);
			2675: out = 16'(-1574);
			2676: out = 16'(-1688);
			2677: out = 16'(-1799);
			2678: out = 16'(-1897);
			2679: out = 16'(-2009);
			2680: out = 16'(-2125);
			2681: out = 16'(-2233);
			2682: out = 16'(-2312);
			2683: out = 16'(-2419);
			2684: out = 16'(-2517);
			2685: out = 16'(-2582);
			2686: out = 16'(-2661);
			2687: out = 16'(-2732);
			2688: out = 16'(-2796);
			2689: out = 16'(-2849);
			2690: out = 16'(-2885);
			2691: out = 16'(-2926);
			2692: out = 16'(-2969);
			2693: out = 16'(-3002);
			2694: out = 16'(-3009);
			2695: out = 16'(-3028);
			2696: out = 16'(-3046);
			2697: out = 16'(-3052);
			2698: out = 16'(-3072);
			2699: out = 16'(-3083);
			2700: out = 16'(-3068);
			2701: out = 16'(-3066);
			2702: out = 16'(-3063);
			2703: out = 16'(-3051);
			2704: out = 16'(-3033);
			2705: out = 16'(-3026);
			2706: out = 16'(-3009);
			2707: out = 16'(-2999);
			2708: out = 16'(-2978);
			2709: out = 16'(-2947);
			2710: out = 16'(-2923);
			2711: out = 16'(-2910);
			2712: out = 16'(-2868);
			2713: out = 16'(-2843);
			2714: out = 16'(-2822);
			2715: out = 16'(-2782);
			2716: out = 16'(-2760);
			2717: out = 16'(-2739);
			2718: out = 16'(-2694);
			2719: out = 16'(-2653);
			2720: out = 16'(-2599);
			2721: out = 16'(-2557);
			2722: out = 16'(-2506);
			2723: out = 16'(-2455);
			2724: out = 16'(-2389);
			2725: out = 16'(-2329);
			2726: out = 16'(-2243);
			2727: out = 16'(-2175);
			2728: out = 16'(-2089);
			2729: out = 16'(-2015);
			2730: out = 16'(-1921);
			2731: out = 16'(-1840);
			2732: out = 16'(-1754);
			2733: out = 16'(-1666);
			2734: out = 16'(-1575);
			2735: out = 16'(-1507);
			2736: out = 16'(-1422);
			2737: out = 16'(-1350);
			2738: out = 16'(-1264);
			2739: out = 16'(-1194);
			2740: out = 16'(-1146);
			2741: out = 16'(-1067);
			2742: out = 16'(-1013);
			2743: out = 16'(-943);
			2744: out = 16'(-892);
			2745: out = 16'(-839);
			2746: out = 16'(-780);
			2747: out = 16'(-734);
			2748: out = 16'(-673);
			2749: out = 16'(-640);
			2750: out = 16'(-589);
			2751: out = 16'(-552);
			2752: out = 16'(-478);
			2753: out = 16'(-408);
			2754: out = 16'(-353);
			2755: out = 16'(-277);
			2756: out = 16'(-230);
			2757: out = 16'(-181);
			2758: out = 16'(-110);
			2759: out = 16'(-79);
			2760: out = 16'(-26);
			2761: out = 16'(12);
			2762: out = 16'(56);
			2763: out = 16'(83);
			2764: out = 16'(140);
			2765: out = 16'(188);
			2766: out = 16'(222);
			2767: out = 16'(268);
			2768: out = 16'(309);
			2769: out = 16'(346);
			2770: out = 16'(388);
			2771: out = 16'(436);
			2772: out = 16'(475);
			2773: out = 16'(518);
			2774: out = 16'(566);
			2775: out = 16'(626);
			2776: out = 16'(682);
			2777: out = 16'(744);
			2778: out = 16'(802);
			2779: out = 16'(888);
			2780: out = 16'(948);
			2781: out = 16'(1038);
			2782: out = 16'(1101);
			2783: out = 16'(1182);
			2784: out = 16'(1251);
			2785: out = 16'(1344);
			2786: out = 16'(1401);
			2787: out = 16'(1476);
			2788: out = 16'(1542);
			2789: out = 16'(1611);
			2790: out = 16'(1675);
			2791: out = 16'(1738);
			2792: out = 16'(1802);
			2793: out = 16'(1844);
			2794: out = 16'(1915);
			2795: out = 16'(1955);
			2796: out = 16'(1991);
			2797: out = 16'(2041);
			2798: out = 16'(2089);
			2799: out = 16'(2124);
			2800: out = 16'(2172);
			2801: out = 16'(2216);
			2802: out = 16'(2254);
			2803: out = 16'(2301);
			2804: out = 16'(2333);
			2805: out = 16'(2363);
			2806: out = 16'(2401);
			2807: out = 16'(2420);
			2808: out = 16'(2452);
			2809: out = 16'(2487);
			2810: out = 16'(2492);
			2811: out = 16'(2507);
			2812: out = 16'(2483);
			2813: out = 16'(2491);
			2814: out = 16'(2490);
			2815: out = 16'(2494);
			2816: out = 16'(2469);
			2817: out = 16'(2480);
			2818: out = 16'(2459);
			2819: out = 16'(2480);
			2820: out = 16'(2491);
			2821: out = 16'(2491);
			2822: out = 16'(2477);
			2823: out = 16'(2483);
			2824: out = 16'(2436);
			2825: out = 16'(2430);
			2826: out = 16'(2440);
			2827: out = 16'(2410);
			2828: out = 16'(2400);
			2829: out = 16'(2352);
			2830: out = 16'(2339);
			2831: out = 16'(2314);
			2832: out = 16'(2279);
			2833: out = 16'(2215);
			2834: out = 16'(2175);
			2835: out = 16'(2137);
			2836: out = 16'(2079);
			2837: out = 16'(2005);
			2838: out = 16'(1938);
			2839: out = 16'(1883);
			2840: out = 16'(1819);
			2841: out = 16'(1750);
			2842: out = 16'(1693);
			2843: out = 16'(1625);
			2844: out = 16'(1565);
			2845: out = 16'(1492);
			2846: out = 16'(1422);
			2847: out = 16'(1369);
			2848: out = 16'(1311);
			2849: out = 16'(1248);
			2850: out = 16'(1193);
			2851: out = 16'(1134);
			2852: out = 16'(1083);
			2853: out = 16'(1031);
			2854: out = 16'(987);
			2855: out = 16'(936);
			2856: out = 16'(893);
			2857: out = 16'(838);
			2858: out = 16'(797);
			2859: out = 16'(751);
			2860: out = 16'(711);
			2861: out = 16'(671);
			2862: out = 16'(637);
			2863: out = 16'(597);
			2864: out = 16'(567);
			2865: out = 16'(531);
			2866: out = 16'(500);
			2867: out = 16'(466);
			2868: out = 16'(441);
			2869: out = 16'(345);
			2870: out = 16'(273);
			2871: out = 16'(197);
			2872: out = 16'(133);
			2873: out = 16'(67);
			2874: out = 16'(4);
			2875: out = 16'(-46);
			2876: out = 16'(-116);
			2877: out = 16'(-154);
			2878: out = 16'(-208);
			2879: out = 16'(-262);
			2880: out = 16'(-304);
			2881: out = 16'(-360);
			2882: out = 16'(-401);
			2883: out = 16'(-443);
			2884: out = 16'(-489);
			2885: out = 16'(-548);
			2886: out = 16'(-575);
			2887: out = 16'(-635);
			2888: out = 16'(-672);
			2889: out = 16'(-728);
			2890: out = 16'(-779);
			2891: out = 16'(-825);
			2892: out = 16'(-884);
			2893: out = 16'(-961);
			2894: out = 16'(-1012);
			2895: out = 16'(-1073);
			2896: out = 16'(-1167);
			2897: out = 16'(-1222);
			2898: out = 16'(-1316);
			2899: out = 16'(-1399);
			2900: out = 16'(-1497);
			2901: out = 16'(-1582);
			2902: out = 16'(-1675);
			2903: out = 16'(-1768);
			2904: out = 16'(-1843);
			2905: out = 16'(-1935);
			2906: out = 16'(-2008);
			2907: out = 16'(-2076);
			2908: out = 16'(-2132);
			2909: out = 16'(-2194);
			2910: out = 16'(-2245);
			2911: out = 16'(-2290);
			2912: out = 16'(-2333);
			2913: out = 16'(-2372);
			2914: out = 16'(-2393);
			2915: out = 16'(-2428);
			2916: out = 16'(-2442);
			2917: out = 16'(-2474);
			2918: out = 16'(-2480);
			2919: out = 16'(-2482);
			2920: out = 16'(-2499);
			2921: out = 16'(-2497);
			2922: out = 16'(-2511);
			2923: out = 16'(-2499);
			2924: out = 16'(-2491);
			2925: out = 16'(-2486);
			2926: out = 16'(-2481);
			2927: out = 16'(-2476);
			2928: out = 16'(-2464);
			2929: out = 16'(-2446);
			2930: out = 16'(-2434);
			2931: out = 16'(-2419);
			2932: out = 16'(-2405);
			2933: out = 16'(-2384);
			2934: out = 16'(-2359);
			2935: out = 16'(-2347);
			2936: out = 16'(-2330);
			2937: out = 16'(-2293);
			2938: out = 16'(-2270);
			2939: out = 16'(-2249);
			2940: out = 16'(-2218);
			2941: out = 16'(-2186);
			2942: out = 16'(-2156);
			2943: out = 16'(-2115);
			2944: out = 16'(-2083);
			2945: out = 16'(-2043);
			2946: out = 16'(-1984);
			2947: out = 16'(-1930);
			2948: out = 16'(-1876);
			2949: out = 16'(-1816);
			2950: out = 16'(-1754);
			2951: out = 16'(-1685);
			2952: out = 16'(-1618);
			2953: out = 16'(-1545);
			2954: out = 16'(-1475);
			2955: out = 16'(-1404);
			2956: out = 16'(-1338);
			2957: out = 16'(-1274);
			2958: out = 16'(-1210);
			2959: out = 16'(-1142);
			2960: out = 16'(-1082);
			2961: out = 16'(-1025);
			2962: out = 16'(-965);
			2963: out = 16'(-910);
			2964: out = 16'(-849);
			2965: out = 16'(-810);
			2966: out = 16'(-761);
			2967: out = 16'(-716);
			2968: out = 16'(-660);
			2969: out = 16'(-630);
			2970: out = 16'(-592);
			2971: out = 16'(-542);
			2972: out = 16'(-510);
			2973: out = 16'(-477);
			2974: out = 16'(-436);
			2975: out = 16'(-380);
			2976: out = 16'(-321);
			2977: out = 16'(-277);
			2978: out = 16'(-226);
			2979: out = 16'(-181);
			2980: out = 16'(-139);
			2981: out = 16'(-102);
			2982: out = 16'(-69);
			2983: out = 16'(-15);
			2984: out = 16'(15);
			2985: out = 16'(46);
			2986: out = 16'(90);
			2987: out = 16'(129);
			2988: out = 16'(151);
			2989: out = 16'(191);
			2990: out = 16'(223);
			2991: out = 16'(253);
			2992: out = 16'(282);
			2993: out = 16'(318);
			2994: out = 16'(359);
			2995: out = 16'(388);
			2996: out = 16'(429);
			2997: out = 16'(467);
			2998: out = 16'(510);
			2999: out = 16'(562);
			3000: out = 16'(613);
			3001: out = 16'(666);
			3002: out = 16'(724);
			3003: out = 16'(780);
			3004: out = 16'(836);
			3005: out = 16'(901);
			3006: out = 16'(960);
			3007: out = 16'(1024);
			3008: out = 16'(1081);
			3009: out = 16'(1156);
			3010: out = 16'(1200);
			3011: out = 16'(1261);
			3012: out = 16'(1312);
			3013: out = 16'(1366);
			3014: out = 16'(1405);
			3015: out = 16'(1452);
			3016: out = 16'(1500);
			3017: out = 16'(1527);
			3018: out = 16'(1586);
			3019: out = 16'(1625);
			3020: out = 16'(1661);
			3021: out = 16'(1690);
			3022: out = 16'(1734);
			3023: out = 16'(1768);
			3024: out = 16'(1791);
			3025: out = 16'(1828);
			3026: out = 16'(1856);
			3027: out = 16'(1886);
			3028: out = 16'(1912);
			3029: out = 16'(1937);
			3030: out = 16'(1977);
			3031: out = 16'(1991);
			3032: out = 16'(2007);
			3033: out = 16'(2027);
			3034: out = 16'(2026);
			3035: out = 16'(2022);
			3036: out = 16'(2017);
			3037: out = 16'(2013);
			3038: out = 16'(2008);
			3039: out = 16'(2009);
			3040: out = 16'(2002);
			3041: out = 16'(2009);
			3042: out = 16'(2009);
			3043: out = 16'(2000);
			3044: out = 16'(1985);
			3045: out = 16'(1986);
			3046: out = 16'(1994);
			3047: out = 16'(1980);
			3048: out = 16'(1969);
			3049: out = 16'(1958);
			3050: out = 16'(1942);
			3051: out = 16'(1924);
			3052: out = 16'(1909);
			3053: out = 16'(1890);
			3054: out = 16'(1856);
			3055: out = 16'(1832);
			3056: out = 16'(1800);
			3057: out = 16'(1745);
			3058: out = 16'(1701);
			3059: out = 16'(1664);
			3060: out = 16'(1613);
			3061: out = 16'(1566);
			3062: out = 16'(1513);
			3063: out = 16'(1462);
			3064: out = 16'(1395);
			3065: out = 16'(1353);
			3066: out = 16'(1299);
			3067: out = 16'(1247);
			3068: out = 16'(1184);
			3069: out = 16'(1142);
			3070: out = 16'(1105);
			3071: out = 16'(1048);
			3072: out = 16'(999);
			3073: out = 16'(944);
			3074: out = 16'(909);
			3075: out = 16'(872);
			3076: out = 16'(830);
			3077: out = 16'(784);
			3078: out = 16'(741);
			3079: out = 16'(706);
			3080: out = 16'(672);
			3081: out = 16'(642);
			3082: out = 16'(605);
			3083: out = 16'(572);
			3084: out = 16'(529);
			3085: out = 16'(515);
			3086: out = 16'(481);
			3087: out = 16'(463);
			3088: out = 16'(442);
			3089: out = 16'(393);
			3090: out = 16'(369);
			3091: out = 16'(332);
			3092: out = 16'(262);
			3093: out = 16'(199);
			3094: out = 16'(156);
			3095: out = 16'(89);
			3096: out = 16'(49);
			3097: out = 16'(-15);
			3098: out = 16'(-52);
			3099: out = 16'(-89);
			3100: out = 16'(-147);
			3101: out = 16'(-192);
			3102: out = 16'(-218);
			3103: out = 16'(-263);
			3104: out = 16'(-299);
			3105: out = 16'(-336);
			3106: out = 16'(-379);
			3107: out = 16'(-417);
			3108: out = 16'(-463);
			3109: out = 16'(-502);
			3110: out = 16'(-526);
			3111: out = 16'(-572);
			3112: out = 16'(-610);
			3113: out = 16'(-655);
			3114: out = 16'(-694);
			3115: out = 16'(-748);
			3116: out = 16'(-795);
			3117: out = 16'(-845);
			3118: out = 16'(-917);
			3119: out = 16'(-978);
			3120: out = 16'(-1033);
			3121: out = 16'(-1090);
			3122: out = 16'(-1188);
			3123: out = 16'(-1252);
			3124: out = 16'(-1312);
			3125: out = 16'(-1389);
			3126: out = 16'(-1459);
			3127: out = 16'(-1529);
			3128: out = 16'(-1599);
			3129: out = 16'(-1654);
			3130: out = 16'(-1709);
			3131: out = 16'(-1761);
			3132: out = 16'(-1802);
			3133: out = 16'(-1835);
			3134: out = 16'(-1880);
			3135: out = 16'(-1910);
			3136: out = 16'(-1945);
			3137: out = 16'(-1960);
			3138: out = 16'(-1994);
			3139: out = 16'(-1992);
			3140: out = 16'(-2017);
			3141: out = 16'(-2022);
			3142: out = 16'(-2024);
			3143: out = 16'(-2041);
			3144: out = 16'(-2040);
			3145: out = 16'(-2041);
			3146: out = 16'(-2039);
			3147: out = 16'(-2031);
			3148: out = 16'(-2031);
			3149: out = 16'(-2021);
			3150: out = 16'(-2025);
			3151: out = 16'(-1995);
			3152: out = 16'(-1991);
			3153: out = 16'(-1983);
			3154: out = 16'(-1963);
			3155: out = 16'(-1946);
			3156: out = 16'(-1936);
			3157: out = 16'(-1915);
			3158: out = 16'(-1898);
			3159: out = 16'(-1885);
			3160: out = 16'(-1861);
			3161: out = 16'(-1847);
			3162: out = 16'(-1819);
			3163: out = 16'(-1795);
			3164: out = 16'(-1768);
			3165: out = 16'(-1748);
			3166: out = 16'(-1716);
			3167: out = 16'(-1679);
			3168: out = 16'(-1642);
			3169: out = 16'(-1608);
			3170: out = 16'(-1563);
			3171: out = 16'(-1513);
			3172: out = 16'(-1471);
			3173: out = 16'(-1406);
			3174: out = 16'(-1351);
			3175: out = 16'(-1299);
			3176: out = 16'(-1246);
			3177: out = 16'(-1187);
			3178: out = 16'(-1133);
			3179: out = 16'(-1081);
			3180: out = 16'(-1021);
			3181: out = 16'(-973);
			3182: out = 16'(-917);
			3183: out = 16'(-880);
			3184: out = 16'(-825);
			3185: out = 16'(-784);
			3186: out = 16'(-738);
			3187: out = 16'(-699);
			3188: out = 16'(-656);
			3189: out = 16'(-606);
			3190: out = 16'(-587);
			3191: out = 16'(-534);
			3192: out = 16'(-502);
			3193: out = 16'(-468);
			3194: out = 16'(-440);
			3195: out = 16'(-413);
			3196: out = 16'(-374);
			3197: out = 16'(-349);
			3198: out = 16'(-310);
			3199: out = 16'(-263);
			3200: out = 16'(-221);
			3201: out = 16'(-183);
			3202: out = 16'(-141);
			3203: out = 16'(-110);
			3204: out = 16'(-69);
			3205: out = 16'(-44);
			3206: out = 16'(-15);
			3207: out = 16'(19);
			3208: out = 16'(36);
			3209: out = 16'(76);
			3210: out = 16'(101);
			3211: out = 16'(120);
			3212: out = 16'(148);
			3213: out = 16'(184);
			3214: out = 16'(204);
			3215: out = 16'(239);
			3216: out = 16'(257);
			3217: out = 16'(283);
			3218: out = 16'(316);
			3219: out = 16'(349);
			3220: out = 16'(381);
			3221: out = 16'(408);
			3222: out = 16'(444);
			3223: out = 16'(493);
			3224: out = 16'(538);
			3225: out = 16'(589);
			3226: out = 16'(644);
			3227: out = 16'(684);
			3228: out = 16'(734);
			3229: out = 16'(793);
			3230: out = 16'(831);
			3231: out = 16'(894);
			3232: out = 16'(943);
			3233: out = 16'(993);
			3234: out = 16'(1028);
			3235: out = 16'(1071);
			3236: out = 16'(1096);
			3237: out = 16'(1144);
			3238: out = 16'(1188);
			3239: out = 16'(1219);
			3240: out = 16'(1249);
			3241: out = 16'(1284);
			3242: out = 16'(1309);
			3243: out = 16'(1348);
			3244: out = 16'(1376);
			3245: out = 16'(1403);
			3246: out = 16'(1422);
			3247: out = 16'(1449);
			3248: out = 16'(1481);
			3249: out = 16'(1503);
			3250: out = 16'(1520);
			3251: out = 16'(1543);
			3252: out = 16'(1575);
			3253: out = 16'(1591);
			3254: out = 16'(1614);
			3255: out = 16'(1620);
			3256: out = 16'(1628);
			3257: out = 16'(1627);
			3258: out = 16'(1634);
			3259: out = 16'(1604);
			3260: out = 16'(1618);
			3261: out = 16'(1620);
			3262: out = 16'(1622);
			3263: out = 16'(1623);
			3264: out = 16'(1612);
			3265: out = 16'(1618);
			3266: out = 16'(1618);
			3267: out = 16'(1611);
			3268: out = 16'(1607);
			3269: out = 16'(1599);
			3270: out = 16'(1607);
			3271: out = 16'(1576);
			3272: out = 16'(1581);
			3273: out = 16'(1570);
			3274: out = 16'(1566);
			3275: out = 16'(1548);
			3276: out = 16'(1518);
			3277: out = 16'(1500);
			3278: out = 16'(1478);
			3279: out = 16'(1435);
			3280: out = 16'(1410);
			3281: out = 16'(1364);
			3282: out = 16'(1332);
			3283: out = 16'(1294);
			3284: out = 16'(1244);
			3285: out = 16'(1204);
			3286: out = 16'(1157);
			3287: out = 16'(1119);
			3288: out = 16'(1059);
			3289: out = 16'(1023);
			3290: out = 16'(989);
			3291: out = 16'(953);
			3292: out = 16'(890);
			3293: out = 16'(862);
			3294: out = 16'(826);
			3295: out = 16'(782);
			3296: out = 16'(738);
			3297: out = 16'(700);
			3298: out = 16'(676);
			3299: out = 16'(634);
			3300: out = 16'(611);
			3301: out = 16'(590);
			3302: out = 16'(552);
			3303: out = 16'(521);
			3304: out = 16'(490);
			3305: out = 16'(458);
			3306: out = 16'(435);
			3307: out = 16'(411);
			3308: out = 16'(392);
			3309: out = 16'(364);
			3310: out = 16'(327);
			3311: out = 16'(309);
			3312: out = 16'(305);
			3313: out = 16'(287);
			3314: out = 16'(226);
			3315: out = 16'(192);
			3316: out = 16'(149);
			3317: out = 16'(87);
			3318: out = 16'(62);
			3319: out = 16'(5);
			3320: out = 16'(-28);
			3321: out = 16'(-64);
			3322: out = 16'(-113);
			3323: out = 16'(-138);
			3324: out = 16'(-169);
			3325: out = 16'(-206);
			3326: out = 16'(-239);
			3327: out = 16'(-270);
			3328: out = 16'(-299);
			3329: out = 16'(-330);
			3330: out = 16'(-351);
			3331: out = 16'(-391);
			3332: out = 16'(-415);
			3333: out = 16'(-445);
			3334: out = 16'(-471);
			3335: out = 16'(-506);
			3336: out = 16'(-553);
			3337: out = 16'(-577);
			3338: out = 16'(-618);
			3339: out = 16'(-663);
			3340: out = 16'(-707);
			3341: out = 16'(-755);
			3342: out = 16'(-795);
			3343: out = 16'(-839);
			3344: out = 16'(-910);
			3345: out = 16'(-971);
			3346: out = 16'(-1035);
			3347: out = 16'(-1085);
			3348: out = 16'(-1134);
			3349: out = 16'(-1197);
			3350: out = 16'(-1245);
			3351: out = 16'(-1306);
			3352: out = 16'(-1358);
			3353: out = 16'(-1395);
			3354: out = 16'(-1438);
			3355: out = 16'(-1463);
			3356: out = 16'(-1504);
			3357: out = 16'(-1532);
			3358: out = 16'(-1551);
			3359: out = 16'(-1577);
			3360: out = 16'(-1592);
			3361: out = 16'(-1608);
			3362: out = 16'(-1630);
			3363: out = 16'(-1638);
			3364: out = 16'(-1637);
			3365: out = 16'(-1643);
			3366: out = 16'(-1654);
			3367: out = 16'(-1647);
			3368: out = 16'(-1648);
			3369: out = 16'(-1653);
			3370: out = 16'(-1650);
			3371: out = 16'(-1637);
			3372: out = 16'(-1638);
			3373: out = 16'(-1624);
			3374: out = 16'(-1615);
			3375: out = 16'(-1618);
			3376: out = 16'(-1603);
			3377: out = 16'(-1590);
			3378: out = 16'(-1574);
			3379: out = 16'(-1567);
			3380: out = 16'(-1560);
			3381: out = 16'(-1535);
			3382: out = 16'(-1513);
			3383: out = 16'(-1504);
			3384: out = 16'(-1486);
			3385: out = 16'(-1469);
			3386: out = 16'(-1454);
			3387: out = 16'(-1437);
			3388: out = 16'(-1415);
			3389: out = 16'(-1391);
			3390: out = 16'(-1354);
			3391: out = 16'(-1329);
			3392: out = 16'(-1298);
			3393: out = 16'(-1263);
			3394: out = 16'(-1216);
			3395: out = 16'(-1182);
			3396: out = 16'(-1143);
			3397: out = 16'(-1099);
			3398: out = 16'(-1046);
			3399: out = 16'(-1003);
			3400: out = 16'(-962);
			3401: out = 16'(-904);
			3402: out = 16'(-868);
			3403: out = 16'(-819);
			3404: out = 16'(-778);
			3405: out = 16'(-743);
			3406: out = 16'(-695);
			3407: out = 16'(-665);
			3408: out = 16'(-634);
			3409: out = 16'(-595);
			3410: out = 16'(-555);
			3411: out = 16'(-517);
			3412: out = 16'(-499);
			3413: out = 16'(-454);
			3414: out = 16'(-438);
			3415: out = 16'(-421);
			3416: out = 16'(-386);
			3417: out = 16'(-351);
			3418: out = 16'(-334);
			3419: out = 16'(-304);
			3420: out = 16'(-281);
			3421: out = 16'(-247);
			3422: out = 16'(-209);
			3423: out = 16'(-178);
			3424: out = 16'(-146);
			3425: out = 16'(-114);
			3426: out = 16'(-89);
			3427: out = 16'(-56);
			3428: out = 16'(-42);
			3429: out = 16'(-10);
			3430: out = 16'(-5);
			3431: out = 16'(27);
			3432: out = 16'(57);
			3433: out = 16'(74);
			3434: out = 16'(100);
			3435: out = 16'(113);
			3436: out = 16'(139);
			3437: out = 16'(164);
			3438: out = 16'(194);
			3439: out = 16'(206);
			3440: out = 16'(230);
			3441: out = 16'(257);
			3442: out = 16'(264);
			3443: out = 16'(306);
			3444: out = 16'(348);
			3445: out = 16'(375);
			3446: out = 16'(410);
			3447: out = 16'(442);
			3448: out = 16'(472);
			3449: out = 16'(517);
			3450: out = 16'(557);
			3451: out = 16'(595);
			3452: out = 16'(640);
			3453: out = 16'(680);
			3454: out = 16'(726);
			3455: out = 16'(752);
			3456: out = 16'(786);
			3457: out = 16'(819);
			3458: out = 16'(860);
			3459: out = 16'(890);
			3460: out = 16'(938);
			3461: out = 16'(959);
			3462: out = 16'(976);
			3463: out = 16'(1010);
			3464: out = 16'(1035);
			3465: out = 16'(1059);
			3466: out = 16'(1085);
			3467: out = 16'(1101);
			3468: out = 16'(1130);
			3469: out = 16'(1150);
			3470: out = 16'(1168);
			3471: out = 16'(1198);
			3472: out = 16'(1211);
			3473: out = 16'(1225);
			3474: out = 16'(1246);
			3475: out = 16'(1247);
			3476: out = 16'(1286);
			3477: out = 16'(1283);
			3478: out = 16'(1311);
			3479: out = 16'(1315);
			3480: out = 16'(1305);
			3481: out = 16'(1311);
			3482: out = 16'(1308);
			3483: out = 16'(1292);
			3484: out = 16'(1292);
			3485: out = 16'(1297);
			3486: out = 16'(1284);
			3487: out = 16'(1298);
			3488: out = 16'(1279);
			3489: out = 16'(1288);
			3490: out = 16'(1286);
			3491: out = 16'(1285);
			3492: out = 16'(1276);
			3493: out = 16'(1274);
			3494: out = 16'(1249);
			3495: out = 16'(1253);
			3496: out = 16'(1247);
			3497: out = 16'(1243);
			3498: out = 16'(1214);
			3499: out = 16'(1194);
			3500: out = 16'(1190);
			3501: out = 16'(1170);
			3502: out = 16'(1149);
			3503: out = 16'(1117);
			3504: out = 16'(1083);
			3505: out = 16'(1047);
			3506: out = 16'(1021);
			3507: out = 16'(974);
			3508: out = 16'(945);
			3509: out = 16'(912);
			3510: out = 16'(880);
			3511: out = 16'(838);
			3512: out = 16'(818);
			3513: out = 16'(772);
			3514: out = 16'(728);
			3515: out = 16'(702);
			3516: out = 16'(681);
			3517: out = 16'(642);
			3518: out = 16'(618);
			3519: out = 16'(597);
			3520: out = 16'(560);
			3521: out = 16'(533);
			3522: out = 16'(504);
			3523: out = 16'(479);
			3524: out = 16'(442);
			3525: out = 16'(430);
			3526: out = 16'(410);
			3527: out = 16'(375);
			3528: out = 16'(358);
			3529: out = 16'(340);
			3530: out = 16'(318);
			3531: out = 16'(303);
			3532: out = 16'(287);
			3533: out = 16'(267);
			3534: out = 16'(245);
			3535: out = 16'(228);
			3536: out = 16'(208);
			3537: out = 16'(174);
			3538: out = 16'(128);
			3539: out = 16'(88);
			3540: out = 16'(46);
			3541: out = 16'(17);
			3542: out = 16'(-13);
			3543: out = 16'(-41);
			3544: out = 16'(-72);
			3545: out = 16'(-93);
			3546: out = 16'(-126);
			3547: out = 16'(-166);
			3548: out = 16'(-174);
			3549: out = 16'(-206);
			3550: out = 16'(-227);
			3551: out = 16'(-252);
			3552: out = 16'(-280);
			3553: out = 16'(-304);
			3554: out = 16'(-334);
			3555: out = 16'(-341);
			3556: out = 16'(-373);
			3557: out = 16'(-410);
			3558: out = 16'(-420);
			3559: out = 16'(-453);
			3560: out = 16'(-480);
			3561: out = 16'(-509);
			3562: out = 16'(-552);
			3563: out = 16'(-585);
			3564: out = 16'(-632);
			3565: out = 16'(-671);
			3566: out = 16'(-717);
			3567: out = 16'(-761);
			3568: out = 16'(-814);
			3569: out = 16'(-856);
			3570: out = 16'(-902);
			3571: out = 16'(-952);
			3572: out = 16'(-991);
			3573: out = 16'(-1038);
			3574: out = 16'(-1074);
			3575: out = 16'(-1105);
			3576: out = 16'(-1146);
			3577: out = 16'(-1177);
			3578: out = 16'(-1197);
			3579: out = 16'(-1227);
			3580: out = 16'(-1241);
			3581: out = 16'(-1261);
			3582: out = 16'(-1270);
			3583: out = 16'(-1288);
			3584: out = 16'(-1304);
			3585: out = 16'(-1316);
			3586: out = 16'(-1331);
			3587: out = 16'(-1341);
			3588: out = 16'(-1336);
			3589: out = 16'(-1342);
			3590: out = 16'(-1343);
			3591: out = 16'(-1329);
			3592: out = 16'(-1331);
			3593: out = 16'(-1327);
			3594: out = 16'(-1320);
			3595: out = 16'(-1319);
			3596: out = 16'(-1321);
			3597: out = 16'(-1308);
			3598: out = 16'(-1303);
			3599: out = 16'(-1294);
			3600: out = 16'(-1271);
			3601: out = 16'(-1263);
			3602: out = 16'(-1255);
			3603: out = 16'(-1247);
			3604: out = 16'(-1239);
			3605: out = 16'(-1226);
			3606: out = 16'(-1219);
			3607: out = 16'(-1201);
			3608: out = 16'(-1179);
			3609: out = 16'(-1166);
			3610: out = 16'(-1157);
			3611: out = 16'(-1137);
			3612: out = 16'(-1118);
			3613: out = 16'(-1086);
			3614: out = 16'(-1074);
			3615: out = 16'(-1044);
			3616: out = 16'(-1011);
			3617: out = 16'(-983);
			3618: out = 16'(-952);
			3619: out = 16'(-919);
			3620: out = 16'(-876);
			3621: out = 16'(-839);
			3622: out = 16'(-802);
			3623: out = 16'(-767);
			3624: out = 16'(-728);
			3625: out = 16'(-704);
			3626: out = 16'(-667);
			3627: out = 16'(-635);
			3628: out = 16'(-598);
			3629: out = 16'(-546);
			3630: out = 16'(-528);
			3631: out = 16'(-504);
			3632: out = 16'(-472);
			3633: out = 16'(-438);
			3634: out = 16'(-412);
			3635: out = 16'(-398);
			3636: out = 16'(-371);
			3637: out = 16'(-342);
			3638: out = 16'(-335);
			3639: out = 16'(-305);
			3640: out = 16'(-281);
			3641: out = 16'(-273);
			3642: out = 16'(-253);
			3643: out = 16'(-223);
			3644: out = 16'(-207);
			3645: out = 16'(-169);
			3646: out = 16'(-144);
			3647: out = 16'(-114);
			3648: out = 16'(-95);
			3649: out = 16'(-69);
			3650: out = 16'(-45);
			3651: out = 16'(-36);
			3652: out = 16'(-10);
			3653: out = 16'(-4);
			3654: out = 16'(27);
			3655: out = 16'(38);
			3656: out = 16'(61);
			3657: out = 16'(87);
			3658: out = 16'(85);
			3659: out = 16'(101);
			3660: out = 16'(128);
			3661: out = 16'(147);
			3662: out = 16'(172);
			3663: out = 16'(182);
			3664: out = 16'(194);
			3665: out = 16'(218);
			3666: out = 16'(247);
			3667: out = 16'(264);
			3668: out = 16'(289);
			3669: out = 16'(321);
			3670: out = 16'(346);
			3671: out = 16'(391);
			3672: out = 16'(418);
			3673: out = 16'(440);
			3674: out = 16'(469);
			3675: out = 16'(510);
			3676: out = 16'(536);
			3677: out = 16'(566);
			3678: out = 16'(610);
			3679: out = 16'(625);
			3680: out = 16'(661);
			3681: out = 16'(681);
			3682: out = 16'(716);
			3683: out = 16'(740);
			3684: out = 16'(771);
			3685: out = 16'(787);
			3686: out = 16'(806);
			3687: out = 16'(829);
			3688: out = 16'(849);
			3689: out = 16'(855);
			3690: out = 16'(878);
			3691: out = 16'(897);
			3692: out = 16'(913);
			3693: out = 16'(925);
			3694: out = 16'(944);
			3695: out = 16'(964);
			3696: out = 16'(973);
			3697: out = 16'(984);
			3698: out = 16'(995);
			3699: out = 16'(1020);
			3700: out = 16'(1039);
			3701: out = 16'(1038);
			3702: out = 16'(1045);
			3703: out = 16'(1038);
			3704: out = 16'(1040);
			3705: out = 16'(1035);
			3706: out = 16'(1035);
			3707: out = 16'(1018);
			3708: out = 16'(1031);
			3709: out = 16'(1019);
			3710: out = 16'(1032);
			3711: out = 16'(1018);
			3712: out = 16'(1023);
			3713: out = 16'(1026);
			3714: out = 16'(1015);
			3715: out = 16'(1022);
			3716: out = 16'(1007);
			3717: out = 16'(1002);
			3718: out = 16'(1002);
			3719: out = 16'(989);
			3720: out = 16'(987);
			3721: out = 16'(979);
			3722: out = 16'(950);
			3723: out = 16'(947);
			3724: out = 16'(927);
			3725: out = 16'(904);
			3726: out = 16'(878);
			3727: out = 16'(850);
			3728: out = 16'(831);
			3729: out = 16'(796);
			3730: out = 16'(774);
			3731: out = 16'(744);
			3732: out = 16'(720);
			3733: out = 16'(699);
			3734: out = 16'(655);
			3735: out = 16'(630);
			3736: out = 16'(614);
			3737: out = 16'(576);
			3738: out = 16'(550);
			3739: out = 16'(537);
			3740: out = 16'(502);
			3741: out = 16'(456);
			3742: out = 16'(459);
			3743: out = 16'(434);
			3744: out = 16'(412);
			3745: out = 16'(379);
			3746: out = 16'(363);
			3747: out = 16'(349);
			3748: out = 16'(330);
			3749: out = 16'(316);
			3750: out = 16'(289);
			3751: out = 16'(269);
			3752: out = 16'(259);
			3753: out = 16'(242);
			3754: out = 16'(219);
			3755: out = 16'(210);
			3756: out = 16'(198);
			3757: out = 16'(186);
			3758: out = 16'(167);
			3759: out = 16'(157);
			3760: out = 16'(128);
			3761: out = 16'(88);
			3762: out = 16'(63);
			3763: out = 16'(38);
			3764: out = 16'(9);
			3765: out = 16'(-18);
			3766: out = 16'(-57);
			3767: out = 16'(-65);
			3768: out = 16'(-99);
			3769: out = 16'(-115);
			3770: out = 16'(-140);
			3771: out = 16'(-162);
			3772: out = 16'(-174);
			3773: out = 16'(-206);
			3774: out = 16'(-209);
			3775: out = 16'(-238);
			3776: out = 16'(-239);
			3777: out = 16'(-269);
			3778: out = 16'(-291);
			3779: out = 16'(-305);
			3780: out = 16'(-327);
			3781: out = 16'(-356);
			3782: out = 16'(-380);
			3783: out = 16'(-410);
			3784: out = 16'(-424);
			3785: out = 16'(-447);
			3786: out = 16'(-492);
			3787: out = 16'(-516);
			3788: out = 16'(-547);
			3789: out = 16'(-583);
			3790: out = 16'(-621);
			3791: out = 16'(-673);
			3792: out = 16'(-701);
			3793: out = 16'(-752);
			3794: out = 16'(-770);
			3795: out = 16'(-805);
			3796: out = 16'(-838);
			3797: out = 16'(-866);
			3798: out = 16'(-896);
			3799: out = 16'(-927);
			3800: out = 16'(-948);
			3801: out = 16'(-969);
			3802: out = 16'(-995);
			3803: out = 16'(-1016);
			3804: out = 16'(-1010);
			3805: out = 16'(-1044);
			3806: out = 16'(-1040);
			3807: out = 16'(-1050);
			3808: out = 16'(-1056);
			3809: out = 16'(-1072);
			3810: out = 16'(-1075);
			3811: out = 16'(-1075);
			3812: out = 16'(-1074);
			3813: out = 16'(-1077);
			3814: out = 16'(-1072);
			3815: out = 16'(-1083);
			3816: out = 16'(-1067);
			3817: out = 16'(-1066);
			3818: out = 16'(-1063);
			3819: out = 16'(-1061);
			3820: out = 16'(-1044);
			3821: out = 16'(-1045);
			3822: out = 16'(-1033);
			3823: out = 16'(-1032);
			3824: out = 16'(-1019);
			3825: out = 16'(-1019);
			3826: out = 16'(-1013);
			3827: out = 16'(-996);
			3828: out = 16'(-991);
			3829: out = 16'(-979);
			3830: out = 16'(-974);
			3831: out = 16'(-944);
			3832: out = 16'(-945);
			3833: out = 16'(-930);
			3834: out = 16'(-913);
			3835: out = 16'(-898);
			3836: out = 16'(-881);
			3837: out = 16'(-851);
			3838: out = 16'(-836);
			3839: out = 16'(-801);
			3840: out = 16'(-779);
			3841: out = 16'(-763);
			3842: out = 16'(-720);
			3843: out = 16'(-711);
			3844: out = 16'(-675);
			3845: out = 16'(-647);
			3846: out = 16'(-612);
			3847: out = 16'(-588);
			3848: out = 16'(-562);
			3849: out = 16'(-531);
			3850: out = 16'(-499);
			3851: out = 16'(-472);
			3852: out = 16'(-448);
			3853: out = 16'(-434);
			3854: out = 16'(-411);
			3855: out = 16'(-386);
			3856: out = 16'(-357);
			3857: out = 16'(-339);
			3858: out = 16'(-322);
			3859: out = 16'(-298);
			3860: out = 16'(-286);
			3861: out = 16'(-270);
			3862: out = 16'(-257);
			3863: out = 16'(-234);
			3864: out = 16'(-222);
			3865: out = 16'(-209);
			3866: out = 16'(-190);
			3867: out = 16'(-163);
			3868: out = 16'(-131);
			3869: out = 16'(-111);
			3870: out = 16'(-97);
			3871: out = 16'(-85);
			3872: out = 16'(-74);
			3873: out = 16'(-41);
			3874: out = 16'(-20);
			3875: out = 16'(-16);
			3876: out = 16'(7);
			3877: out = 16'(20);
			3878: out = 16'(27);
			3879: out = 16'(41);
			3880: out = 16'(54);
			3881: out = 16'(68);
			3882: out = 16'(87);
			3883: out = 16'(103);
			3884: out = 16'(117);
			3885: out = 16'(128);
			3886: out = 16'(136);
			3887: out = 16'(171);
			3888: out = 16'(188);
			3889: out = 16'(208);
			3890: out = 16'(220);
			3891: out = 16'(237);
			3892: out = 16'(261);
			3893: out = 16'(281);
			3894: out = 16'(298);
			3895: out = 16'(332);
			3896: out = 16'(372);
			3897: out = 16'(397);
			3898: out = 16'(420);
			3899: out = 16'(443);
			3900: out = 16'(459);
			3901: out = 16'(490);
			3902: out = 16'(517);
			3903: out = 16'(529);
			3904: out = 16'(545);
			3905: out = 16'(560);
			3906: out = 16'(589);
			3907: out = 16'(609);
			3908: out = 16'(631);
			3909: out = 16'(642);
			3910: out = 16'(655);
			3911: out = 16'(667);
			3912: out = 16'(684);
			3913: out = 16'(712);
			3914: out = 16'(727);
			3915: out = 16'(729);
			3916: out = 16'(744);
			3917: out = 16'(762);
			3918: out = 16'(764);
			3919: out = 16'(778);
			3920: out = 16'(789);
			3921: out = 16'(807);
			3922: out = 16'(813);
			3923: out = 16'(819);
			3924: out = 16'(811);
			3925: out = 16'(810);
			3926: out = 16'(807);
			3927: out = 16'(813);
			3928: out = 16'(818);
			3929: out = 16'(812);
			3930: out = 16'(805);
			3931: out = 16'(801);
			3932: out = 16'(805);
			3933: out = 16'(811);
			3934: out = 16'(801);
			3935: out = 16'(793);
			3936: out = 16'(789);
			3937: out = 16'(797);
			3938: out = 16'(796);
			3939: out = 16'(782);
			3940: out = 16'(778);
			3941: out = 16'(785);
			3942: out = 16'(774);
			3943: out = 16'(770);
			3944: out = 16'(749);
			3945: out = 16'(747);
			3946: out = 16'(734);
			3947: out = 16'(714);
			3948: out = 16'(693);
			3949: out = 16'(679);
			3950: out = 16'(668);
			3951: out = 16'(634);
			3952: out = 16'(617);
			3953: out = 16'(596);
			3954: out = 16'(572);
			3955: out = 16'(542);
			3956: out = 16'(531);
			3957: out = 16'(515);
			3958: out = 16'(490);
			3959: out = 16'(466);
			3960: out = 16'(441);
			3961: out = 16'(430);
			3962: out = 16'(399);
			3963: out = 16'(386);
			3964: out = 16'(363);
			3965: out = 16'(345);
			3966: out = 16'(327);
			3967: out = 16'(306);
			3968: out = 16'(285);
			3969: out = 16'(267);
			3970: out = 16'(257);
			3971: out = 16'(250);
			3972: out = 16'(227);
			3973: out = 16'(208);
			3974: out = 16'(209);
			3975: out = 16'(187);
			3976: out = 16'(180);
			3977: out = 16'(164);
			3978: out = 16'(160);
			3979: out = 16'(133);
			3980: out = 16'(128);
			3981: out = 16'(129);
			3982: out = 16'(104);
			3983: out = 16'(74);
			3984: out = 16'(51);
			3985: out = 16'(30);
			3986: out = 16'(15);
			3987: out = 16'(-9);
			3988: out = 16'(-32);
			3989: out = 16'(-50);
			3990: out = 16'(-68);
			3991: out = 16'(-81);
			3992: out = 16'(-97);
			3993: out = 16'(-113);
			3994: out = 16'(-140);
			3995: out = 16'(-154);
			3996: out = 16'(-167);
			3997: out = 16'(-179);
			3998: out = 16'(-192);
			3999: out = 16'(-205);
			4000: out = 16'(-221);
			4001: out = 16'(-246);
			4002: out = 16'(-268);
			4003: out = 16'(-278);
			4004: out = 16'(-301);
			4005: out = 16'(-318);
			4006: out = 16'(-336);
			4007: out = 16'(-348);
			4008: out = 16'(-370);
			4009: out = 16'(-405);
			4010: out = 16'(-424);
			4011: out = 16'(-452);
			4012: out = 16'(-481);
			4013: out = 16'(-507);
			4014: out = 16'(-539);
			4015: out = 16'(-581);
			4016: out = 16'(-609);
			4017: out = 16'(-632);
			4018: out = 16'(-660);
			4019: out = 16'(-683);
			4020: out = 16'(-706);
			4021: out = 16'(-723);
			4022: out = 16'(-748);
			4023: out = 16'(-774);
			4024: out = 16'(-786);
			4025: out = 16'(-794);
			4026: out = 16'(-819);
			4027: out = 16'(-826);
			4028: out = 16'(-837);
			4029: out = 16'(-836);
			4030: out = 16'(-857);
			4031: out = 16'(-847);
			4032: out = 16'(-851);
			4033: out = 16'(-855);
			4034: out = 16'(-867);
			4035: out = 16'(-867);
			4036: out = 16'(-867);
			4037: out = 16'(-866);
			4038: out = 16'(-864);
			4039: out = 16'(-843);
			4040: out = 16'(-846);
			4041: out = 16'(-846);
			4042: out = 16'(-846);
			4043: out = 16'(-842);
			4044: out = 16'(-836);
			4045: out = 16'(-841);
			4046: out = 16'(-842);
			4047: out = 16'(-825);
			4048: out = 16'(-812);
			4049: out = 16'(-801);
			4050: out = 16'(-806);
			4051: out = 16'(-794);
			4052: out = 16'(-784);
			4053: out = 16'(-770);
			4054: out = 16'(-765);
			4055: out = 16'(-744);
			4056: out = 16'(-742);
			4057: out = 16'(-725);
			4058: out = 16'(-717);
			4059: out = 16'(-703);
			4060: out = 16'(-683);
			4061: out = 16'(-667);
			4062: out = 16'(-648);
			4063: out = 16'(-640);
			4064: out = 16'(-599);
			4065: out = 16'(-584);
			4066: out = 16'(-557);
			4067: out = 16'(-527);
			4068: out = 16'(-515);
			4069: out = 16'(-483);
			4070: out = 16'(-460);
			4071: out = 16'(-443);
			4072: out = 16'(-418);
			4073: out = 16'(-401);
			4074: out = 16'(-386);
			4075: out = 16'(-365);
			4076: out = 16'(-347);
			4077: out = 16'(-317);
			4078: out = 16'(-302);
			4079: out = 16'(-298);
			4080: out = 16'(-280);
			4081: out = 16'(-255);
			4082: out = 16'(-247);
			4083: out = 16'(-238);
			4084: out = 16'(-210);
			4085: out = 16'(-203);
			4086: out = 16'(-184);
			4087: out = 16'(-181);
			4088: out = 16'(-162);
			4089: out = 16'(-147);
			4090: out = 16'(-133);
			4091: out = 16'(-108);
			4092: out = 16'(-95);
			4093: out = 16'(-74);
			4094: out = 16'(-67);
			4095: out = 16'(-51);
			4096: out = 16'(-38);
			4097: out = 16'(-24);
			4098: out = 16'(-16);
			4099: out = 16'(-4);
			4100: out = 16'(9);
			4101: out = 16'(20);
			4102: out = 16'(32);
			4103: out = 16'(38);
			4104: out = 16'(57);
			4105: out = 16'(70);
			4106: out = 16'(85);
			4107: out = 16'(89);
			4108: out = 16'(101);
			4109: out = 16'(111);
			4110: out = 16'(127);
			4111: out = 16'(131);
			4112: out = 16'(143);
			4113: out = 16'(172);
			4114: out = 16'(190);
			4115: out = 16'(219);
			4116: out = 16'(229);
			4117: out = 16'(242);
			4118: out = 16'(264);
			4119: out = 16'(282);
			4120: out = 16'(309);
			4121: out = 16'(328);
			4122: out = 16'(342);
			4123: out = 16'(367);
			4124: out = 16'(397);
			4125: out = 16'(404);
			4126: out = 16'(432);
			4127: out = 16'(429);
			4128: out = 16'(456);
			4129: out = 16'(457);
			4130: out = 16'(474);
			4131: out = 16'(495);
			4132: out = 16'(507);
			4133: out = 16'(530);
			4134: out = 16'(529);
			4135: out = 16'(547);
			4136: out = 16'(557);
			4137: out = 16'(561);
			4138: out = 16'(572);
			4139: out = 16'(581);
			4140: out = 16'(587);
			4141: out = 16'(605);
			4142: out = 16'(602);
			4143: out = 16'(620);
			4144: out = 16'(620);
			4145: out = 16'(633);
			4146: out = 16'(646);
			4147: out = 16'(646);
			4148: out = 16'(640);
			4149: out = 16'(634);
			4150: out = 16'(623);
			4151: out = 16'(632);
			4152: out = 16'(634);
			4153: out = 16'(638);
			4154: out = 16'(625);
			4155: out = 16'(633);
			4156: out = 16'(623);
			4157: out = 16'(623);
			4158: out = 16'(631);
			4159: out = 16'(614);
			4160: out = 16'(614);
			4161: out = 16'(619);
			4162: out = 16'(610);
			4163: out = 16'(619);
			4164: out = 16'(610);
			4165: out = 16'(602);
			4166: out = 16'(598);
			4167: out = 16'(598);
			4168: out = 16'(583);
			4169: out = 16'(558);
			4170: out = 16'(549);
			4171: out = 16'(543);
			4172: out = 16'(526);
			4173: out = 16'(505);
			4174: out = 16'(477);
			4175: out = 16'(477);
			4176: out = 16'(454);
			4177: out = 16'(445);
			4178: out = 16'(425);
			4179: out = 16'(404);
			4180: out = 16'(392);
			4181: out = 16'(363);
			4182: out = 16'(347);
			4183: out = 16'(333);
			4184: out = 16'(312);
			4185: out = 16'(314);
			4186: out = 16'(296);
			4187: out = 16'(267);
			4188: out = 16'(255);
			4189: out = 16'(245);
			4190: out = 16'(231);
			4191: out = 16'(220);
			4192: out = 16'(202);
			4193: out = 16'(185);
			4194: out = 16'(176);
			4195: out = 16'(173);
			4196: out = 16'(161);
			4197: out = 16'(160);
			4198: out = 16'(134);
			4199: out = 16'(124);
			4200: out = 16'(121);
			4201: out = 16'(110);
			4202: out = 16'(92);
			4203: out = 16'(97);
			4204: out = 16'(88);
			4205: out = 16'(67);
			4206: out = 16'(50);
			4207: out = 16'(31);
			4208: out = 16'(3);
			4209: out = 16'(-7);
			4210: out = 16'(-16);
			4211: out = 16'(-38);
			4212: out = 16'(-53);
			4213: out = 16'(-75);
			4214: out = 16'(-85);
			4215: out = 16'(-102);
			4216: out = 16'(-123);
			4217: out = 16'(-127);
			4218: out = 16'(-132);
			4219: out = 16'(-148);
			4220: out = 16'(-173);
			4221: out = 16'(-181);
			4222: out = 16'(-181);
			4223: out = 16'(-199);
			4224: out = 16'(-205);
			4225: out = 16'(-210);
			4226: out = 16'(-235);
			4227: out = 16'(-249);
			4228: out = 16'(-261);
			4229: out = 16'(-283);
			4230: out = 16'(-292);
			4231: out = 16'(-320);
			4232: out = 16'(-337);
			4233: out = 16'(-359);
			4234: out = 16'(-379);
			4235: out = 16'(-396);
			4236: out = 16'(-415);
			4237: out = 16'(-440);
			4238: out = 16'(-458);
			4239: out = 16'(-484);
			4240: out = 16'(-518);
			4241: out = 16'(-527);
			4242: out = 16'(-554);
			4243: out = 16'(-559);
			4244: out = 16'(-590);
			4245: out = 16'(-605);
			4246: out = 16'(-618);
			4247: out = 16'(-629);
			4248: out = 16'(-642);
			4249: out = 16'(-645);
			4250: out = 16'(-658);
			4251: out = 16'(-665);
			4252: out = 16'(-675);
			4253: out = 16'(-677);
			4254: out = 16'(-681);
			4255: out = 16'(-681);
			4256: out = 16'(-688);
			4257: out = 16'(-690);
			4258: out = 16'(-688);
			4259: out = 16'(-687);
			4260: out = 16'(-684);
			4261: out = 16'(-684);
			4262: out = 16'(-681);
			4263: out = 16'(-679);
			4264: out = 16'(-679);
			4265: out = 16'(-663);
			4266: out = 16'(-670);
			4267: out = 16'(-666);
			4268: out = 16'(-668);
			4269: out = 16'(-656);
			4270: out = 16'(-656);
			4271: out = 16'(-645);
			4272: out = 16'(-646);
			4273: out = 16'(-633);
			4274: out = 16'(-629);
			4275: out = 16'(-610);
			4276: out = 16'(-617);
			4277: out = 16'(-610);
			4278: out = 16'(-602);
			4279: out = 16'(-583);
			4280: out = 16'(-576);
			4281: out = 16'(-560);
			4282: out = 16'(-548);
			4283: out = 16'(-540);
			4284: out = 16'(-516);
			4285: out = 16'(-509);
			4286: out = 16'(-494);
			4287: out = 16'(-476);
			4288: out = 16'(-463);
			4289: out = 16'(-438);
			4290: out = 16'(-432);
			4291: out = 16'(-397);
			4292: out = 16'(-381);
			4293: out = 16'(-369);
			4294: out = 16'(-356);
			4295: out = 16'(-330);
			4296: out = 16'(-327);
			4297: out = 16'(-308);
			4298: out = 16'(-294);
			4299: out = 16'(-276);
			4300: out = 16'(-262);
			4301: out = 16'(-232);
			4302: out = 16'(-239);
			4303: out = 16'(-219);
			4304: out = 16'(-208);
			4305: out = 16'(-193);
			4306: out = 16'(-180);
			4307: out = 16'(-184);
			4308: out = 16'(-170);
			4309: out = 16'(-154);
			4310: out = 16'(-147);
			4311: out = 16'(-131);
			4312: out = 16'(-128);
			4313: out = 16'(-105);
			4314: out = 16'(-95);
			4315: out = 16'(-76);
			4316: out = 16'(-78);
			4317: out = 16'(-53);
			4318: out = 16'(-40);
			4319: out = 16'(-41);
			4320: out = 16'(-21);
			4321: out = 16'(-22);
			4322: out = 16'(-8);
			4323: out = 16'(-6);
			4324: out = 16'(13);
			4325: out = 16'(21);
			4326: out = 16'(34);
			4327: out = 16'(38);
			4328: out = 16'(54);
			4329: out = 16'(56);
			4330: out = 16'(67);
			4331: out = 16'(67);
			4332: out = 16'(79);
			4333: out = 16'(96);
			4334: out = 16'(103);
			4335: out = 16'(113);
			4336: out = 16'(125);
			4337: out = 16'(134);
			4338: out = 16'(158);
			4339: out = 16'(176);
			4340: out = 16'(194);
			4341: out = 16'(202);
			4342: out = 16'(221);
			4343: out = 16'(228);
			4344: out = 16'(255);
			4345: out = 16'(276);
			4346: out = 16'(278);
			4347: out = 16'(306);
			4348: out = 16'(315);
			4349: out = 16'(326);
			4350: out = 16'(333);
			4351: out = 16'(340);
			4352: out = 16'(364);
			4353: out = 16'(373);
			4354: out = 16'(384);
			4355: out = 16'(386);
			4356: out = 16'(400);
			4357: out = 16'(413);
			4358: out = 16'(418);
			4359: out = 16'(422);
			4360: out = 16'(444);
			4361: out = 16'(450);
			4362: out = 16'(450);
			4363: out = 16'(474);
			4364: out = 16'(467);
			4365: out = 16'(486);
			4366: out = 16'(483);
			4367: out = 16'(489);
			4368: out = 16'(489);
			4369: out = 16'(482);
			4370: out = 16'(493);
			4371: out = 16'(500);
			4372: out = 16'(501);
			4373: out = 16'(493);
			4374: out = 16'(486);
			4375: out = 16'(490);
			4376: out = 16'(482);
			4377: out = 16'(482);
			4378: out = 16'(475);
			4379: out = 16'(476);
			4380: out = 16'(470);
			4381: out = 16'(468);
			4382: out = 16'(479);
			4383: out = 16'(462);
			4384: out = 16'(482);
			4385: out = 16'(472);
			4386: out = 16'(465);
			4387: out = 16'(463);
			4388: out = 16'(458);
			4389: out = 16'(447);
			4390: out = 16'(444);
			4391: out = 16'(436);
			4392: out = 16'(417);
			4393: out = 16'(411);
			4394: out = 16'(405);
			4395: out = 16'(391);
			4396: out = 16'(377);
			4397: out = 16'(362);
			4398: out = 16'(352);
			4399: out = 16'(341);
			4400: out = 16'(327);
			4401: out = 16'(305);
			4402: out = 16'(289);
			4403: out = 16'(286);
			4404: out = 16'(277);
			4405: out = 16'(253);
			4406: out = 16'(241);
			4407: out = 16'(223);
			4408: out = 16'(220);
			4409: out = 16'(197);
			4410: out = 16'(193);
			4411: out = 16'(186);
			4412: out = 16'(170);
			4413: out = 16'(161);
			4414: out = 16'(149);
			4415: out = 16'(139);
			4416: out = 16'(120);
			4417: out = 16'(124);
			4418: out = 16'(119);
			4419: out = 16'(93);
			4420: out = 16'(98);
			4421: out = 16'(88);
			4422: out = 16'(80);
			4423: out = 16'(74);
			4424: out = 16'(65);
			4425: out = 16'(53);
			4426: out = 16'(51);
			4427: out = 16'(44);
			4428: out = 16'(36);
			4429: out = 16'(14);
			4430: out = 16'(5);
			4431: out = 16'(-5);
			4432: out = 16'(-21);
			4433: out = 16'(-32);
			4434: out = 16'(-48);
			4435: out = 16'(-60);
			4436: out = 16'(-63);
			4437: out = 16'(-76);
			4438: out = 16'(-81);
			4439: out = 16'(-97);
			4440: out = 16'(-104);
			4441: out = 16'(-111);
			4442: out = 16'(-131);
			4443: out = 16'(-133);
			4444: out = 16'(-155);
			4445: out = 16'(-156);
			4446: out = 16'(-169);
			4447: out = 16'(-182);
			4448: out = 16'(-183);
			4449: out = 16'(-196);
			4450: out = 16'(-206);
			4451: out = 16'(-214);
			4452: out = 16'(-229);
			4453: out = 16'(-247);
			4454: out = 16'(-255);
			4455: out = 16'(-261);
			4456: out = 16'(-298);
			4457: out = 16'(-310);
			4458: out = 16'(-314);
			4459: out = 16'(-348);
			4460: out = 16'(-365);
			4461: out = 16'(-379);
			4462: out = 16'(-391);
			4463: out = 16'(-410);
			4464: out = 16'(-424);
			4465: out = 16'(-445);
			4466: out = 16'(-468);
			4467: out = 16'(-462);
			4468: out = 16'(-472);
			4469: out = 16'(-483);
			4470: out = 16'(-503);
			4471: out = 16'(-505);
			4472: out = 16'(-518);
			4473: out = 16'(-526);
			4474: out = 16'(-526);
			4475: out = 16'(-540);
			4476: out = 16'(-531);
			4477: out = 16'(-538);
			4478: out = 16'(-540);
			4479: out = 16'(-543);
			4480: out = 16'(-533);
			4481: out = 16'(-553);
			4482: out = 16'(-539);
			4483: out = 16'(-540);
			4484: out = 16'(-545);
			4485: out = 16'(-537);
			4486: out = 16'(-538);
			4487: out = 16'(-534);
			4488: out = 16'(-531);
			4489: out = 16'(-528);
			4490: out = 16'(-519);
			4491: out = 16'(-518);
			4492: out = 16'(-527);
			4493: out = 16'(-516);
			4494: out = 16'(-507);
			4495: out = 16'(-515);
			4496: out = 16'(-519);
			4497: out = 16'(-501);
			4498: out = 16'(-496);
			4499: out = 16'(-487);
			4500: out = 16'(-486);
			4501: out = 16'(-470);
			4502: out = 16'(-467);
			4503: out = 16'(-460);
			4504: out = 16'(-454);
			4505: out = 16'(-433);
			4506: out = 16'(-432);
			4507: out = 16'(-413);
			4508: out = 16'(-397);
			4509: out = 16'(-399);
			4510: out = 16'(-369);
			4511: out = 16'(-369);
			4512: out = 16'(-350);
			4513: out = 16'(-332);
			4514: out = 16'(-329);
			4515: out = 16'(-298);
			4516: out = 16'(-297);
			4517: out = 16'(-275);
			4518: out = 16'(-269);
			4519: out = 16'(-247);
			4520: out = 16'(-241);
			4521: out = 16'(-220);
			4522: out = 16'(-214);
			4523: out = 16'(-217);
			4524: out = 16'(-195);
			4525: out = 16'(-183);
			4526: out = 16'(-183);
			4527: out = 16'(-162);
			4528: out = 16'(-150);
			4529: out = 16'(-150);
			4530: out = 16'(-143);
			4531: out = 16'(-137);
			4532: out = 16'(-134);
			4533: out = 16'(-120);
			4534: out = 16'(-120);
			4535: out = 16'(-95);
			4536: out = 16'(-98);
			4537: out = 16'(-75);
			4538: out = 16'(-73);
			4539: out = 16'(-52);
			4540: out = 16'(-44);
			4541: out = 16'(-36);
			4542: out = 16'(-36);
			4543: out = 16'(-24);
			4544: out = 16'(-25);
			4545: out = 16'(-15);
			4546: out = 16'(-1);
			4547: out = 16'(2);
			4548: out = 16'(4);
			4549: out = 16'(21);
			4550: out = 16'(19);
			4551: out = 16'(32);
			4552: out = 16'(36);
			4553: out = 16'(42);
			4554: out = 16'(43);
			4555: out = 16'(51);
			4556: out = 16'(62);
			4557: out = 16'(79);
			4558: out = 16'(86);
			4559: out = 16'(111);
			4560: out = 16'(116);
			4561: out = 16'(128);
			4562: out = 16'(136);
			4563: out = 16'(143);
			4564: out = 16'(155);
			4565: out = 16'(174);
			4566: out = 16'(179);
			4567: out = 16'(203);
			4568: out = 16'(211);
			4569: out = 16'(218);
			4570: out = 16'(232);
			4571: out = 16'(241);
			4572: out = 16'(253);
			4573: out = 16'(262);
			4574: out = 16'(277);
			4575: out = 16'(283);
			4576: out = 16'(283);
			4577: out = 16'(294);
			4578: out = 16'(291);
			4579: out = 16'(306);
			4580: out = 16'(312);
			4581: out = 16'(322);
			4582: out = 16'(322);
			4583: out = 16'(327);
			4584: out = 16'(340);
			4585: out = 16'(338);
			4586: out = 16'(347);
			4587: out = 16'(348);
			4588: out = 16'(361);
			4589: out = 16'(367);
			4590: out = 16'(369);
			4591: out = 16'(380);
			4592: out = 16'(380);
			4593: out = 16'(364);
			4594: out = 16'(367);
			4595: out = 16'(363);
			4596: out = 16'(374);
			4597: out = 16'(372);
			4598: out = 16'(374);
			4599: out = 16'(373);
			4600: out = 16'(348);
			4601: out = 16'(358);
			4602: out = 16'(359);
			4603: out = 16'(364);
			4604: out = 16'(363);
			4605: out = 16'(352);
			4606: out = 16'(361);
			4607: out = 16'(361);
			4608: out = 16'(351);
			4609: out = 16'(357);
			4610: out = 16'(342);
			4611: out = 16'(341);
			4612: out = 16'(330);
			4613: out = 16'(333);
			4614: out = 16'(317);
			4615: out = 16'(311);
			4616: out = 16'(308);
			4617: out = 16'(306);
			4618: out = 16'(281);
			4619: out = 16'(288);
			4620: out = 16'(269);
			4621: out = 16'(256);
			4622: out = 16'(235);
			4623: out = 16'(232);
			4624: out = 16'(219);
			4625: out = 16'(210);
			4626: out = 16'(202);
			4627: out = 16'(187);
			4628: out = 16'(171);
			4629: out = 16'(178);
			4630: out = 16'(167);
			4631: out = 16'(150);
			4632: out = 16'(143);
			4633: out = 16'(133);
			4634: out = 16'(131);
			4635: out = 16'(112);
			4636: out = 16'(119);
			4637: out = 16'(100);
			4638: out = 16'(97);
			4639: out = 16'(85);
			4640: out = 16'(83);
			4641: out = 16'(81);
			4642: out = 16'(80);
			4643: out = 16'(68);
			4644: out = 16'(63);
			4645: out = 16'(52);
			4646: out = 16'(48);
			4647: out = 16'(48);
			4648: out = 16'(36);
			4649: out = 16'(36);
			4650: out = 16'(30);
			4651: out = 16'(6);
			4652: out = 16'(2);
			4653: out = 16'(-5);
			4654: out = 16'(-16);
			4655: out = 16'(-24);
			4656: out = 16'(-42);
			4657: out = 16'(-54);
			4658: out = 16'(-55);
			4659: out = 16'(-67);
			4660: out = 16'(-83);
			4661: out = 16'(-83);
			4662: out = 16'(-86);
			4663: out = 16'(-109);
			4664: out = 16'(-109);
			4665: out = 16'(-116);
			4666: out = 16'(-110);
			4667: out = 16'(-128);
			4668: out = 16'(-134);
			4669: out = 16'(-151);
			4670: out = 16'(-144);
			4671: out = 16'(-159);
			4672: out = 16'(-166);
			4673: out = 16'(-166);
			4674: out = 16'(-183);
			4675: out = 16'(-192);
			4676: out = 16'(-196);
			4677: out = 16'(-203);
			4678: out = 16'(-217);
			4679: out = 16'(-234);
			4680: out = 16'(-249);
			4681: out = 16'(-256);
			4682: out = 16'(-273);
			4683: out = 16'(-289);
			4684: out = 16'(-299);
			4685: out = 16'(-313);
			4686: out = 16'(-336);
			4687: out = 16'(-342);
			4688: out = 16'(-360);
			4689: out = 16'(-359);
			4690: out = 16'(-367);
			4691: out = 16'(-380);
			4692: out = 16'(-386);
			4693: out = 16'(-396);
			4694: out = 16'(-407);
			4695: out = 16'(-394);
			4696: out = 16'(-403);
			4697: out = 16'(-407);
			4698: out = 16'(-422);
			4699: out = 16'(-417);
			4700: out = 16'(-415);
			4701: out = 16'(-427);
			4702: out = 16'(-425);
			4703: out = 16'(-423);
			4704: out = 16'(-411);
			4705: out = 16'(-420);
			4706: out = 16'(-428);
			4707: out = 16'(-427);
			4708: out = 16'(-419);
			4709: out = 16'(-416);
			4710: out = 16'(-421);
			4711: out = 16'(-422);
			4712: out = 16'(-415);
			4713: out = 16'(-419);
			4714: out = 16'(-408);
			4715: out = 16'(-411);
			4716: out = 16'(-407);
			4717: out = 16'(-397);
			4718: out = 16'(-400);
			4719: out = 16'(-399);
			4720: out = 16'(-382);
			4721: out = 16'(-388);
			4722: out = 16'(-381);
			4723: out = 16'(-377);
			4724: out = 16'(-377);
			4725: out = 16'(-365);
			4726: out = 16'(-363);
			4727: out = 16'(-356);
			4728: out = 16'(-356);
			4729: out = 16'(-332);
			4730: out = 16'(-322);
			4731: out = 16'(-316);
			4732: out = 16'(-304);
			4733: out = 16'(-293);
			4734: out = 16'(-278);
			4735: out = 16'(-275);
			4736: out = 16'(-256);
			4737: out = 16'(-252);
			4738: out = 16'(-250);
			4739: out = 16'(-232);
			4740: out = 16'(-219);
			4741: out = 16'(-210);
			4742: out = 16'(-200);
			4743: out = 16'(-205);
			4744: out = 16'(-191);
			4745: out = 16'(-176);
			4746: out = 16'(-179);
			4747: out = 16'(-172);
			4748: out = 16'(-159);
			4749: out = 16'(-144);
			4750: out = 16'(-141);
			4751: out = 16'(-132);
			4752: out = 16'(-119);
			4753: out = 16'(-110);
			4754: out = 16'(-120);
			4755: out = 16'(-113);
			4756: out = 16'(-102);
			4757: out = 16'(-88);
			4758: out = 16'(-90);
			4759: out = 16'(-66);
			4760: out = 16'(-63);
			4761: out = 16'(-51);
			4762: out = 16'(-51);
			4763: out = 16'(-39);
			4764: out = 16'(-46);
			4765: out = 16'(-25);
			4766: out = 16'(-27);
			4767: out = 16'(-18);
			4768: out = 16'(-19);
			4769: out = 16'(-8);
			4770: out = 16'(1);
			4771: out = 16'(-2);
			4772: out = 16'(2);
			4773: out = 16'(16);
			4774: out = 16'(22);
			4775: out = 16'(33);
			4776: out = 16'(27);
			4777: out = 16'(21);
			4778: out = 16'(44);
			4779: out = 16'(38);
			4780: out = 16'(52);
			4781: out = 16'(49);
			4782: out = 16'(72);
			4783: out = 16'(79);
			4784: out = 16'(80);
			4785: out = 16'(96);
			4786: out = 16'(105);
			4787: out = 16'(112);
			4788: out = 16'(124);
			4789: out = 16'(127);
			4790: out = 16'(135);
			4791: out = 16'(154);
			4792: out = 16'(163);
			4793: out = 16'(170);
			4794: out = 16'(172);
			4795: out = 16'(186);
			4796: out = 16'(190);
			4797: out = 16'(200);
			4798: out = 16'(203);
			4799: out = 16'(208);
			4800: out = 16'(220);
			4801: out = 16'(227);
			4802: out = 16'(216);
			4803: out = 16'(240);
			4804: out = 16'(247);
			4805: out = 16'(255);
			4806: out = 16'(256);
			4807: out = 16'(255);
			4808: out = 16'(252);
			4809: out = 16'(269);
			4810: out = 16'(263);
			4811: out = 16'(273);
			4812: out = 16'(273);
			4813: out = 16'(270);
			4814: out = 16'(275);
			4815: out = 16'(282);
			4816: out = 16'(278);
			4817: out = 16'(275);
			4818: out = 16'(255);
			4819: out = 16'(267);
			4820: out = 16'(267);
			4821: out = 16'(274);
			4822: out = 16'(262);
			4823: out = 16'(261);
			4824: out = 16'(254);
			4825: out = 16'(267);
			4826: out = 16'(256);
			4827: out = 16'(268);
			4828: out = 16'(253);
			4829: out = 16'(261);
			4830: out = 16'(251);
			4831: out = 16'(265);
			4832: out = 16'(250);
			4833: out = 16'(246);
			4834: out = 16'(252);
			4835: out = 16'(237);
			4836: out = 16'(240);
			4837: out = 16'(238);
			4838: out = 16'(222);
			4839: out = 16'(223);
			4840: out = 16'(203);
			4841: out = 16'(194);
			4842: out = 16'(207);
			4843: out = 16'(183);
			4844: out = 16'(184);
			4845: out = 16'(175);
			4846: out = 16'(161);
			4847: out = 16'(157);
			4848: out = 16'(158);
			4849: out = 16'(136);
			4850: out = 16'(139);
			4851: out = 16'(128);
			4852: out = 16'(116);
			4853: out = 16'(115);
			4854: out = 16'(107);
			4855: out = 16'(89);
			4856: out = 16'(86);
			4857: out = 16'(79);
			4858: out = 16'(68);
			4859: out = 16'(84);
			4860: out = 16'(73);
			4861: out = 16'(60);
			4862: out = 16'(49);
			4863: out = 16'(41);
			4864: out = 16'(42);
			4865: out = 16'(37);
			4866: out = 16'(41);
			4867: out = 16'(37);
			4868: out = 16'(29);
			4869: out = 16'(16);
			4870: out = 16'(25);
			4871: out = 16'(25);
			4872: out = 16'(9);
			4873: out = 16'(2);
			4874: out = 16'(1);
			4875: out = 16'(-16);
			4876: out = 16'(-30);
			4877: out = 16'(-41);
			4878: out = 16'(-38);
			4879: out = 16'(-29);
			4880: out = 16'(-49);
			4881: out = 16'(-53);
			4882: out = 16'(-57);
			4883: out = 16'(-61);
			4884: out = 16'(-77);
			4885: out = 16'(-72);
			4886: out = 16'(-80);
			4887: out = 16'(-96);
			4888: out = 16'(-105);
			4889: out = 16'(-104);
			4890: out = 16'(-113);
			4891: out = 16'(-122);
			4892: out = 16'(-117);
			4893: out = 16'(-127);
			4894: out = 16'(-120);
			4895: out = 16'(-132);
			4896: out = 16'(-137);
			4897: out = 16'(-143);
			4898: out = 16'(-156);
			4899: out = 16'(-163);
			4900: out = 16'(-175);
			4901: out = 16'(-174);
			4902: out = 16'(-193);
			4903: out = 16'(-187);
			4904: out = 16'(-215);
			4905: out = 16'(-226);
			4906: out = 16'(-239);
			4907: out = 16'(-243);
			4908: out = 16'(-250);
			4909: out = 16'(-254);
			4910: out = 16'(-271);
			4911: out = 16'(-282);
			4912: out = 16'(-279);
			4913: out = 16'(-279);
			4914: out = 16'(-286);
			4915: out = 16'(-300);
			4916: out = 16'(-305);
			4917: out = 16'(-312);
			4918: out = 16'(-316);
			4919: out = 16'(-324);
			4920: out = 16'(-313);
			4921: out = 16'(-322);
			4922: out = 16'(-322);
			4923: out = 16'(-333);
			4924: out = 16'(-323);
			4925: out = 16'(-333);
			4926: out = 16'(-328);
			4927: out = 16'(-326);
			4928: out = 16'(-323);
			4929: out = 16'(-318);
			4930: out = 16'(-327);
			4931: out = 16'(-313);
			4932: out = 16'(-321);
			4933: out = 16'(-330);
			4934: out = 16'(-320);
			4935: out = 16'(-328);
			4936: out = 16'(-321);
			4937: out = 16'(-321);
			4938: out = 16'(-309);
			4939: out = 16'(-316);
			4940: out = 16'(-309);
			4941: out = 16'(-305);
			4942: out = 16'(-310);
			4943: out = 16'(-309);
			4944: out = 16'(-316);
			4945: out = 16'(-299);
			4946: out = 16'(-298);
			4947: out = 16'(-296);
			4948: out = 16'(-293);
			4949: out = 16'(-285);
			4950: out = 16'(-283);
			4951: out = 16'(-266);
			4952: out = 16'(-262);
			4953: out = 16'(-268);
			4954: out = 16'(-250);
			4955: out = 16'(-241);
			4956: out = 16'(-219);
			4957: out = 16'(-227);
			4958: out = 16'(-212);
			4959: out = 16'(-207);
			4960: out = 16'(-203);
			4961: out = 16'(-190);
			4962: out = 16'(-179);
			4963: out = 16'(-175);
			4964: out = 16'(-171);
			4965: out = 16'(-150);
			4966: out = 16'(-162);
			4967: out = 16'(-156);
			4968: out = 16'(-135);
			4969: out = 16'(-146);
			4970: out = 16'(-131);
			4971: out = 16'(-119);
			4972: out = 16'(-121);
			4973: out = 16'(-116);
			4974: out = 16'(-103);
			4975: out = 16'(-104);
			4976: out = 16'(-105);
			4977: out = 16'(-104);
			4978: out = 16'(-88);
			4979: out = 16'(-85);
			4980: out = 16'(-79);
			4981: out = 16'(-70);
			4982: out = 16'(-61);
			4983: out = 16'(-48);
			4984: out = 16'(-46);
			4985: out = 16'(-49);
			4986: out = 16'(-36);
			4987: out = 16'(-37);
			4988: out = 16'(-31);
			4989: out = 16'(-21);
			4990: out = 16'(-25);
			4991: out = 16'(-20);
			4992: out = 16'(-18);
			4993: out = 16'(-20);
			4994: out = 16'(-9);
			4995: out = 16'(-13);
			4996: out = 16'(1);
			4997: out = 16'(3);
			4998: out = 16'(14);
			4999: out = 16'(14);
			5000: out = 16'(13);
			5001: out = 16'(28);
			5002: out = 16'(28);
			5003: out = 16'(30);
			5004: out = 16'(43);
			5005: out = 16'(50);
			5006: out = 16'(53);
			5007: out = 16'(66);
			5008: out = 16'(69);
			5009: out = 16'(77);
			5010: out = 16'(83);
			5011: out = 16'(86);
			5012: out = 16'(95);
			5013: out = 16'(100);
			5014: out = 16'(98);
			5015: out = 16'(113);
			5016: out = 16'(122);
			5017: out = 16'(136);
			5018: out = 16'(139);
			5019: out = 16'(134);
			5020: out = 16'(143);
			5021: out = 16'(146);
			5022: out = 16'(157);
			5023: out = 16'(156);
			5024: out = 16'(155);
			5025: out = 16'(166);
			5026: out = 16'(167);
			5027: out = 16'(174);
			5028: out = 16'(182);
			5029: out = 16'(164);
			5030: out = 16'(182);
			5031: out = 16'(179);
			5032: out = 16'(188);
			5033: out = 16'(191);
			5034: out = 16'(194);
			5035: out = 16'(198);
			5036: out = 16'(199);
			5037: out = 16'(199);
			5038: out = 16'(188);
			5039: out = 16'(183);
			5040: out = 16'(190);
			5041: out = 16'(199);
			5042: out = 16'(194);
			5043: out = 16'(179);
			5044: out = 16'(198);
			5045: out = 16'(179);
			5046: out = 16'(192);
			5047: out = 16'(183);
			5048: out = 16'(187);
			5049: out = 16'(195);
			5050: out = 16'(173);
			5051: out = 16'(185);
			5052: out = 16'(183);
			5053: out = 16'(185);
			5054: out = 16'(183);
			5055: out = 16'(176);
			5056: out = 16'(162);
			5057: out = 16'(164);
			5058: out = 16'(164);
			5059: out = 16'(172);
			5060: out = 16'(149);
			5061: out = 16'(154);
			5062: out = 16'(148);
			5063: out = 16'(143);
			5064: out = 16'(139);
			5065: out = 16'(140);
			5066: out = 16'(119);
			5067: out = 16'(116);
			5068: out = 16'(114);
			5069: out = 16'(102);
			5070: out = 16'(107);
			5071: out = 16'(98);
			5072: out = 16'(98);
			5073: out = 16'(91);
			5074: out = 16'(76);
			5075: out = 16'(75);
			5076: out = 16'(63);
			5077: out = 16'(70);
			5078: out = 16'(62);
			5079: out = 16'(62);
			5080: out = 16'(50);
			5081: out = 16'(38);
			5082: out = 16'(33);
			5083: out = 16'(44);
			5084: out = 16'(40);
			5085: out = 16'(24);
			5086: out = 16'(26);
			5087: out = 16'(28);
			5088: out = 16'(15);
			5089: out = 16'(12);
			5090: out = 16'(12);
			5091: out = 16'(8);
			5092: out = 16'(6);
			5093: out = 16'(8);
			5094: out = 16'(10);
			5095: out = 16'(-14);
			5096: out = 16'(-8);
			5097: out = 16'(-4);
			5098: out = 16'(-21);
			5099: out = 16'(-27);
			5100: out = 16'(-37);
			5101: out = 16'(-45);
			5102: out = 16'(-42);
			5103: out = 16'(-54);
			5104: out = 16'(-49);
			5105: out = 16'(-43);
			5106: out = 16'(-69);
			5107: out = 16'(-64);
			5108: out = 16'(-77);
			5109: out = 16'(-78);
			5110: out = 16'(-74);
			5111: out = 16'(-75);
			5112: out = 16'(-86);
			5113: out = 16'(-83);
			5114: out = 16'(-100);
			5115: out = 16'(-101);
			5116: out = 16'(-101);
			5117: out = 16'(-104);
			5118: out = 16'(-103);
			5119: out = 16'(-112);
			5120: out = 16'(-122);
			5121: out = 16'(-120);
			5122: out = 16'(-132);
			5123: out = 16'(-139);
			5124: out = 16'(-137);
			5125: out = 16'(-160);
			5126: out = 16'(-152);
			5127: out = 16'(-159);
			5128: out = 16'(-167);
			5129: out = 16'(-173);
			5130: out = 16'(-185);
			5131: out = 16'(-197);
			5132: out = 16'(-200);
			5133: out = 16'(-207);
			5134: out = 16'(-207);
			5135: out = 16'(-222);
			5136: out = 16'(-222);
			5137: out = 16'(-225);
			5138: out = 16'(-233);
			5139: out = 16'(-233);
			5140: out = 16'(-235);
			5141: out = 16'(-233);
			5142: out = 16'(-241);
			5143: out = 16'(-250);
			5144: out = 16'(-253);
			5145: out = 16'(-245);
			5146: out = 16'(-245);
			5147: out = 16'(-254);
			5148: out = 16'(-252);
			5149: out = 16'(-251);
			5150: out = 16'(-261);
			5151: out = 16'(-253);
			5152: out = 16'(-257);
			5153: out = 16'(-250);
			5154: out = 16'(-251);
			5155: out = 16'(-253);
			5156: out = 16'(-255);
			5157: out = 16'(-255);
			5158: out = 16'(-243);
			5159: out = 16'(-256);
			5160: out = 16'(-252);
			5161: out = 16'(-245);
			5162: out = 16'(-240);
			5163: out = 16'(-238);
			5164: out = 16'(-241);
			5165: out = 16'(-242);
			5166: out = 16'(-233);
			5167: out = 16'(-233);
			5168: out = 16'(-223);
			5169: out = 16'(-230);
			5170: out = 16'(-210);
			5171: out = 16'(-214);
			5172: out = 16'(-207);
			5173: out = 16'(-214);
			5174: out = 16'(-209);
			5175: out = 16'(-196);
			5176: out = 16'(-184);
			5177: out = 16'(-194);
			5178: out = 16'(-186);
			5179: out = 16'(-180);
			5180: out = 16'(-176);
			5181: out = 16'(-176);
			5182: out = 16'(-161);
			5183: out = 16'(-164);
			5184: out = 16'(-143);
			5185: out = 16'(-136);
			5186: out = 16'(-129);
			5187: out = 16'(-137);
			5188: out = 16'(-117);
			5189: out = 16'(-133);
			5190: out = 16'(-121);
			5191: out = 16'(-115);
			5192: out = 16'(-119);
			5193: out = 16'(-111);
			5194: out = 16'(-101);
			5195: out = 16'(-97);
			5196: out = 16'(-85);
			5197: out = 16'(-83);
			5198: out = 16'(-81);
			5199: out = 16'(-80);
			5200: out = 16'(-80);
			5201: out = 16'(-77);
			5202: out = 16'(-66);
			5203: out = 16'(-56);
			5204: out = 16'(-52);
			5205: out = 16'(-60);
			5206: out = 16'(-51);
			5207: out = 16'(-52);
			5208: out = 16'(-45);
			5209: out = 16'(-42);
			5210: out = 16'(-31);
			5211: out = 16'(-30);
			5212: out = 16'(-28);
			5213: out = 16'(-21);
			5214: out = 16'(-26);
			5215: out = 16'(-19);
			5216: out = 16'(-21);
			5217: out = 16'(-9);
			5218: out = 16'(-10);
			5219: out = 16'(-9);
			5220: out = 16'(-8);
			5221: out = 16'(0);
			5222: out = 16'(2);
			5223: out = 16'(10);
			5224: out = 16'(7);
			5225: out = 16'(6);
			5226: out = 16'(12);
			5227: out = 16'(22);
			5228: out = 16'(26);
			5229: out = 16'(29);
			5230: out = 16'(37);
			5231: out = 16'(38);
			5232: out = 16'(49);
			5233: out = 16'(54);
			5234: out = 16'(64);
			5235: out = 16'(58);
			5236: out = 16'(64);
			5237: out = 16'(68);
			5238: out = 16'(74);
			5239: out = 16'(81);
			5240: out = 16'(85);
			5241: out = 16'(90);
			5242: out = 16'(90);
			5243: out = 16'(102);
			5244: out = 16'(97);
			5245: out = 16'(107);
			5246: out = 16'(108);
			5247: out = 16'(108);
			5248: out = 16'(115);
			5249: out = 16'(113);
			5250: out = 16'(123);
			5251: out = 16'(121);
			5252: out = 16'(117);
			5253: out = 16'(116);
			5254: out = 16'(128);
			5255: out = 16'(133);
			5256: out = 16'(133);
			5257: out = 16'(128);
			5258: out = 16'(133);
			5259: out = 16'(134);
			5260: out = 16'(132);
			5261: out = 16'(141);
			5262: out = 16'(127);
			5263: out = 16'(127);
			5264: out = 16'(121);
			5265: out = 16'(125);
			5266: out = 16'(135);
			5267: out = 16'(132);
			5268: out = 16'(128);
			5269: out = 16'(132);
			5270: out = 16'(124);
			5271: out = 16'(124);
			5272: out = 16'(117);
			5273: out = 16'(122);
			5274: out = 16'(122);
			5275: out = 16'(121);
			5276: out = 16'(122);
			5277: out = 16'(121);
			5278: out = 16'(117);
			5279: out = 16'(112);
			5280: out = 16'(105);
			5281: out = 16'(109);
			5282: out = 16'(98);
			5283: out = 16'(103);
			5284: out = 16'(87);
			5285: out = 16'(99);
			5286: out = 16'(97);
			5287: out = 16'(97);
			5288: out = 16'(92);
			5289: out = 16'(79);
			5290: out = 16'(72);
			5291: out = 16'(65);
			5292: out = 16'(66);
			5293: out = 16'(51);
			5294: out = 16'(48);
			5295: out = 16'(49);
			5296: out = 16'(36);
			5297: out = 16'(49);
			5298: out = 16'(37);
			5299: out = 16'(36);
			5300: out = 16'(28);
			5301: out = 16'(15);
			5302: out = 16'(20);
			5303: out = 16'(24);
			5304: out = 16'(15);
			5305: out = 16'(19);
			5306: out = 16'(5);
			5307: out = 16'(13);
			5308: out = 16'(4);
			5309: out = 16'(5);
			5310: out = 16'(2);
			5311: out = 16'(-12);
			5312: out = 16'(0);
			5313: out = 16'(-6);
			5314: out = 16'(-10);
			5315: out = 16'(-19);
			5316: out = 16'(-12);
			5317: out = 16'(-14);
			5318: out = 16'(-21);
			5319: out = 16'(-24);
			5320: out = 16'(-24);
			5321: out = 16'(-27);
			5322: out = 16'(-37);
			5323: out = 16'(-38);
			5324: out = 16'(-40);
			5325: out = 16'(-44);
			5326: out = 16'(-58);
			5327: out = 16'(-58);
			5328: out = 16'(-56);
			5329: out = 16'(-54);
			5330: out = 16'(-58);
			5331: out = 16'(-66);
			5332: out = 16'(-79);
			5333: out = 16'(-72);
			5334: out = 16'(-75);
			5335: out = 16'(-67);
			5336: out = 16'(-76);
			5337: out = 16'(-77);
			5338: out = 16'(-83);
			5339: out = 16'(-79);
			5340: out = 16'(-86);
			5341: out = 16'(-91);
			5342: out = 16'(-95);
			5343: out = 16'(-100);
			5344: out = 16'(-99);
			5345: out = 16'(-107);
			5346: out = 16'(-110);
			5347: out = 16'(-115);
			5348: out = 16'(-119);
			5349: out = 16'(-128);
			5350: out = 16'(-128);
			5351: out = 16'(-140);
			5352: out = 16'(-139);
			5353: out = 16'(-148);
			5354: out = 16'(-149);
			5355: out = 16'(-164);
			5356: out = 16'(-160);
			5357: out = 16'(-167);
			5358: out = 16'(-166);
			5359: out = 16'(-174);
			5360: out = 16'(-166);
			5361: out = 16'(-172);
			5362: out = 16'(-184);
			5363: out = 16'(-163);
			5364: out = 16'(-181);
			5365: out = 16'(-181);
			5366: out = 16'(-181);
			5367: out = 16'(-191);
			5368: out = 16'(-190);
			5369: out = 16'(-192);
			5370: out = 16'(-190);
			5371: out = 16'(-191);
			5372: out = 16'(-187);
			5373: out = 16'(-186);
			5374: out = 16'(-184);
			5375: out = 16'(-182);
			5376: out = 16'(-190);
			5377: out = 16'(-185);
			5378: out = 16'(-180);
			5379: out = 16'(-179);
			5380: out = 16'(-182);
			5381: out = 16'(-191);
			5382: out = 16'(-191);
			5383: out = 16'(-194);
			5384: out = 16'(-182);
			5385: out = 16'(-187);
			5386: out = 16'(-181);
			5387: out = 16'(-184);
			5388: out = 16'(-194);
			5389: out = 16'(-178);
			5390: out = 16'(-184);
			5391: out = 16'(-178);
			5392: out = 16'(-163);
			5393: out = 16'(-179);
			5394: out = 16'(-175);
			5395: out = 16'(-164);
			5396: out = 16'(-159);
			5397: out = 16'(-167);
			5398: out = 16'(-161);
			5399: out = 16'(-155);
			5400: out = 16'(-158);
			5401: out = 16'(-150);
			5402: out = 16'(-143);
			5403: out = 16'(-137);
			5404: out = 16'(-132);
			5405: out = 16'(-124);
			5406: out = 16'(-127);
			5407: out = 16'(-116);
			5408: out = 16'(-105);
			5409: out = 16'(-101);
			5410: out = 16'(-108);
			5411: out = 16'(-100);
			5412: out = 16'(-95);
			5413: out = 16'(-98);
			5414: out = 16'(-85);
			5415: out = 16'(-96);
			5416: out = 16'(-86);
			5417: out = 16'(-87);
			5418: out = 16'(-76);
			5419: out = 16'(-81);
			5420: out = 16'(-77);
			5421: out = 16'(-79);
			5422: out = 16'(-68);
			5423: out = 16'(-77);
			5424: out = 16'(-66);
			5425: out = 16'(-63);
			5426: out = 16'(-60);
			5427: out = 16'(-46);
			5428: out = 16'(-49);
			5429: out = 16'(-42);
			5430: out = 16'(-43);
			5431: out = 16'(-54);
			5432: out = 16'(-37);
			5433: out = 16'(-33);
			5434: out = 16'(-37);
			5435: out = 16'(-38);
			5436: out = 16'(-28);
			5437: out = 16'(-27);
			5438: out = 16'(-24);
			5439: out = 16'(-20);
			5440: out = 16'(-22);
			5441: out = 16'(-24);
			5442: out = 16'(-17);
			5443: out = 16'(-14);
			5444: out = 16'(-2);
			5445: out = 16'(-6);
			5446: out = 16'(-12);
			default: out = 0;
		endcase
	end
endmodule
