module snare_lookup(index, out);
	input logic unsigned [11:0] index;
	output logic signed [15:0] out;
	always_comb begin
		case(index)
			0: out = 16'(18770);
			1: out = 16'(16727);
			2: out = 16'(16);
			3: out = 16'(-21435);
			4: out = 16'(2);
			5: out = 16'(23562);
			6: out = 16'(13);
			7: out = 16'(-52);
			8: out = 16'(7171);
			9: out = 16'(2183);
			10: out = 16'(-5407);
			11: out = 16'(-9265);
			12: out = 16'(1518);
			13: out = 16'(6871);
			14: out = 16'(-4366);
			15: out = 16'(-10684);
			16: out = 16'(-5174);
			17: out = 16'(19084);
			18: out = 16'(-8681);
			19: out = 16'(-7718);
			20: out = 16'(-11558);
			21: out = 16'(22781);
			22: out = 16'(1547);
			23: out = 16'(1475);
			24: out = 16'(-11965);
			25: out = 16'(8095);
			26: out = 16'(12069);
			27: out = 16'(-5930);
			28: out = 16'(21052);
			29: out = 16'(-14769);
			30: out = 16'(30798);
			31: out = 16'(21219);
			32: out = 16'(30918);
			33: out = 16'(28162);
			34: out = 16'(30695);
			35: out = 16'(30600);
			36: out = 16'(30557);
			37: out = 16'(30421);
			38: out = 16'(30364);
			39: out = 16'(30222);
			40: out = 16'(30118);
			41: out = 16'(30066);
			42: out = 16'(29918);
			43: out = 16'(26620);
			44: out = 16'(9283);
			45: out = 16'(-7249);
			46: out = 16'(-7541);
			47: out = 16'(-14923);
			48: out = 16'(-25236);
			49: out = 16'(-31114);
			50: out = 16'(-30870);
			51: out = 16'(-26714);
			52: out = 16'(-30997);
			53: out = 16'(-30693);
			54: out = 16'(-30399);
			55: out = 16'(-30972);
			56: out = 16'(-30718);
			57: out = 16'(-28153);
			58: out = 16'(-30378);
			59: out = 16'(-24247);
			60: out = 16'(-6742);
			61: out = 16'(-5105);
			62: out = 16'(-597);
			63: out = 16'(874);
			64: out = 16'(28876);
			65: out = 16'(17035);
			66: out = 16'(30894);
			67: out = 16'(18741);
			68: out = 16'(31049);
			69: out = 16'(30672);
			70: out = 16'(29874);
			71: out = 16'(30366);
			72: out = 16'(29949);
			73: out = 16'(30543);
			74: out = 16'(28273);
			75: out = 16'(22155);
			76: out = 16'(18665);
			77: out = 16'(945);
			78: out = 16'(3700);
			79: out = 16'(-782);
			80: out = 16'(11605);
			81: out = 16'(6661);
			82: out = 16'(-5079);
			83: out = 16'(-9182);
			84: out = 16'(9792);
			85: out = 16'(7102);
			86: out = 16'(-35);
			87: out = 16'(-13159);
			88: out = 16'(12526);
			89: out = 16'(-1022);
			90: out = 16'(16283);
			91: out = 16'(-1713);
			92: out = 16'(-1111);
			93: out = 16'(14412);
			94: out = 16'(-1358);
			95: out = 16'(-13815);
			96: out = 16'(396);
			97: out = 16'(-32765);
			98: out = 16'(-14964);
			99: out = 16'(1723);
			100: out = 16'(-22260);
			101: out = 16'(-29749);
			102: out = 16'(-29064);
			103: out = 16'(-27936);
			104: out = 16'(-30966);
			105: out = 16'(-29694);
			106: out = 16'(-19788);
			107: out = 16'(-30024);
			108: out = 16'(-30245);
			109: out = 16'(-18594);
			110: out = 16'(-30593);
			111: out = 16'(-29460);
			112: out = 16'(-30528);
			113: out = 16'(-29078);
			114: out = 16'(-30506);
			115: out = 16'(-9507);
			116: out = 16'(-29409);
			117: out = 16'(-30307);
			118: out = 16'(-17672);
			119: out = 16'(-10843);
			120: out = 16'(-12737);
			121: out = 16'(-20699);
			122: out = 16'(2611);
			123: out = 16'(-4679);
			124: out = 16'(3589);
			125: out = 16'(1156);
			126: out = 16'(14380);
			127: out = 16'(9843);
			128: out = 16'(23271);
			129: out = 16'(19789);
			130: out = 16'(31498);
			131: out = 16'(28838);
			132: out = 16'(27106);
			133: out = 16'(27318);
			134: out = 16'(30860);
			135: out = 16'(30724);
			136: out = 16'(30672);
			137: out = 16'(30578);
			138: out = 16'(30649);
			139: out = 16'(30919);
			140: out = 16'(21298);
			141: out = 16'(30716);
			142: out = 16'(29611);
			143: out = 16'(29403);
			144: out = 16'(30107);
			145: out = 16'(30081);
			146: out = 16'(23283);
			147: out = 16'(19088);
			148: out = 16'(24879);
			149: out = 16'(9585);
			150: out = 16'(15219);
			151: out = 16'(6589);
			152: out = 16'(10244);
			153: out = 16'(15590);
			154: out = 16'(9658);
			155: out = 16'(-2812);
			156: out = 16'(3153);
			157: out = 16'(-4328);
			158: out = 16'(-491);
			159: out = 16'(-10437);
			160: out = 16'(-14276);
			161: out = 16'(-32257);
			162: out = 16'(-25517);
			163: out = 16'(-18036);
			164: out = 16'(-31525);
			165: out = 16'(-27097);
			166: out = 16'(-31682);
			167: out = 16'(-28460);
			168: out = 16'(-31135);
			169: out = 16'(-31009);
			170: out = 16'(-30867);
			171: out = 16'(-30717);
			172: out = 16'(-30641);
			173: out = 16'(-30504);
			174: out = 16'(-28026);
			175: out = 16'(-30064);
			176: out = 16'(-29917);
			177: out = 16'(-30281);
			178: out = 16'(-30152);
			179: out = 16'(-26486);
			180: out = 16'(-29834);
			181: out = 16'(-29799);
			182: out = 16'(-30651);
			183: out = 16'(-26047);
			184: out = 16'(-18019);
			185: out = 16'(-16674);
			186: out = 16'(-9414);
			187: out = 16'(-278);
			188: out = 16'(-208);
			189: out = 16'(6470);
			190: out = 16'(13010);
			191: out = 16'(9059);
			192: out = 16'(22820);
			193: out = 16'(25046);
			194: out = 16'(9415);
			195: out = 16'(18157);
			196: out = 16'(23314);
			197: out = 16'(18343);
			198: out = 16'(21753);
			199: out = 16'(22808);
			200: out = 16'(18243);
			201: out = 16'(31230);
			202: out = 16'(19048);
			203: out = 16'(31176);
			204: out = 16'(28509);
			205: out = 16'(15475);
			206: out = 16'(23050);
			207: out = 16'(21405);
			208: out = 16'(6916);
			209: out = 16'(2957);
			210: out = 16'(20172);
			211: out = 16'(17661);
			212: out = 16'(26416);
			213: out = 16'(10576);
			214: out = 16'(11733);
			215: out = 16'(10716);
			216: out = 16'(13685);
			217: out = 16'(-2396);
			218: out = 16'(8098);
			219: out = 16'(10050);
			220: out = 16'(-9944);
			221: out = 16'(-11667);
			222: out = 16'(17990);
			223: out = 16'(-19215);
			224: out = 16'(-3966);
			225: out = 16'(1129);
			226: out = 16'(-15400);
			227: out = 16'(-14431);
			228: out = 16'(5558);
			229: out = 16'(-3915);
			230: out = 16'(-12082);
			231: out = 16'(-9438);
			232: out = 16'(1367);
			233: out = 16'(-11488);
			234: out = 16'(-19585);
			235: out = 16'(1921);
			236: out = 16'(-13368);
			237: out = 16'(-14597);
			238: out = 16'(-16361);
			239: out = 16'(-23802);
			240: out = 16'(-335);
			241: out = 16'(-17204);
			242: out = 16'(-13480);
			243: out = 16'(-19297);
			244: out = 16'(-21497);
			245: out = 16'(-14748);
			246: out = 16'(-14815);
			247: out = 16'(-220);
			248: out = 16'(-17930);
			249: out = 16'(-12572);
			250: out = 16'(-8447);
			251: out = 16'(1906);
			252: out = 16'(-14169);
			253: out = 16'(-18963);
			254: out = 16'(7758);
			255: out = 16'(-27055);
			256: out = 16'(-20767);
			257: out = 16'(-7164);
			258: out = 16'(-5336);
			259: out = 16'(-12856);
			260: out = 16'(-16243);
			261: out = 16'(-10502);
			262: out = 16'(-10212);
			263: out = 16'(-8632);
			264: out = 16'(-10683);
			265: out = 16'(-1326);
			266: out = 16'(-13394);
			267: out = 16'(358);
			268: out = 16'(15720);
			269: out = 16'(-10751);
			270: out = 16'(6355);
			271: out = 16'(-10340);
			272: out = 16'(-5591);
			273: out = 16'(1514);
			274: out = 16'(-148);
			275: out = 16'(13578);
			276: out = 16'(6946);
			277: out = 16'(5666);
			278: out = 16'(1658);
			279: out = 16'(5872);
			280: out = 16'(944);
			281: out = 16'(11848);
			282: out = 16'(-5582);
			283: out = 16'(11537);
			284: out = 16'(3296);
			285: out = 16'(6651);
			286: out = 16'(-4833);
			287: out = 16'(9942);
			288: out = 16'(-1483);
			289: out = 16'(13056);
			290: out = 16'(5425);
			291: out = 16'(14555);
			292: out = 16'(-1549);
			293: out = 16'(4719);
			294: out = 16'(18279);
			295: out = 16'(20229);
			296: out = 16'(347);
			297: out = 16'(-2260);
			298: out = 16'(28062);
			299: out = 16'(-12553);
			300: out = 16'(11723);
			301: out = 16'(22485);
			302: out = 16'(4322);
			303: out = 16'(10961);
			304: out = 16'(15485);
			305: out = 16'(16964);
			306: out = 16'(-3859);
			307: out = 16'(17968);
			308: out = 16'(3734);
			309: out = 16'(11956);
			310: out = 16'(15259);
			311: out = 16'(4783);
			312: out = 16'(-7888);
			313: out = 16'(6230);
			314: out = 16'(10208);
			315: out = 16'(2689);
			316: out = 16'(2311);
			317: out = 16'(13419);
			318: out = 16'(-6346);
			319: out = 16'(14569);
			320: out = 16'(-20218);
			321: out = 16'(11509);
			322: out = 16'(5037);
			323: out = 16'(-10771);
			324: out = 16'(1221);
			325: out = 16'(5100);
			326: out = 16'(-2054);
			327: out = 16'(-15423);
			328: out = 16'(-13533);
			329: out = 16'(110);
			330: out = 16'(-20329);
			331: out = 16'(-12594);
			332: out = 16'(-4328);
			333: out = 16'(-19143);
			334: out = 16'(-12507);
			335: out = 16'(-16545);
			336: out = 16'(-8458);
			337: out = 16'(-20542);
			338: out = 16'(-12650);
			339: out = 16'(-9857);
			340: out = 16'(-19195);
			341: out = 16'(-17254);
			342: out = 16'(-22035);
			343: out = 16'(-11863);
			344: out = 16'(-29567);
			345: out = 16'(-11764);
			346: out = 16'(-14306);
			347: out = 16'(-27548);
			348: out = 16'(-30155);
			349: out = 16'(-9422);
			350: out = 16'(-17330);
			351: out = 16'(-14370);
			352: out = 16'(-9558);
			353: out = 16'(-12521);
			354: out = 16'(-20146);
			355: out = 16'(-17904);
			356: out = 16'(-23080);
			357: out = 16'(-11154);
			358: out = 16'(1716);
			359: out = 16'(7422);
			360: out = 16'(4015);
			361: out = 16'(4466);
			362: out = 16'(14273);
			363: out = 16'(-491);
			364: out = 16'(13164);
			365: out = 16'(-3798);
			366: out = 16'(23083);
			367: out = 16'(-522);
			368: out = 16'(2247);
			369: out = 16'(18325);
			370: out = 16'(20098);
			371: out = 16'(12196);
			372: out = 16'(8442);
			373: out = 16'(24693);
			374: out = 16'(4683);
			375: out = 16'(19988);
			376: out = 16'(-4137);
			377: out = 16'(9094);
			378: out = 16'(8892);
			379: out = 16'(26070);
			380: out = 16'(-3723);
			381: out = 16'(-113);
			382: out = 16'(27262);
			383: out = 16'(4403);
			384: out = 16'(1617);
			385: out = 16'(16241);
			386: out = 16'(-1137);
			387: out = 16'(9262);
			388: out = 16'(12847);
			389: out = 16'(24281);
			390: out = 16'(13562);
			391: out = 16'(388);
			392: out = 16'(-2087);
			393: out = 16'(11443);
			394: out = 16'(17247);
			395: out = 16'(-7728);
			396: out = 16'(9820);
			397: out = 16'(5599);
			398: out = 16'(7905);
			399: out = 16'(18197);
			400: out = 16'(1820);
			401: out = 16'(-3524);
			402: out = 16'(9381);
			403: out = 16'(-13897);
			404: out = 16'(330);
			405: out = 16'(-13190);
			406: out = 16'(-446);
			407: out = 16'(-22495);
			408: out = 16'(6691);
			409: out = 16'(-8529);
			410: out = 16'(-19118);
			411: out = 16'(-2879);
			412: out = 16'(-6180);
			413: out = 16'(4852);
			414: out = 16'(-12973);
			415: out = 16'(-9442);
			416: out = 16'(-3340);
			417: out = 16'(-11512);
			418: out = 16'(-2701);
			419: out = 16'(639);
			420: out = 16'(-13499);
			421: out = 16'(-12242);
			422: out = 16'(4341);
			423: out = 16'(-15255);
			424: out = 16'(-17008);
			425: out = 16'(-8507);
			426: out = 16'(-11461);
			427: out = 16'(-310);
			428: out = 16'(-13521);
			429: out = 16'(-10350);
			430: out = 16'(-4942);
			431: out = 16'(-15904);
			432: out = 16'(11704);
			433: out = 16'(2258);
			434: out = 16'(-7036);
			435: out = 16'(-9413);
			436: out = 16'(-2625);
			437: out = 16'(-13502);
			438: out = 16'(-18154);
			439: out = 16'(9011);
			440: out = 16'(-7822);
			441: out = 16'(-21185);
			442: out = 16'(-3846);
			443: out = 16'(3692);
			444: out = 16'(-3121);
			445: out = 16'(3162);
			446: out = 16'(-16272);
			447: out = 16'(10981);
			448: out = 16'(1967);
			449: out = 16'(6030);
			450: out = 16'(-5996);
			451: out = 16'(17746);
			452: out = 16'(10715);
			453: out = 16'(-1947);
			454: out = 16'(9717);
			455: out = 16'(4253);
			456: out = 16'(2352);
			457: out = 16'(8141);
			458: out = 16'(-3395);
			459: out = 16'(12969);
			460: out = 16'(-3219);
			461: out = 16'(18733);
			462: out = 16'(22745);
			463: out = 16'(11689);
			464: out = 16'(485);
			465: out = 16'(3867);
			466: out = 16'(17432);
			467: out = 16'(-10602);
			468: out = 16'(10032);
			469: out = 16'(15629);
			470: out = 16'(-5881);
			471: out = 16'(2996);
			472: out = 16'(-11228);
			473: out = 16'(26984);
			474: out = 16'(1396);
			475: out = 16'(-4421);
			476: out = 16'(773);
			477: out = 16'(788);
			478: out = 16'(2973);
			479: out = 16'(13025);
			480: out = 16'(4436);
			481: out = 16'(18119);
			482: out = 16'(2426);
			483: out = 16'(1986);
			484: out = 16'(15520);
			485: out = 16'(-5944);
			486: out = 16'(-15474);
			487: out = 16'(11048);
			488: out = 16'(-15374);
			489: out = 16'(16);
			490: out = 16'(14351);
			491: out = 16'(2332);
			492: out = 16'(5183);
			493: out = 16'(2014);
			494: out = 16'(4381);
			495: out = 16'(-15282);
			496: out = 16'(2823);
			497: out = 16'(5763);
			498: out = 16'(-262);
			499: out = 16'(5216);
			500: out = 16'(217);
			501: out = 16'(-4668);
			502: out = 16'(-8326);
			503: out = 16'(-7257);
			504: out = 16'(3321);
			505: out = 16'(-464);
			506: out = 16'(-13599);
			507: out = 16'(-10683);
			508: out = 16'(-12786);
			509: out = 16'(7983);
			510: out = 16'(-10266);
			511: out = 16'(-4557);
			512: out = 16'(2252);
			513: out = 16'(-7970);
			514: out = 16'(-12228);
			515: out = 16'(-1070);
			516: out = 16'(1759);
			517: out = 16'(-9468);
			518: out = 16'(985);
			519: out = 16'(-12860);
			520: out = 16'(-7906);
			521: out = 16'(-16538);
			522: out = 16'(-6847);
			523: out = 16'(-3882);
			524: out = 16'(-11561);
			525: out = 16'(-10818);
			526: out = 16'(-16795);
			527: out = 16'(-6781);
			528: out = 16'(-10541);
			529: out = 16'(-15642);
			530: out = 16'(-8367);
			531: out = 16'(-3960);
			532: out = 16'(-9723);
			533: out = 16'(-1043);
			534: out = 16'(-13867);
			535: out = 16'(-9242);
			536: out = 16'(-8076);
			537: out = 16'(-4760);
			538: out = 16'(-4133);
			539: out = 16'(9146);
			540: out = 16'(-3671);
			541: out = 16'(-8797);
			542: out = 16'(-7086);
			543: out = 16'(3708);
			544: out = 16'(9571);
			545: out = 16'(-4379);
			546: out = 16'(13447);
			547: out = 16'(-3361);
			548: out = 16'(-2642);
			549: out = 16'(15937);
			550: out = 16'(-1705);
			551: out = 16'(4148);
			552: out = 16'(2239);
			553: out = 16'(-2662);
			554: out = 16'(5794);
			555: out = 16'(3265);
			556: out = 16'(7572);
			557: out = 16'(5633);
			558: out = 16'(11165);
			559: out = 16'(14392);
			560: out = 16'(2789);
			561: out = 16'(8155);
			562: out = 16'(794);
			563: out = 16'(14619);
			564: out = 16'(21077);
			565: out = 16'(6369);
			566: out = 16'(11230);
			567: out = 16'(12726);
			568: out = 16'(5679);
			569: out = 16'(16053);
			570: out = 16'(3638);
			571: out = 16'(9149);
			572: out = 16'(-2392);
			573: out = 16'(14084);
			574: out = 16'(13985);
			575: out = 16'(13495);
			576: out = 16'(1415);
			577: out = 16'(4334);
			578: out = 16'(8994);
			579: out = 16'(9708);
			580: out = 16'(5681);
			581: out = 16'(-685);
			582: out = 16'(8597);
			583: out = 16'(-11309);
			584: out = 16'(11311);
			585: out = 16'(-1384);
			586: out = 16'(-1271);
			587: out = 16'(-586);
			588: out = 16'(-449);
			589: out = 16'(3252);
			590: out = 16'(9040);
			591: out = 16'(8060);
			592: out = 16'(-7123);
			593: out = 16'(4130);
			594: out = 16'(-9372);
			595: out = 16'(-6630);
			596: out = 16'(-5331);
			597: out = 16'(-1089);
			598: out = 16'(4754);
			599: out = 16'(6674);
			600: out = 16'(-2822);
			601: out = 16'(-3751);
			602: out = 16'(-9550);
			603: out = 16'(-20642);
			604: out = 16'(-4561);
			605: out = 16'(8676);
			606: out = 16'(-6684);
			607: out = 16'(-6450);
			608: out = 16'(-5507);
			609: out = 16'(-4826);
			610: out = 16'(-4996);
			611: out = 16'(-25989);
			612: out = 16'(-3405);
			613: out = 16'(-901);
			614: out = 16'(-4031);
			615: out = 16'(-5724);
			616: out = 16'(-4069);
			617: out = 16'(829);
			618: out = 16'(-4565);
			619: out = 16'(-10570);
			620: out = 16'(-243);
			621: out = 16'(-3251);
			622: out = 16'(-1322);
			623: out = 16'(-20853);
			624: out = 16'(4430);
			625: out = 16'(9441);
			626: out = 16'(-7861);
			627: out = 16'(6224);
			628: out = 16'(-5172);
			629: out = 16'(3281);
			630: out = 16'(4021);
			631: out = 16'(-5683);
			632: out = 16'(4190);
			633: out = 16'(6189);
			634: out = 16'(2283);
			635: out = 16'(8661);
			636: out = 16'(3020);
			637: out = 16'(8856);
			638: out = 16'(6425);
			639: out = 16'(8220);
			640: out = 16'(-3271);
			641: out = 16'(3268);
			642: out = 16'(6198);
			643: out = 16'(2786);
			644: out = 16'(-4075);
			645: out = 16'(2315);
			646: out = 16'(-1956);
			647: out = 16'(-2415);
			648: out = 16'(4286);
			649: out = 16'(-6525);
			650: out = 16'(5681);
			651: out = 16'(21060);
			652: out = 16'(8723);
			653: out = 16'(-2165);
			654: out = 16'(-8121);
			655: out = 16'(15900);
			656: out = 16'(3367);
			657: out = 16'(8216);
			658: out = 16'(8196);
			659: out = 16'(-2053);
			660: out = 16'(-1534);
			661: out = 16'(-6082);
			662: out = 16'(11905);
			663: out = 16'(-2489);
			664: out = 16'(-5934);
			665: out = 16'(12642);
			666: out = 16'(-11071);
			667: out = 16'(11386);
			668: out = 16'(-3803);
			669: out = 16'(3752);
			670: out = 16'(11799);
			671: out = 16'(-2638);
			672: out = 16'(1366);
			673: out = 16'(7846);
			674: out = 16'(-1070);
			675: out = 16'(-4983);
			676: out = 16'(5426);
			677: out = 16'(4566);
			678: out = 16'(-1917);
			679: out = 16'(-3262);
			680: out = 16'(12855);
			681: out = 16'(-3737);
			682: out = 16'(-3444);
			683: out = 16'(-757);
			684: out = 16'(-4808);
			685: out = 16'(-4646);
			686: out = 16'(2828);
			687: out = 16'(-3643);
			688: out = 16'(-4613);
			689: out = 16'(8965);
			690: out = 16'(-4053);
			691: out = 16'(2882);
			692: out = 16'(-3139);
			693: out = 16'(-18772);
			694: out = 16'(-1470);
			695: out = 16'(7507);
			696: out = 16'(2899);
			697: out = 16'(-9511);
			698: out = 16'(-4724);
			699: out = 16'(-3408);
			700: out = 16'(1101);
			701: out = 16'(6810);
			702: out = 16'(-6971);
			703: out = 16'(-3100);
			704: out = 16'(-5757);
			705: out = 16'(4506);
			706: out = 16'(-14518);
			707: out = 16'(-7484);
			708: out = 16'(-7593);
			709: out = 16'(-10965);
			710: out = 16'(16490);
			711: out = 16'(-12738);
			712: out = 16'(4616);
			713: out = 16'(1312);
			714: out = 16'(-18183);
			715: out = 16'(10007);
			716: out = 16'(-432);
			717: out = 16'(3829);
			718: out = 16'(-8285);
			719: out = 16'(1324);
			720: out = 16'(-606);
			721: out = 16'(-3432);
			722: out = 16'(-6971);
			723: out = 16'(-2299);
			724: out = 16'(6000);
			725: out = 16'(-9698);
			726: out = 16'(-145);
			727: out = 16'(5564);
			728: out = 16'(3647);
			729: out = 16'(-6675);
			730: out = 16'(-6807);
			731: out = 16'(-6742);
			732: out = 16'(-684);
			733: out = 16'(-1899);
			734: out = 16'(1287);
			735: out = 16'(15406);
			736: out = 16'(-5845);
			737: out = 16'(6321);
			738: out = 16'(8217);
			739: out = 16'(-11143);
			740: out = 16'(872);
			741: out = 16'(11785);
			742: out = 16'(-1901);
			743: out = 16'(-2311);
			744: out = 16'(-471);
			745: out = 16'(800);
			746: out = 16'(2500);
			747: out = 16'(-6597);
			748: out = 16'(11929);
			749: out = 16'(-10365);
			750: out = 16'(2863);
			751: out = 16'(-2745);
			752: out = 16'(10889);
			753: out = 16'(19673);
			754: out = 16'(-7392);
			755: out = 16'(9268);
			756: out = 16'(-215);
			757: out = 16'(-5079);
			758: out = 16'(12451);
			759: out = 16'(23236);
			760: out = 16'(124);
			761: out = 16'(1223);
			762: out = 16'(1647);
			763: out = 16'(10603);
			764: out = 16'(-621);
			765: out = 16'(10899);
			766: out = 16'(12101);
			767: out = 16'(-8003);
			768: out = 16'(-183);
			769: out = 16'(-2325);
			770: out = 16'(-1664);
			771: out = 16'(-1322);
			772: out = 16'(-581);
			773: out = 16'(-6103);
			774: out = 16'(7657);
			775: out = 16'(7361);
			776: out = 16'(-4285);
			777: out = 16'(8175);
			778: out = 16'(1824);
			779: out = 16'(-14907);
			780: out = 16'(-455);
			781: out = 16'(11993);
			782: out = 16'(-11674);
			783: out = 16'(1627);
			784: out = 16'(-4730);
			785: out = 16'(-8705);
			786: out = 16'(10542);
			787: out = 16'(2401);
			788: out = 16'(-10119);
			789: out = 16'(-2458);
			790: out = 16'(-11612);
			791: out = 16'(6754);
			792: out = 16'(10661);
			793: out = 16'(-14867);
			794: out = 16'(-2477);
			795: out = 16'(3656);
			796: out = 16'(-7357);
			797: out = 16'(-17651);
			798: out = 16'(9754);
			799: out = 16'(-10021);
			800: out = 16'(10170);
			801: out = 16'(9465);
			802: out = 16'(-8069);
			803: out = 16'(-12784);
			804: out = 16'(770);
			805: out = 16'(-3258);
			806: out = 16'(3204);
			807: out = 16'(-5143);
			808: out = 16'(-1934);
			809: out = 16'(-2117);
			810: out = 16'(-751);
			811: out = 16'(-7530);
			812: out = 16'(-3167);
			813: out = 16'(-9928);
			814: out = 16'(-3360);
			815: out = 16'(1910);
			816: out = 16'(4368);
			817: out = 16'(2747);
			818: out = 16'(1893);
			819: out = 16'(3140);
			820: out = 16'(4027);
			821: out = 16'(-6838);
			822: out = 16'(14326);
			823: out = 16'(12206);
			824: out = 16'(-10076);
			825: out = 16'(-7260);
			826: out = 16'(10626);
			827: out = 16'(-5391);
			828: out = 16'(-602);
			829: out = 16'(-2188);
			830: out = 16'(-2346);
			831: out = 16'(12531);
			832: out = 16'(-8609);
			833: out = 16'(4845);
			834: out = 16'(-16043);
			835: out = 16'(-795);
			836: out = 16'(15005);
			837: out = 16'(2101);
			838: out = 16'(435);
			839: out = 16'(5231);
			840: out = 16'(4263);
			841: out = 16'(-11712);
			842: out = 16'(-2164);
			843: out = 16'(9053);
			844: out = 16'(-7588);
			845: out = 16'(9684);
			846: out = 16'(8236);
			847: out = 16'(-9038);
			848: out = 16'(6674);
			849: out = 16'(-3396);
			850: out = 16'(-354);
			851: out = 16'(3924);
			852: out = 16'(3500);
			853: out = 16'(-186);
			854: out = 16'(-14617);
			855: out = 16'(-1649);
			856: out = 16'(1532);
			857: out = 16'(3985);
			858: out = 16'(-15463);
			859: out = 16'(1549);
			860: out = 16'(-2635);
			861: out = 16'(3460);
			862: out = 16'(8452);
			863: out = 16'(-6787);
			864: out = 16'(-2815);
			865: out = 16'(-10314);
			866: out = 16'(12774);
			867: out = 16'(-1418);
			868: out = 16'(-6818);
			869: out = 16'(-7011);
			870: out = 16'(-10556);
			871: out = 16'(1056);
			872: out = 16'(-5992);
			873: out = 16'(-6513);
			874: out = 16'(1154);
			875: out = 16'(1731);
			876: out = 16'(-7169);
			877: out = 16'(3064);
			878: out = 16'(8924);
			879: out = 16'(-936);
			880: out = 16'(1885);
			881: out = 16'(-2000);
			882: out = 16'(10294);
			883: out = 16'(-20069);
			884: out = 16'(684);
			885: out = 16'(14427);
			886: out = 16'(2892);
			887: out = 16'(3846);
			888: out = 16'(-497);
			889: out = 16'(-7742);
			890: out = 16'(131);
			891: out = 16'(-3077);
			892: out = 16'(2074);
			893: out = 16'(3086);
			894: out = 16'(-258);
			895: out = 16'(-806);
			896: out = 16'(6660);
			897: out = 16'(-4599);
			898: out = 16'(-11319);
			899: out = 16'(2201);
			900: out = 16'(-10208);
			901: out = 16'(19575);
			902: out = 16'(-333);
			903: out = 16'(105);
			904: out = 16'(-9941);
			905: out = 16'(3286);
			906: out = 16'(-10188);
			907: out = 16'(-260);
			908: out = 16'(11334);
			909: out = 16'(-2326);
			910: out = 16'(-1712);
			911: out = 16'(11495);
			912: out = 16'(-6542);
			913: out = 16'(-1518);
			914: out = 16'(-9201);
			915: out = 16'(5759);
			916: out = 16'(-1452);
			917: out = 16'(2380);
			918: out = 16'(-689);
			919: out = 16'(3928);
			920: out = 16'(-582);
			921: out = 16'(-3403);
			922: out = 16'(15161);
			923: out = 16'(-1398);
			924: out = 16'(10468);
			925: out = 16'(-1388);
			926: out = 16'(-4435);
			927: out = 16'(-4296);
			928: out = 16'(8362);
			929: out = 16'(3147);
			930: out = 16'(4432);
			931: out = 16'(-2432);
			932: out = 16'(13922);
			933: out = 16'(11558);
			934: out = 16'(3165);
			935: out = 16'(3599);
			936: out = 16'(-740);
			937: out = 16'(8936);
			938: out = 16'(693);
			939: out = 16'(6179);
			940: out = 16'(-8425);
			941: out = 16'(14117);
			942: out = 16'(-1376);
			943: out = 16'(6597);
			944: out = 16'(-5458);
			945: out = 16'(-1768);
			946: out = 16'(-8767);
			947: out = 16'(2588);
			948: out = 16'(-12771);
			949: out = 16'(11214);
			950: out = 16'(10290);
			951: out = 16'(-359);
			952: out = 16'(446);
			953: out = 16'(-5560);
			954: out = 16'(8490);
			955: out = 16'(-5647);
			956: out = 16'(-3670);
			957: out = 16'(-14522);
			958: out = 16'(14405);
			959: out = 16'(3123);
			960: out = 16'(-7464);
			961: out = 16'(-6426);
			962: out = 16'(-3388);
			963: out = 16'(8848);
			964: out = 16'(12486);
			965: out = 16'(299);
			966: out = 16'(-14177);
			967: out = 16'(2690);
			968: out = 16'(-9190);
			969: out = 16'(6426);
			970: out = 16'(632);
			971: out = 16'(12286);
			972: out = 16'(-2404);
			973: out = 16'(-259);
			974: out = 16'(3991);
			975: out = 16'(-5970);
			976: out = 16'(-6677);
			977: out = 16'(-5342);
			978: out = 16'(-2128);
			979: out = 16'(-4355);
			980: out = 16'(3975);
			981: out = 16'(-502);
			982: out = 16'(1597);
			983: out = 16'(-909);
			984: out = 16'(-945);
			985: out = 16'(2333);
			986: out = 16'(-5834);
			987: out = 16'(-16005);
			988: out = 16'(19352);
			989: out = 16'(-6496);
			990: out = 16'(-3973);
			991: out = 16'(-6964);
			992: out = 16'(-484);
			993: out = 16'(1300);
			994: out = 16'(2160);
			995: out = 16'(-2250);
			996: out = 16'(-4792);
			997: out = 16'(1716);
			998: out = 16'(2095);
			999: out = 16'(-5767);
			1000: out = 16'(1190);
			1001: out = 16'(-5922);
			1002: out = 16'(-625);
			1003: out = 16'(6051);
			1004: out = 16'(2244);
			1005: out = 16'(11318);
			1006: out = 16'(-6974);
			1007: out = 16'(-6496);
			1008: out = 16'(-4080);
			1009: out = 16'(-4000);
			1010: out = 16'(-14713);
			1011: out = 16'(2313);
			1012: out = 16'(1532);
			1013: out = 16'(-6203);
			1014: out = 16'(11053);
			1015: out = 16'(4560);
			1016: out = 16'(-1398);
			1017: out = 16'(4297);
			1018: out = 16'(2198);
			1019: out = 16'(7050);
			1020: out = 16'(-184);
			1021: out = 16'(-4682);
			1022: out = 16'(-2685);
			1023: out = 16'(629);
			1024: out = 16'(4551);
			1025: out = 16'(4592);
			1026: out = 16'(7361);
			1027: out = 16'(-5536);
			1028: out = 16'(-3722);
			1029: out = 16'(-4066);
			1030: out = 16'(8879);
			1031: out = 16'(-7085);
			1032: out = 16'(5467);
			1033: out = 16'(419);
			1034: out = 16'(-178);
			1035: out = 16'(-8101);
			1036: out = 16'(2900);
			1037: out = 16'(-7688);
			1038: out = 16'(-12509);
			1039: out = 16'(1643);
			1040: out = 16'(3063);
			1041: out = 16'(1914);
			1042: out = 16'(-178);
			1043: out = 16'(-448);
			1044: out = 16'(-11147);
			1045: out = 16'(-9766);
			1046: out = 16'(-243);
			1047: out = 16'(9471);
			1048: out = 16'(-7627);
			1049: out = 16'(-4957);
			1050: out = 16'(2886);
			1051: out = 16'(5423);
			1052: out = 16'(4375);
			1053: out = 16'(7131);
			1054: out = 16'(-15223);
			1055: out = 16'(5981);
			1056: out = 16'(-5344);
			1057: out = 16'(1158);
			1058: out = 16'(8567);
			1059: out = 16'(-932);
			1060: out = 16'(5476);
			1061: out = 16'(1317);
			1062: out = 16'(3454);
			1063: out = 16'(5924);
			1064: out = 16'(-13283);
			1065: out = 16'(-944);
			1066: out = 16'(-708);
			1067: out = 16'(-5018);
			1068: out = 16'(-3577);
			1069: out = 16'(-3821);
			1070: out = 16'(-14715);
			1071: out = 16'(9750);
			1072: out = 16'(2711);
			1073: out = 16'(9399);
			1074: out = 16'(-238);
			1075: out = 16'(-2521);
			1076: out = 16'(445);
			1077: out = 16'(-5855);
			1078: out = 16'(-11273);
			1079: out = 16'(5215);
			1080: out = 16'(-6098);
			1081: out = 16'(928);
			1082: out = 16'(-12997);
			1083: out = 16'(6398);
			1084: out = 16'(-1234);
			1085: out = 16'(-3608);
			1086: out = 16'(4100);
			1087: out = 16'(-3634);
			1088: out = 16'(685);
			1089: out = 16'(-10080);
			1090: out = 16'(9219);
			1091: out = 16'(8081);
			1092: out = 16'(-9073);
			1093: out = 16'(-6588);
			1094: out = 16'(9405);
			1095: out = 16'(2825);
			1096: out = 16'(7374);
			1097: out = 16'(-6665);
			1098: out = 16'(1713);
			1099: out = 16'(-1419);
			1100: out = 16'(7321);
			1101: out = 16'(-9836);
			1102: out = 16'(-3792);
			1103: out = 16'(-3063);
			1104: out = 16'(6277);
			1105: out = 16'(1362);
			1106: out = 16'(3672);
			1107: out = 16'(2770);
			1108: out = 16'(32);
			1109: out = 16'(6975);
			1110: out = 16'(4122);
			1111: out = 16'(34);
			1112: out = 16'(-875);
			1113: out = 16'(8989);
			1114: out = 16'(-719);
			1115: out = 16'(-8337);
			1116: out = 16'(-142);
			1117: out = 16'(-5932);
			1118: out = 16'(8506);
			1119: out = 16'(-170);
			1120: out = 16'(-5120);
			1121: out = 16'(1404);
			1122: out = 16'(-9065);
			1123: out = 16'(-2553);
			1124: out = 16'(-8811);
			1125: out = 16'(1768);
			1126: out = 16'(-8636);
			1127: out = 16'(337);
			1128: out = 16'(6451);
			1129: out = 16'(10190);
			1130: out = 16'(523);
			1131: out = 16'(277);
			1132: out = 16'(1348);
			1133: out = 16'(-3677);
			1134: out = 16'(3418);
			1135: out = 16'(-6001);
			1136: out = 16'(3224);
			1137: out = 16'(-9454);
			1138: out = 16'(5877);
			1139: out = 16'(-6318);
			1140: out = 16'(525);
			1141: out = 16'(-1320);
			1142: out = 16'(-342);
			1143: out = 16'(11775);
			1144: out = 16'(-3122);
			1145: out = 16'(-5131);
			1146: out = 16'(7194);
			1147: out = 16'(-11433);
			1148: out = 16'(9141);
			1149: out = 16'(-5327);
			1150: out = 16'(-4340);
			1151: out = 16'(12056);
			1152: out = 16'(2471);
			1153: out = 16'(-2426);
			1154: out = 16'(2594);
			1155: out = 16'(-12847);
			1156: out = 16'(-3877);
			1157: out = 16'(14591);
			1158: out = 16'(-1474);
			1159: out = 16'(-3397);
			1160: out = 16'(-13233);
			1161: out = 16'(7131);
			1162: out = 16'(-8941);
			1163: out = 16'(-9199);
			1164: out = 16'(-6178);
			1165: out = 16'(1784);
			1166: out = 16'(-3646);
			1167: out = 16'(1405);
			1168: out = 16'(10399);
			1169: out = 16'(-5176);
			1170: out = 16'(-1749);
			1171: out = 16'(10720);
			1172: out = 16'(6708);
			1173: out = 16'(-655);
			1174: out = 16'(3258);
			1175: out = 16'(-11623);
			1176: out = 16'(12633);
			1177: out = 16'(8259);
			1178: out = 16'(-6284);
			1179: out = 16'(-8418);
			1180: out = 16'(2443);
			1181: out = 16'(433);
			1182: out = 16'(-9348);
			1183: out = 16'(-358);
			1184: out = 16'(-740);
			1185: out = 16'(6298);
			1186: out = 16'(6821);
			1187: out = 16'(-891);
			1188: out = 16'(4835);
			1189: out = 16'(-6556);
			1190: out = 16'(-4006);
			1191: out = 16'(1215);
			1192: out = 16'(3025);
			1193: out = 16'(5683);
			1194: out = 16'(-920);
			1195: out = 16'(-309);
			1196: out = 16'(1994);
			1197: out = 16'(-15305);
			1198: out = 16'(12000);
			1199: out = 16'(12393);
			1200: out = 16'(-2379);
			1201: out = 16'(-8327);
			1202: out = 16'(4886);
			1203: out = 16'(-508);
			1204: out = 16'(-9562);
			1205: out = 16'(4992);
			1206: out = 16'(1772);
			1207: out = 16'(2937);
			1208: out = 16'(-7589);
			1209: out = 16'(5929);
			1210: out = 16'(2634);
			1211: out = 16'(-11395);
			1212: out = 16'(12);
			1213: out = 16'(4673);
			1214: out = 16'(4592);
			1215: out = 16'(-759);
			1216: out = 16'(7204);
			1217: out = 16'(-15096);
			1218: out = 16'(3026);
			1219: out = 16'(-829);
			1220: out = 16'(-5785);
			1221: out = 16'(-2180);
			1222: out = 16'(1984);
			1223: out = 16'(7542);
			1224: out = 16'(874);
			1225: out = 16'(-8120);
			1226: out = 16'(-4112);
			1227: out = 16'(11535);
			1228: out = 16'(-4232);
			1229: out = 16'(-6309);
			1230: out = 16'(5406);
			1231: out = 16'(10575);
			1232: out = 16'(-579);
			1233: out = 16'(-56);
			1234: out = 16'(3745);
			1235: out = 16'(-7041);
			1236: out = 16'(1557);
			1237: out = 16'(-2478);
			1238: out = 16'(-5024);
			1239: out = 16'(3296);
			1240: out = 16'(7833);
			1241: out = 16'(-2776);
			1242: out = 16'(1588);
			1243: out = 16'(-5379);
			1244: out = 16'(-3017);
			1245: out = 16'(-4920);
			1246: out = 16'(3894);
			1247: out = 16'(-8919);
			1248: out = 16'(4058);
			1249: out = 16'(-1349);
			1250: out = 16'(11571);
			1251: out = 16'(-1519);
			1252: out = 16'(7857);
			1253: out = 16'(5340);
			1254: out = 16'(-2808);
			1255: out = 16'(-4354);
			1256: out = 16'(-8464);
			1257: out = 16'(5027);
			1258: out = 16'(8354);
			1259: out = 16'(-1550);
			1260: out = 16'(-3958);
			1261: out = 16'(1425);
			1262: out = 16'(1808);
			1263: out = 16'(-4934);
			1264: out = 16'(-2288);
			1265: out = 16'(-10906);
			1266: out = 16'(3792);
			1267: out = 16'(972);
			1268: out = 16'(-932);
			1269: out = 16'(-1611);
			1270: out = 16'(-3960);
			1271: out = 16'(8789);
			1272: out = 16'(3328);
			1273: out = 16'(-3866);
			1274: out = 16'(-2708);
			1275: out = 16'(-6229);
			1276: out = 16'(3783);
			1277: out = 16'(-5976);
			1278: out = 16'(-2127);
			1279: out = 16'(4610);
			1280: out = 16'(-4418);
			1281: out = 16'(5932);
			1282: out = 16'(-4601);
			1283: out = 16'(-1012);
			1284: out = 16'(-7968);
			1285: out = 16'(2015);
			1286: out = 16'(7309);
			1287: out = 16'(-1480);
			1288: out = 16'(-2119);
			1289: out = 16'(-1448);
			1290: out = 16'(-6293);
			1291: out = 16'(-4391);
			1292: out = 16'(3498);
			1293: out = 16'(4559);
			1294: out = 16'(-8285);
			1295: out = 16'(11337);
			1296: out = 16'(-8722);
			1297: out = 16'(-2046);
			1298: out = 16'(12276);
			1299: out = 16'(6083);
			1300: out = 16'(3625);
			1301: out = 16'(-926);
			1302: out = 16'(-77);
			1303: out = 16'(-3705);
			1304: out = 16'(3304);
			1305: out = 16'(-2006);
			1306: out = 16'(5442);
			1307: out = 16'(-6528);
			1308: out = 16'(13203);
			1309: out = 16'(5550);
			1310: out = 16'(-4246);
			1311: out = 16'(-4608);
			1312: out = 16'(5960);
			1313: out = 16'(-2823);
			1314: out = 16'(1442);
			1315: out = 16'(-1229);
			1316: out = 16'(-795);
			1317: out = 16'(-337);
			1318: out = 16'(2926);
			1319: out = 16'(-668);
			1320: out = 16'(-842);
			1321: out = 16'(-7212);
			1322: out = 16'(2639);
			1323: out = 16'(-7508);
			1324: out = 16'(13702);
			1325: out = 16'(4881);
			1326: out = 16'(-9201);
			1327: out = 16'(1901);
			1328: out = 16'(-6820);
			1329: out = 16'(584);
			1330: out = 16'(-2463);
			1331: out = 16'(-12488);
			1332: out = 16'(-1893);
			1333: out = 16'(2082);
			1334: out = 16'(-3052);
			1335: out = 16'(-8489);
			1336: out = 16'(7289);
			1337: out = 16'(-8309);
			1338: out = 16'(6587);
			1339: out = 16'(-3130);
			1340: out = 16'(-15586);
			1341: out = 16'(3556);
			1342: out = 16'(10727);
			1343: out = 16'(-3583);
			1344: out = 16'(-8903);
			1345: out = 16'(1196);
			1346: out = 16'(2284);
			1347: out = 16'(-5510);
			1348: out = 16'(8870);
			1349: out = 16'(-8654);
			1350: out = 16'(-3968);
			1351: out = 16'(3951);
			1352: out = 16'(5664);
			1353: out = 16'(-5935);
			1354: out = 16'(-5227);
			1355: out = 16'(3653);
			1356: out = 16'(-216);
			1357: out = 16'(-4855);
			1358: out = 16'(-4640);
			1359: out = 16'(-1084);
			1360: out = 16'(205);
			1361: out = 16'(-6314);
			1362: out = 16'(-1582);
			1363: out = 16'(3683);
			1364: out = 16'(1436);
			1365: out = 16'(-16063);
			1366: out = 16'(9166);
			1367: out = 16'(2533);
			1368: out = 16'(-2563);
			1369: out = 16'(-3056);
			1370: out = 16'(4694);
			1371: out = 16'(-9587);
			1372: out = 16'(5358);
			1373: out = 16'(-6133);
			1374: out = 16'(-4016);
			1375: out = 16'(5428);
			1376: out = 16'(-2278);
			1377: out = 16'(-1997);
			1378: out = 16'(-452);
			1379: out = 16'(-1011);
			1380: out = 16'(-7733);
			1381: out = 16'(9256);
			1382: out = 16'(6144);
			1383: out = 16'(-2466);
			1384: out = 16'(9249);
			1385: out = 16'(-3350);
			1386: out = 16'(3229);
			1387: out = 16'(-1006);
			1388: out = 16'(-2214);
			1389: out = 16'(-6688);
			1390: out = 16'(-1091);
			1391: out = 16'(8102);
			1392: out = 16'(-1379);
			1393: out = 16'(972);
			1394: out = 16'(-4097);
			1395: out = 16'(-814);
			1396: out = 16'(-14777);
			1397: out = 16'(10807);
			1398: out = 16'(-537);
			1399: out = 16'(8444);
			1400: out = 16'(9949);
			1401: out = 16'(-1310);
			1402: out = 16'(7287);
			1403: out = 16'(-7456);
			1404: out = 16'(-6737);
			1405: out = 16'(9934);
			1406: out = 16'(-811);
			1407: out = 16'(2770);
			1408: out = 16'(1407);
			1409: out = 16'(2543);
			1410: out = 16'(-4447);
			1411: out = 16'(-3704);
			1412: out = 16'(-17129);
			1413: out = 16'(11324);
			1414: out = 16'(-4482);
			1415: out = 16'(-9190);
			1416: out = 16'(6503);
			1417: out = 16'(1795);
			1418: out = 16'(-594);
			1419: out = 16'(6667);
			1420: out = 16'(-2868);
			1421: out = 16'(-217);
			1422: out = 16'(835);
			1423: out = 16'(-13570);
			1424: out = 16'(8354);
			1425: out = 16'(-838);
			1426: out = 16'(2140);
			1427: out = 16'(1105);
			1428: out = 16'(1762);
			1429: out = 16'(-4631);
			1430: out = 16'(1725);
			1431: out = 16'(43);
			1432: out = 16'(7254);
			1433: out = 16'(1071);
			1434: out = 16'(-4662);
			1435: out = 16'(-4390);
			1436: out = 16'(5654);
			1437: out = 16'(-8753);
			1438: out = 16'(673);
			1439: out = 16'(-3568);
			1440: out = 16'(4411);
			1441: out = 16'(-12881);
			1442: out = 16'(-5516);
			1443: out = 16'(1386);
			1444: out = 16'(696);
			1445: out = 16'(7321);
			1446: out = 16'(-11174);
			1447: out = 16'(11460);
			1448: out = 16'(2368);
			1449: out = 16'(-10143);
			1450: out = 16'(577);
			1451: out = 16'(2089);
			1452: out = 16'(5790);
			1453: out = 16'(-4760);
			1454: out = 16'(-6136);
			1455: out = 16'(4955);
			1456: out = 16'(-2889);
			1457: out = 16'(2823);
			1458: out = 16'(9366);
			1459: out = 16'(1126);
			1460: out = 16'(-470);
			1461: out = 16'(-1030);
			1462: out = 16'(2569);
			1463: out = 16'(807);
			1464: out = 16'(-1045);
			1465: out = 16'(-5982);
			1466: out = 16'(-2531);
			1467: out = 16'(7904);
			1468: out = 16'(10418);
			1469: out = 16'(3507);
			1470: out = 16'(-4847);
			1471: out = 16'(-3814);
			1472: out = 16'(-1155);
			1473: out = 16'(725);
			1474: out = 16'(-699);
			1475: out = 16'(8673);
			1476: out = 16'(-6179);
			1477: out = 16'(-6079);
			1478: out = 16'(1956);
			1479: out = 16'(5260);
			1480: out = 16'(-5529);
			1481: out = 16'(10578);
			1482: out = 16'(-629);
			1483: out = 16'(4681);
			1484: out = 16'(774);
			1485: out = 16'(1970);
			1486: out = 16'(-1621);
			1487: out = 16'(14015);
			1488: out = 16'(1158);
			1489: out = 16'(-1373);
			1490: out = 16'(950);
			1491: out = 16'(-7512);
			1492: out = 16'(9420);
			1493: out = 16'(1840);
			1494: out = 16'(1365);
			1495: out = 16'(-4098);
			1496: out = 16'(4732);
			1497: out = 16'(2768);
			1498: out = 16'(1455);
			1499: out = 16'(-3762);
			1500: out = 16'(-2745);
			1501: out = 16'(5447);
			1502: out = 16'(-681);
			1503: out = 16'(-5624);
			1504: out = 16'(-6181);
			1505: out = 16'(8008);
			1506: out = 16'(-3123);
			1507: out = 16'(-2514);
			1508: out = 16'(-2340);
			1509: out = 16'(-1365);
			1510: out = 16'(-1143);
			1511: out = 16'(-5221);
			1512: out = 16'(9505);
			1513: out = 16'(-989);
			1514: out = 16'(-5702);
			1515: out = 16'(-3570);
			1516: out = 16'(4165);
			1517: out = 16'(1675);
			1518: out = 16'(-210);
			1519: out = 16'(-11308);
			1520: out = 16'(187);
			1521: out = 16'(-2893);
			1522: out = 16'(-179);
			1523: out = 16'(1200);
			1524: out = 16'(2371);
			1525: out = 16'(-10485);
			1526: out = 16'(-1331);
			1527: out = 16'(-1598);
			1528: out = 16'(-1635);
			1529: out = 16'(978);
			1530: out = 16'(-5140);
			1531: out = 16'(6661);
			1532: out = 16'(-1628);
			1533: out = 16'(-2922);
			1534: out = 16'(5497);
			1535: out = 16'(-8614);
			1536: out = 16'(-4590);
			1537: out = 16'(1049);
			1538: out = 16'(-4273);
			1539: out = 16'(-8174);
			1540: out = 16'(3819);
			1541: out = 16'(3286);
			1542: out = 16'(1427);
			1543: out = 16'(3649);
			1544: out = 16'(-5133);
			1545: out = 16'(-3975);
			1546: out = 16'(4544);
			1547: out = 16'(-5042);
			1548: out = 16'(4206);
			1549: out = 16'(9193);
			1550: out = 16'(-4595);
			1551: out = 16'(754);
			1552: out = 16'(2316);
			1553: out = 16'(-3630);
			1554: out = 16'(3607);
			1555: out = 16'(1443);
			1556: out = 16'(-6678);
			1557: out = 16'(-682);
			1558: out = 16'(237);
			1559: out = 16'(-2095);
			1560: out = 16'(-3321);
			1561: out = 16'(-1744);
			1562: out = 16'(3452);
			1563: out = 16'(-2503);
			1564: out = 16'(694);
			1565: out = 16'(7239);
			1566: out = 16'(-8698);
			1567: out = 16'(2944);
			1568: out = 16'(-1085);
			1569: out = 16'(-1620);
			1570: out = 16'(-2568);
			1571: out = 16'(7782);
			1572: out = 16'(4978);
			1573: out = 16'(847);
			1574: out = 16'(4454);
			1575: out = 16'(-1583);
			1576: out = 16'(-6343);
			1577: out = 16'(1723);
			1578: out = 16'(-2831);
			1579: out = 16'(5234);
			1580: out = 16'(3413);
			1581: out = 16'(1456);
			1582: out = 16'(-5174);
			1583: out = 16'(-1919);
			1584: out = 16'(3052);
			1585: out = 16'(-8233);
			1586: out = 16'(2488);
			1587: out = 16'(2663);
			1588: out = 16'(1349);
			1589: out = 16'(-5545);
			1590: out = 16'(6032);
			1591: out = 16'(-702);
			1592: out = 16'(1818);
			1593: out = 16'(5921);
			1594: out = 16'(686);
			1595: out = 16'(193);
			1596: out = 16'(-2970);
			1597: out = 16'(1890);
			1598: out = 16'(3332);
			1599: out = 16'(4721);
			1600: out = 16'(-4302);
			1601: out = 16'(-4341);
			1602: out = 16'(1376);
			1603: out = 16'(-4942);
			1604: out = 16'(9785);
			1605: out = 16'(5483);
			1606: out = 16'(-989);
			1607: out = 16'(-6863);
			1608: out = 16'(1287);
			1609: out = 16'(840);
			1610: out = 16'(-4048);
			1611: out = 16'(-1432);
			1612: out = 16'(5782);
			1613: out = 16'(-2372);
			1614: out = 16'(-6639);
			1615: out = 16'(1912);
			1616: out = 16'(-9104);
			1617: out = 16'(4883);
			1618: out = 16'(466);
			1619: out = 16'(4475);
			1620: out = 16'(3370);
			1621: out = 16'(4121);
			1622: out = 16'(-1220);
			1623: out = 16'(3679);
			1624: out = 16'(617);
			1625: out = 16'(-4431);
			1626: out = 16'(-356);
			1627: out = 16'(-6889);
			1628: out = 16'(6305);
			1629: out = 16'(447);
			1630: out = 16'(4188);
			1631: out = 16'(324);
			1632: out = 16'(-5699);
			1633: out = 16'(-5647);
			1634: out = 16'(981);
			1635: out = 16'(267);
			1636: out = 16'(1748);
			1637: out = 16'(-3041);
			1638: out = 16'(-5134);
			1639: out = 16'(4851);
			1640: out = 16'(811);
			1641: out = 16'(1915);
			1642: out = 16'(-6374);
			1643: out = 16'(129);
			1644: out = 16'(1251);
			1645: out = 16'(-5720);
			1646: out = 16'(7870);
			1647: out = 16'(5936);
			1648: out = 16'(-3949);
			1649: out = 16'(-5680);
			1650: out = 16'(2239);
			1651: out = 16'(-2436);
			1652: out = 16'(5038);
			1653: out = 16'(839);
			1654: out = 16'(-550);
			1655: out = 16'(-11524);
			1656: out = 16'(7693);
			1657: out = 16'(684);
			1658: out = 16'(-1796);
			1659: out = 16'(-10781);
			1660: out = 16'(6813);
			1661: out = 16'(241);
			1662: out = 16'(-2235);
			1663: out = 16'(4812);
			1664: out = 16'(1061);
			1665: out = 16'(-2284);
			1666: out = 16'(5309);
			1667: out = 16'(-2291);
			1668: out = 16'(865);
			1669: out = 16'(-172);
			1670: out = 16'(-2098);
			1671: out = 16'(-1220);
			1672: out = 16'(-9107);
			1673: out = 16'(3388);
			1674: out = 16'(291);
			1675: out = 16'(8106);
			1676: out = 16'(875);
			1677: out = 16'(4358);
			1678: out = 16'(2573);
			1679: out = 16'(-1288);
			1680: out = 16'(2951);
			1681: out = 16'(8376);
			1682: out = 16'(1666);
			1683: out = 16'(5504);
			1684: out = 16'(-3651);
			1685: out = 16'(1434);
			1686: out = 16'(-10966);
			1687: out = 16'(4008);
			1688: out = 16'(-1206);
			1689: out = 16'(6383);
			1690: out = 16'(5445);
			1691: out = 16'(3854);
			1692: out = 16'(591);
			1693: out = 16'(-4253);
			1694: out = 16'(-1291);
			1695: out = 16'(6455);
			1696: out = 16'(-8926);
			1697: out = 16'(-3059);
			1698: out = 16'(-1048);
			1699: out = 16'(2631);
			1700: out = 16'(2701);
			1701: out = 16'(-4120);
			1702: out = 16'(-856);
			1703: out = 16'(2891);
			1704: out = 16'(2992);
			1705: out = 16'(-2373);
			1706: out = 16'(359);
			1707: out = 16'(3877);
			1708: out = 16'(-3842);
			1709: out = 16'(-7916);
			1710: out = 16'(2471);
			1711: out = 16'(8654);
			1712: out = 16'(-2359);
			1713: out = 16'(-3144);
			1714: out = 16'(-9715);
			1715: out = 16'(7676);
			1716: out = 16'(-7770);
			1717: out = 16'(2140);
			1718: out = 16'(1198);
			1719: out = 16'(-2450);
			1720: out = 16'(-1861);
			1721: out = 16'(-8855);
			1722: out = 16'(8436);
			1723: out = 16'(-1785);
			1724: out = 16'(253);
			1725: out = 16'(-2884);
			1726: out = 16'(-659);
			1727: out = 16'(-6465);
			1728: out = 16'(-344);
			1729: out = 16'(-3899);
			1730: out = 16'(4131);
			1731: out = 16'(-974);
			1732: out = 16'(-2097);
			1733: out = 16'(1618);
			1734: out = 16'(3164);
			1735: out = 16'(-462);
			1736: out = 16'(2318);
			1737: out = 16'(-1358);
			1738: out = 16'(1079);
			1739: out = 16'(-1066);
			1740: out = 16'(3188);
			1741: out = 16'(-573);
			1742: out = 16'(-1581);
			1743: out = 16'(4805);
			1744: out = 16'(-4800);
			1745: out = 16'(-6504);
			1746: out = 16'(9968);
			1747: out = 16'(6310);
			1748: out = 16'(-337);
			1749: out = 16'(853);
			1750: out = 16'(-7688);
			1751: out = 16'(2006);
			1752: out = 16'(-472);
			1753: out = 16'(-6182);
			1754: out = 16'(1871);
			1755: out = 16'(4399);
			1756: out = 16'(-1488);
			1757: out = 16'(2848);
			1758: out = 16'(-1985);
			1759: out = 16'(-2201);
			1760: out = 16'(-784);
			1761: out = 16'(-583);
			1762: out = 16'(-4230);
			1763: out = 16'(1031);
			1764: out = 16'(444);
			1765: out = 16'(4106);
			1766: out = 16'(5852);
			1767: out = 16'(863);
			1768: out = 16'(1149);
			1769: out = 16'(1395);
			1770: out = 16'(-1801);
			1771: out = 16'(4241);
			1772: out = 16'(-88);
			1773: out = 16'(2823);
			1774: out = 16'(-1037);
			1775: out = 16'(-1526);
			1776: out = 16'(-2134);
			1777: out = 16'(1379);
			1778: out = 16'(-4034);
			1779: out = 16'(2212);
			1780: out = 16'(-7904);
			1781: out = 16'(765);
			1782: out = 16'(-3482);
			1783: out = 16'(-10114);
			1784: out = 16'(2412);
			1785: out = 16'(7762);
			1786: out = 16'(1680);
			1787: out = 16'(1258);
			1788: out = 16'(-2241);
			1789: out = 16'(414);
			1790: out = 16'(-5557);
			1791: out = 16'(79);
			1792: out = 16'(329);
			1793: out = 16'(-4165);
			1794: out = 16'(1861);
			1795: out = 16'(3504);
			1796: out = 16'(-6513);
			1797: out = 16'(632);
			1798: out = 16'(4831);
			1799: out = 16'(538);
			1800: out = 16'(3357);
			1801: out = 16'(1006);
			1802: out = 16'(1944);
			1803: out = 16'(3377);
			1804: out = 16'(-5732);
			1805: out = 16'(-1472);
			1806: out = 16'(925);
			1807: out = 16'(-2768);
			1808: out = 16'(-575);
			1809: out = 16'(-6971);
			1810: out = 16'(1033);
			1811: out = 16'(-1553);
			1812: out = 16'(-3692);
			1813: out = 16'(3086);
			1814: out = 16'(-561);
			1815: out = 16'(820);
			1816: out = 16'(-1373);
			1817: out = 16'(-5327);
			1818: out = 16'(3962);
			1819: out = 16'(3558);
			1820: out = 16'(-1119);
			1821: out = 16'(-5429);
			1822: out = 16'(-500);
			1823: out = 16'(4956);
			1824: out = 16'(-3564);
			1825: out = 16'(5435);
			1826: out = 16'(-638);
			1827: out = 16'(-192);
			1828: out = 16'(-2618);
			1829: out = 16'(3392);
			1830: out = 16'(482);
			1831: out = 16'(1632);
			1832: out = 16'(3066);
			1833: out = 16'(-3045);
			1834: out = 16'(1023);
			1835: out = 16'(3456);
			1836: out = 16'(1944);
			1837: out = 16'(-2875);
			1838: out = 16'(-3937);
			1839: out = 16'(-3260);
			1840: out = 16'(4431);
			1841: out = 16'(-8108);
			1842: out = 16'(-8715);
			1843: out = 16'(6755);
			1844: out = 16'(-5925);
			1845: out = 16'(4695);
			1846: out = 16'(4577);
			1847: out = 16'(2615);
			1848: out = 16'(-371);
			1849: out = 16'(-1837);
			1850: out = 16'(2743);
			1851: out = 16'(4223);
			1852: out = 16'(40);
			1853: out = 16'(-395);
			1854: out = 16'(2749);
			1855: out = 16'(-2955);
			1856: out = 16'(2939);
			1857: out = 16'(-4101);
			1858: out = 16'(5358);
			1859: out = 16'(-4952);
			1860: out = 16'(-2904);
			1861: out = 16'(6696);
			1862: out = 16'(-4035);
			1863: out = 16'(-934);
			1864: out = 16'(-955);
			1865: out = 16'(4493);
			1866: out = 16'(-3752);
			1867: out = 16'(-742);
			1868: out = 16'(1932);
			1869: out = 16'(-4391);
			1870: out = 16'(-499);
			1871: out = 16'(-7854);
			1872: out = 16'(3499);
			1873: out = 16'(6078);
			1874: out = 16'(-2715);
			1875: out = 16'(-1666);
			1876: out = 16'(-189);
			1877: out = 16'(-257);
			1878: out = 16'(182);
			1879: out = 16'(-1934);
			1880: out = 16'(556);
			1881: out = 16'(1329);
			1882: out = 16'(809);
			1883: out = 16'(-557);
			1884: out = 16'(-1274);
			1885: out = 16'(-3919);
			1886: out = 16'(-981);
			1887: out = 16'(4628);
			1888: out = 16'(5507);
			1889: out = 16'(1612);
			1890: out = 16'(-3313);
			1891: out = 16'(6770);
			1892: out = 16'(2329);
			1893: out = 16'(-3351);
			1894: out = 16'(1969);
			1895: out = 16'(-4170);
			1896: out = 16'(1276);
			1897: out = 16'(-562);
			1898: out = 16'(-3213);
			1899: out = 16'(4204);
			1900: out = 16'(-4756);
			1901: out = 16'(-3777);
			1902: out = 16'(-743);
			1903: out = 16'(781);
			1904: out = 16'(381);
			1905: out = 16'(2991);
			1906: out = 16'(-1033);
			1907: out = 16'(2218);
			1908: out = 16'(377);
			1909: out = 16'(3507);
			1910: out = 16'(-533);
			1911: out = 16'(-2856);
			1912: out = 16'(-2902);
			1913: out = 16'(2167);
			1914: out = 16'(-9783);
			1915: out = 16'(-1447);
			1916: out = 16'(-970);
			1917: out = 16'(4249);
			1918: out = 16'(-7121);
			1919: out = 16'(2781);
			1920: out = 16'(3182);
			1921: out = 16'(-4825);
			1922: out = 16'(4126);
			1923: out = 16'(495);
			1924: out = 16'(4371);
			1925: out = 16'(-4134);
			1926: out = 16'(3488);
			1927: out = 16'(-28);
			1928: out = 16'(-2410);
			1929: out = 16'(1677);
			1930: out = 16'(435);
			1931: out = 16'(-3010);
			1932: out = 16'(599);
			1933: out = 16'(-986);
			1934: out = 16'(2079);
			1935: out = 16'(-1095);
			1936: out = 16'(-2040);
			1937: out = 16'(2938);
			1938: out = 16'(-1358);
			1939: out = 16'(5926);
			1940: out = 16'(-164);
			1941: out = 16'(2344);
			1942: out = 16'(178);
			1943: out = 16'(2211);
			1944: out = 16'(-4436);
			1945: out = 16'(2648);
			1946: out = 16'(931);
			1947: out = 16'(3050);
			1948: out = 16'(1225);
			1949: out = 16'(190);
			1950: out = 16'(-6875);
			1951: out = 16'(1651);
			1952: out = 16'(2284);
			1953: out = 16'(-3366);
			1954: out = 16'(4610);
			1955: out = 16'(-2694);
			1956: out = 16'(-1946);
			1957: out = 16'(-893);
			1958: out = 16'(-1240);
			1959: out = 16'(68);
			1960: out = 16'(-3641);
			1961: out = 16'(-4579);
			1962: out = 16'(-1695);
			1963: out = 16'(2831);
			1964: out = 16'(-9117);
			1965: out = 16'(229);
			1966: out = 16'(4528);
			1967: out = 16'(4597);
			1968: out = 16'(-1743);
			1969: out = 16'(-236);
			1970: out = 16'(-631);
			1971: out = 16'(-142);
			1972: out = 16'(-5752);
			1973: out = 16'(726);
			1974: out = 16'(5770);
			1975: out = 16'(-1523);
			1976: out = 16'(404);
			1977: out = 16'(-1073);
			1978: out = 16'(186);
			1979: out = 16'(442);
			1980: out = 16'(5044);
			1981: out = 16'(210);
			1982: out = 16'(-2589);
			1983: out = 16'(-3367);
			1984: out = 16'(492);
			1985: out = 16'(496);
			1986: out = 16'(1283);
			1987: out = 16'(3077);
			1988: out = 16'(-1116);
			1989: out = 16'(416);
			1990: out = 16'(904);
			1991: out = 16'(414);
			1992: out = 16'(-242);
			1993: out = 16'(-3103);
			1994: out = 16'(4160);
			1995: out = 16'(128);
			1996: out = 16'(-1110);
			1997: out = 16'(-1411);
			1998: out = 16'(2578);
			1999: out = 16'(46);
			2000: out = 16'(1931);
			2001: out = 16'(-6255);
			2002: out = 16'(23);
			2003: out = 16'(901);
			2004: out = 16'(2595);
			2005: out = 16'(-190);
			2006: out = 16'(-5799);
			2007: out = 16'(4181);
			2008: out = 16'(-170);
			2009: out = 16'(-3059);
			2010: out = 16'(215);
			2011: out = 16'(1829);
			2012: out = 16'(-2783);
			2013: out = 16'(7133);
			2014: out = 16'(-284);
			2015: out = 16'(-5983);
			2016: out = 16'(1733);
			2017: out = 16'(-2346);
			2018: out = 16'(1337);
			2019: out = 16'(3215);
			2020: out = 16'(-810);
			2021: out = 16'(1165);
			2022: out = 16'(-3631);
			2023: out = 16'(-2210);
			2024: out = 16'(1321);
			2025: out = 16'(2824);
			2026: out = 16'(2357);
			2027: out = 16'(1898);
			2028: out = 16'(-3602);
			2029: out = 16'(204);
			2030: out = 16'(-2040);
			2031: out = 16'(-553);
			2032: out = 16'(128);
			2033: out = 16'(4583);
			2034: out = 16'(256);
			2035: out = 16'(-1769);
			2036: out = 16'(-4458);
			2037: out = 16'(4598);
			2038: out = 16'(3185);
			2039: out = 16'(-781);
			2040: out = 16'(2227);
			2041: out = 16'(-2291);
			2042: out = 16'(-863);
			2043: out = 16'(-3281);
			2044: out = 16'(722);
			2045: out = 16'(-2125);
			2046: out = 16'(-918);
			2047: out = 16'(2062);
			2048: out = 16'(-3395);
			2049: out = 16'(2490);
			2050: out = 16'(3043);
			2051: out = 16'(1869);
			2052: out = 16'(-5444);
			2053: out = 16'(-1072);
			2054: out = 16'(1513);
			2055: out = 16'(-3500);
			2056: out = 16'(-80);
			2057: out = 16'(3220);
			2058: out = 16'(2803);
			2059: out = 16'(1055);
			2060: out = 16'(3147);
			2061: out = 16'(-3156);
			2062: out = 16'(-3323);
			2063: out = 16'(4566);
			2064: out = 16'(-448);
			2065: out = 16'(2824);
			2066: out = 16'(-4528);
			2067: out = 16'(3701);
			2068: out = 16'(1102);
			2069: out = 16'(-6100);
			2070: out = 16'(-1034);
			2071: out = 16'(133);
			2072: out = 16'(-309);
			2073: out = 16'(-2048);
			2074: out = 16'(1406);
			2075: out = 16'(-3081);
			2076: out = 16'(-622);
			2077: out = 16'(5612);
			2078: out = 16'(-188);
			2079: out = 16'(-460);
			2080: out = 16'(-2153);
			2081: out = 16'(-2891);
			2082: out = 16'(2905);
			2083: out = 16'(-3526);
			2084: out = 16'(2885);
			2085: out = 16'(-1221);
			2086: out = 16'(2498);
			2087: out = 16'(-1990);
			2088: out = 16'(-2588);
			2089: out = 16'(1399);
			2090: out = 16'(319);
			2091: out = 16'(344);
			2092: out = 16'(-1541);
			2093: out = 16'(361);
			2094: out = 16'(1508);
			2095: out = 16'(1786);
			2096: out = 16'(-2487);
			2097: out = 16'(820);
			2098: out = 16'(-3110);
			2099: out = 16'(653);
			2100: out = 16'(-4645);
			2101: out = 16'(181);
			2102: out = 16'(205);
			2103: out = 16'(-1043);
			2104: out = 16'(2543);
			2105: out = 16'(1573);
			2106: out = 16'(-67);
			2107: out = 16'(-127);
			2108: out = 16'(2219);
			2109: out = 16'(-607);
			2110: out = 16'(-1849);
			2111: out = 16'(-857);
			2112: out = 16'(3260);
			2113: out = 16'(-1186);
			2114: out = 16'(127);
			2115: out = 16'(-220);
			2116: out = 16'(2213);
			2117: out = 16'(-1457);
			2118: out = 16'(2384);
			2119: out = 16'(-4853);
			2120: out = 16'(-2585);
			2121: out = 16'(1897);
			2122: out = 16'(-1282);
			2123: out = 16'(807);
			2124: out = 16'(-2226);
			2125: out = 16'(231);
			2126: out = 16'(680);
			2127: out = 16'(272);
			2128: out = 16'(-2963);
			2129: out = 16'(-2029);
			2130: out = 16'(1);
			2131: out = 16'(334);
			2132: out = 16'(-2801);
			2133: out = 16'(-226);
			2134: out = 16'(378);
			2135: out = 16'(-4834);
			2136: out = 16'(2248);
			2137: out = 16'(2255);
			2138: out = 16'(3694);
			2139: out = 16'(-1768);
			2140: out = 16'(-3069);
			2141: out = 16'(610);
			2142: out = 16'(608);
			2143: out = 16'(2370);
			2144: out = 16'(4602);
			2145: out = 16'(-2348);
			2146: out = 16'(908);
			2147: out = 16'(-7114);
			2148: out = 16'(2909);
			2149: out = 16'(-2028);
			2150: out = 16'(3941);
			2151: out = 16'(2069);
			2152: out = 16'(-146);
			2153: out = 16'(-2574);
			2154: out = 16'(479);
			2155: out = 16'(-707);
			2156: out = 16'(285);
			2157: out = 16'(1498);
			2158: out = 16'(-4253);
			2159: out = 16'(-6268);
			2160: out = 16'(2287);
			2161: out = 16'(415);
			2162: out = 16'(-448);
			2163: out = 16'(-1148);
			2164: out = 16'(-2141);
			2165: out = 16'(2323);
			2166: out = 16'(-3316);
			2167: out = 16'(-403);
			2168: out = 16'(-2778);
			2169: out = 16'(4349);
			2170: out = 16'(936);
			2171: out = 16'(971);
			2172: out = 16'(-1926);
			2173: out = 16'(1446);
			2174: out = 16'(-3258);
			2175: out = 16'(2821);
			2176: out = 16'(-3519);
			2177: out = 16'(2602);
			2178: out = 16'(1638);
			2179: out = 16'(-608);
			2180: out = 16'(-4816);
			2181: out = 16'(4151);
			2182: out = 16'(2425);
			2183: out = 16'(-1516);
			2184: out = 16'(1860);
			2185: out = 16'(145);
			2186: out = 16'(1872);
			2187: out = 16'(-2012);
			2188: out = 16'(3844);
			2189: out = 16'(1251);
			2190: out = 16'(-3443);
			2191: out = 16'(1225);
			2192: out = 16'(1365);
			2193: out = 16'(2304);
			2194: out = 16'(-469);
			2195: out = 16'(-432);
			2196: out = 16'(-2553);
			2197: out = 16'(1434);
			2198: out = 16'(1569);
			2199: out = 16'(2314);
			2200: out = 16'(-1259);
			2201: out = 16'(-168);
			2202: out = 16'(-2646);
			2203: out = 16'(3389);
			2204: out = 16'(-2110);
			2205: out = 16'(1125);
			2206: out = 16'(958);
			2207: out = 16'(-2297);
			2208: out = 16'(-3511);
			2209: out = 16'(256);
			2210: out = 16'(1913);
			2211: out = 16'(-797);
			2212: out = 16'(-2230);
			2213: out = 16'(-1171);
			2214: out = 16'(2144);
			2215: out = 16'(-597);
			2216: out = 16'(2122);
			2217: out = 16'(-824);
			2218: out = 16'(2549);
			2219: out = 16'(-459);
			2220: out = 16'(-6055);
			2221: out = 16'(4067);
			2222: out = 16'(-2471);
			2223: out = 16'(-1131);
			2224: out = 16'(3618);
			2225: out = 16'(-944);
			2226: out = 16'(529);
			2227: out = 16'(-3856);
			2228: out = 16'(-1120);
			2229: out = 16'(869);
			2230: out = 16'(396);
			2231: out = 16'(243);
			2232: out = 16'(1445);
			2233: out = 16'(-1667);
			2234: out = 16'(1943);
			2235: out = 16'(-1106);
			2236: out = 16'(569);
			2237: out = 16'(-594);
			2238: out = 16'(2551);
			2239: out = 16'(796);
			2240: out = 16'(-2725);
			2241: out = 16'(-1909);
			2242: out = 16'(2991);
			2243: out = 16'(-418);
			2244: out = 16'(2899);
			2245: out = 16'(-905);
			2246: out = 16'(-748);
			2247: out = 16'(1651);
			2248: out = 16'(-2102);
			2249: out = 16'(2684);
			2250: out = 16'(265);
			2251: out = 16'(2190);
			2252: out = 16'(1882);
			2253: out = 16'(-2789);
			2254: out = 16'(-46);
			2255: out = 16'(1417);
			2256: out = 16'(904);
			2257: out = 16'(1311);
			2258: out = 16'(607);
			2259: out = 16'(-574);
			2260: out = 16'(-4645);
			2261: out = 16'(3519);
			2262: out = 16'(3312);
			2263: out = 16'(1082);
			2264: out = 16'(597);
			2265: out = 16'(-960);
			2266: out = 16'(-767);
			2267: out = 16'(675);
			2268: out = 16'(-2036);
			2269: out = 16'(-792);
			2270: out = 16'(3448);
			2271: out = 16'(2357);
			2272: out = 16'(-266);
			2273: out = 16'(-1929);
			2274: out = 16'(862);
			2275: out = 16'(-1347);
			2276: out = 16'(79);
			2277: out = 16'(-4597);
			2278: out = 16'(-70);
			2279: out = 16'(597);
			2280: out = 16'(-2237);
			2281: out = 16'(4557);
			2282: out = 16'(-675);
			2283: out = 16'(2322);
			2284: out = 16'(1658);
			2285: out = 16'(-971);
			2286: out = 16'(897);
			2287: out = 16'(-2710);
			2288: out = 16'(-251);
			2289: out = 16'(-493);
			2290: out = 16'(1171);
			2291: out = 16'(508);
			2292: out = 16'(-231);
			2293: out = 16'(-393);
			2294: out = 16'(-1459);
			2295: out = 16'(76);
			2296: out = 16'(3782);
			2297: out = 16'(1526);
			2298: out = 16'(-684);
			2299: out = 16'(-1837);
			2300: out = 16'(936);
			2301: out = 16'(-616);
			2302: out = 16'(473);
			2303: out = 16'(2234);
			2304: out = 16'(-1388);
			2305: out = 16'(-830);
			2306: out = 16'(2222);
			2307: out = 16'(844);
			2308: out = 16'(-2075);
			2309: out = 16'(-3696);
			2310: out = 16'(4944);
			2311: out = 16'(-1478);
			2312: out = 16'(1318);
			2313: out = 16'(875);
			2314: out = 16'(-2598);
			2315: out = 16'(4229);
			2316: out = 16'(-1368);
			2317: out = 16'(663);
			2318: out = 16'(1117);
			2319: out = 16'(-1309);
			2320: out = 16'(668);
			2321: out = 16'(-1296);
			2322: out = 16'(-538);
			2323: out = 16'(-332);
			2324: out = 16'(2479);
			2325: out = 16'(-3111);
			2326: out = 16'(-757);
			2327: out = 16'(2427);
			2328: out = 16'(-1598);
			2329: out = 16'(1798);
			2330: out = 16'(914);
			2331: out = 16'(2288);
			2332: out = 16'(-970);
			2333: out = 16'(-1090);
			2334: out = 16'(-2541);
			2335: out = 16'(1289);
			2336: out = 16'(571);
			2337: out = 16'(533);
			2338: out = 16'(438);
			2339: out = 16'(904);
			2340: out = 16'(1287);
			2341: out = 16'(-1688);
			2342: out = 16'(22);
			2343: out = 16'(-678);
			2344: out = 16'(263);
			2345: out = 16'(-3420);
			2346: out = 16'(-778);
			2347: out = 16'(2613);
			2348: out = 16'(-1915);
			2349: out = 16'(-633);
			2350: out = 16'(833);
			2351: out = 16'(1266);
			2352: out = 16'(-3038);
			2353: out = 16'(-7);
			2354: out = 16'(2274);
			2355: out = 16'(-595);
			2356: out = 16'(713);
			2357: out = 16'(-503);
			2358: out = 16'(223);
			2359: out = 16'(-990);
			2360: out = 16'(-1219);
			2361: out = 16'(704);
			2362: out = 16'(-361);
			2363: out = 16'(-118);
			2364: out = 16'(-3197);
			2365: out = 16'(2399);
			2366: out = 16'(233);
			2367: out = 16'(1260);
			2368: out = 16'(-949);
			2369: out = 16'(-1987);
			2370: out = 16'(-146);
			2371: out = 16'(-2348);
			2372: out = 16'(234);
			2373: out = 16'(-798);
			2374: out = 16'(665);
			2375: out = 16'(-1727);
			2376: out = 16'(-3560);
			2377: out = 16'(2770);
			2378: out = 16'(757);
			2379: out = 16'(973);
			2380: out = 16'(-1732);
			2381: out = 16'(1082);
			2382: out = 16'(772);
			2383: out = 16'(589);
			2384: out = 16'(-683);
			2385: out = 16'(-614);
			2386: out = 16'(-76);
			2387: out = 16'(1844);
			2388: out = 16'(-419);
			2389: out = 16'(243);
			2390: out = 16'(-4558);
			2391: out = 16'(1387);
			2392: out = 16'(-4732);
			2393: out = 16'(2441);
			2394: out = 16'(240);
			2395: out = 16'(-2473);
			2396: out = 16'(-876);
			2397: out = 16'(1632);
			2398: out = 16'(-2704);
			2399: out = 16'(-397);
			2400: out = 16'(498);
			2401: out = 16'(-1349);
			2402: out = 16'(-572);
			2403: out = 16'(1782);
			2404: out = 16'(729);
			2405: out = 16'(561);
			2406: out = 16'(-2417);
			2407: out = 16'(-7);
			2408: out = 16'(2814);
			2409: out = 16'(166);
			2410: out = 16'(-539);
			2411: out = 16'(-2014);
			2412: out = 16'(884);
			2413: out = 16'(-1014);
			2414: out = 16'(-763);
			2415: out = 16'(-216);
			2416: out = 16'(4232);
			2417: out = 16'(650);
			2418: out = 16'(1035);
			2419: out = 16'(-2252);
			2420: out = 16'(-159);
			2421: out = 16'(1023);
			2422: out = 16'(1067);
			2423: out = 16'(341);
			2424: out = 16'(-796);
			2425: out = 16'(-2143);
			2426: out = 16'(193);
			2427: out = 16'(288);
			2428: out = 16'(-1466);
			2429: out = 16'(-1652);
			2430: out = 16'(402);
			2431: out = 16'(-47);
			2432: out = 16'(-1617);
			2433: out = 16'(395);
			2434: out = 16'(-2049);
			2435: out = 16'(2403);
			2436: out = 16'(-4598);
			2437: out = 16'(-255);
			2438: out = 16'(365);
			2439: out = 16'(-2009);
			2440: out = 16'(-3631);
			2441: out = 16'(1600);
			2442: out = 16'(-5161);
			2443: out = 16'(803);
			2444: out = 16'(2009);
			2445: out = 16'(-2498);
			2446: out = 16'(2673);
			2447: out = 16'(-1193);
			2448: out = 16'(-1865);
			2449: out = 16'(-688);
			2450: out = 16'(645);
			2451: out = 16'(-375);
			2452: out = 16'(1146);
			2453: out = 16'(1361);
			2454: out = 16'(-887);
			2455: out = 16'(1608);
			2456: out = 16'(-1348);
			2457: out = 16'(-2121);
			2458: out = 16'(1372);
			2459: out = 16'(-2182);
			2460: out = 16'(-1310);
			2461: out = 16'(-213);
			2462: out = 16'(-122);
			2463: out = 16'(518);
			2464: out = 16'(1591);
			2465: out = 16'(1631);
			2466: out = 16'(-1734);
			2467: out = 16'(1049);
			2468: out = 16'(-82);
			2469: out = 16'(298);
			2470: out = 16'(114);
			2471: out = 16'(-205);
			2472: out = 16'(-1318);
			2473: out = 16'(-1758);
			2474: out = 16'(1307);
			2475: out = 16'(3030);
			2476: out = 16'(1080);
			2477: out = 16'(-251);
			2478: out = 16'(-1367);
			2479: out = 16'(-755);
			2480: out = 16'(-715);
			2481: out = 16'(2551);
			2482: out = 16'(1297);
			2483: out = 16'(-1525);
			2484: out = 16'(-1466);
			2485: out = 16'(2259);
			2486: out = 16'(-1136);
			2487: out = 16'(455);
			2488: out = 16'(-428);
			2489: out = 16'(709);
			2490: out = 16'(-414);
			2491: out = 16'(-174);
			2492: out = 16'(-2200);
			2493: out = 16'(1267);
			2494: out = 16'(27);
			2495: out = 16'(1067);
			2496: out = 16'(1714);
			2497: out = 16'(-1018);
			2498: out = 16'(21);
			2499: out = 16'(-1809);
			2500: out = 16'(1015);
			2501: out = 16'(-1828);
			2502: out = 16'(1409);
			2503: out = 16'(356);
			2504: out = 16'(-2268);
			2505: out = 16'(-1820);
			2506: out = 16'(302);
			2507: out = 16'(1642);
			2508: out = 16'(-3);
			2509: out = 16'(704);
			2510: out = 16'(367);
			2511: out = 16'(570);
			2512: out = 16'(511);
			2513: out = 16'(-95);
			2514: out = 16'(-1688);
			2515: out = 16'(2207);
			2516: out = 16'(-2101);
			2517: out = 16'(449);
			2518: out = 16'(1069);
			2519: out = 16'(-2526);
			2520: out = 16'(-1961);
			2521: out = 16'(897);
			2522: out = 16'(371);
			2523: out = 16'(699);
			2524: out = 16'(1534);
			2525: out = 16'(-21);
			2526: out = 16'(-1441);
			2527: out = 16'(-1481);
			2528: out = 16'(1624);
			2529: out = 16'(59);
			2530: out = 16'(-569);
			2531: out = 16'(468);
			2532: out = 16'(359);
			2533: out = 16'(704);
			2534: out = 16'(904);
			2535: out = 16'(-795);
			2536: out = 16'(1502);
			2537: out = 16'(88);
			2538: out = 16'(872);
			2539: out = 16'(831);
			2540: out = 16'(-113);
			2541: out = 16'(-1333);
			2542: out = 16'(3661);
			2543: out = 16'(-887);
			2544: out = 16'(1467);
			2545: out = 16'(-1300);
			2546: out = 16'(-38);
			2547: out = 16'(-1835);
			2548: out = 16'(610);
			2549: out = 16'(120);
			2550: out = 16'(-310);
			2551: out = 16'(-1982);
			2552: out = 16'(1616);
			2553: out = 16'(-60);
			2554: out = 16'(-810);
			2555: out = 16'(2287);
			2556: out = 16'(-770);
			2557: out = 16'(-1154);
			2558: out = 16'(641);
			2559: out = 16'(27);
			2560: out = 16'(1115);
			2561: out = 16'(1618);
			2562: out = 16'(-1808);
			2563: out = 16'(-765);
			2564: out = 16'(2205);
			2565: out = 16'(-885);
			2566: out = 16'(-1252);
			2567: out = 16'(2147);
			2568: out = 16'(-2009);
			2569: out = 16'(-1168);
			2570: out = 16'(1658);
			2571: out = 16'(-1422);
			2572: out = 16'(2067);
			2573: out = 16'(568);
			2574: out = 16'(-1082);
			2575: out = 16'(-1218);
			2576: out = 16'(73);
			2577: out = 16'(758);
			2578: out = 16'(1491);
			2579: out = 16'(-996);
			2580: out = 16'(-2133);
			2581: out = 16'(-1686);
			2582: out = 16'(-1);
			2583: out = 16'(-224);
			2584: out = 16'(-120);
			2585: out = 16'(143);
			2586: out = 16'(131);
			2587: out = 16'(-635);
			2588: out = 16'(-1045);
			2589: out = 16'(-1140);
			2590: out = 16'(609);
			2591: out = 16'(246);
			2592: out = 16'(-1349);
			2593: out = 16'(-47);
			2594: out = 16'(544);
			2595: out = 16'(-970);
			2596: out = 16'(-234);
			2597: out = 16'(-2518);
			2598: out = 16'(1617);
			2599: out = 16'(945);
			2600: out = 16'(-1546);
			2601: out = 16'(1);
			2602: out = 16'(-1026);
			2603: out = 16'(-391);
			2604: out = 16'(-293);
			2605: out = 16'(-1280);
			2606: out = 16'(-764);
			2607: out = 16'(951);
			2608: out = 16'(-1092);
			2609: out = 16'(1298);
			2610: out = 16'(1405);
			2611: out = 16'(778);
			2612: out = 16'(20);
			2613: out = 16'(475);
			2614: out = 16'(-269);
			2615: out = 16'(631);
			2616: out = 16'(1160);
			2617: out = 16'(-118);
			2618: out = 16'(-1476);
			2619: out = 16'(530);
			2620: out = 16'(-272);
			2621: out = 16'(-380);
			2622: out = 16'(404);
			2623: out = 16'(-82);
			2624: out = 16'(542);
			2625: out = 16'(361);
			2626: out = 16'(489);
			2627: out = 16'(-619);
			2628: out = 16'(649);
			2629: out = 16'(-14);
			2630: out = 16'(738);
			2631: out = 16'(299);
			2632: out = 16'(-234);
			2633: out = 16'(770);
			2634: out = 16'(495);
			2635: out = 16'(-2068);
			2636: out = 16'(-139);
			2637: out = 16'(173);
			2638: out = 16'(-127);
			2639: out = 16'(-1561);
			2640: out = 16'(-421);
			2641: out = 16'(968);
			2642: out = 16'(294);
			2643: out = 16'(735);
			2644: out = 16'(-1130);
			2645: out = 16'(-609);
			2646: out = 16'(365);
			2647: out = 16'(-1676);
			2648: out = 16'(-787);
			2649: out = 16'(-556);
			2650: out = 16'(562);
			2651: out = 16'(-152);
			2652: out = 16'(493);
			2653: out = 16'(582);
			2654: out = 16'(74);
			2655: out = 16'(909);
			2656: out = 16'(-1134);
			2657: out = 16'(-547);
			2658: out = 16'(-1907);
			2659: out = 16'(2062);
			2660: out = 16'(1920);
			2661: out = 16'(669);
			2662: out = 16'(-544);
			2663: out = 16'(793);
			2664: out = 16'(-1233);
			2665: out = 16'(666);
			2666: out = 16'(295);
			2667: out = 16'(328);
			2668: out = 16'(784);
			2669: out = 16'(-549);
			2670: out = 16'(-443);
			2671: out = 16'(-297);
			2672: out = 16'(761);
			2673: out = 16'(806);
			2674: out = 16'(-301);
			2675: out = 16'(-289);
			2676: out = 16'(-112);
			2677: out = 16'(-42);
			2678: out = 16'(-454);
			2679: out = 16'(870);
			2680: out = 16'(-1013);
			2681: out = 16'(-444);
			2682: out = 16'(1363);
			2683: out = 16'(1095);
			2684: out = 16'(-112);
			2685: out = 16'(1307);
			2686: out = 16'(-1503);
			2687: out = 16'(-1531);
			2688: out = 16'(1469);
			2689: out = 16'(-119);
			2690: out = 16'(956);
			2691: out = 16'(-1109);
			2692: out = 16'(-666);
			2693: out = 16'(-663);
			2694: out = 16'(1060);
			2695: out = 16'(-385);
			2696: out = 16'(111);
			2697: out = 16'(-316);
			2698: out = 16'(-1084);
			2699: out = 16'(789);
			2700: out = 16'(-722);
			2701: out = 16'(104);
			2702: out = 16'(1398);
			2703: out = 16'(-1858);
			2704: out = 16'(666);
			2705: out = 16'(2);
			2706: out = 16'(1161);
			2707: out = 16'(1174);
			2708: out = 16'(267);
			2709: out = 16'(-272);
			2710: out = 16'(-228);
			2711: out = 16'(-298);
			2712: out = 16'(1326);
			2713: out = 16'(-270);
			2714: out = 16'(-616);
			2715: out = 16'(455);
			2716: out = 16'(-1355);
			2717: out = 16'(-205);
			2718: out = 16'(353);
			2719: out = 16'(523);
			2720: out = 16'(-817);
			2721: out = 16'(215);
			2722: out = 16'(-479);
			2723: out = 16'(-74);
			2724: out = 16'(-792);
			2725: out = 16'(-796);
			2726: out = 16'(428);
			2727: out = 16'(-712);
			2728: out = 16'(-966);
			2729: out = 16'(-1258);
			2730: out = 16'(654);
			2731: out = 16'(-1017);
			2732: out = 16'(-289);
			2733: out = 16'(-2437);
			2734: out = 16'(1389);
			2735: out = 16'(-418);
			2736: out = 16'(-1523);
			2737: out = 16'(85);
			2738: out = 16'(-301);
			2739: out = 16'(320);
			2740: out = 16'(-262);
			2741: out = 16'(133);
			2742: out = 16'(742);
			2743: out = 16'(420);
			2744: out = 16'(-469);
			2745: out = 16'(-631);
			2746: out = 16'(1025);
			2747: out = 16'(-189);
			2748: out = 16'(-62);
			2749: out = 16'(41);
			2750: out = 16'(-907);
			2751: out = 16'(816);
			2752: out = 16'(191);
			2753: out = 16'(-711);
			2754: out = 16'(-1583);
			2755: out = 16'(-706);
			2756: out = 16'(658);
			2757: out = 16'(800);
			2758: out = 16'(-342);
			2759: out = 16'(455);
			2760: out = 16'(481);
			2761: out = 16'(-276);
			2762: out = 16'(-7);
			2763: out = 16'(-213);
			2764: out = 16'(-786);
			2765: out = 16'(497);
			2766: out = 16'(-935);
			2767: out = 16'(-733);
			2768: out = 16'(567);
			2769: out = 16'(532);
			2770: out = 16'(486);
			2771: out = 16'(-912);
			2772: out = 16'(-1537);
			2773: out = 16'(2022);
			2774: out = 16'(500);
			2775: out = 16'(737);
			2776: out = 16'(-1348);
			2777: out = 16'(823);
			2778: out = 16'(38);
			2779: out = 16'(167);
			2780: out = 16'(-825);
			2781: out = 16'(730);
			2782: out = 16'(-1841);
			2783: out = 16'(-711);
			2784: out = 16'(1084);
			2785: out = 16'(-1510);
			2786: out = 16'(-387);
			2787: out = 16'(545);
			2788: out = 16'(144);
			2789: out = 16'(782);
			2790: out = 16'(-506);
			2791: out = 16'(108);
			2792: out = 16'(630);
			2793: out = 16'(-1857);
			2794: out = 16'(374);
			2795: out = 16'(147);
			2796: out = 16'(-467);
			2797: out = 16'(-691);
			2798: out = 16'(472);
			2799: out = 16'(-115);
			2800: out = 16'(-923);
			2801: out = 16'(-1493);
			2802: out = 16'(640);
			2803: out = 16'(-483);
			2804: out = 16'(-48);
			2805: out = 16'(749);
			2806: out = 16'(-73);
			2807: out = 16'(-101);
			2808: out = 16'(570);
			2809: out = 16'(-112);
			2810: out = 16'(-267);
			2811: out = 16'(-1331);
			2812: out = 16'(1118);
			2813: out = 16'(-1065);
			2814: out = 16'(257);
			2815: out = 16'(1317);
			2816: out = 16'(-77);
			2817: out = 16'(-509);
			2818: out = 16'(255);
			2819: out = 16'(44);
			2820: out = 16'(-385);
			2821: out = 16'(-59);
			2822: out = 16'(202);
			2823: out = 16'(220);
			2824: out = 16'(-686);
			2825: out = 16'(379);
			2826: out = 16'(-230);
			2827: out = 16'(224);
			2828: out = 16'(542);
			2829: out = 16'(-215);
			2830: out = 16'(414);
			2831: out = 16'(-667);
			2832: out = 16'(-972);
			2833: out = 16'(1427);
			2834: out = 16'(-613);
			2835: out = 16'(61);
			2836: out = 16'(-127);
			2837: out = 16'(246);
			2838: out = 16'(258);
			2839: out = 16'(-243);
			2840: out = 16'(-518);
			2841: out = 16'(218);
			2842: out = 16'(-18);
			2843: out = 16'(917);
			2844: out = 16'(398);
			2845: out = 16'(384);
			2846: out = 16'(-179);
			2847: out = 16'(312);
			2848: out = 16'(-273);
			2849: out = 16'(-31);
			2850: out = 16'(542);
			2851: out = 16'(-666);
			2852: out = 16'(163);
			2853: out = 16'(-128);
			2854: out = 16'(69);
			2855: out = 16'(789);
			2856: out = 16'(-54);
			2857: out = 16'(93);
			2858: out = 16'(-496);
			2859: out = 16'(456);
			2860: out = 16'(-58);
			2861: out = 16'(264);
			2862: out = 16'(278);
			2863: out = 16'(-54);
			2864: out = 16'(-798);
			2865: out = 16'(-690);
			2866: out = 16'(850);
			2867: out = 16'(-1300);
			2868: out = 16'(-53);
			2869: out = 16'(-354);
			2870: out = 16'(778);
			2871: out = 16'(467);
			2872: out = 16'(-336);
			2873: out = 16'(-360);
			2874: out = 16'(-251);
			2875: out = 16'(362);
			2876: out = 16'(-753);
			2877: out = 16'(-781);
			2878: out = 16'(731);
			2879: out = 16'(-642);
			2880: out = 16'(-246);
			2881: out = 16'(-210);
			2882: out = 16'(-247);
			2883: out = 16'(422);
			2884: out = 16'(412);
			2885: out = 16'(-836);
			2886: out = 16'(269);
			2887: out = 16'(-607);
			2888: out = 16'(337);
			2889: out = 16'(-367);
			2890: out = 16'(293);
			2891: out = 16'(374);
			2892: out = 16'(-655);
			2893: out = 16'(-493);
			2894: out = 16'(-240);
			2895: out = 16'(331);
			2896: out = 16'(-382);
			2897: out = 16'(523);
			2898: out = 16'(266);
			2899: out = 16'(259);
			2900: out = 16'(-382);
			2901: out = 16'(445);
			2902: out = 16'(-97);
			2903: out = 16'(-236);
			2904: out = 16'(113);
			2905: out = 16'(-299);
			2906: out = 16'(-30);
			2907: out = 16'(-293);
			2908: out = 16'(394);
			2909: out = 16'(-564);
			2910: out = 16'(40);
			2911: out = 16'(402);
			2912: out = 16'(180);
			2913: out = 16'(-439);
			2914: out = 16'(-47);
			2915: out = 16'(-709);
			2916: out = 16'(510);
			2917: out = 16'(-187);
			2918: out = 16'(-10);
			2919: out = 16'(-12);
			2920: out = 16'(-211);
			2921: out = 16'(-228);
			2922: out = 16'(-231);
			2923: out = 16'(469);
			2924: out = 16'(-562);
			2925: out = 16'(48);
			2926: out = 16'(-211);
			2927: out = 16'(-101);
			2928: out = 16'(294);
			2929: out = 16'(-140);
			2930: out = 16'(66);
			2931: out = 16'(553);
			2932: out = 16'(-24);
			2933: out = 16'(665);
			2934: out = 16'(-66);
			2935: out = 16'(-203);
			2936: out = 16'(-299);
			default: out = 0;
		endcase
	end
endmodule
