module kick_lookup(index, out);
	input logic unsigned [10:0] index;
	output logic signed [15:0] out;
	always_comb begin
		case(index)
			0: out = 16'(0);
			1: out = 16'(3069);
			2: out = 16'(6789);
			3: out = 16'(9756);
			4: out = 16'(32112);
			5: out = 16'(31670);
			6: out = 16'(22038);
			7: out = 16'(-6732);
			8: out = 16'(-28912);
			9: out = 16'(-32262);
			10: out = 16'(-31750);
			11: out = 16'(-25403);
			12: out = 16'(-3197);
			13: out = 16'(20281);
			14: out = 16'(32481);
			15: out = 16'(31999);
			16: out = 16'(22692);
			17: out = 16'(8592);
			18: out = 16'(-14380);
			19: out = 16'(-29308);
			20: out = 16'(-31885);
			21: out = 16'(-31144);
			22: out = 16'(-23476);
			23: out = 16'(-11318);
			24: out = 16'(5527);
			25: out = 16'(20041);
			26: out = 16'(32429);
			27: out = 16'(32289);
			28: out = 16'(26841);
			29: out = 16'(18304);
			30: out = 16'(6280);
			31: out = 16'(-8205);
			32: out = 16'(-22653);
			33: out = 16'(-30874);
			34: out = 16'(-31388);
			35: out = 16'(-26401);
			36: out = 16'(-21378);
			37: out = 16'(-12879);
			38: out = 16'(-4659);
			39: out = 16'(7214);
			40: out = 16'(15761);
			41: out = 16'(25025);
			42: out = 16'(31368);
			43: out = 16'(29331);
			44: out = 16'(23742);
			45: out = 16'(15591);
			46: out = 16'(9865);
			47: out = 16'(2968);
			48: out = 16'(-8893);
			49: out = 16'(-19162);
			50: out = 16'(-24208);
			51: out = 16'(-28007);
			52: out = 16'(-28503);
			53: out = 16'(-24537);
			54: out = 16'(-18451);
			55: out = 16'(-14245);
			56: out = 16'(-7969);
			57: out = 16'(-3386);
			58: out = 16'(3190);
			59: out = 16'(11344);
			60: out = 16'(17468);
			61: out = 16'(22175);
			62: out = 16'(26295);
			63: out = 16'(27597);
			64: out = 16'(24352);
			65: out = 16'(19807);
			66: out = 16'(15304);
			67: out = 16'(10087);
			68: out = 16'(5519);
			69: out = 16'(990);
			70: out = 16'(-4602);
			71: out = 16'(-12017);
			72: out = 16'(-17874);
			73: out = 16'(-21737);
			74: out = 16'(-23589);
			75: out = 16'(-24291);
			76: out = 16'(-24087);
			77: out = 16'(-21100);
			78: out = 16'(-16648);
			79: out = 16'(-12911);
			80: out = 16'(-9520);
			81: out = 16'(-5521);
			82: out = 16'(-2043);
			83: out = 16'(1268);
			84: out = 16'(5665);
			85: out = 16'(10601);
			86: out = 16'(14695);
			87: out = 16'(17852);
			88: out = 16'(20370);
			89: out = 16'(22242);
			90: out = 16'(23334);
			91: out = 16'(21656);
			92: out = 16'(18323);
			93: out = 16'(14779);
			94: out = 16'(11575);
			95: out = 16'(9014);
			96: out = 16'(6198);
			97: out = 16'(2711);
			98: out = 16'(-176);
			99: out = 16'(-2950);
			100: out = 16'(-6363);
			101: out = 16'(-10989);
			102: out = 16'(-15320);
			103: out = 16'(-18278);
			104: out = 16'(-19959);
			105: out = 16'(-20712);
			106: out = 16'(-20830);
			107: out = 16'(-20376);
			108: out = 16'(-19056);
			109: out = 16'(-16254);
			110: out = 16'(-12921);
			111: out = 16'(-9971);
			112: out = 16'(-7504);
			113: out = 16'(-4873);
			114: out = 16'(-2301);
			115: out = 16'(-138);
			116: out = 16'(1957);
			117: out = 16'(4705);
			118: out = 16'(8220);
			119: out = 16'(11473);
			120: out = 16'(14067);
			121: out = 16'(16101);
			122: out = 16'(17700);
			123: out = 16'(19012);
			124: out = 16'(19194);
			125: out = 16'(18788);
			126: out = 16'(17613);
			127: out = 16'(15428);
			128: out = 16'(12829);
			129: out = 16'(10281);
			130: out = 16'(8107);
			131: out = 16'(6314);
			132: out = 16'(4807);
			133: out = 16'(2192);
			134: out = 16'(-83);
			135: out = 16'(-2060);
			136: out = 16'(-4083);
			137: out = 16'(-6529);
			138: out = 16'(-9830);
			139: out = 16'(-13321);
			140: out = 16'(-15863);
			141: out = 16'(-17403);
			142: out = 16'(-18170);
			143: out = 16'(-18320);
			144: out = 16'(-18129);
			145: out = 16'(-17531);
			146: out = 16'(-16523);
			147: out = 16'(-14576);
			148: out = 16'(-11887);
			149: out = 16'(-9260);
			150: out = 16'(-6974);
			151: out = 16'(-5153);
			152: out = 16'(-3133);
			153: out = 16'(-1169);
			154: out = 16'(463);
			155: out = 16'(1861);
			156: out = 16'(3575);
			157: out = 16'(5830);
			158: out = 16'(8421);
			159: out = 16'(10652);
			160: out = 16'(12383);
			161: out = 16'(13746);
			162: out = 16'(14772);
			163: out = 16'(15484);
			164: out = 16'(15240);
			165: out = 16'(14895);
			166: out = 16'(14477);
			167: out = 16'(13333);
			168: out = 16'(11476);
			169: out = 16'(9437);
			170: out = 16'(7538);
			171: out = 16'(5866);
			172: out = 16'(4529);
			173: out = 16'(3386);
			174: out = 16'(1963);
			175: out = 16'(67);
			176: out = 16'(-1450);
			177: out = 16'(-2819);
			178: out = 16'(-4250);
			179: out = 16'(-6132);
			180: out = 16'(-8654);
			181: out = 16'(-11197);
			182: out = 16'(-13045);
			183: out = 16'(-14109);
			184: out = 16'(-14633);
			185: out = 16'(-14705);
			186: out = 16'(-14502);
			187: out = 16'(-14035);
			188: out = 16'(-13332);
			189: out = 16'(-12132);
			190: out = 16'(-10251);
			191: out = 16'(-8120);
			192: out = 16'(-6220);
			193: out = 16'(-4616);
			194: out = 16'(-3323);
			195: out = 16'(-1756);
			196: out = 16'(-330);
			197: out = 16'(820);
			198: out = 16'(1888);
			199: out = 16'(3117);
			200: out = 16'(4855);
			201: out = 16'(6826);
			202: out = 16'(8561);
			203: out = 16'(9937);
			204: out = 16'(11019);
			205: out = 16'(11856);
			206: out = 16'(12489);
			207: out = 16'(12246);
			208: out = 16'(12012);
			209: out = 16'(11835);
			210: out = 16'(11213);
			211: out = 16'(10108);
			212: out = 16'(8547);
			213: out = 16'(6974);
			214: out = 16'(5528);
			215: out = 16'(4280);
			216: out = 16'(3286);
			217: out = 16'(2446);
			218: out = 16'(1058);
			219: out = 16'(-358);
			220: out = 16'(-1546);
			221: out = 16'(-2607);
			222: out = 16'(-3787);
			223: out = 16'(-5346);
			224: out = 16'(-7381);
			225: out = 16'(-9402);
			226: out = 16'(-10818);
			227: out = 16'(-11649);
			228: out = 16'(-12014);
			229: out = 16'(-12039);
			230: out = 16'(-11825);
			231: out = 16'(-11420);
			232: out = 16'(-10837);
			233: out = 16'(-9919);
			234: out = 16'(-8404);
			235: out = 16'(-6718);
			236: out = 16'(-5129);
			237: out = 16'(-3805);
			238: out = 16'(-2738);
			239: out = 16'(-1552);
			240: out = 16'(-348);
			241: out = 16'(574);
			242: out = 16'(1436);
			243: out = 16'(2338);
			244: out = 16'(3618);
			245: out = 16'(5201);
			246: out = 16'(6692);
			247: out = 16'(7894);
			248: out = 16'(8843);
			249: out = 16'(9597);
			250: out = 16'(10182);
			251: out = 16'(10157);
			252: out = 16'(10031);
			253: out = 16'(9915);
			254: out = 16'(9529);
			255: out = 16'(8716);
			256: out = 16'(7519);
			257: out = 16'(6240);
			258: out = 16'(4988);
			259: out = 16'(3910);
			260: out = 16'(3038);
			261: out = 16'(2266);
			262: out = 16'(1493);
			263: out = 16'(202);
			264: out = 16'(-886);
			265: out = 16'(-1800);
			266: out = 16'(-2705);
			267: out = 16'(-3820);
			268: out = 16'(-5342);
			269: out = 16'(-7128);
			270: out = 16'(-8515);
			271: out = 16'(-9400);
			272: out = 16'(-9860);
			273: out = 16'(-9961);
			274: out = 16'(-9847);
			275: out = 16'(-9566);
			276: out = 16'(-9143);
			277: out = 16'(-8521);
			278: out = 16'(-7497);
			279: out = 16'(-6121);
			280: out = 16'(-4766);
			281: out = 16'(-3577);
			282: out = 16'(-2596);
			283: out = 16'(-1813);
			284: out = 16'(-680);
			285: out = 16'(163);
			286: out = 16'(880);
			287: out = 16'(1590);
			288: out = 16'(2467);
			289: out = 16'(3651);
			290: out = 16'(4944);
			291: out = 16'(6017);
			292: out = 16'(6891);
			293: out = 16'(7575);
			294: out = 16'(8149);
			295: out = 16'(8405);
			296: out = 16'(8332);
			297: out = 16'(8238);
			298: out = 16'(8080);
			299: out = 16'(7637);
			300: out = 16'(6826);
			301: out = 16'(5748);
			302: out = 16'(4656);
			303: out = 16'(3713);
			304: out = 16'(2889);
			305: out = 16'(2192);
			306: out = 16'(1660);
			307: out = 16'(670);
			308: out = 16'(-326);
			309: out = 16'(-1107);
			310: out = 16'(-1844);
			311: out = 16'(-2678);
			312: out = 16'(-3772);
			313: out = 16'(-5187);
			314: out = 16'(-6554);
			315: out = 16'(-7486);
			316: out = 16'(-8027);
			317: out = 16'(-8220);
			318: out = 16'(-8207);
			319: out = 16'(-8005);
			320: out = 16'(-7702);
			321: out = 16'(-7256);
			322: out = 16'(-6578);
			323: out = 16'(-5578);
			324: out = 16'(-4416);
			325: out = 16'(-3345);
			326: out = 16'(-2459);
			327: out = 16'(-1778);
			328: out = 16'(-978);
			329: out = 16'(-203);
			330: out = 16'(423);
			331: out = 16'(975);
			332: out = 16'(1608);
			333: out = 16'(2440);
			334: out = 16'(3499);
			335: out = 16'(4489);
			336: out = 16'(5312);
			337: out = 16'(5942);
			338: out = 16'(6468);
			339: out = 16'(6896);
			340: out = 16'(6889);
			341: out = 16'(6833);
			342: out = 16'(6741);
			343: out = 16'(6505);
			344: out = 16'(6012);
			345: out = 16'(5214);
			346: out = 16'(4332);
			347: out = 16'(3466);
			348: out = 16'(2737);
			349: out = 16'(2123);
			350: out = 16'(1607);
			351: out = 16'(1087);
			352: out = 16'(135);
			353: out = 16'(-576);
			354: out = 16'(-1222);
			355: out = 16'(-1860);
			356: out = 16'(-2614);
			357: out = 16'(-3640);
			358: out = 16'(-4836);
			359: out = 16'(-5814);
			360: out = 16'(-6427);
			361: out = 16'(-6705);
			362: out = 16'(-6782);
			363: out = 16'(-6681);
			364: out = 16'(-6474);
			365: out = 16'(-6176);
			366: out = 16'(-5745);
			367: out = 16'(-5046);
			368: out = 16'(-4131);
			369: out = 16'(-3197);
			370: out = 16'(-2398);
			371: out = 16'(-1750);
			372: out = 16'(-1219);
			373: out = 16'(-482);
			374: out = 16'(79);
			375: out = 16'(559);
			376: out = 16'(1035);
			377: out = 16'(1600);
			378: out = 16'(2370);
			379: out = 16'(3245);
			380: out = 16'(3988);
			381: out = 16'(4577);
			382: out = 16'(5066);
			383: out = 16'(5456);
			384: out = 16'(5694);
			385: out = 16'(5633);
			386: out = 16'(5592);
			387: out = 16'(5504);
			388: out = 16'(5240);
			389: out = 16'(4684);
			390: out = 16'(3945);
			391: out = 16'(3244);
			392: out = 16'(2584);
			393: out = 16'(2021);
			394: out = 16'(1536);
			395: out = 16'(1175);
			396: out = 16'(529);
			397: out = 16'(-151);
			398: out = 16'(-709);
			399: out = 16'(-1226);
			400: out = 16'(-1765);
			401: out = 16'(-2501);
			402: out = 16'(-3470);
			403: out = 16'(-4393);
			404: out = 16'(-5067);
			405: out = 16'(-5425);
			406: out = 16'(-5581);
			407: out = 16'(-5563);
			408: out = 16'(-5421);
			409: out = 16'(-5204);
			410: out = 16'(-4907);
			411: out = 16'(-4487);
			412: out = 16'(-3813);
			413: out = 16'(-3027);
			414: out = 16'(-2302);
			415: out = 16'(-1703);
			416: out = 16'(-1221);
			417: out = 16'(-704);
			418: out = 16'(-176);
			419: out = 16'(231);
			420: out = 16'(614);
			421: out = 16'(1011);
			422: out = 16'(1552);
			423: out = 16'(2240);
			424: out = 16'(2906);
			425: out = 16'(3458);
			426: out = 16'(3917);
			427: out = 16'(4255);
			428: out = 16'(4584);
			429: out = 16'(4642);
			430: out = 16'(4587);
			431: out = 16'(4554);
			432: out = 16'(4445);
			433: out = 16'(4140);
			434: out = 16'(3601);
			435: out = 16'(3013);
			436: out = 16'(2435);
			437: out = 16'(1923);
			438: out = 16'(1483);
			439: out = 16'(1125);
			440: out = 16'(811);
			441: out = 16'(154);
			442: out = 16'(-356);
			443: out = 16'(-798);
			444: out = 16'(-1221);
			445: out = 16'(-1717);
			446: out = 16'(-2384);
			447: out = 16'(-3214);
			448: out = 16'(-3890);
			449: out = 16'(-4343);
			450: out = 16'(-4523);
			451: out = 16'(-4590);
			452: out = 16'(-4507);
			453: out = 16'(-4370);
			454: out = 16'(-4172);
			455: out = 16'(-3886);
			456: out = 16'(-3442);
			457: out = 16'(-2836);
			458: out = 16'(-2211);
			459: out = 16'(-1650);
			460: out = 16'(-1205);
			461: out = 16'(-854);
			462: out = 16'(-372);
			463: out = 16'(5);
			464: out = 16'(316);
			465: out = 16'(622);
			466: out = 16'(980);
			467: out = 16'(1475);
			468: out = 16'(2067);
			469: out = 16'(2574);
			470: out = 16'(2984);
			471: out = 16'(3326);
			472: out = 16'(3600);
			473: out = 16'(3813);
			474: out = 16'(3775);
			475: out = 16'(3728);
			476: out = 16'(3686);
			477: out = 16'(3529);
			478: out = 16'(3201);
			479: out = 16'(2751);
			480: out = 16'(2262);
			481: out = 16'(1792);
			482: out = 16'(1402);
			483: out = 16'(1086);
			484: out = 16'(817);
			485: out = 16'(409);
			486: out = 16'(-62);
			487: out = 16'(-456);
			488: out = 16'(-793);
			489: out = 16'(-1166);
			490: out = 16'(-1637);
			491: out = 16'(-2258);
			492: out = 16'(-2907);
			493: out = 16'(-3371);
			494: out = 16'(-3640);
			495: out = 16'(-3736);
			496: out = 16'(-3731);
			497: out = 16'(-3652);
			498: out = 16'(-3501);
			499: out = 16'(-3308);
			500: out = 16'(-3030);
			501: out = 16'(-2606);
			502: out = 16'(-2085);
			503: out = 16'(-1604);
			504: out = 16'(-1188);
			505: out = 16'(-854);
			506: out = 16'(-531);
			507: out = 16'(-166);
			508: out = 16'(124);
			509: out = 16'(371);
			510: out = 16'(640);
			511: out = 16'(986);
			512: out = 16'(1426);
			513: out = 16'(1871);
			514: out = 16'(2257);
			515: out = 16'(2554);
			516: out = 16'(2815);
			517: out = 16'(3009);
			518: out = 16'(3079);
			519: out = 16'(3050);
			520: out = 16'(3013);
			521: out = 16'(2951);
			522: out = 16'(2763);
			523: out = 16'(2430);
			524: out = 16'(2034);
			525: out = 16'(1639);
			526: out = 16'(1294);
			527: out = 16'(1010);
			528: out = 16'(771);
			529: out = 16'(567);
			530: out = 16'(128);
			531: out = 16'(-227);
			532: out = 16'(-519);
			533: out = 16'(-797);
			534: out = 16'(-1134);
			535: out = 16'(-1574);
			536: out = 16'(-2125);
			537: out = 16'(-2582);
			538: out = 16'(-2885);
			539: out = 16'(-3028);
			540: out = 16'(-3068);
			541: out = 16'(-3026);
			542: out = 16'(-2923);
			543: out = 16'(-2782);
			544: out = 16'(-2599);
			545: out = 16'(-2329);
			546: out = 16'(-1921);
			547: out = 16'(-1507);
			548: out = 16'(-1146);
			549: out = 16'(-839);
			550: out = 16'(-589);
			551: out = 16'(-277);
			552: out = 16'(-26);
			553: out = 16'(188);
			554: out = 16'(388);
			555: out = 16'(626);
			556: out = 16'(948);
			557: out = 16'(1344);
			558: out = 16'(1675);
			559: out = 16'(1955);
			560: out = 16'(2172);
			561: out = 16'(2363);
			562: out = 16'(2492);
			563: out = 16'(2494);
			564: out = 16'(2491);
			565: out = 16'(2430);
			566: out = 16'(2339);
			567: out = 16'(2137);
			568: out = 16'(1819);
			569: out = 16'(1492);
			570: out = 16'(1193);
			571: out = 16'(936);
			572: out = 16'(711);
			573: out = 16'(531);
			574: out = 16'(273);
			575: out = 16'(-46);
			576: out = 16'(-304);
			577: out = 16'(-548);
			578: out = 16'(-779);
			579: out = 16'(-1073);
			580: out = 16'(-1497);
			581: out = 16'(-1935);
			582: out = 16'(-2245);
			583: out = 16'(-2428);
			584: out = 16'(-2499);
			585: out = 16'(-2486);
			586: out = 16'(-2434);
			587: out = 16'(-2347);
			588: out = 16'(-2218);
			589: out = 16'(-2043);
			590: out = 16'(-1754);
			591: out = 16'(-1404);
			592: out = 16'(-1082);
			593: out = 16'(-810);
			594: out = 16'(-592);
			595: out = 16'(-380);
			596: out = 16'(-139);
			597: out = 16'(46);
			598: out = 16'(223);
			599: out = 16'(388);
			600: out = 16'(613);
			601: out = 16'(901);
			602: out = 16'(1200);
			603: out = 16'(1452);
			604: out = 16'(1661);
			605: out = 16'(1828);
			606: out = 16'(1977);
			607: out = 16'(2022);
			608: out = 16'(2002);
			609: out = 16'(1986);
			610: out = 16'(1942);
			611: out = 16'(1832);
			612: out = 16'(1613);
			613: out = 16'(1353);
			614: out = 16'(1105);
			615: out = 16'(872);
			616: out = 16'(672);
			617: out = 16'(515);
			618: out = 16'(369);
			619: out = 16'(89);
			620: out = 16'(-147);
			621: out = 16'(-336);
			622: out = 16'(-526);
			623: out = 16'(-748);
			624: out = 16'(-1033);
			625: out = 16'(-1389);
			626: out = 16'(-1709);
			627: out = 16'(-1910);
			628: out = 16'(-2017);
			629: out = 16'(-2041);
			630: out = 16'(-2025);
			631: out = 16'(-1946);
			632: out = 16'(-1861);
			633: out = 16'(-1748);
			634: out = 16'(-1563);
			635: out = 16'(-1299);
			636: out = 16'(-1021);
			637: out = 16'(-784);
			638: out = 16'(-587);
			639: out = 16'(-413);
			640: out = 16'(-221);
			641: out = 16'(-44);
			642: out = 16'(101);
			643: out = 16'(239);
			644: out = 16'(381);
			645: out = 16'(589);
			646: out = 16'(831);
			647: out = 16'(1071);
			648: out = 16'(1249);
			649: out = 16'(1403);
			650: out = 16'(1520);
			651: out = 16'(1620);
			652: out = 16'(1618);
			653: out = 16'(1618);
			654: out = 16'(1607);
			655: out = 16'(1548);
			656: out = 16'(1410);
			657: out = 16'(1204);
			658: out = 16'(989);
			659: out = 16'(782);
			660: out = 16'(611);
			661: out = 16'(458);
			662: out = 16'(327);
			663: out = 16'(192);
			664: out = 16'(-28);
			665: out = 16'(-206);
			666: out = 16'(-351);
			667: out = 16'(-506);
			668: out = 16'(-707);
			669: out = 16'(-971);
			670: out = 16'(-1245);
			671: out = 16'(-1463);
			672: out = 16'(-1592);
			673: out = 16'(-1643);
			674: out = 16'(-1650);
			675: out = 16'(-1618);
			676: out = 16'(-1560);
			677: out = 16'(-1469);
			678: out = 16'(-1354);
			679: out = 16'(-1182);
			680: out = 16'(-962);
			681: out = 16'(-743);
			682: out = 16'(-555);
			683: out = 16'(-421);
			684: out = 16'(-281);
			685: out = 16'(-114);
			686: out = 16'(-5);
			687: out = 16'(113);
			688: out = 16'(230);
			689: out = 16'(375);
			690: out = 16'(557);
			691: out = 16'(752);
			692: out = 16'(938);
			693: out = 16'(1059);
			694: out = 16'(1168);
			695: out = 16'(1247);
			696: out = 16'(1305);
			697: out = 16'(1297);
			698: out = 16'(1286);
			699: out = 16'(1253);
			700: out = 16'(1190);
			701: out = 16'(1047);
			702: out = 16'(880);
			703: out = 16'(702);
			704: out = 16'(560);
			705: out = 16'(430);
			706: out = 16'(318);
			707: out = 16'(228);
			708: out = 16'(46);
			709: out = 16'(-93);
			710: out = 16'(-227);
			711: out = 16'(-341);
			712: out = 16'(-480);
			713: out = 16'(-671);
			714: out = 16'(-902);
			715: out = 16'(-1105);
			716: out = 16'(-1241);
			717: out = 16'(-1316);
			718: out = 16'(-1343);
			719: out = 16'(-1319);
			720: out = 16'(-1271);
			721: out = 16'(-1226);
			722: out = 16'(-1157);
			723: out = 16'(-1044);
			724: out = 16'(-876);
			725: out = 16'(-704);
			726: out = 16'(-528);
			727: out = 16'(-398);
			728: out = 16'(-281);
			729: out = 16'(-169);
			730: out = 16'(-45);
			731: out = 16'(38);
			732: out = 16'(128);
			733: out = 16'(218);
			734: out = 16'(346);
			735: out = 16'(510);
			736: out = 16'(661);
			737: out = 16'(787);
			738: out = 16'(878);
			739: out = 16'(964);
			740: out = 16'(1039);
			741: out = 16'(1035);
			742: out = 16'(1032);
			743: out = 16'(1022);
			744: out = 16'(987);
			745: out = 16'(904);
			746: out = 16'(774);
			747: out = 16'(630);
			748: out = 16'(502);
			749: out = 16'(379);
			750: out = 16'(289);
			751: out = 16'(210);
			752: out = 16'(128);
			753: out = 16'(-18);
			754: out = 16'(-140);
			755: out = 16'(-238);
			756: out = 16'(-327);
			757: out = 16'(-447);
			758: out = 16'(-621);
			759: out = 16'(-805);
			760: out = 16'(-948);
			761: out = 16'(-1044);
			762: out = 16'(-1075);
			763: out = 16'(-1083);
			764: out = 16'(-1044);
			765: out = 16'(-1019);
			766: out = 16'(-974);
			767: out = 16'(-898);
			768: out = 16'(-779);
			769: out = 16'(-647);
			770: out = 16'(-499);
			771: out = 16'(-386);
			772: out = 16'(-286);
			773: out = 16'(-209);
			774: out = 16'(-97);
			775: out = 16'(-16);
			776: out = 16'(54);
			777: out = 16'(128);
			778: out = 16'(220);
			779: out = 16'(332);
			780: out = 16'(459);
			781: out = 16'(560);
			782: out = 16'(655);
			783: out = 16'(729);
			784: out = 16'(789);
			785: out = 16'(810);
			786: out = 16'(805);
			787: out = 16'(793);
			788: out = 16'(778);
			789: out = 16'(747);
			790: out = 16'(668);
			791: out = 16'(542);
			792: out = 16'(441);
			793: out = 16'(345);
			794: out = 16'(257);
			795: out = 16'(187);
			796: out = 16'(128);
			797: out = 16'(30);
			798: out = 16'(-68);
			799: out = 16'(-154);
			800: out = 16'(-221);
			801: out = 16'(-318);
			802: out = 16'(-424);
			803: out = 16'(-581);
			804: out = 16'(-706);
			805: out = 16'(-794);
			806: out = 16'(-857);
			807: out = 16'(-867);
			808: out = 16'(-846);
			809: out = 16'(-841);
			810: out = 16'(-806);
			811: out = 16'(-744);
			812: out = 16'(-683);
			813: out = 16'(-584);
			814: out = 16'(-460);
			815: out = 16'(-365);
			816: out = 16'(-280);
			817: out = 16'(-203);
			818: out = 16'(-133);
			819: out = 16'(-51);
			820: out = 16'(9);
			821: out = 16'(70);
			822: out = 16'(127);
			823: out = 16'(219);
			824: out = 16'(309);
			825: out = 16'(404);
			826: out = 16'(474);
			827: out = 16'(547);
			828: out = 16'(587);
			829: out = 16'(633);
			830: out = 16'(623);
			831: out = 16'(633);
			832: out = 16'(614);
			833: out = 16'(602);
			834: out = 16'(549);
			835: out = 16'(477);
			836: out = 16'(392);
			837: out = 16'(314);
			838: out = 16'(231);
			839: out = 16'(173);
			840: out = 16'(121);
			841: out = 16'(67);
			842: out = 16'(-16);
			843: out = 16'(-102);
			844: out = 16'(-173);
			845: out = 16'(-210);
			846: out = 16'(-292);
			847: out = 16'(-396);
			848: out = 16'(-518);
			849: out = 16'(-605);
			850: out = 16'(-658);
			851: out = 16'(-681);
			852: out = 16'(-684);
			853: out = 16'(-663);
			854: out = 16'(-656);
			855: out = 16'(-610);
			856: out = 16'(-576);
			857: out = 16'(-509);
			858: out = 16'(-432);
			859: out = 16'(-330);
			860: out = 16'(-262);
			861: out = 16'(-193);
			862: out = 16'(-147);
			863: out = 16'(-76);
			864: out = 16'(-21);
			865: out = 16'(21);
			866: out = 16'(67);
			867: out = 16'(113);
			868: out = 16'(194);
			869: out = 16'(276);
			870: out = 16'(333);
			871: out = 16'(386);
			872: out = 16'(444);
			873: out = 16'(486);
			874: out = 16'(493);
			875: out = 16'(490);
			876: out = 16'(470);
			877: out = 16'(472);
			878: out = 16'(444);
			879: out = 16'(391);
			880: out = 16'(327);
			881: out = 16'(253);
			882: out = 16'(193);
			883: out = 16'(139);
			884: out = 16'(98);
			885: out = 16'(53);
			886: out = 16'(5);
			887: out = 16'(-60);
			888: out = 16'(-104);
			889: out = 16'(-156);
			890: out = 16'(-206);
			891: out = 16'(-261);
			892: out = 16'(-365);
			893: out = 16'(-445);
			894: out = 16'(-503);
			895: out = 16'(-540);
			896: out = 16'(-533);
			897: out = 16'(-537);
			898: out = 16'(-519);
			899: out = 16'(-515);
			900: out = 16'(-486);
			901: out = 16'(-433);
			902: out = 16'(-369);
			903: out = 16'(-298);
			904: out = 16'(-241);
			905: out = 16'(-183);
			906: out = 16'(-143);
			907: out = 16'(-95);
			908: out = 16'(-44);
			909: out = 16'(-15);
			910: out = 16'(19);
			911: out = 16'(51);
			912: out = 16'(116);
			913: out = 16'(174);
			914: out = 16'(232);
			915: out = 16'(283);
			916: out = 16'(312);
			917: out = 16'(338);
			918: out = 16'(369);
			919: out = 16'(363);
			920: out = 16'(348);
			921: out = 16'(352);
			922: out = 16'(342);
			923: out = 16'(311);
			924: out = 16'(269);
			925: out = 16'(210);
			926: out = 16'(167);
			927: out = 16'(112);
			928: out = 16'(83);
			929: out = 16'(52);
			930: out = 16'(30);
			931: out = 16'(-24);
			932: out = 16'(-83);
			933: out = 16'(-116);
			934: out = 16'(-144);
			935: out = 16'(-192);
			936: out = 16'(-249);
			937: out = 16'(-313);
			938: out = 16'(-367);
			939: out = 16'(-394);
			940: out = 16'(-415);
			941: out = 16'(-420);
			942: out = 16'(-421);
			943: out = 16'(-411);
			944: out = 16'(-382);
			945: out = 16'(-365);
			946: out = 16'(-322);
			947: out = 16'(-275);
			948: out = 16'(-219);
			949: out = 16'(-176);
			950: out = 16'(-141);
			951: out = 16'(-113);
			952: out = 16'(-63);
			953: out = 16'(-25);
			954: out = 16'(1);
			955: out = 16'(33);
			956: out = 16'(52);
			957: out = 16'(96);
			958: out = 16'(135);
			959: out = 16'(186);
			960: out = 16'(220);
			961: out = 16'(255);
			962: out = 16'(263);
			963: out = 16'(282);
			964: out = 16'(267);
			965: out = 16'(267);
			966: out = 16'(251);
			967: out = 16'(237);
			968: out = 16'(203);
			969: out = 16'(175);
			970: out = 16'(139);
			971: out = 16'(89);
			972: out = 16'(73);
			973: out = 16'(37);
			974: out = 16'(25);
			975: out = 16'(-16);
			976: out = 16'(-49);
			977: out = 16'(-72);
			978: out = 16'(-113);
			979: out = 16'(-132);
			980: out = 16'(-175);
			981: out = 16'(-226);
			982: out = 16'(-271);
			983: out = 16'(-300);
			984: out = 16'(-313);
			985: out = 16'(-333);
			986: out = 16'(-327);
			987: out = 16'(-328);
			988: out = 16'(-309);
			989: out = 16'(-299);
			990: out = 16'(-283);
			991: out = 16'(-241);
			992: out = 16'(-203);
			993: out = 16'(-150);
			994: out = 16'(-131);
			995: out = 16'(-104);
			996: out = 16'(-79);
			997: out = 16'(-49);
			998: out = 16'(-25);
			999: out = 16'(-13);
			1000: out = 16'(13);
			1001: out = 16'(50);
			1002: out = 16'(83);
			1003: out = 16'(113);
			1004: out = 16'(143);
			1005: out = 16'(166);
			1006: out = 16'(182);
			1007: out = 16'(198);
			1008: out = 16'(190);
			1009: out = 16'(179);
			1010: out = 16'(173);
			1011: out = 16'(176);
			1012: out = 16'(149);
			1013: out = 16'(140);
			1014: out = 16'(107);
			1015: out = 16'(75);
			1016: out = 16'(50);
			1017: out = 16'(24);
			1018: out = 16'(12);
			1019: out = 16'(-14);
			1020: out = 16'(-37);
			1021: out = 16'(-43);
			1022: out = 16'(-74);
			1023: out = 16'(-101);
			1024: out = 16'(-122);
			1025: out = 16'(-160);
			1026: out = 16'(-185);
			1027: out = 16'(-222);
			1028: out = 16'(-235);
			1029: out = 16'(-245);
			1030: out = 16'(-261);
			1031: out = 16'(-253);
			1032: out = 16'(-252);
			1033: out = 16'(-242);
			1034: out = 16'(-210);
			1035: out = 16'(-196);
			1036: out = 16'(-176);
			1037: out = 16'(-136);
			1038: out = 16'(-121);
			1039: out = 16'(-97);
			1040: out = 16'(-80);
			1041: out = 16'(-60);
			1042: out = 16'(-31);
			1043: out = 16'(-19);
			1044: out = 16'(-8);
			1045: out = 16'(6);
			1046: out = 16'(37);
			1047: out = 16'(58);
			1048: out = 16'(85);
			1049: out = 16'(107);
			1050: out = 16'(123);
			1051: out = 16'(133);
			1052: out = 16'(132);
			1053: out = 16'(125);
			1054: out = 16'(124);
			1055: out = 16'(121);
			1056: out = 16'(105);
			1057: out = 16'(99);
			1058: out = 16'(72);
			1059: out = 16'(49);
			1060: out = 16'(28);
			1061: out = 16'(19);
			1062: out = 16'(2);
			1063: out = 16'(-19);
			1064: out = 16'(-24);
			1065: out = 16'(-44);
			1066: out = 16'(-58);
			1067: out = 16'(-67);
			1068: out = 16'(-86);
			1069: out = 16'(-107);
			1070: out = 16'(-128);
			1071: out = 16'(-164);
			1072: out = 16'(-166);
			1073: out = 16'(-181);
			1074: out = 16'(-190);
			1075: out = 16'(-182);
			1076: out = 16'(-182);
			1077: out = 16'(-187);
			1078: out = 16'(-184);
			1079: out = 16'(-164);
			1080: out = 16'(-158);
			1081: out = 16'(-124);
			1082: out = 16'(-108);
			1083: out = 16'(-96);
			1084: out = 16'(-77);
			1085: out = 16'(-63);
			1086: out = 16'(-43);
			1087: out = 16'(-38);
			1088: out = 16'(-22);
			1089: out = 16'(-6);
			default: out = 0;
		endcase
	end
endmodule
