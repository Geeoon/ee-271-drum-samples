module snare_lookup(index, out);
	input logic unsigned [10:0] index;
	output logic signed [15:0] out;
	always_comb begin
		case(index)
			0: out = 16'(18770);
			1: out = 16'(23562);
			2: out = 16'(-5407);
			3: out = 16'(-10684);
			4: out = 16'(-11558);
			5: out = 16'(8095);
			6: out = 16'(30798);
			7: out = 16'(30600);
			8: out = 16'(30118);
			9: out = 16'(-7249);
			10: out = 16'(-30870);
			11: out = 16'(-30972);
			12: out = 16'(-6742);
			13: out = 16'(17035);
			14: out = 16'(29874);
			15: out = 16'(22155);
			16: out = 16'(11605);
			17: out = 16'(7102);
			18: out = 16'(16283);
			19: out = 16'(-13815);
			20: out = 16'(-22260);
			21: out = 16'(-29694);
			22: out = 16'(-30593);
			23: out = 16'(-9507);
			24: out = 16'(-12737);
			25: out = 16'(1156);
			26: out = 16'(31498);
			27: out = 16'(30724);
			28: out = 16'(21298);
			29: out = 16'(30081);
			30: out = 16'(15219);
			31: out = 16'(-2812);
			32: out = 16'(-14276);
			33: out = 16'(-27097);
			34: out = 16'(-30867);
			35: out = 16'(-30064);
			36: out = 16'(-29834);
			37: out = 16'(-16674);
			38: out = 16'(13010);
			39: out = 16'(18157);
			40: out = 16'(18243);
			41: out = 16'(15475);
			42: out = 16'(20172);
			43: out = 16'(10716);
			44: out = 16'(-9944);
			45: out = 16'(1129);
			46: out = 16'(-12082);
			47: out = 16'(1921);
			48: out = 16'(-335);
			49: out = 16'(-14748);
			50: out = 16'(-8447);
			51: out = 16'(-27055);
			52: out = 16'(-16243);
			53: out = 16'(-1326);
			54: out = 16'(6355);
			55: out = 16'(13578);
			56: out = 16'(944);
			57: out = 16'(6651);
			58: out = 16'(5425);
			59: out = 16'(20229);
			60: out = 16'(11723);
			61: out = 16'(16964);
			62: out = 16'(15259);
			63: out = 16'(2689);
			64: out = 16'(-20218);
			65: out = 16'(5100);
			66: out = 16'(-20329);
			67: out = 16'(-16545);
			68: out = 16'(-19195);
			69: out = 16'(-11764);
			70: out = 16'(-17330);
			71: out = 16'(-17904);
			72: out = 16'(4015);
			73: out = 16'(-3798);
			74: out = 16'(20098);
			75: out = 16'(19988);
			76: out = 16'(-3723);
			77: out = 16'(16241);
			78: out = 16'(13562);
			79: out = 16'(-7728);
			80: out = 16'(1820);
			81: out = 16'(-13190);
			82: out = 16'(-19118);
			83: out = 16'(-9442);
			84: out = 16'(-13499);
			85: out = 16'(-8507);
			86: out = 16'(-4942);
			87: out = 16'(-9413);
			88: out = 16'(-7822);
			89: out = 16'(3162);
			90: out = 16'(-5996);
			91: out = 16'(4253);
			92: out = 16'(-3219);
			93: out = 16'(3867);
			94: out = 16'(-5881);
			95: out = 16'(-4421);
			96: out = 16'(4436);
			97: out = 16'(-5944);
			98: out = 16'(14351);
			99: out = 16'(-15282);
			100: out = 16'(217);
			101: out = 16'(-464);
			102: out = 16'(-10266);
			103: out = 16'(-1070);
			104: out = 16'(-7906);
			105: out = 16'(-10818);
			106: out = 16'(-8367);
			107: out = 16'(-9242);
			108: out = 16'(-3671);
			109: out = 16'(-4379);
			110: out = 16'(-1705);
			111: out = 16'(3265);
			112: out = 16'(2789);
			113: out = 16'(6369);
			114: out = 16'(3638);
			115: out = 16'(13495);
			116: out = 16'(5681);
			117: out = 16'(-1384);
			118: out = 16'(9040);
			119: out = 16'(-6630);
			120: out = 16'(-2822);
			121: out = 16'(8676);
			122: out = 16'(-4996);
			123: out = 16'(-5724);
			124: out = 16'(-243);
			125: out = 16'(9441);
			126: out = 16'(4021);
			127: out = 16'(8661);
			128: out = 16'(-3271);
			129: out = 16'(2315);
			130: out = 16'(5681);
			131: out = 16'(15900);
			132: out = 16'(-1534);
			133: out = 16'(12642);
			134: out = 16'(11799);
			135: out = 16'(-4983);
			136: out = 16'(12855);
			137: out = 16'(-4646);
			138: out = 16'(-4053);
			139: out = 16'(7507);
			140: out = 16'(1101);
			141: out = 16'(4506);
			142: out = 16'(16490);
			143: out = 16'(10007);
			144: out = 16'(-606);
			145: out = 16'(-9698);
			146: out = 16'(-6807);
			147: out = 16'(15406);
			148: out = 16'(872);
			149: out = 16'(800);
			150: out = 16'(2863);
			151: out = 16'(9268);
			152: out = 16'(124);
			153: out = 16'(10899);
			154: out = 16'(-1664);
			155: out = 16'(7361);
			156: out = 16'(-455);
			157: out = 16'(-8705);
			158: out = 16'(-11612);
			159: out = 16'(3656);
			160: out = 16'(10170);
			161: out = 16'(-3258);
			162: out = 16'(-751);
			163: out = 16'(1910);
			164: out = 16'(4027);
			165: out = 16'(-7260);
			166: out = 16'(-2346);
			167: out = 16'(-795);
			168: out = 16'(4263);
			169: out = 16'(9684);
			170: out = 16'(-354);
			171: out = 16'(-1649);
			172: out = 16'(-2635);
			173: out = 16'(-10314);
			174: out = 16'(-10556);
			175: out = 16'(1731);
			176: out = 16'(1885);
			177: out = 16'(14427);
			178: out = 16'(131);
			179: out = 16'(-806);
			180: out = 16'(-10208);
			181: out = 16'(3286);
			182: out = 16'(-1712);
			183: out = 16'(5759);
			184: out = 16'(-582);
			185: out = 16'(-1388);
			186: out = 16'(4432);
			187: out = 16'(3599);
			188: out = 16'(-8425);
			189: out = 16'(-1768);
			190: out = 16'(10290);
			191: out = 16'(-5647);
			192: out = 16'(-7464);
			193: out = 16'(299);
			194: out = 16'(632);
			195: out = 16'(-5970);
			196: out = 16'(3975);
			197: out = 16'(2333);
			198: out = 16'(-3973);
			199: out = 16'(-2250);
			200: out = 16'(1190);
			201: out = 16'(11318);
			202: out = 16'(-14713);
			203: out = 16'(4560);
			204: out = 16'(-184);
			205: out = 16'(4592);
			206: out = 16'(8879);
			207: out = 16'(-8101);
			208: out = 16'(3063);
			209: out = 16'(-9766);
			210: out = 16'(2886);
			211: out = 16'(5981);
			212: out = 16'(5476);
			213: out = 16'(-944);
			214: out = 16'(-14715);
			215: out = 16'(-2521);
			216: out = 16'(-6098);
			217: out = 16'(-3608);
			218: out = 16'(9219);
			219: out = 16'(2825);
			220: out = 16'(7321);
			221: out = 16'(1362);
			222: out = 16'(4122);
			223: out = 16'(-8337);
			224: out = 16'(-5120);
			225: out = 16'(1768);
			226: out = 16'(523);
			227: out = 16'(-6001);
			228: out = 16'(525);
			229: out = 16'(-5131);
			230: out = 16'(-4340);
			231: out = 16'(-12847);
			232: out = 16'(-13233);
			233: out = 16'(1784);
			234: out = 16'(-1749);
			235: out = 16'(-11623);
			236: out = 16'(2443);
			237: out = 16'(6298);
			238: out = 16'(-4006);
			239: out = 16'(-309);
			240: out = 16'(-2379);
			241: out = 16'(4992);
			242: out = 16'(2634);
			243: out = 16'(-759);
			244: out = 16'(-5785);
			245: out = 16'(-8120);
			246: out = 16'(5406);
			247: out = 16'(-7041);
			248: out = 16'(7833);
			249: out = 16'(-4920);
			250: out = 16'(11571);
			251: out = 16'(-4354);
			252: out = 16'(-3958);
			253: out = 16'(-10906);
			254: out = 16'(-3960);
			255: out = 16'(-6229);
			256: out = 16'(-4418);
			257: out = 16'(2015);
			258: out = 16'(-6293);
			259: out = 16'(11337);
			260: out = 16'(3625);
			261: out = 16'(-2006);
			262: out = 16'(-4246);
			263: out = 16'(-1229);
			264: out = 16'(-842);
			265: out = 16'(4881);
			266: out = 16'(-2463);
			267: out = 16'(-8489);
			268: out = 16'(-15586);
			269: out = 16'(1196);
			270: out = 16'(-3968);
			271: out = 16'(3653);
			272: out = 16'(205);
			273: out = 16'(-16063);
			274: out = 16'(4694);
			275: out = 16'(5428);
			276: out = 16'(-7733);
			277: out = 16'(-3350);
			278: out = 16'(-1091);
			279: out = 16'(-814);
			280: out = 16'(9949);
			281: out = 16'(9934);
			282: out = 16'(-4447);
			283: out = 16'(-9190);
			284: out = 16'(-2868);
			285: out = 16'(-838);
			286: out = 16'(1725);
			287: out = 16'(-4390);
			288: out = 16'(4411);
			289: out = 16'(7321);
			290: out = 16'(577);
			291: out = 16'(4955);
			292: out = 16'(-470);
			293: out = 16'(-5982);
			294: out = 16'(-4847);
			295: out = 16'(8673);
			296: out = 16'(-5529);
			297: out = 16'(1970);
			298: out = 16'(950);
			299: out = 16'(-4098);
			300: out = 16'(-2745);
			301: out = 16'(8008);
			302: out = 16'(-1143);
			303: out = 16'(-3570);
			304: out = 16'(187);
			305: out = 16'(-10485);
			306: out = 16'(-5140);
			307: out = 16'(-8614);
			308: out = 16'(3819);
			309: out = 16'(-3975);
			310: out = 16'(-4595);
			311: out = 16'(1443);
			312: out = 16'(-3321);
			313: out = 16'(7239);
			314: out = 16'(-2568);
			315: out = 16'(-1583);
			316: out = 16'(3413);
			317: out = 16'(-8233);
			318: out = 16'(6032);
			319: out = 16'(193);
			320: out = 16'(-4302);
			321: out = 16'(5483);
			322: out = 16'(-4048);
			323: out = 16'(1912);
			324: out = 16'(3370);
			325: out = 16'(-4431);
			326: out = 16'(4188);
			327: out = 16'(267);
			328: out = 16'(811);
			329: out = 16'(-5720);
			330: out = 16'(2239);
			331: out = 16'(-11524);
			332: out = 16'(6813);
			333: out = 16'(-2284);
			334: out = 16'(-2098);
			335: out = 16'(8106);
			336: out = 16'(2951);
			337: out = 16'(1434);
			338: out = 16'(5445);
			339: out = 16'(6455);
			340: out = 16'(2701);
			341: out = 16'(-2373);
			342: out = 16'(2471);
			343: out = 16'(7676);
			344: out = 16'(-1861);
			345: out = 16'(-2884);
			346: out = 16'(4131);
			347: out = 16'(-462);
			348: out = 16'(3188);
			349: out = 16'(-6504);
			350: out = 16'(-7688);
			351: out = 16'(4399);
			352: out = 16'(-784);
			353: out = 16'(4106);
			354: out = 16'(-1801);
			355: out = 16'(-1526);
			356: out = 16'(-7904);
			357: out = 16'(7762);
			358: out = 16'(-5557);
			359: out = 16'(3504);
			360: out = 16'(3357);
			361: out = 16'(-1472);
			362: out = 16'(1033);
			363: out = 16'(820);
			364: out = 16'(-1119);
			365: out = 16'(5435);
			366: out = 16'(482);
			367: out = 16'(3456);
			368: out = 16'(4431);
			369: out = 16'(4695);
			370: out = 16'(2743);
			371: out = 16'(-2955);
			372: out = 16'(-2904);
			373: out = 16'(4493);
			374: out = 16'(-499);
			375: out = 16'(-1666);
			376: out = 16'(556);
			377: out = 16'(-3919);
			378: out = 16'(-3313);
			379: out = 16'(-4170);
			380: out = 16'(-4756);
			381: out = 16'(2991);
			382: out = 16'(-533);
			383: out = 16'(-1447);
			384: out = 16'(3182);
			385: out = 16'(-4134);
			386: out = 16'(435);
			387: out = 16'(-1095);
			388: out = 16'(-164);
			389: out = 16'(2648);
			390: out = 16'(-6875);
			391: out = 16'(-2694);
			392: out = 16'(-3641);
			393: out = 16'(229);
			394: out = 16'(-631);
			395: out = 16'(-1523);
			396: out = 16'(5044);
			397: out = 16'(496);
			398: out = 16'(904);
			399: out = 16'(128);
			400: out = 16'(1931);
			401: out = 16'(-190);
			402: out = 16'(215);
			403: out = 16'(-5983);
			404: out = 16'(-810);
			405: out = 16'(2824);
			406: out = 16'(-2040);
			407: out = 16'(-1769);
			408: out = 16'(2227);
			409: out = 16'(-2125);
			410: out = 16'(3043);
			411: out = 16'(-3500);
			412: out = 16'(3147);
			413: out = 16'(2824);
			414: out = 16'(-1034);
			415: out = 16'(-3081);
			416: out = 16'(-2153);
			417: out = 16'(-1221);
			418: out = 16'(319);
			419: out = 16'(1786);
			420: out = 16'(-4645);
			421: out = 16'(1573);
			422: out = 16'(-1849);
			423: out = 16'(-220);
			424: out = 16'(-2585);
			425: out = 16'(231);
			426: out = 16'(1);
			427: out = 16'(-4834);
			428: out = 16'(-3069);
			429: out = 16'(-2348);
			430: out = 16'(3941);
			431: out = 16'(-707);
			432: out = 16'(2287);
			433: out = 16'(2323);
			434: out = 16'(936);
			435: out = 16'(2821);
			436: out = 16'(-4816);
			437: out = 16'(145);
			438: out = 16'(-3443);
			439: out = 16'(-432);
			440: out = 16'(-1259);
			441: out = 16'(1125);
			442: out = 16'(1913);
			443: out = 16'(-597);
			444: out = 16'(-6055);
			445: out = 16'(-944);
			446: out = 16'(396);
			447: out = 16'(-1106);
			448: out = 16'(-2725);
			449: out = 16'(-905);
			450: out = 16'(265);
			451: out = 16'(1417);
			452: out = 16'(-4645);
			453: out = 16'(-960);
			454: out = 16'(3448);
			455: out = 16'(-1347);
			456: out = 16'(-2237);
			457: out = 16'(-971);
			458: out = 16'(1171);
			459: out = 16'(76);
			460: out = 16'(936);
			461: out = 16'(-830);
			462: out = 16'(4944);
			463: out = 16'(4229);
			464: out = 16'(668);
			465: out = 16'(-3111);
			466: out = 16'(914);
			467: out = 16'(1289);
			468: out = 16'(1287);
			469: out = 16'(-3420);
			470: out = 16'(833);
			471: out = 16'(-595);
			472: out = 16'(-1219);
			473: out = 16'(2399);
			474: out = 16'(-146);
			475: out = 16'(-1727);
			476: out = 16'(-1732);
			477: out = 16'(-614);
			478: out = 16'(-4558);
			479: out = 16'(-2473);
			480: out = 16'(498);
			481: out = 16'(561);
			482: out = 16'(-539);
			483: out = 16'(-216);
			484: out = 16'(-159);
			485: out = 16'(-2143);
			486: out = 16'(402);
			487: out = 16'(2403);
			488: out = 16'(-3631);
			489: out = 16'(-2498);
			490: out = 16'(645);
			491: out = 16'(1608);
			492: out = 16'(-1310);
			493: out = 16'(1631);
			494: out = 16'(114);
			495: out = 16'(3030);
			496: out = 16'(-715);
			497: out = 16'(2259);
			498: out = 16'(-414);
			499: out = 16'(1067);
			500: out = 16'(1015);
			501: out = 16'(-1820);
			502: out = 16'(367);
			503: out = 16'(2207);
			504: out = 16'(-1961);
			505: out = 16'(-21);
			506: out = 16'(-569);
			507: out = 16'(-795);
			508: out = 16'(-113);
			509: out = 16'(-1300);
			510: out = 16'(-310);
			511: out = 16'(2287);
			512: out = 16'(1115);
			513: out = 16'(-885);
			514: out = 16'(1658);
			515: out = 16'(-1218);
			516: out = 16'(-2133);
			517: out = 16'(143);
			518: out = 16'(609);
			519: out = 16'(-970);
			520: out = 16'(-1546);
			521: out = 16'(-1280);
			522: out = 16'(1405);
			523: out = 16'(631);
			524: out = 16'(-272);
			525: out = 16'(361);
			526: out = 16'(738);
			527: out = 16'(-2068);
			528: out = 16'(-421);
			529: out = 16'(-609);
			530: out = 16'(562);
			531: out = 16'(909);
			532: out = 16'(1920);
			533: out = 16'(666);
			534: out = 16'(-443);
			535: out = 16'(-289);
			536: out = 16'(-1013);
			537: out = 16'(1307);
			538: out = 16'(956);
			539: out = 16'(-385);
			540: out = 16'(-722);
			541: out = 16'(2);
			542: out = 16'(-228);
			543: out = 16'(455);
			544: out = 16'(-817);
			545: out = 16'(-796);
			546: out = 16'(654);
			547: out = 16'(-418);
			548: out = 16'(-262);
			549: out = 16'(-631);
			550: out = 16'(-907);
			551: out = 16'(-706);
			552: out = 16'(481);
			553: out = 16'(497);
			554: out = 16'(486);
			555: out = 16'(737);
			556: out = 16'(-825);
			557: out = 16'(-1510);
			558: out = 16'(-506);
			559: out = 16'(147);
			560: out = 16'(-923);
			561: out = 16'(749);
			562: out = 16'(-267);
			563: out = 16'(1317);
			564: out = 16'(-385);
			565: out = 16'(379);
			566: out = 16'(414);
			567: out = 16'(61);
			568: out = 16'(-518);
			569: out = 16'(384);
			570: out = 16'(542);
			571: out = 16'(789);
			572: out = 16'(-58);
			573: out = 16'(-690);
			574: out = 16'(778);
			575: out = 16'(362);
			576: out = 16'(-246);
			577: out = 16'(-836);
			578: out = 16'(293);
			579: out = 16'(331);
			580: out = 16'(-382);
			581: out = 16'(-299);
			582: out = 16'(40);
			583: out = 16'(-709);
			584: out = 16'(-211);
			585: out = 16'(48);
			586: out = 16'(66);
			587: out = 16'(-203);
			default: out = 0;
		endcase
	end
endmodule
