module closed_hihat_lookup(index, out);
	input logic unsigned [12:0] index;
	output logic signed [23:0] out;
	always_comb begin
		case(index)
			0: out = 24'(0);
			1: out = 24'(0);
			2: out = 24'(128);
			3: out = 24'(-476);
			4: out = 24'(232);
			5: out = 24'(-612);
			6: out = 24'(368);
			7: out = 24'(-760);
			8: out = 24'(544);
			9: out = 24'(-984);
			10: out = 24'(800);
			11: out = 24'(-1276);
			12: out = 24'(1188);
			13: out = 24'(-1932);
			14: out = 24'(2188);
			15: out = 24'(-3512);
			16: out = 24'(5228);
			17: out = 24'(-14560);
			18: out = 24'(41252);
			19: out = 24'(112940);
			20: out = 24'(-31780);
			21: out = 24'(-59212);
			22: out = 24'(-42624);
			23: out = 24'(67588);
			24: out = 24'(46124);
			25: out = 24'(101904);
			26: out = 24'(72372);
			27: out = 24'(-96064);
			28: out = 24'(-128932);
			29: out = 24'(-75892);
			30: out = 24'(87560);
			31: out = 24'(131064);
			32: out = 24'(10640);
			33: out = 24'(-107096);
			34: out = 24'(11020);
			35: out = 24'(77636);
			36: out = 24'(75056);
			37: out = 24'(8508);
			38: out = 24'(-92360);
			39: out = 24'(-26264);
			40: out = 24'(100120);
			41: out = 24'(53540);
			42: out = 24'(-15544);
			43: out = 24'(-86164);
			44: out = 24'(-25480);
			45: out = 24'(-76668);
			46: out = 24'(54444);
			47: out = 24'(116332);
			48: out = 24'(41532);
			49: out = 24'(-86876);
			50: out = 24'(-106452);
			51: out = 24'(11400);
			52: out = 24'(105200);
			53: out = 24'(87008);
			54: out = 24'(-15560);
			55: out = 24'(-108880);
			56: out = 24'(-121568);
			57: out = 24'(-72672);
			58: out = 24'(41324);
			59: out = 24'(50168);
			60: out = 24'(113684);
			61: out = 24'(103800);
			62: out = 24'(-8452);
			63: out = 24'(-116484);
			64: out = 24'(-84512);
			65: out = 24'(39388);
			66: out = 24'(9828);
			67: out = 24'(-76324);
			68: out = 24'(-85324);
			69: out = 24'(82424);
			70: out = 24'(89440);
			71: out = 24'(26264);
			72: out = 24'(-79912);
			73: out = 24'(-88608);
			74: out = 24'(-10676);
			75: out = 24'(25572);
			76: out = 24'(-131068);
			77: out = 24'(42980);
			78: out = 24'(124572);
			79: out = 24'(111000);
			80: out = 24'(-86532);
			81: out = 24'(-87048);
			82: out = 24'(16236);
			83: out = 24'(119872);
			84: out = 24'(30280);
			85: out = 24'(45472);
			86: out = 24'(100700);
			87: out = 24'(8788);
			88: out = 24'(-90452);
			89: out = 24'(-118312);
			90: out = 24'(-3276);
			91: out = 24'(90796);
			92: out = 24'(106864);
			93: out = 24'(62912);
			94: out = 24'(-64444);
			95: out = 24'(-109460);
			96: out = 24'(-116676);
			97: out = 24'(-111372);
			98: out = 24'(-66124);
			99: out = 24'(24588);
			100: out = 24'(73540);
			101: out = 24'(36152);
			102: out = 24'(-10720);
			103: out = 24'(-23732);
			104: out = 24'(-20772);
			105: out = 24'(83060);
			106: out = 24'(-9500);
			107: out = 24'(-125884);
			108: out = 24'(-119148);
			109: out = 24'(-42280);
			110: out = 24'(93804);
			111: out = 24'(47436);
			112: out = 24'(-66960);
			113: out = 24'(-118488);
			114: out = 24'(-45392);
			115: out = 24'(-127136);
			116: out = 24'(18784);
			117: out = 24'(12772);
			118: out = 24'(-111616);
			119: out = 24'(-123988);
			120: out = 24'(-10096);
			121: out = 24'(94900);
			122: out = 24'(-90320);
			123: out = 24'(-90172);
			124: out = 24'(-84900);
			125: out = 24'(-45044);
			126: out = 24'(-75920);
			127: out = 24'(-83868);
			128: out = 24'(-78056);
			129: out = 24'(76596);
			130: out = 24'(-61156);
			131: out = 24'(-101228);
			132: out = 24'(-11532);
			133: out = 24'(-34192);
			134: out = 24'(-74860);
			135: out = 24'(-112044);
			136: out = 24'(-99276);
			137: out = 24'(-31380);
			138: out = 24'(12088);
			139: out = 24'(-7792);
			140: out = 24'(-101824);
			141: out = 24'(-84384);
			142: out = 24'(-20972);
			143: out = 24'(-103548);
			144: out = 24'(-3028);
			145: out = 24'(55480);
			146: out = 24'(43692);
			147: out = 24'(-49452);
			148: out = 24'(-94792);
			149: out = 24'(-12376);
			150: out = 24'(126304);
			151: out = 24'(116908);
			152: out = 24'(108376);
			153: out = 24'(-492);
			154: out = 24'(-107464);
			155: out = 24'(-119360);
			156: out = 24'(-96916);
			157: out = 24'(29960);
			158: out = 24'(116832);
			159: out = 24'(104108);
			160: out = 24'(51300);
			161: out = 24'(-27976);
			162: out = 24'(-9288);
			163: out = 24'(44716);
			164: out = 24'(69212);
			165: out = 24'(9584);
			166: out = 24'(-76944);
			167: out = 24'(-119636);
			168: out = 24'(-89472);
			169: out = 24'(-52768);
			170: out = 24'(484);
			171: out = 24'(67560);
			172: out = 24'(20628);
			173: out = 24'(-63852);
			174: out = 24'(-93652);
			175: out = 24'(96720);
			176: out = 24'(127924);
			177: out = 24'(100888);
			178: out = 24'(26768);
			179: out = 24'(-52820);
			180: out = 24'(-69844);
			181: out = 24'(-1512);
			182: out = 24'(109456);
			183: out = 24'(121604);
			184: out = 24'(121436);
			185: out = 24'(119076);
			186: out = 24'(107112);
			187: out = 24'(28456);
			188: out = 24'(-53108);
			189: out = 24'(-117296);
			190: out = 24'(-44816);
			191: out = 24'(61104);
			192: out = 24'(119152);
			193: out = 24'(-23644);
			194: out = 24'(-63720);
			195: out = 24'(-1808);
			196: out = 24'(105428);
			197: out = 24'(62444);
			198: out = 24'(-11676);
			199: out = 24'(-72500);
			200: out = 24'(19424);
			201: out = 24'(45260);
			202: out = 24'(54684);
			203: out = 24'(113492);
			204: out = 24'(122624);
			205: out = 24'(36848);
			206: out = 24'(-115656);
			207: out = 24'(-90208);
			208: out = 24'(35064);
			209: out = 24'(131064);
			210: out = 24'(112716);
			211: out = 24'(108092);
			212: out = 24'(59008);
			213: out = 24'(-8400);
			214: out = 24'(-97928);
			215: out = 24'(-124916);
			216: out = 24'(-77240);
			217: out = 24'(102744);
			218: out = 24'(129884);
			219: out = 24'(60208);
			220: out = 24'(-83796);
			221: out = 24'(46004);
			222: out = 24'(97572);
			223: out = 24'(73216);
			224: out = 24'(-103568);
			225: out = 24'(-61028);
			226: out = 24'(-38328);
			227: out = 24'(-81760);
			228: out = 24'(81944);
			229: out = 24'(60224);
			230: out = 24'(18920);
			231: out = 24'(23116);
			232: out = 24'(91320);
			233: out = 24'(84952);
			234: out = 24'(4928);
			235: out = 24'(-61976);
			236: out = 24'(-19932);
			237: out = 24'(62364);
			238: out = 24'(-11080);
			239: out = 24'(46296);
			240: out = 24'(6940);
			241: out = 24'(-29720);
			242: out = 24'(-67760);
			243: out = 24'(42204);
			244: out = 24'(102592);
			245: out = 24'(19356);
			246: out = 24'(-25628);
			247: out = 24'(-83172);
			248: out = 24'(-96092);
			249: out = 24'(97836);
			250: out = 24'(48040);
			251: out = 24'(-71652);
			252: out = 24'(-120796);
			253: out = 24'(-67840);
			254: out = 24'(17844);
			255: out = 24'(27068);
			256: out = 24'(-122264);
			257: out = 24'(-5524);
			258: out = 24'(128120);
			259: out = 24'(40028);
			260: out = 24'(-81944);
			261: out = 24'(-127416);
			262: out = 24'(-37088);
			263: out = 24'(90376);
			264: out = 24'(129776);
			265: out = 24'(74140);
			266: out = 24'(-7268);
			267: out = 24'(-10100);
			268: out = 24'(52920);
			269: out = 24'(102640);
			270: out = 24'(82096);
			271: out = 24'(54092);
			272: out = 24'(18028);
			273: out = 24'(-44568);
			274: out = 24'(81100);
			275: out = 24'(77292);
			276: out = 24'(24340);
			277: out = 24'(-11372);
			278: out = 24'(42072);
			279: out = 24'(31732);
			280: out = 24'(-112256);
			281: out = 24'(14024);
			282: out = 24'(66952);
			283: out = 24'(54256);
			284: out = 24'(-61004);
			285: out = 24'(-111584);
			286: out = 24'(-86800);
			287: out = 24'(16520);
			288: out = 24'(-72724);
			289: out = 24'(-104300);
			290: out = 24'(-83640);
			291: out = 24'(-73656);
			292: out = 24'(37628);
			293: out = 24'(50312);
			294: out = 24'(-63700);
			295: out = 24'(-26984);
			296: out = 24'(-43384);
			297: out = 24'(-77892);
			298: out = 24'(-119388);
			299: out = 24'(-111492);
			300: out = 24'(-101576);
			301: out = 24'(-52744);
			302: out = 24'(2472);
			303: out = 24'(42472);
			304: out = 24'(20416);
			305: out = 24'(-33372);
			306: out = 24'(-107604);
			307: out = 24'(-85708);
			308: out = 24'(7940);
			309: out = 24'(-33180);
			310: out = 24'(-90064);
			311: out = 24'(-73900);
			312: out = 24'(114512);
			313: out = 24'(67564);
			314: out = 24'(-16256);
			315: out = 24'(-102700);
			316: out = 24'(-17256);
			317: out = 24'(67308);
			318: out = 24'(77820);
			319: out = 24'(-90244);
			320: out = 24'(-23736);
			321: out = 24'(65640);
			322: out = 24'(111044);
			323: out = 24'(-102280);
			324: out = 24'(-64724);
			325: out = 24'(81756);
			326: out = 24'(120192);
			327: out = 24'(109116);
			328: out = 24'(67968);
			329: out = 24'(17888);
			330: out = 24'(48428);
			331: out = 24'(-14712);
			332: out = 24'(-70488);
			333: out = 24'(-64420);
			334: out = 24'(62316);
			335: out = 24'(114340);
			336: out = 24'(66048);
			337: out = 24'(80168);
			338: out = 24'(14636);
			339: out = 24'(8236);
			340: out = 24'(56908);
			341: out = 24'(37204);
			342: out = 24'(-4812);
			343: out = 24'(-30332);
			344: out = 24'(-31712);
			345: out = 24'(68484);
			346: out = 24'(115200);
			347: out = 24'(61312);
			348: out = 24'(52252);
			349: out = 24'(71276);
			350: out = 24'(96656);
			351: out = 24'(-88188);
			352: out = 24'(-41000);
			353: out = 24'(35264);
			354: out = 24'(64520);
			355: out = 24'(19092);
			356: out = 24'(-33644);
			357: out = 24'(-57164);
			358: out = 24'(-4580);
			359: out = 24'(24780);
			360: out = 24'(61600);
			361: out = 24'(116336);
			362: out = 24'(-13232);
			363: out = 24'(-26188);
			364: out = 24'(29672);
			365: out = 24'(38752);
			366: out = 24'(71308);
			367: out = 24'(29496);
			368: out = 24'(-85208);
			369: out = 24'(12068);
			370: out = 24'(50700);
			371: out = 24'(50480);
			372: out = 24'(-2492);
			373: out = 24'(44212);
			374: out = 24'(64436);
			375: out = 24'(11968);
			376: out = 24'(-95108);
			377: out = 24'(-123636);
			378: out = 24'(-93828);
			379: out = 24'(46844);
			380: out = 24'(81328);
			381: out = 24'(73408);
			382: out = 24'(56740);
			383: out = 24'(-44736);
			384: out = 24'(-62868);
			385: out = 24'(-18268);
			386: out = 24'(11216);
			387: out = 24'(11808);
			388: out = 24'(-24792);
			389: out = 24'(-36788);
			390: out = 24'(-84292);
			391: out = 24'(-35712);
			392: out = 24'(21228);
			393: out = 24'(100256);
			394: out = 24'(-42548);
			395: out = 24'(-65552);
			396: out = 24'(47324);
			397: out = 24'(-63060);
			398: out = 24'(-110908);
			399: out = 24'(-110332);
			400: out = 24'(-59628);
			401: out = 24'(88012);
			402: out = 24'(97148);
			403: out = 24'(13500);
			404: out = 24'(-111120);
			405: out = 24'(-54012);
			406: out = 24'(58064);
			407: out = 24'(52004);
			408: out = 24'(-25252);
			409: out = 24'(-96408);
			410: out = 24'(-114392);
			411: out = 24'(56896);
			412: out = 24'(1056);
			413: out = 24'(-113376);
			414: out = 24'(-116324);
			415: out = 24'(30608);
			416: out = 24'(118076);
			417: out = 24'(47888);
			418: out = 24'(9092);
			419: out = 24'(-79360);
			420: out = 24'(-104132);
			421: out = 24'(-36604);
			422: out = 24'(-96560);
			423: out = 24'(-80088);
			424: out = 24'(35768);
			425: out = 24'(69872);
			426: out = 24'(79548);
			427: out = 24'(30776);
			428: out = 24'(-29352);
			429: out = 24'(-56628);
			430: out = 24'(-37412);
			431: out = 24'(4196);
			432: out = 24'(14836);
			433: out = 24'(48008);
			434: out = 24'(34556);
			435: out = 24'(-66484);
			436: out = 24'(-17648);
			437: out = 24'(63288);
			438: out = 24'(120648);
			439: out = 24'(-20776);
			440: out = 24'(-6512);
			441: out = 24'(12572);
			442: out = 24'(6656);
			443: out = 24'(-95080);
			444: out = 24'(-94876);
			445: out = 24'(-2664);
			446: out = 24'(20232);
			447: out = 24'(3896);
			448: out = 24'(10840);
			449: out = 24'(131064);
			450: out = 24'(-32116);
			451: out = 24'(-12204);
			452: out = 24'(71296);
			453: out = 24'(120308);
			454: out = 24'(-4332);
			455: out = 24'(-92864);
			456: out = 24'(-14104);
			457: out = 24'(34024);
			458: out = 24'(79072);
			459: out = 24'(69752);
			460: out = 24'(100364);
			461: out = 24'(68916);
			462: out = 24'(53780);
			463: out = 24'(1040);
			464: out = 24'(80096);
			465: out = 24'(18068);
			466: out = 24'(-46236);
			467: out = 24'(-3632);
			468: out = 24'(84876);
			469: out = 24'(114480);
			470: out = 24'(69084);
			471: out = 24'(9660);
			472: out = 24'(-8240);
			473: out = 24'(1328);
			474: out = 24'(-36600);
			475: out = 24'(-94328);
			476: out = 24'(-113124);
			477: out = 24'(-32516);
			478: out = 24'(29452);
			479: out = 24'(68400);
			480: out = 24'(34932);
			481: out = 24'(-41892);
			482: out = 24'(-64104);
			483: out = 24'(-11652);
			484: out = 24'(48020);
			485: out = 24'(14640);
			486: out = 24'(-12520);
			487: out = 24'(-14808);
			488: out = 24'(-51668);
			489: out = 24'(27804);
			490: out = 24'(28540);
			491: out = 24'(-4336);
			492: out = 24'(-101056);
			493: out = 24'(-13508);
			494: out = 24'(98560);
			495: out = 24'(120780);
			496: out = 24'(-31964);
			497: out = 24'(-91792);
			498: out = 24'(-4196);
			499: out = 24'(-65884);
			500: out = 24'(-83592);
			501: out = 24'(-103476);
			502: out = 24'(-58656);
			503: out = 24'(-2688);
			504: out = 24'(11376);
			505: out = 24'(-38936);
			506: out = 24'(-32684);
			507: out = 24'(8676);
			508: out = 24'(42640);
			509: out = 24'(-95820);
			510: out = 24'(33936);
			511: out = 24'(-6868);
			512: out = 24'(-118088);
			513: out = 24'(-85672);
			514: out = 24'(9544);
			515: out = 24'(99420);
			516: out = 24'(80980);
			517: out = 24'(45760);
			518: out = 24'(-63008);
			519: out = 24'(-115464);
			520: out = 24'(-106728);
			521: out = 24'(-10936);
			522: out = 24'(37444);
			523: out = 24'(-12488);
			524: out = 24'(12696);
			525: out = 24'(59720);
			526: out = 24'(100872);
			527: out = 24'(-48872);
			528: out = 24'(-31904);
			529: out = 24'(19304);
			530: out = 24'(101392);
			531: out = 24'(10688);
			532: out = 24'(-24920);
			533: out = 24'(-42460);
			534: out = 24'(80264);
			535: out = 24'(-36928);
			536: out = 24'(-53880);
			537: out = 24'(114432);
			538: out = 24'(82140);
			539: out = 24'(59856);
			540: out = 24'(1980);
			541: out = 24'(-28040);
			542: out = 24'(-33944);
			543: out = 24'(-15952);
			544: out = 24'(-24128);
			545: out = 24'(16208);
			546: out = 24'(24804);
			547: out = 24'(32964);
			548: out = 24'(16376);
			549: out = 24'(49632);
			550: out = 24'(68516);
			551: out = 24'(71820);
			552: out = 24'(-14976);
			553: out = 24'(-21820);
			554: out = 24'(16408);
			555: out = 24'(168);
			556: out = 24'(48308);
			557: out = 24'(50660);
			558: out = 24'(27004);
			559: out = 24'(-42056);
			560: out = 24'(-34588);
			561: out = 24'(25736);
			562: out = 24'(94244);
			563: out = 24'(52704);
			564: out = 24'(19560);
			565: out = 24'(32560);
			566: out = 24'(-4124);
			567: out = 24'(25328);
			568: out = 24'(54560);
			569: out = 24'(72024);
			570: out = 24'(6300);
			571: out = 24'(-3592);
			572: out = 24'(68316);
			573: out = 24'(-62540);
			574: out = 24'(-9624);
			575: out = 24'(48992);
			576: out = 24'(1324);
			577: out = 24'(33180);
			578: out = 24'(16572);
			579: out = 24'(-52176);
			580: out = 24'(-18240);
			581: out = 24'(-80092);
			582: out = 24'(-91256);
			583: out = 24'(29588);
			584: out = 24'(71996);
			585: out = 24'(60104);
			586: out = 24'(21696);
			587: out = 24'(-72216);
			588: out = 24'(-30684);
			589: out = 24'(22076);
			590: out = 24'(-29320);
			591: out = 24'(-15420);
			592: out = 24'(72);
			593: out = 24'(10820);
			594: out = 24'(-2600);
			595: out = 24'(-72340);
			596: out = 24'(-87716);
			597: out = 24'(46648);
			598: out = 24'(72068);
			599: out = 24'(30928);
			600: out = 24'(-71020);
			601: out = 24'(-48908);
			602: out = 24'(-83004);
			603: out = 24'(-101572);
			604: out = 24'(-93372);
			605: out = 24'(-5496);
			606: out = 24'(75324);
			607: out = 24'(87624);
			608: out = 24'(93812);
			609: out = 24'(-43156);
			610: out = 24'(-108904);
			611: out = 24'(-9808);
			612: out = 24'(78148);
			613: out = 24'(49312);
			614: out = 24'(-44176);
			615: out = 24'(1116);
			616: out = 24'(46312);
			617: out = 24'(74472);
			618: out = 24'(-7692);
			619: out = 24'(54516);
			620: out = 24'(2444);
			621: out = 24'(-66324);
			622: out = 24'(-10488);
			623: out = 24'(7192);
			624: out = 24'(34224);
			625: out = 24'(42204);
			626: out = 24'(44176);
			627: out = 24'(10820);
			628: out = 24'(6872);
			629: out = 24'(66624);
			630: out = 24'(74216);
			631: out = 24'(8528);
			632: out = 24'(-91044);
			633: out = 24'(-103448);
			634: out = 24'(488);
			635: out = 24'(84728);
			636: out = 24'(32440);
			637: out = 24'(-58664);
			638: out = 24'(-87868);
			639: out = 24'(10944);
			640: out = 24'(-3928);
			641: out = 24'(-32768);
			642: out = 24'(-76872);
			643: out = 24'(-96816);
			644: out = 24'(-32744);
			645: out = 24'(24544);
			646: out = 24'(43652);
			647: out = 24'(-41512);
			648: out = 24'(5876);
			649: out = 24'(56436);
			650: out = 24'(-101812);
			651: out = 24'(-104876);
			652: out = 24'(-45280);
			653: out = 24'(63564);
			654: out = 24'(26712);
			655: out = 24'(-31772);
			656: out = 24'(-94324);
			657: out = 24'(-23752);
			658: out = 24'(3116);
			659: out = 24'(39236);
			660: out = 24'(38768);
			661: out = 24'(-51656);
			662: out = 24'(-86092);
			663: out = 24'(-60760);
			664: out = 24'(-43048);
			665: out = 24'(29012);
			666: out = 24'(60772);
			667: out = 24'(62196);
			668: out = 24'(55740);
			669: out = 24'(23060);
			670: out = 24'(-32156);
			671: out = 24'(-101392);
			672: out = 24'(-73556);
			673: out = 24'(-5832);
			674: out = 24'(34604);
			675: out = 24'(30044);
			676: out = 24'(5412);
			677: out = 24'(-17724);
			678: out = 24'(-94032);
			679: out = 24'(39148);
			680: out = 24'(55044);
			681: out = 24'(-42584);
			682: out = 24'(-69056);
			683: out = 24'(-70500);
			684: out = 24'(-9284);
			685: out = 24'(7416);
			686: out = 24'(59288);
			687: out = 24'(17764);
			688: out = 24'(-37284);
			689: out = 24'(33284);
			690: out = 24'(53896);
			691: out = 24'(39876);
			692: out = 24'(28472);
			693: out = 24'(-82092);
			694: out = 24'(-82300);
			695: out = 24'(25104);
			696: out = 24'(76660);
			697: out = 24'(77264);
			698: out = 24'(30020);
			699: out = 24'(-2184);
			700: out = 24'(-78660);
			701: out = 24'(-80480);
			702: out = 24'(-17016);
			703: out = 24'(39284);
			704: out = 24'(75640);
			705: out = 24'(48280);
			706: out = 24'(-38772);
			707: out = 24'(-98536);
			708: out = 24'(-71388);
			709: out = 24'(45316);
			710: out = 24'(24456);
			711: out = 24'(94492);
			712: out = 24'(54900);
			713: out = 24'(-54132);
			714: out = 24'(-95676);
			715: out = 24'(-38204);
			716: out = 24'(50796);
			717: out = 24'(74440);
			718: out = 24'(51504);
			719: out = 24'(34744);
			720: out = 24'(19776);
			721: out = 24'(96168);
			722: out = 24'(28916);
			723: out = 24'(-76436);
			724: out = 24'(-113740);
			725: out = 24'(-4464);
			726: out = 24'(87676);
			727: out = 24'(63524);
			728: out = 24'(-37864);
			729: out = 24'(-67040);
			730: out = 24'(112);
			731: out = 24'(50876);
			732: out = 24'(14256);
			733: out = 24'(-54480);
			734: out = 24'(-65180);
			735: out = 24'(-24740);
			736: out = 24'(57652);
			737: out = 24'(64404);
			738: out = 24'(-86076);
			739: out = 24'(-118308);
			740: out = 24'(-89456);
			741: out = 24'(4612);
			742: out = 24'(55936);
			743: out = 24'(93052);
			744: out = 24'(57036);
			745: out = 24'(-73128);
			746: out = 24'(-108428);
			747: out = 24'(-47820);
			748: out = 24'(49852);
			749: out = 24'(24072);
			750: out = 24'(-22260);
			751: out = 24'(-31100);
			752: out = 24'(80592);
			753: out = 24'(34472);
			754: out = 24'(-32416);
			755: out = 24'(-85164);
			756: out = 24'(-54136);
			757: out = 24'(34196);
			758: out = 24'(69736);
			759: out = 24'(17736);
			760: out = 24'(-53480);
			761: out = 24'(-48572);
			762: out = 24'(41996);
			763: out = 24'(71612);
			764: out = 24'(62564);
			765: out = 24'(16396);
			766: out = 24'(-63792);
			767: out = 24'(24772);
			768: out = 24'(67400);
			769: out = 24'(49868);
			770: out = 24'(-54692);
			771: out = 24'(1184);
			772: out = 24'(72988);
			773: out = 24'(10128);
			774: out = 24'(2928);
			775: out = 24'(-47028);
			776: out = 24'(-63988);
			777: out = 24'(-816);
			778: out = 24'(42388);
			779: out = 24'(31416);
			780: out = 24'(-63440);
			781: out = 24'(-16548);
			782: out = 24'(-45540);
			783: out = 24'(-115020);
			784: out = 24'(-36592);
			785: out = 24'(9996);
			786: out = 24'(54776);
			787: out = 24'(76244);
			788: out = 24'(59916);
			789: out = 24'(39972);
			790: out = 24'(21736);
			791: out = 24'(-28224);
			792: out = 24'(-31692);
			793: out = 24'(-31504);
			794: out = 24'(-63932);
			795: out = 24'(52308);
			796: out = 24'(72360);
			797: out = 24'(31984);
			798: out = 24'(-13340);
			799: out = 24'(-7940);
			800: out = 24'(42276);
			801: out = 24'(91484);
			802: out = 24'(23220);
			803: out = 24'(-21368);
			804: out = 24'(-23796);
			805: out = 24'(47248);
			806: out = 24'(50168);
			807: out = 24'(18492);
			808: out = 24'(-43796);
			809: out = 24'(792);
			810: out = 24'(21992);
			811: out = 24'(39228);
			812: out = 24'(54436);
			813: out = 24'(59560);
			814: out = 24'(45024);
			815: out = 24'(29680);
			816: out = 24'(5600);
			817: out = 24'(19488);
			818: out = 24'(34032);
			819: out = 24'(47676);
			820: out = 24'(-6172);
			821: out = 24'(-2248);
			822: out = 24'(71812);
			823: out = 24'(51464);
			824: out = 24'(664);
			825: out = 24'(-69880);
			826: out = 24'(4188);
			827: out = 24'(-11020);
			828: out = 24'(37432);
			829: out = 24'(77708);
			830: out = 24'(28200);
			831: out = 24'(-55204);
			832: out = 24'(-104424);
			833: out = 24'(-35184);
			834: out = 24'(40996);
			835: out = 24'(74448);
			836: out = 24'(56732);
			837: out = 24'(-52696);
			838: out = 24'(-52132);
			839: out = 24'(12568);
			840: out = 24'(932);
			841: out = 24'(56328);
			842: out = 24'(35908);
			843: out = 24'(-7944);
			844: out = 24'(5128);
			845: out = 24'(33632);
			846: out = 24'(25696);
			847: out = 24'(-103784);
			848: out = 24'(-82656);
			849: out = 24'(-36556);
			850: out = 24'(23864);
			851: out = 24'(-7072);
			852: out = 24'(36440);
			853: out = 24'(55472);
			854: out = 24'(13356);
			855: out = 24'(-46236);
			856: out = 24'(-64372);
			857: out = 24'(-4172);
			858: out = 24'(-76160);
			859: out = 24'(12384);
			860: out = 24'(71392);
			861: out = 24'(-6572);
			862: out = 24'(9384);
			863: out = 24'(-24368);
			864: out = 24'(-58336);
			865: out = 24'(-60644);
			866: out = 24'(-11052);
			867: out = 24'(31220);
			868: out = 24'(14588);
			869: out = 24'(37288);
			870: out = 24'(38548);
			871: out = 24'(32784);
			872: out = 24'(-33972);
			873: out = 24'(-42588);
			874: out = 24'(-33960);
			875: out = 24'(-10684);
			876: out = 24'(-29844);
			877: out = 24'(-20000);
			878: out = 24'(8980);
			879: out = 24'(6864);
			880: out = 24'(28408);
			881: out = 24'(17212);
			882: out = 24'(-72616);
			883: out = 24'(-29252);
			884: out = 24'(-11324);
			885: out = 24'(6220);
			886: out = 24'(-62216);
			887: out = 24'(8092);
			888: out = 24'(48220);
			889: out = 24'(25984);
			890: out = 24'(-71948);
			891: out = 24'(-84064);
			892: out = 24'(-3088);
			893: out = 24'(32840);
			894: out = 24'(49520);
			895: out = 24'(32184);
			896: out = 24'(21244);
			897: out = 24'(-9072);
			898: out = 24'(-15604);
			899: out = 24'(-6932);
			900: out = 24'(-13480);
			901: out = 24'(9040);
			902: out = 24'(-11544);
			903: out = 24'(-79688);
			904: out = 24'(-2152);
			905: out = 24'(60824);
			906: out = 24'(66372);
			907: out = 24'(8624);
			908: out = 24'(-76252);
			909: out = 24'(-89788);
			910: out = 24'(13308);
			911: out = 24'(61384);
			912: out = 24'(47504);
			913: out = 24'(-23164);
			914: out = 24'(-74696);
			915: out = 24'(-88512);
			916: out = 24'(-59428);
			917: out = 24'(-49112);
			918: out = 24'(31148);
			919: out = 24'(22120);
			920: out = 24'(-8344);
			921: out = 24'(-33796);
			922: out = 24'(-46472);
			923: out = 24'(-49964);
			924: out = 24'(-28600);
			925: out = 24'(-48236);
			926: out = 24'(-3308);
			927: out = 24'(43760);
			928: out = 24'(62504);
			929: out = 24'(-10892);
			930: out = 24'(-77836);
			931: out = 24'(-96208);
			932: out = 24'(-8644);
			933: out = 24'(34488);
			934: out = 24'(12684);
			935: out = 24'(-91508);
			936: out = 24'(-54676);
			937: out = 24'(-9412);
			938: out = 24'(6108);
			939: out = 24'(75632);
			940: out = 24'(58152);
			941: out = 24'(36404);
			942: out = 24'(59652);
			943: out = 24'(-17632);
			944: out = 24'(-78512);
			945: out = 24'(-104912);
			946: out = 24'(21496);
			947: out = 24'(57848);
			948: out = 24'(47632);
			949: out = 24'(8672);
			950: out = 24'(29520);
			951: out = 24'(18780);
			952: out = 24'(-16348);
			953: out = 24'(-32640);
			954: out = 24'(-18364);
			955: out = 24'(1080);
			956: out = 24'(-33712);
			957: out = 24'(31408);
			958: out = 24'(44764);
			959: out = 24'(26496);
			960: out = 24'(-312);
			961: out = 24'(-8896);
			962: out = 24'(6252);
			963: out = 24'(42028);
			964: out = 24'(1164);
			965: out = 24'(34720);
			966: out = 24'(104360);
			967: out = 24'(-65504);
			968: out = 24'(15424);
			969: out = 24'(49876);
			970: out = 24'(3408);
			971: out = 24'(-17628);
			972: out = 24'(13948);
			973: out = 24'(58968);
			974: out = 24'(55192);
			975: out = 24'(2880);
			976: out = 24'(-23236);
			977: out = 24'(13520);
			978: out = 24'(40136);
			979: out = 24'(20692);
			980: out = 24'(-29848);
			981: out = 24'(-87924);
			982: out = 24'(-25124);
			983: out = 24'(45176);
			984: out = 24'(42372);
			985: out = 24'(12280);
			986: out = 24'(-11852);
			987: out = 24'(-2396);
			988: out = 24'(41388);
			989: out = 24'(-9116);
			990: out = 24'(-17056);
			991: out = 24'(72304);
			992: out = 24'(6544);
			993: out = 24'(-20960);
			994: out = 24'(-49116);
			995: out = 24'(115176);
			996: out = 24'(-49700);
			997: out = 24'(-91812);
			998: out = 24'(32320);
			999: out = 24'(71328);
			1000: out = 24'(70844);
			1001: out = 24'(21948);
			1002: out = 24'(-68588);
			1003: out = 24'(-42116);
			1004: out = 24'(-2364);
			1005: out = 24'(-4108);
			1006: out = 24'(-43652);
			1007: out = 24'(-67380);
			1008: out = 24'(-44504);
			1009: out = 24'(19940);
			1010: out = 24'(24700);
			1011: out = 24'(60);
			1012: out = 24'(-42796);
			1013: out = 24'(-44844);
			1014: out = 24'(-46484);
			1015: out = 24'(-24972);
			1016: out = 24'(-1480);
			1017: out = 24'(40252);
			1018: out = 24'(40516);
			1019: out = 24'(26524);
			1020: out = 24'(-39036);
			1021: out = 24'(7880);
			1022: out = 24'(34844);
			1023: out = 24'(-110028);
			1024: out = 24'(-69104);
			1025: out = 24'(-2436);
			1026: out = 24'(70204);
			1027: out = 24'(58300);
			1028: out = 24'(31340);
			1029: out = 24'(-21240);
			1030: out = 24'(-39132);
			1031: out = 24'(-16648);
			1032: out = 24'(34004);
			1033: out = 24'(40352);
			1034: out = 24'(61576);
			1035: out = 24'(1788);
			1036: out = 24'(-31272);
			1037: out = 24'(-51860);
			1038: out = 24'(51964);
			1039: out = 24'(46584);
			1040: out = 24'(-19076);
			1041: out = 24'(-68864);
			1042: out = 24'(-11040);
			1043: out = 24'(56064);
			1044: out = 24'(43016);
			1045: out = 24'(-29764);
			1046: out = 24'(-40220);
			1047: out = 24'(34616);
			1048: out = 24'(-52124);
			1049: out = 24'(-6308);
			1050: out = 24'(16480);
			1051: out = 24'(-356);
			1052: out = 24'(-13108);
			1053: out = 24'(-40500);
			1054: out = 24'(-62216);
			1055: out = 24'(-10412);
			1056: out = 24'(18404);
			1057: out = 24'(30108);
			1058: out = 24'(20004);
			1059: out = 24'(48);
			1060: out = 24'(892);
			1061: out = 24'(21320);
			1062: out = 24'(17704);
			1063: out = 24'(24396);
			1064: out = 24'(21424);
			1065: out = 24'(19772);
			1066: out = 24'(14672);
			1067: out = 24'(19476);
			1068: out = 24'(23788);
			1069: out = 24'(-13916);
			1070: out = 24'(31960);
			1071: out = 24'(63360);
			1072: out = 24'(36020);
			1073: out = 24'(9400);
			1074: out = 24'(-24172);
			1075: out = 24'(-21296);
			1076: out = 24'(-67792);
			1077: out = 24'(28760);
			1078: out = 24'(51788);
			1079: out = 24'(-21516);
			1080: out = 24'(164);
			1081: out = 24'(40156);
			1082: out = 24'(71992);
			1083: out = 24'(-32144);
			1084: out = 24'(-26340);
			1085: out = 24'(-18688);
			1086: out = 24'(8632);
			1087: out = 24'(-42448);
			1088: out = 24'(-38084);
			1089: out = 24'(-6788);
			1090: out = 24'(40352);
			1091: out = 24'(15792);
			1092: out = 24'(14632);
			1093: out = 24'(70496);
			1094: out = 24'(-46552);
			1095: out = 24'(-2624);
			1096: out = 24'(66464);
			1097: out = 24'(45632);
			1098: out = 24'(18628);
			1099: out = 24'(4048);
			1100: out = 24'(49708);
			1101: out = 24'(-62888);
			1102: out = 24'(-39828);
			1103: out = 24'(21236);
			1104: out = 24'(87540);
			1105: out = 24'(2172);
			1106: out = 24'(-56496);
			1107: out = 24'(-44612);
			1108: out = 24'(31248);
			1109: out = 24'(72324);
			1110: out = 24'(57028);
			1111: out = 24'(20680);
			1112: out = 24'(-37400);
			1113: out = 24'(-65748);
			1114: out = 24'(-55656);
			1115: out = 24'(4780);
			1116: out = 24'(35792);
			1117: out = 24'(34020);
			1118: out = 24'(-12416);
			1119: out = 24'(-16856);
			1120: out = 24'(-37276);
			1121: out = 24'(-50808);
			1122: out = 24'(6964);
			1123: out = 24'(35900);
			1124: out = 24'(33900);
			1125: out = 24'(26140);
			1126: out = 24'(-49700);
			1127: out = 24'(-32864);
			1128: out = 24'(61828);
			1129: out = 24'(-65640);
			1130: out = 24'(-29296);
			1131: out = 24'(-8464);
			1132: out = 24'(-49152);
			1133: out = 24'(-20112);
			1134: out = 24'(16752);
			1135: out = 24'(36008);
			1136: out = 24'(16308);
			1137: out = 24'(-45932);
			1138: out = 24'(-86416);
			1139: out = 24'(-3732);
			1140: out = 24'(-51220);
			1141: out = 24'(-2496);
			1142: out = 24'(64676);
			1143: out = 24'(-32196);
			1144: out = 24'(-49888);
			1145: out = 24'(-58552);
			1146: out = 24'(-28224);
			1147: out = 24'(-13752);
			1148: out = 24'(12540);
			1149: out = 24'(13528);
			1150: out = 24'(55244);
			1151: out = 24'(-4508);
			1152: out = 24'(-16556);
			1153: out = 24'(33072);
			1154: out = 24'(58232);
			1155: out = 24'(-13120);
			1156: out = 24'(-122384);
			1157: out = 24'(-53928);
			1158: out = 24'(-17224);
			1159: out = 24'(11272);
			1160: out = 24'(-17800);
			1161: out = 24'(49584);
			1162: out = 24'(68588);
			1163: out = 24'(61436);
			1164: out = 24'(-95128);
			1165: out = 24'(-40280);
			1166: out = 24'(32996);
			1167: out = 24'(48644);
			1168: out = 24'(29188);
			1169: out = 24'(-10260);
			1170: out = 24'(-31732);
			1171: out = 24'(-8640);
			1172: out = 24'(22112);
			1173: out = 24'(29736);
			1174: out = 24'(-3060);
			1175: out = 24'(43996);
			1176: out = 24'(31244);
			1177: out = 24'(15864);
			1178: out = 24'(31796);
			1179: out = 24'(37700);
			1180: out = 24'(17412);
			1181: out = 24'(-41144);
			1182: out = 24'(21028);
			1183: out = 24'(-6000);
			1184: out = 24'(-54412);
			1185: out = 24'(-33896);
			1186: out = 24'(-34424);
			1187: out = 24'(5268);
			1188: out = 24'(36476);
			1189: out = 24'(25044);
			1190: out = 24'(-33008);
			1191: out = 24'(-80988);
			1192: out = 24'(-51008);
			1193: out = 24'(-10496);
			1194: out = 24'(36796);
			1195: out = 24'(68420);
			1196: out = 24'(-15304);
			1197: out = 24'(-11588);
			1198: out = 24'(16960);
			1199: out = 24'(58124);
			1200: out = 24'(-38556);
			1201: out = 24'(-61536);
			1202: out = 24'(28472);
			1203: out = 24'(-31256);
			1204: out = 24'(25300);
			1205: out = 24'(54944);
			1206: out = 24'(23192);
			1207: out = 24'(7172);
			1208: out = 24'(-26108);
			1209: out = 24'(-57140);
			1210: out = 24'(-24996);
			1211: out = 24'(8080);
			1212: out = 24'(30416);
			1213: out = 24'(13044);
			1214: out = 24'(17500);
			1215: out = 24'(-1488);
			1216: out = 24'(-20128);
			1217: out = 24'(-9452);
			1218: out = 24'(1032);
			1219: out = 24'(724);
			1220: out = 24'(-14748);
			1221: out = 24'(-1244);
			1222: out = 24'(27536);
			1223: out = 24'(55944);
			1224: out = 24'(27996);
			1225: out = 24'(22496);
			1226: out = 24'(-1420);
			1227: out = 24'(-52444);
			1228: out = 24'(9908);
			1229: out = 24'(47880);
			1230: out = 24'(40388);
			1231: out = 24'(-14108);
			1232: out = 24'(-11084);
			1233: out = 24'(31012);
			1234: out = 24'(45676);
			1235: out = 24'(42424);
			1236: out = 24'(-35384);
			1237: out = 24'(-106876);
			1238: out = 24'(-53736);
			1239: out = 24'(28592);
			1240: out = 24'(66144);
			1241: out = 24'(52940);
			1242: out = 24'(-38472);
			1243: out = 24'(-46472);
			1244: out = 24'(14644);
			1245: out = 24'(48080);
			1246: out = 24'(21704);
			1247: out = 24'(-10172);
			1248: out = 24'(10868);
			1249: out = 24'(41244);
			1250: out = 24'(32380);
			1251: out = 24'(-15656);
			1252: out = 24'(62724);
			1253: out = 24'(-41380);
			1254: out = 24'(-71024);
			1255: out = 24'(13044);
			1256: out = 24'(-7700);
			1257: out = 24'(8032);
			1258: out = 24'(17600);
			1259: out = 24'(43856);
			1260: out = 24'(-15312);
			1261: out = 24'(-47568);
			1262: out = 24'(-12124);
			1263: out = 24'(-37464);
			1264: out = 24'(-24368);
			1265: out = 24'(-9244);
			1266: out = 24'(62020);
			1267: out = 24'(-17432);
			1268: out = 24'(-59676);
			1269: out = 24'(-42992);
			1270: out = 24'(-39352);
			1271: out = 24'(-32760);
			1272: out = 24'(-14080);
			1273: out = 24'(37208);
			1274: out = 24'(49132);
			1275: out = 24'(9716);
			1276: out = 24'(-73272);
			1277: out = 24'(-77748);
			1278: out = 24'(-17880);
			1279: out = 24'(45764);
			1280: out = 24'(-74808);
			1281: out = 24'(-7280);
			1282: out = 24'(25368);
			1283: out = 24'(62656);
			1284: out = 24'(-66784);
			1285: out = 24'(-13516);
			1286: out = 24'(59312);
			1287: out = 24'(49264);
			1288: out = 24'(-19560);
			1289: out = 24'(-66724);
			1290: out = 24'(-39672);
			1291: out = 24'(19332);
			1292: out = 24'(32804);
			1293: out = 24'(10368);
			1294: out = 24'(29864);
			1295: out = 24'(-9440);
			1296: out = 24'(8132);
			1297: out = 24'(51916);
			1298: out = 24'(23444);
			1299: out = 24'(34780);
			1300: out = 24'(35512);
			1301: out = 24'(9312);
			1302: out = 24'(16244);
			1303: out = 24'(25900);
			1304: out = 24'(31140);
			1305: out = 24'(15660);
			1306: out = 24'(-14688);
			1307: out = 24'(-30708);
			1308: out = 24'(9752);
			1309: out = 24'(30828);
			1310: out = 24'(52108);
			1311: out = 24'(44152);
			1312: out = 24'(33816);
			1313: out = 24'(-2820);
			1314: out = 24'(-29000);
			1315: out = 24'(-58512);
			1316: out = 24'(19148);
			1317: out = 24'(48536);
			1318: out = 24'(29488);
			1319: out = 24'(-42712);
			1320: out = 24'(-57004);
			1321: out = 24'(-28792);
			1322: out = 24'(28188);
			1323: out = 24'(-4740);
			1324: out = 24'(3516);
			1325: out = 24'(35392);
			1326: out = 24'(14024);
			1327: out = 24'(14284);
			1328: out = 24'(5424);
			1329: out = 24'(3100);
			1330: out = 24'(-3192);
			1331: out = 24'(9588);
			1332: out = 24'(24296);
			1333: out = 24'(5704);
			1334: out = 24'(-15144);
			1335: out = 24'(-32320);
			1336: out = 24'(6120);
			1337: out = 24'(-50032);
			1338: out = 24'(-13360);
			1339: out = 24'(41836);
			1340: out = 24'(35268);
			1341: out = 24'(-5296);
			1342: out = 24'(-39836);
			1343: out = 24'(-36680);
			1344: out = 24'(-5440);
			1345: out = 24'(-3092);
			1346: out = 24'(-24932);
			1347: out = 24'(-53396);
			1348: out = 24'(-9084);
			1349: out = 24'(36072);
			1350: out = 24'(36804);
			1351: out = 24'(-16936);
			1352: out = 24'(-33152);
			1353: out = 24'(-4952);
			1354: out = 24'(-16180);
			1355: out = 24'(19240);
			1356: out = 24'(22008);
			1357: out = 24'(11172);
			1358: out = 24'(-2284);
			1359: out = 24'(2392);
			1360: out = 24'(7428);
			1361: out = 24'(448);
			1362: out = 24'(6040);
			1363: out = 24'(15504);
			1364: out = 24'(18848);
			1365: out = 24'(36840);
			1366: out = 24'(28304);
			1367: out = 24'(3440);
			1368: out = 24'(-86724);
			1369: out = 24'(-37664);
			1370: out = 24'(17420);
			1371: out = 24'(41444);
			1372: out = 24'(-1280);
			1373: out = 24'(-3220);
			1374: out = 24'(10556);
			1375: out = 24'(11516);
			1376: out = 24'(22064);
			1377: out = 24'(31436);
			1378: out = 24'(33252);
			1379: out = 24'(21600);
			1380: out = 24'(-4060);
			1381: out = 24'(-14252);
			1382: out = 24'(6968);
			1383: out = 24'(4556);
			1384: out = 24'(-7104);
			1385: out = 24'(-10368);
			1386: out = 24'(-97060);
			1387: out = 24'(-43040);
			1388: out = 24'(40060);
			1389: out = 24'(48264);
			1390: out = 24'(1952);
			1391: out = 24'(-32268);
			1392: out = 24'(-12248);
			1393: out = 24'(-27008);
			1394: out = 24'(-18252);
			1395: out = 24'(-12920);
			1396: out = 24'(56824);
			1397: out = 24'(-52052);
			1398: out = 24'(-55704);
			1399: out = 24'(27872);
			1400: out = 24'(-11996);
			1401: out = 24'(39864);
			1402: out = 24'(32708);
			1403: out = 24'(-88420);
			1404: out = 24'(-36916);
			1405: out = 24'(-11144);
			1406: out = 24'(-11908);
			1407: out = 24'(18920);
			1408: out = 24'(15596);
			1409: out = 24'(4340);
			1410: out = 24'(-56032);
			1411: out = 24'(42400);
			1412: out = 24'(41328);
			1413: out = 24'(-14088);
			1414: out = 24'(-76780);
			1415: out = 24'(-65144);
			1416: out = 24'(-1272);
			1417: out = 24'(53816);
			1418: out = 24'(16692);
			1419: out = 24'(-13012);
			1420: out = 24'(-23392);
			1421: out = 24'(-1300);
			1422: out = 24'(-11964);
			1423: out = 24'(-23128);
			1424: out = 24'(-18392);
			1425: out = 24'(7596);
			1426: out = 24'(10208);
			1427: out = 24'(-5592);
			1428: out = 24'(10568);
			1429: out = 24'(1436);
			1430: out = 24'(1940);
			1431: out = 24'(3108);
			1432: out = 24'(15480);
			1433: out = 24'(11960);
			1434: out = 24'(9472);
			1435: out = 24'(46300);
			1436: out = 24'(12180);
			1437: out = 24'(-5244);
			1438: out = 24'(19188);
			1439: out = 24'(-20744);
			1440: out = 24'(552);
			1441: out = 24'(28624);
			1442: out = 24'(8984);
			1443: out = 24'(11604);
			1444: out = 24'(-836);
			1445: out = 24'(-19104);
			1446: out = 24'(7124);
			1447: out = 24'(9564);
			1448: out = 24'(6956);
			1449: out = 24'(43612);
			1450: out = 24'(3704);
			1451: out = 24'(-24380);
			1452: out = 24'(-36072);
			1453: out = 24'(12468);
			1454: out = 24'(5668);
			1455: out = 24'(-16548);
			1456: out = 24'(29876);
			1457: out = 24'(-16052);
			1458: out = 24'(-31072);
			1459: out = 24'(-21828);
			1460: out = 24'(28288);
			1461: out = 24'(29132);
			1462: out = 24'(15328);
			1463: out = 24'(13912);
			1464: out = 24'(608);
			1465: out = 24'(-18364);
			1466: out = 24'(-36308);
			1467: out = 24'(-7728);
			1468: out = 24'(12348);
			1469: out = 24'(16796);
			1470: out = 24'(4616);
			1471: out = 24'(-9384);
			1472: out = 24'(-3480);
			1473: out = 24'(14716);
			1474: out = 24'(2048);
			1475: out = 24'(-3996);
			1476: out = 24'(-2140);
			1477: out = 24'(10032);
			1478: out = 24'(17172);
			1479: out = 24'(21352);
			1480: out = 24'(30892);
			1481: out = 24'(-17784);
			1482: out = 24'(20864);
			1483: out = 24'(37920);
			1484: out = 24'(-28060);
			1485: out = 24'(-8940);
			1486: out = 24'(2632);
			1487: out = 24'(9612);
			1488: out = 24'(39816);
			1489: out = 24'(-11732);
			1490: out = 24'(-52920);
			1491: out = 24'(-3712);
			1492: out = 24'(14076);
			1493: out = 24'(30844);
			1494: out = 24'(9112);
			1495: out = 24'(-18748);
			1496: out = 24'(-28832);
			1497: out = 24'(-8128);
			1498: out = 24'(-19232);
			1499: out = 24'(53468);
			1500: out = 24'(43280);
			1501: out = 24'(8696);
			1502: out = 24'(-81840);
			1503: out = 24'(-54540);
			1504: out = 24'(-2624);
			1505: out = 24'(38736);
			1506: out = 24'(-24784);
			1507: out = 24'(-12720);
			1508: out = 24'(35968);
			1509: out = 24'(19000);
			1510: out = 24'(-14996);
			1511: out = 24'(-47840);
			1512: out = 24'(-35364);
			1513: out = 24'(16128);
			1514: out = 24'(42196);
			1515: out = 24'(30692);
			1516: out = 24'(-30412);
			1517: out = 24'(-864);
			1518: out = 24'(11808);
			1519: out = 24'(-50812);
			1520: out = 24'(-26140);
			1521: out = 24'(-8960);
			1522: out = 24'(25820);
			1523: out = 24'(37160);
			1524: out = 24'(28296);
			1525: out = 24'(-6540);
			1526: out = 24'(-30040);
			1527: out = 24'(-32320);
			1528: out = 24'(1704);
			1529: out = 24'(24660);
			1530: out = 24'(1536);
			1531: out = 24'(-13928);
			1532: out = 24'(-6392);
			1533: out = 24'(33736);
			1534: out = 24'(23812);
			1535: out = 24'(7280);
			1536: out = 24'(-31204);
			1537: out = 24'(-42588);
			1538: out = 24'(-57656);
			1539: out = 24'(-22312);
			1540: out = 24'(21512);
			1541: out = 24'(35392);
			1542: out = 24'(-8204);
			1543: out = 24'(-44604);
			1544: out = 24'(-1704);
			1545: out = 24'(30464);
			1546: out = 24'(27120);
			1547: out = 24'(-19204);
			1548: out = 24'(-15680);
			1549: out = 24'(-1708);
			1550: out = 24'(19596);
			1551: out = 24'(6032);
			1552: out = 24'(-5860);
			1553: out = 24'(-9788);
			1554: out = 24'(13668);
			1555: out = 24'(-30420);
			1556: out = 24'(-32828);
			1557: out = 24'(-25256);
			1558: out = 24'(-5736);
			1559: out = 24'(17520);
			1560: out = 24'(23896);
			1561: out = 24'(-1412);
			1562: out = 24'(26888);
			1563: out = 24'(9052);
			1564: out = 24'(6560);
			1565: out = 24'(12928);
			1566: out = 24'(35348);
			1567: out = 24'(16860);
			1568: out = 24'(-15336);
			1569: out = 24'(5708);
			1570: out = 24'(20944);
			1571: out = 24'(21988);
			1572: out = 24'(35004);
			1573: out = 24'(-24948);
			1574: out = 24'(-7192);
			1575: out = 24'(49188);
			1576: out = 24'(-1964);
			1577: out = 24'(-39424);
			1578: out = 24'(-52852);
			1579: out = 24'(6320);
			1580: out = 24'(33940);
			1581: out = 24'(27388);
			1582: out = 24'(-13652);
			1583: out = 24'(-81944);
			1584: out = 24'(-36940);
			1585: out = 24'(42520);
			1586: out = 24'(25332);
			1587: out = 24'(41388);
			1588: out = 24'(-5600);
			1589: out = 24'(-36044);
			1590: out = 24'(-30992);
			1591: out = 24'(24040);
			1592: out = 24'(49532);
			1593: out = 24'(32904);
			1594: out = 24'(-22616);
			1595: out = 24'(-56804);
			1596: out = 24'(-49488);
			1597: out = 24'(24052);
			1598: out = 24'(40480);
			1599: out = 24'(36888);
			1600: out = 24'(19584);
			1601: out = 24'(13048);
			1602: out = 24'(-25432);
			1603: out = 24'(-63796);
			1604: out = 24'(-11644);
			1605: out = 24'(22668);
			1606: out = 24'(39820);
			1607: out = 24'(17096);
			1608: out = 24'(-13212);
			1609: out = 24'(-49464);
			1610: out = 24'(-53868);
			1611: out = 24'(20052);
			1612: out = 24'(6220);
			1613: out = 24'(-18168);
			1614: out = 24'(-5604);
			1615: out = 24'(-53856);
			1616: out = 24'(-35660);
			1617: out = 24'(2252);
			1618: out = 24'(22460);
			1619: out = 24'(-1880);
			1620: out = 24'(-21424);
			1621: out = 24'(-7288);
			1622: out = 24'(7236);
			1623: out = 24'(20604);
			1624: out = 24'(13056);
			1625: out = 24'(288);
			1626: out = 24'(-19288);
			1627: out = 24'(-1260);
			1628: out = 24'(50124);
			1629: out = 24'(-37144);
			1630: out = 24'(-60376);
			1631: out = 24'(-41672);
			1632: out = 24'(22472);
			1633: out = 24'(13732);
			1634: out = 24'(-6344);
			1635: out = 24'(-22568);
			1636: out = 24'(-12948);
			1637: out = 24'(-1896);
			1638: out = 24'(4144);
			1639: out = 24'(-7780);
			1640: out = 24'(8824);
			1641: out = 24'(19652);
			1642: out = 24'(20776);
			1643: out = 24'(4140);
			1644: out = 24'(-5984);
			1645: out = 24'(-12960);
			1646: out = 24'(-18440);
			1647: out = 24'(-7100);
			1648: out = 24'(17300);
			1649: out = 24'(36480);
			1650: out = 24'(-8608);
			1651: out = 24'(-32580);
			1652: out = 24'(-30644);
			1653: out = 24'(16288);
			1654: out = 24'(13788);
			1655: out = 24'(13280);
			1656: out = 24'(19396);
			1657: out = 24'(20448);
			1658: out = 24'(32160);
			1659: out = 24'(16832);
			1660: out = 24'(-58424);
			1661: out = 24'(-36172);
			1662: out = 24'(-564);
			1663: out = 24'(27696);
			1664: out = 24'(23432);
			1665: out = 24'(22188);
			1666: out = 24'(20288);
			1667: out = 24'(2364);
			1668: out = 24'(14620);
			1669: out = 24'(19248);
			1670: out = 24'(30236);
			1671: out = 24'(-71148);
			1672: out = 24'(-33764);
			1673: out = 24'(17008);
			1674: out = 24'(39340);
			1675: out = 24'(-36776);
			1676: out = 24'(-65720);
			1677: out = 24'(-37892);
			1678: out = 24'(36384);
			1679: out = 24'(1152);
			1680: out = 24'(-30364);
			1681: out = 24'(27052);
			1682: out = 24'(15712);
			1683: out = 24'(11872);
			1684: out = 24'(-12988);
			1685: out = 24'(-4276);
			1686: out = 24'(2096);
			1687: out = 24'(23552);
			1688: out = 24'(27008);
			1689: out = 24'(13160);
			1690: out = 24'(-13768);
			1691: out = 24'(-23652);
			1692: out = 24'(-14316);
			1693: out = 24'(18444);
			1694: out = 24'(33716);
			1695: out = 24'(20716);
			1696: out = 24'(4256);
			1697: out = 24'(-17672);
			1698: out = 24'(-29572);
			1699: out = 24'(-20728);
			1700: out = 24'(2376);
			1701: out = 24'(22380);
			1702: out = 24'(18808);
			1703: out = 24'(32864);
			1704: out = 24'(-1536);
			1705: out = 24'(-46664);
			1706: out = 24'(-35704);
			1707: out = 24'(-20888);
			1708: out = 24'(11624);
			1709: out = 24'(26360);
			1710: out = 24'(35284);
			1711: out = 24'(13060);
			1712: out = 24'(-3876);
			1713: out = 24'(-1852);
			1714: out = 24'(18764);
			1715: out = 24'(16700);
			1716: out = 24'(-11928);
			1717: out = 24'(-18140);
			1718: out = 24'(-8824);
			1719: out = 24'(3936);
			1720: out = 24'(-42740);
			1721: out = 24'(2420);
			1722: out = 24'(36876);
			1723: out = 24'(37252);
			1724: out = 24'(25488);
			1725: out = 24'(-24296);
			1726: out = 24'(-51644);
			1727: out = 24'(38212);
			1728: out = 24'(14040);
			1729: out = 24'(-14144);
			1730: out = 24'(-51692);
			1731: out = 24'(20184);
			1732: out = 24'(34752);
			1733: out = 24'(28740);
			1734: out = 24'(6576);
			1735: out = 24'(4388);
			1736: out = 24'(7940);
			1737: out = 24'(22224);
			1738: out = 24'(-29604);
			1739: out = 24'(-20752);
			1740: out = 24'(-1392);
			1741: out = 24'(12312);
			1742: out = 24'(-20812);
			1743: out = 24'(-22596);
			1744: out = 24'(17160);
			1745: out = 24'(22608);
			1746: out = 24'(25692);
			1747: out = 24'(15208);
			1748: out = 24'(36608);
			1749: out = 24'(-5896);
			1750: out = 24'(2928);
			1751: out = 24'(40192);
			1752: out = 24'(-5732);
			1753: out = 24'(4288);
			1754: out = 24'(3736);
			1755: out = 24'(-45404);
			1756: out = 24'(-9216);
			1757: out = 24'(5480);
			1758: out = 24'(-2544);
			1759: out = 24'(-6884);
			1760: out = 24'(-21788);
			1761: out = 24'(-19448);
			1762: out = 24'(17096);
			1763: out = 24'(-1036);
			1764: out = 24'(1352);
			1765: out = 24'(16132);
			1766: out = 24'(-7820);
			1767: out = 24'(-3164);
			1768: out = 24'(-6820);
			1769: out = 24'(-22604);
			1770: out = 24'(8644);
			1771: out = 24'(34432);
			1772: out = 24'(33664);
			1773: out = 24'(6296);
			1774: out = 24'(-32708);
			1775: out = 24'(-38452);
			1776: out = 24'(13384);
			1777: out = 24'(2772);
			1778: out = 24'(-3868);
			1779: out = 24'(-9048);
			1780: out = 24'(-864);
			1781: out = 24'(7768);
			1782: out = 24'(7956);
			1783: out = 24'(1560);
			1784: out = 24'(-1472);
			1785: out = 24'(9280);
			1786: out = 24'(16264);
			1787: out = 24'(4540);
			1788: out = 24'(-11652);
			1789: out = 24'(-10668);
			1790: out = 24'(1312);
			1791: out = 24'(37804);
			1792: out = 24'(2004);
			1793: out = 24'(-56736);
			1794: out = 24'(2120);
			1795: out = 24'(13904);
			1796: out = 24'(9664);
			1797: out = 24'(-54872);
			1798: out = 24'(5164);
			1799: out = 24'(2664);
			1800: out = 24'(-4448);
			1801: out = 24'(12360);
			1802: out = 24'(26996);
			1803: out = 24'(2768);
			1804: out = 24'(-78304);
			1805: out = 24'(-22928);
			1806: out = 24'(-3636);
			1807: out = 24'(11784);
			1808: out = 24'(39072);
			1809: out = 24'(27696);
			1810: out = 24'(-1084);
			1811: out = 24'(-32180);
			1812: out = 24'(-34068);
			1813: out = 24'(-8864);
			1814: out = 24'(16204);
			1815: out = 24'(416);
			1816: out = 24'(-9900);
			1817: out = 24'(-24300);
			1818: out = 24'(-20884);
			1819: out = 24'(-8288);
			1820: out = 24'(4824);
			1821: out = 24'(-3276);
			1822: out = 24'(-19764);
			1823: out = 24'(-28324);
			1824: out = 24'(-212);
			1825: out = 24'(38744);
			1826: out = 24'(7768);
			1827: out = 24'(1984);
			1828: out = 24'(1552);
			1829: out = 24'(-55664);
			1830: out = 24'(14796);
			1831: out = 24'(38508);
			1832: out = 24'(26996);
			1833: out = 24'(-29960);
			1834: out = 24'(-18544);
			1835: out = 24'(5040);
			1836: out = 24'(11724);
			1837: out = 24'(-13504);
			1838: out = 24'(2060);
			1839: out = 24'(34576);
			1840: out = 24'(12984);
			1841: out = 24'(-48004);
			1842: out = 24'(-75576);
			1843: out = 24'(29484);
			1844: out = 24'(35540);
			1845: out = 24'(10732);
			1846: out = 24'(-50652);
			1847: out = 24'(-32284);
			1848: out = 24'(-13800);
			1849: out = 24'(18256);
			1850: out = 24'(33156);
			1851: out = 24'(8228);
			1852: out = 24'(1640);
			1853: out = 24'(22464);
			1854: out = 24'(33424);
			1855: out = 24'(23368);
			1856: out = 24'(-124);
			1857: out = 24'(-13616);
			1858: out = 24'(-2584);
			1859: out = 24'(5208);
			1860: out = 24'(520);
			1861: out = 24'(-11360);
			1862: out = 24'(-496);
			1863: out = 24'(14448);
			1864: out = 24'(18024);
			1865: out = 24'(-16564);
			1866: out = 24'(-11264);
			1867: out = 24'(25960);
			1868: out = 24'(-66740);
			1869: out = 24'(-6756);
			1870: out = 24'(34448);
			1871: out = 24'(20416);
			1872: out = 24'(-10516);
			1873: out = 24'(-27732);
			1874: out = 24'(-10840);
			1875: out = 24'(14668);
			1876: out = 24'(25456);
			1877: out = 24'(9088);
			1878: out = 24'(-13516);
			1879: out = 24'(-7660);
			1880: out = 24'(13096);
			1881: out = 24'(22524);
			1882: out = 24'(13576);
			1883: out = 24'(-11832);
			1884: out = 24'(-9712);
			1885: out = 24'(28108);
			1886: out = 24'(-2304);
			1887: out = 24'(-20632);
			1888: out = 24'(-26736);
			1889: out = 24'(14708);
			1890: out = 24'(20476);
			1891: out = 24'(18688);
			1892: out = 24'(6804);
			1893: out = 24'(9828);
			1894: out = 24'(-3996);
			1895: out = 24'(-17408);
			1896: out = 24'(17400);
			1897: out = 24'(484);
			1898: out = 24'(7612);
			1899: out = 24'(20800);
			1900: out = 24'(16388);
			1901: out = 24'(-32096);
			1902: out = 24'(-71008);
			1903: out = 24'(1584);
			1904: out = 24'(26980);
			1905: out = 24'(44640);
			1906: out = 24'(30952);
			1907: out = 24'(13008);
			1908: out = 24'(-10772);
			1909: out = 24'(-18224);
			1910: out = 24'(-19604);
			1911: out = 24'(3604);
			1912: out = 24'(13804);
			1913: out = 24'(10092);
			1914: out = 24'(8520);
			1915: out = 24'(4308);
			1916: out = 24'(2260);
			1917: out = 24'(-2424);
			1918: out = 24'(-3460);
			1919: out = 24'(-2216);
			1920: out = 24'(7552);
			1921: out = 24'(7928);
			1922: out = 24'(19176);
			1923: out = 24'(21168);
			1924: out = 24'(23740);
			1925: out = 24'(-5788);
			1926: out = 24'(-3112);
			1927: out = 24'(23400);
			1928: out = 24'(18372);
			1929: out = 24'(11880);
			1930: out = 24'(4504);
			1931: out = 24'(16616);
			1932: out = 24'(15804);
			1933: out = 24'(11156);
			1934: out = 24'(-2724);
			1935: out = 24'(472);
			1936: out = 24'(5216);
			1937: out = 24'(8348);
			1938: out = 24'(-20404);
			1939: out = 24'(-10432);
			1940: out = 24'(-15152);
			1941: out = 24'(-9240);
			1942: out = 24'(460);
			1943: out = 24'(29724);
			1944: out = 24'(21332);
			1945: out = 24'(-40504);
			1946: out = 24'(-55448);
			1947: out = 24'(-32032);
			1948: out = 24'(22600);
			1949: out = 24'(18636);
			1950: out = 24'(27664);
			1951: out = 24'(17236);
			1952: out = 24'(13304);
			1953: out = 24'(-19312);
			1954: out = 24'(-26448);
			1955: out = 24'(-20284);
			1956: out = 24'(-2312);
			1957: out = 24'(6864);
			1958: out = 24'(15076);
			1959: out = 24'(11100);
			1960: out = 24'(10844);
			1961: out = 24'(-6500);
			1962: out = 24'(-17588);
			1963: out = 24'(-22620);
			1964: out = 24'(1500);
			1965: out = 24'(5928);
			1966: out = 24'(-13076);
			1967: out = 24'(-34340);
			1968: out = 24'(-16472);
			1969: out = 24'(17836);
			1970: out = 24'(4412);
			1971: out = 24'(-5848);
			1972: out = 24'(-12004);
			1973: out = 24'(9024);
			1974: out = 24'(8788);
			1975: out = 24'(9596);
			1976: out = 24'(884);
			1977: out = 24'(2432);
			1978: out = 24'(-12232);
			1979: out = 24'(-24176);
			1980: out = 24'(-30256);
			1981: out = 24'(-7088);
			1982: out = 24'(8988);
			1983: out = 24'(12568);
			1984: out = 24'(32472);
			1985: out = 24'(2216);
			1986: out = 24'(468);
			1987: out = 24'(28036);
			1988: out = 24'(18936);
			1989: out = 24'(1468);
			1990: out = 24'(-21452);
			1991: out = 24'(-48088);
			1992: out = 24'(-7504);
			1993: out = 24'(21844);
			1994: out = 24'(9884);
			1995: out = 24'(13100);
			1996: out = 24'(-2352);
			1997: out = 24'(-9420);
			1998: out = 24'(1424);
			1999: out = 24'(-10180);
			2000: out = 24'(-9748);
			2001: out = 24'(8204);
			2002: out = 24'(-2240);
			2003: out = 24'(10788);
			2004: out = 24'(24264);
			2005: out = 24'(15716);
			2006: out = 24'(8132);
			2007: out = 24'(-22576);
			2008: out = 24'(-53488);
			2009: out = 24'(-35804);
			2010: out = 24'(7840);
			2011: out = 24'(32636);
			2012: out = 24'(4060);
			2013: out = 24'(-6804);
			2014: out = 24'(-3924);
			2015: out = 24'(17196);
			2016: out = 24'(-19640);
			2017: out = 24'(-30392);
			2018: out = 24'(-23580);
			2019: out = 24'(24664);
			2020: out = 24'(8228);
			2021: out = 24'(-8864);
			2022: out = 24'(-28588);
			2023: out = 24'(-11100);
			2024: out = 24'(-4480);
			2025: out = 24'(972);
			2026: out = 24'(-12040);
			2027: out = 24'(16896);
			2028: out = 24'(6912);
			2029: out = 24'(-29448);
			2030: out = 24'(26996);
			2031: out = 24'(1876);
			2032: out = 24'(-23512);
			2033: out = 24'(-32084);
			2034: out = 24'(8);
			2035: out = 24'(12868);
			2036: out = 24'(1012);
			2037: out = 24'(27024);
			2038: out = 24'(6564);
			2039: out = 24'(-13060);
			2040: out = 24'(-33040);
			2041: out = 24'(4476);
			2042: out = 24'(23364);
			2043: out = 24'(17604);
			2044: out = 24'(-16156);
			2045: out = 24'(-33896);
			2046: out = 24'(-32596);
			2047: out = 24'(-8928);
			2048: out = 24'(2912);
			2049: out = 24'(16);
			2050: out = 24'(-19116);
			2051: out = 24'(24400);
			2052: out = 24'(-14112);
			2053: out = 24'(-24192);
			2054: out = 24'(13748);
			2055: out = 24'(32576);
			2056: out = 24'(19984);
			2057: out = 24'(-16416);
			2058: out = 24'(-15296);
			2059: out = 24'(-23636);
			2060: out = 24'(-6528);
			2061: out = 24'(22624);
			2062: out = 24'(17224);
			2063: out = 24'(1448);
			2064: out = 24'(-19608);
			2065: out = 24'(10652);
			2066: out = 24'(-20816);
			2067: out = 24'(-17440);
			2068: out = 24'(29576);
			2069: out = 24'(19292);
			2070: out = 24'(1604);
			2071: out = 24'(-24224);
			2072: out = 24'(-22436);
			2073: out = 24'(6596);
			2074: out = 24'(32608);
			2075: out = 24'(15656);
			2076: out = 24'(26376);
			2077: out = 24'(-13220);
			2078: out = 24'(-45916);
			2079: out = 24'(-45508);
			2080: out = 24'(2528);
			2081: out = 24'(34876);
			2082: out = 24'(24836);
			2083: out = 24'(10256);
			2084: out = 24'(-9588);
			2085: out = 24'(-4488);
			2086: out = 24'(25944);
			2087: out = 24'(27084);
			2088: out = 24'(3464);
			2089: out = 24'(-31600);
			2090: out = 24'(-15408);
			2091: out = 24'(-5456);
			2092: out = 24'(4776);
			2093: out = 24'(32024);
			2094: out = 24'(-1048);
			2095: out = 24'(-11444);
			2096: out = 24'(6960);
			2097: out = 24'(-5796);
			2098: out = 24'(620);
			2099: out = 24'(4560);
			2100: out = 24'(7604);
			2101: out = 24'(5052);
			2102: out = 24'(12416);
			2103: out = 24'(27280);
			2104: out = 24'(-9680);
			2105: out = 24'(-5132);
			2106: out = 24'(5344);
			2107: out = 24'(11340);
			2108: out = 24'(6984);
			2109: out = 24'(7320);
			2110: out = 24'(8156);
			2111: out = 24'(1680);
			2112: out = 24'(-6932);
			2113: out = 24'(-12672);
			2114: out = 24'(-32588);
			2115: out = 24'(14020);
			2116: out = 24'(15808);
			2117: out = 24'(-14620);
			2118: out = 24'(-16268);
			2119: out = 24'(3184);
			2120: out = 24'(20588);
			2121: out = 24'(-23676);
			2122: out = 24'(11860);
			2123: out = 24'(15960);
			2124: out = 24'(19836);
			2125: out = 24'(2976);
			2126: out = 24'(22904);
			2127: out = 24'(22252);
			2128: out = 24'(-5344);
			2129: out = 24'(-18144);
			2130: out = 24'(-1504);
			2131: out = 24'(29148);
			2132: out = 24'(6384);
			2133: out = 24'(7536);
			2134: out = 24'(-4908);
			2135: out = 24'(-36340);
			2136: out = 24'(-1244);
			2137: out = 24'(17340);
			2138: out = 24'(22520);
			2139: out = 24'(10016);
			2140: out = 24'(14084);
			2141: out = 24'(1804);
			2142: out = 24'(-34460);
			2143: out = 24'(-27628);
			2144: out = 24'(-6952);
			2145: out = 24'(15812);
			2146: out = 24'(16904);
			2147: out = 24'(-7820);
			2148: out = 24'(-23064);
			2149: out = 24'(6276);
			2150: out = 24'(-18456);
			2151: out = 24'(-12296);
			2152: out = 24'(-3124);
			2153: out = 24'(19528);
			2154: out = 24'(2160);
			2155: out = 24'(-4184);
			2156: out = 24'(11252);
			2157: out = 24'(-17124);
			2158: out = 24'(-28588);
			2159: out = 24'(-22916);
			2160: out = 24'(31384);
			2161: out = 24'(19528);
			2162: out = 24'(13308);
			2163: out = 24'(23844);
			2164: out = 24'(-8376);
			2165: out = 24'(-8496);
			2166: out = 24'(-1892);
			2167: out = 24'(-28192);
			2168: out = 24'(-15568);
			2169: out = 24'(-3252);
			2170: out = 24'(10468);
			2171: out = 24'(1020);
			2172: out = 24'(14612);
			2173: out = 24'(19216);
			2174: out = 24'(-38856);
			2175: out = 24'(-12596);
			2176: out = 24'(13224);
			2177: out = 24'(19140);
			2178: out = 24'(26372);
			2179: out = 24'(5552);
			2180: out = 24'(-13528);
			2181: out = 24'(-15936);
			2182: out = 24'(4744);
			2183: out = 24'(13156);
			2184: out = 24'(-1228);
			2185: out = 24'(11832);
			2186: out = 24'(592);
			2187: out = 24'(-9452);
			2188: out = 24'(444);
			2189: out = 24'(944);
			2190: out = 24'(11432);
			2191: out = 24'(16852);
			2192: out = 24'(19328);
			2193: out = 24'(-16108);
			2194: out = 24'(-45824);
			2195: out = 24'(-12832);
			2196: out = 24'(8484);
			2197: out = 24'(28384);
			2198: out = 24'(18248);
			2199: out = 24'(16828);
			2200: out = 24'(-21076);
			2201: out = 24'(-48924);
			2202: out = 24'(-56616);
			2203: out = 24'(-16000);
			2204: out = 24'(7016);
			2205: out = 24'(1732);
			2206: out = 24'(31268);
			2207: out = 24'(11892);
			2208: out = 24'(-7444);
			2209: out = 24'(2620);
			2210: out = 24'(-30324);
			2211: out = 24'(-36824);
			2212: out = 24'(-21280);
			2213: out = 24'(-17488);
			2214: out = 24'(-9116);
			2215: out = 24'(1464);
			2216: out = 24'(26564);
			2217: out = 24'(1196);
			2218: out = 24'(-17096);
			2219: out = 24'(-24768);
			2220: out = 24'(-12956);
			2221: out = 24'(9124);
			2222: out = 24'(28272);
			2223: out = 24'(28888);
			2224: out = 24'(-4872);
			2225: out = 24'(-45468);
			2226: out = 24'(-63896);
			2227: out = 24'(-21468);
			2228: out = 24'(21604);
			2229: out = 24'(34384);
			2230: out = 24'(7128);
			2231: out = 24'(6184);
			2232: out = 24'(5272);
			2233: out = 24'(8468);
			2234: out = 24'(-11528);
			2235: out = 24'(-12912);
			2236: out = 24'(-8704);
			2237: out = 24'(3948);
			2238: out = 24'(-7284);
			2239: out = 24'(-10396);
			2240: out = 24'(-6108);
			2241: out = 24'(-4100);
			2242: out = 24'(9916);
			2243: out = 24'(6548);
			2244: out = 24'(-27444);
			2245: out = 24'(-23632);
			2246: out = 24'(-13292);
			2247: out = 24'(9028);
			2248: out = 24'(-23128);
			2249: out = 24'(11376);
			2250: out = 24'(15944);
			2251: out = 24'(-16812);
			2252: out = 24'(5168);
			2253: out = 24'(10480);
			2254: out = 24'(3416);
			2255: out = 24'(26496);
			2256: out = 24'(-26552);
			2257: out = 24'(-34000);
			2258: out = 24'(33716);
			2259: out = 24'(13204);
			2260: out = 24'(10204);
			2261: out = 24'(-4648);
			2262: out = 24'(-4888);
			2263: out = 24'(-10252);
			2264: out = 24'(-9920);
			2265: out = 24'(-19932);
			2266: out = 24'(17736);
			2267: out = 24'(17176);
			2268: out = 24'(10068);
			2269: out = 24'(20396);
			2270: out = 24'(7096);
			2271: out = 24'(-1232);
			2272: out = 24'(2324);
			2273: out = 24'(-10016);
			2274: out = 24'(1016);
			2275: out = 24'(13432);
			2276: out = 24'(12916);
			2277: out = 24'(11148);
			2278: out = 24'(4332);
			2279: out = 24'(-6180);
			2280: out = 24'(-7064);
			2281: out = 24'(-4028);
			2282: out = 24'(10364);
			2283: out = 24'(19000);
			2284: out = 24'(25612);
			2285: out = 24'(5416);
			2286: out = 24'(-19320);
			2287: out = 24'(-23200);
			2288: out = 24'(2024);
			2289: out = 24'(23464);
			2290: out = 24'(32228);
			2291: out = 24'(-15068);
			2292: out = 24'(-27996);
			2293: out = 24'(-20);
			2294: out = 24'(3020);
			2295: out = 24'(-2832);
			2296: out = 24'(-10048);
			2297: out = 24'(17840);
			2298: out = 24'(27280);
			2299: out = 24'(28156);
			2300: out = 24'(7500);
			2301: out = 24'(4144);
			2302: out = 24'(-1736);
			2303: out = 24'(-2356);
			2304: out = 24'(-35416);
			2305: out = 24'(76);
			2306: out = 24'(13684);
			2307: out = 24'(20796);
			2308: out = 24'(-23248);
			2309: out = 24'(-4632);
			2310: out = 24'(15152);
			2311: out = 24'(31056);
			2312: out = 24'(-13696);
			2313: out = 24'(-15588);
			2314: out = 24'(12216);
			2315: out = 24'(32876);
			2316: out = 24'(13200);
			2317: out = 24'(-17308);
			2318: out = 24'(-35356);
			2319: out = 24'(-8248);
			2320: out = 24'(10112);
			2321: out = 24'(10608);
			2322: out = 24'(1312);
			2323: out = 24'(5404);
			2324: out = 24'(4300);
			2325: out = 24'(-10636);
			2326: out = 24'(-10132);
			2327: out = 24'(7620);
			2328: out = 24'(26188);
			2329: out = 24'(-1280);
			2330: out = 24'(-11512);
			2331: out = 24'(-7168);
			2332: out = 24'(26340);
			2333: out = 24'(-11736);
			2334: out = 24'(-33632);
			2335: out = 24'(-38920);
			2336: out = 24'(26492);
			2337: out = 24'(30008);
			2338: out = 24'(25992);
			2339: out = 24'(9892);
			2340: out = 24'(7920);
			2341: out = 24'(-4760);
			2342: out = 24'(-15724);
			2343: out = 24'(-45856);
			2344: out = 24'(-12160);
			2345: out = 24'(16052);
			2346: out = 24'(14688);
			2347: out = 24'(2980);
			2348: out = 24'(-12540);
			2349: out = 24'(-14008);
			2350: out = 24'(-4152);
			2351: out = 24'(10240);
			2352: out = 24'(14036);
			2353: out = 24'(9552);
			2354: out = 24'(-5376);
			2355: out = 24'(-4972);
			2356: out = 24'(2692);
			2357: out = 24'(1040);
			2358: out = 24'(-1016);
			2359: out = 24'(-8688);
			2360: out = 24'(-12072);
			2361: out = 24'(-17408);
			2362: out = 24'(-3856);
			2363: out = 24'(6144);
			2364: out = 24'(-19100);
			2365: out = 24'(1556);
			2366: out = 24'(16652);
			2367: out = 24'(19948);
			2368: out = 24'(564);
			2369: out = 24'(-16336);
			2370: out = 24'(-20816);
			2371: out = 24'(5452);
			2372: out = 24'(-3516);
			2373: out = 24'(-8860);
			2374: out = 24'(-7908);
			2375: out = 24'(18380);
			2376: out = 24'(20328);
			2377: out = 24'(3404);
			2378: out = 24'(-30124);
			2379: out = 24'(-30772);
			2380: out = 24'(-12368);
			2381: out = 24'(13792);
			2382: out = 24'(18400);
			2383: out = 24'(7688);
			2384: out = 24'(-14368);
			2385: out = 24'(-20704);
			2386: out = 24'(-21556);
			2387: out = 24'(2660);
			2388: out = 24'(20400);
			2389: out = 24'(8684);
			2390: out = 24'(-22300);
			2391: out = 24'(-33496);
			2392: out = 24'(7836);
			2393: out = 24'(18416);
			2394: out = 24'(8536);
			2395: out = 24'(-24664);
			2396: out = 24'(-3060);
			2397: out = 24'(-12780);
			2398: out = 24'(-11668);
			2399: out = 24'(3300);
			2400: out = 24'(-11496);
			2401: out = 24'(-16908);
			2402: out = 24'(-5300);
			2403: out = 24'(-4688);
			2404: out = 24'(18220);
			2405: out = 24'(21768);
			2406: out = 24'(-4744);
			2407: out = 24'(912);
			2408: out = 24'(1844);
			2409: out = 24'(1572);
			2410: out = 24'(9684);
			2411: out = 24'(-6256);
			2412: out = 24'(-18208);
			2413: out = 24'(-5068);
			2414: out = 24'(-4828);
			2415: out = 24'(6888);
			2416: out = 24'(11900);
			2417: out = 24'(4732);
			2418: out = 24'(-8476);
			2419: out = 24'(-16260);
			2420: out = 24'(-15420);
			2421: out = 24'(13612);
			2422: out = 24'(21892);
			2423: out = 24'(12096);
			2424: out = 24'(18780);
			2425: out = 24'(-2904);
			2426: out = 24'(-12516);
			2427: out = 24'(-5532);
			2428: out = 24'(6788);
			2429: out = 24'(7296);
			2430: out = 24'(-3840);
			2431: out = 24'(-7696);
			2432: out = 24'(-9248);
			2433: out = 24'(4856);
			2434: out = 24'(22524);
			2435: out = 24'(15356);
			2436: out = 24'(1008);
			2437: out = 24'(-7304);
			2438: out = 24'(9960);
			2439: out = 24'(11144);
			2440: out = 24'(204);
			2441: out = 24'(-22084);
			2442: out = 24'(5208);
			2443: out = 24'(15452);
			2444: out = 24'(15868);
			2445: out = 24'(27720);
			2446: out = 24'(4692);
			2447: out = 24'(-3020);
			2448: out = 24'(4624);
			2449: out = 24'(-364);
			2450: out = 24'(-12528);
			2451: out = 24'(-21580);
			2452: out = 24'(-8008);
			2453: out = 24'(10560);
			2454: out = 24'(13100);
			2455: out = 24'(-9588);
			2456: out = 24'(-460);
			2457: out = 24'(2280);
			2458: out = 24'(7848);
			2459: out = 24'(-18888);
			2460: out = 24'(7260);
			2461: out = 24'(11844);
			2462: out = 24'(756);
			2463: out = 24'(16524);
			2464: out = 24'(4060);
			2465: out = 24'(-16372);
			2466: out = 24'(-4992);
			2467: out = 24'(-23896);
			2468: out = 24'(-4648);
			2469: out = 24'(25940);
			2470: out = 24'(20724);
			2471: out = 24'(-8220);
			2472: out = 24'(-37536);
			2473: out = 24'(-42856);
			2474: out = 24'(4512);
			2475: out = 24'(33904);
			2476: out = 24'(23328);
			2477: out = 24'(-13288);
			2478: out = 24'(-22816);
			2479: out = 24'(-5880);
			2480: out = 24'(-1296);
			2481: out = 24'(24652);
			2482: out = 24'(17564);
			2483: out = 24'(-2172);
			2484: out = 24'(-23924);
			2485: out = 24'(-13812);
			2486: out = 24'(9060);
			2487: out = 24'(16988);
			2488: out = 24'(20476);
			2489: out = 24'(-2912);
			2490: out = 24'(-30080);
			2491: out = 24'(17372);
			2492: out = 24'(19428);
			2493: out = 24'(12008);
			2494: out = 24'(-2604);
			2495: out = 24'(-4792);
			2496: out = 24'(-10736);
			2497: out = 24'(-13596);
			2498: out = 24'(14116);
			2499: out = 24'(16800);
			2500: out = 24'(10124);
			2501: out = 24'(-9408);
			2502: out = 24'(10692);
			2503: out = 24'(7832);
			2504: out = 24'(-6352);
			2505: out = 24'(19232);
			2506: out = 24'(6092);
			2507: out = 24'(-744);
			2508: out = 24'(348);
			2509: out = 24'(2484);
			2510: out = 24'(-5052);
			2511: out = 24'(-11760);
			2512: out = 24'(15096);
			2513: out = 24'(12868);
			2514: out = 24'(6140);
			2515: out = 24'(-1612);
			2516: out = 24'(4344);
			2517: out = 24'(9292);
			2518: out = 24'(4036);
			2519: out = 24'(-37668);
			2520: out = 24'(-23240);
			2521: out = 24'(7964);
			2522: out = 24'(20964);
			2523: out = 24'(21000);
			2524: out = 24'(-14952);
			2525: out = 24'(-44176);
			2526: out = 24'(-14052);
			2527: out = 24'(8844);
			2528: out = 24'(17284);
			2529: out = 24'(6952);
			2530: out = 24'(-92);
			2531: out = 24'(6116);
			2532: out = 24'(14864);
			2533: out = 24'(10268);
			2534: out = 24'(-6476);
			2535: out = 24'(-9064);
			2536: out = 24'(11744);
			2537: out = 24'(14616);
			2538: out = 24'(12708);
			2539: out = 24'(1384);
			2540: out = 24'(-15208);
			2541: out = 24'(3020);
			2542: out = 24'(14888);
			2543: out = 24'(7264);
			2544: out = 24'(-8576);
			2545: out = 24'(-5976);
			2546: out = 24'(8760);
			2547: out = 24'(-5488);
			2548: out = 24'(1480);
			2549: out = 24'(-4720);
			2550: out = 24'(-2788);
			2551: out = 24'(-14516);
			2552: out = 24'(2188);
			2553: out = 24'(11244);
			2554: out = 24'(10480);
			2555: out = 24'(-13628);
			2556: out = 24'(-16376);
			2557: out = 24'(-1416);
			2558: out = 24'(5092);
			2559: out = 24'(-6804);
			2560: out = 24'(-14492);
			2561: out = 24'(5808);
			2562: out = 24'(13936);
			2563: out = 24'(5208);
			2564: out = 24'(-20368);
			2565: out = 24'(-28300);
			2566: out = 24'(-15028);
			2567: out = 24'(8080);
			2568: out = 24'(2432);
			2569: out = 24'(18812);
			2570: out = 24'(3340);
			2571: out = 24'(-28148);
			2572: out = 24'(-11448);
			2573: out = 24'(-26792);
			2574: out = 24'(-21232);
			2575: out = 24'(29920);
			2576: out = 24'(10388);
			2577: out = 24'(-12972);
			2578: out = 24'(-39956);
			2579: out = 24'(-4956);
			2580: out = 24'(2408);
			2581: out = 24'(11372);
			2582: out = 24'(17004);
			2583: out = 24'(9176);
			2584: out = 24'(-5824);
			2585: out = 24'(-16020);
			2586: out = 24'(-11080);
			2587: out = 24'(5264);
			2588: out = 24'(8948);
			2589: out = 24'(-22060);
			2590: out = 24'(12084);
			2591: out = 24'(15892);
			2592: out = 24'(5168);
			2593: out = 24'(4092);
			2594: out = 24'(-3148);
			2595: out = 24'(-7360);
			2596: out = 24'(-12980);
			2597: out = 24'(4900);
			2598: out = 24'(11008);
			2599: out = 24'(7764);
			2600: out = 24'(-2900);
			2601: out = 24'(-4052);
			2602: out = 24'(392);
			2603: out = 24'(6404);
			2604: out = 24'(4024);
			2605: out = 24'(-2652);
			2606: out = 24'(-10392);
			2607: out = 24'(-3068);
			2608: out = 24'(-1632);
			2609: out = 24'(5248);
			2610: out = 24'(8916);
			2611: out = 24'(14192);
			2612: out = 24'(6784);
			2613: out = 24'(444);
			2614: out = 24'(768);
			2615: out = 24'(3216);
			2616: out = 24'(6360);
			2617: out = 24'(20148);
			2618: out = 24'(-29144);
			2619: out = 24'(-25100);
			2620: out = 24'(780);
			2621: out = 24'(25696);
			2622: out = 24'(-3920);
			2623: out = 24'(-22524);
			2624: out = 24'(-3388);
			2625: out = 24'(4236);
			2626: out = 24'(12496);
			2627: out = 24'(5572);
			2628: out = 24'(16);
			2629: out = 24'(4192);
			2630: out = 24'(14244);
			2631: out = 24'(12436);
			2632: out = 24'(-7644);
			2633: out = 24'(-9952);
			2634: out = 24'(2756);
			2635: out = 24'(-40532);
			2636: out = 24'(10096);
			2637: out = 24'(17840);
			2638: out = 24'(-508);
			2639: out = 24'(-27420);
			2640: out = 24'(-4912);
			2641: out = 24'(17292);
			2642: out = 24'(-18288);
			2643: out = 24'(-24376);
			2644: out = 24'(-14152);
			2645: out = 24'(17820);
			2646: out = 24'(19496);
			2647: out = 24'(4384);
			2648: out = 24'(-16056);
			2649: out = 24'(5112);
			2650: out = 24'(6784);
			2651: out = 24'(17176);
			2652: out = 24'(14120);
			2653: out = 24'(-4352);
			2654: out = 24'(-17904);
			2655: out = 24'(-11536);
			2656: out = 24'(13292);
			2657: out = 24'(7292);
			2658: out = 24'(-8304);
			2659: out = 24'(-21788);
			2660: out = 24'(5852);
			2661: out = 24'(14624);
			2662: out = 24'(8800);
			2663: out = 24'(-15588);
			2664: out = 24'(-10152);
			2665: out = 24'(-3304);
			2666: out = 24'(2492);
			2667: out = 24'(3880);
			2668: out = 24'(3428);
			2669: out = 24'(1980);
			2670: out = 24'(1948);
			2671: out = 24'(1944);
			2672: out = 24'(2604);
			2673: out = 24'(1900);
			2674: out = 24'(2704);
			2675: out = 24'(232);
			2676: out = 24'(2880);
			2677: out = 24'(14496);
			2678: out = 24'(5576);
			2679: out = 24'(-5968);
			2680: out = 24'(-15752);
			2681: out = 24'(17096);
			2682: out = 24'(6508);
			2683: out = 24'(-8852);
			2684: out = 24'(-17896);
			2685: out = 24'(-7056);
			2686: out = 24'(-2420);
			2687: out = 24'(-7708);
			2688: out = 24'(22244);
			2689: out = 24'(-3748);
			2690: out = 24'(-22404);
			2691: out = 24'(-12296);
			2692: out = 24'(1812);
			2693: out = 24'(13840);
			2694: out = 24'(9028);
			2695: out = 24'(-1596);
			2696: out = 24'(-19632);
			2697: out = 24'(-14904);
			2698: out = 24'(19060);
			2699: out = 24'(6196);
			2700: out = 24'(-4840);
			2701: out = 24'(-14644);
			2702: out = 24'(25344);
			2703: out = 24'(5616);
			2704: out = 24'(-14440);
			2705: out = 24'(-35332);
			2706: out = 24'(5780);
			2707: out = 24'(21036);
			2708: out = 24'(18252);
			2709: out = 24'(-20684);
			2710: out = 24'(-556);
			2711: out = 24'(10828);
			2712: out = 24'(148);
			2713: out = 24'(4536);
			2714: out = 24'(12104);
			2715: out = 24'(16388);
			2716: out = 24'(-16804);
			2717: out = 24'(-11604);
			2718: out = 24'(-2512);
			2719: out = 24'(4824);
			2720: out = 24'(12064);
			2721: out = 24'(184);
			2722: out = 24'(-14160);
			2723: out = 24'(-12856);
			2724: out = 24'(4512);
			2725: out = 24'(10584);
			2726: out = 24'(-7872);
			2727: out = 24'(6512);
			2728: out = 24'(5496);
			2729: out = 24'(5568);
			2730: out = 24'(-11672);
			2731: out = 24'(-4940);
			2732: out = 24'(-252);
			2733: out = 24'(12680);
			2734: out = 24'(12484);
			2735: out = 24'(17336);
			2736: out = 24'(6184);
			2737: out = 24'(2348);
			2738: out = 24'(-31716);
			2739: out = 24'(-17996);
			2740: out = 24'(24984);
			2741: out = 24'(18436);
			2742: out = 24'(-1416);
			2743: out = 24'(-23492);
			2744: out = 24'(-21036);
			2745: out = 24'(5668);
			2746: out = 24'(20144);
			2747: out = 24'(12176);
			2748: out = 24'(556);
			2749: out = 24'(488);
			2750: out = 24'(1400);
			2751: out = 24'(-19072);
			2752: out = 24'(-4652);
			2753: out = 24'(5816);
			2754: out = 24'(6012);
			2755: out = 24'(23008);
			2756: out = 24'(-17916);
			2757: out = 24'(-46860);
			2758: out = 24'(-5380);
			2759: out = 24'(5932);
			2760: out = 24'(17580);
			2761: out = 24'(7592);
			2762: out = 24'(-972);
			2763: out = 24'(-10828);
			2764: out = 24'(-7036);
			2765: out = 24'(-6184);
			2766: out = 24'(9820);
			2767: out = 24'(4564);
			2768: out = 24'(-5832);
			2769: out = 24'(13220);
			2770: out = 24'(11884);
			2771: out = 24'(9376);
			2772: out = 24'(11988);
			2773: out = 24'(-572);
			2774: out = 24'(-4456);
			2775: out = 24'(-2728);
			2776: out = 24'(12556);
			2777: out = 24'(5548);
			2778: out = 24'(-4164);
			2779: out = 24'(-12036);
			2780: out = 24'(2940);
			2781: out = 24'(8676);
			2782: out = 24'(4584);
			2783: out = 24'(-17100);
			2784: out = 24'(-2536);
			2785: out = 24'(11984);
			2786: out = 24'(2252);
			2787: out = 24'(8492);
			2788: out = 24'(-11764);
			2789: out = 24'(-25456);
			2790: out = 24'(9236);
			2791: out = 24'(16372);
			2792: out = 24'(8112);
			2793: out = 24'(-24268);
			2794: out = 24'(5812);
			2795: out = 24'(-856);
			2796: out = 24'(-14548);
			2797: out = 24'(10224);
			2798: out = 24'(-1952);
			2799: out = 24'(-7316);
			2800: out = 24'(-7080);
			2801: out = 24'(4892);
			2802: out = 24'(-2408);
			2803: out = 24'(-13788);
			2804: out = 24'(10396);
			2805: out = 24'(6964);
			2806: out = 24'(-548);
			2807: out = 24'(-30796);
			2808: out = 24'(13408);
			2809: out = 24'(-3140);
			2810: out = 24'(-23280);
			2811: out = 24'(-14928);
			2812: out = 24'(6704);
			2813: out = 24'(9840);
			2814: out = 24'(-9900);
			2815: out = 24'(-11000);
			2816: out = 24'(-852);
			2817: out = 24'(8400);
			2818: out = 24'(-17184);
			2819: out = 24'(-12992);
			2820: out = 24'(-5744);
			2821: out = 24'(2172);
			2822: out = 24'(1260);
			2823: out = 24'(-15004);
			2824: out = 24'(-21708);
			2825: out = 24'(18472);
			2826: out = 24'(5752);
			2827: out = 24'(-10892);
			2828: out = 24'(-26368);
			2829: out = 24'(-27872);
			2830: out = 24'(-1688);
			2831: out = 24'(23060);
			2832: out = 24'(14396);
			2833: out = 24'(3740);
			2834: out = 24'(-6080);
			2835: out = 24'(1520);
			2836: out = 24'(828);
			2837: out = 24'(8364);
			2838: out = 24'(7004);
			2839: out = 24'(4120);
			2840: out = 24'(-4056);
			2841: out = 24'(-844);
			2842: out = 24'(7936);
			2843: out = 24'(4724);
			2844: out = 24'(3052);
			2845: out = 24'(-2860);
			2846: out = 24'(-12632);
			2847: out = 24'(-7816);
			2848: out = 24'(684);
			2849: out = 24'(7044);
			2850: out = 24'(2720);
			2851: out = 24'(-5392);
			2852: out = 24'(-6488);
			2853: out = 24'(15488);
			2854: out = 24'(-2256);
			2855: out = 24'(-7436);
			2856: out = 24'(-6268);
			2857: out = 24'(6768);
			2858: out = 24'(-1608);
			2859: out = 24'(-8044);
			2860: out = 24'(5196);
			2861: out = 24'(4812);
			2862: out = 24'(9392);
			2863: out = 24'(8176);
			2864: out = 24'(8804);
			2865: out = 24'(2120);
			2866: out = 24'(36);
			2867: out = 24'(-2808);
			2868: out = 24'(7152);
			2869: out = 24'(5560);
			2870: out = 24'(2324);
			2871: out = 24'(-948);
			2872: out = 24'(4240);
			2873: out = 24'(4328);
			2874: out = 24'(7464);
			2875: out = 24'(-13260);
			2876: out = 24'(-2636);
			2877: out = 24'(13012);
			2878: out = 24'(-9016);
			2879: out = 24'(-23824);
			2880: out = 24'(-21168);
			2881: out = 24'(10056);
			2882: out = 24'(19100);
			2883: out = 24'(5372);
			2884: out = 24'(-20256);
			2885: out = 24'(13672);
			2886: out = 24'(5104);
			2887: out = 24'(828);
			2888: out = 24'(-11772);
			2889: out = 24'(12624);
			2890: out = 24'(7112);
			2891: out = 24'(-6488);
			2892: out = 24'(2504);
			2893: out = 24'(-1228);
			2894: out = 24'(4676);
			2895: out = 24'(12816);
			2896: out = 24'(9656);
			2897: out = 24'(-1612);
			2898: out = 24'(-7324);
			2899: out = 24'(14268);
			2900: out = 24'(15396);
			2901: out = 24'(7380);
			2902: out = 24'(-9988);
			2903: out = 24'(-1160);
			2904: out = 24'(4860);
			2905: out = 24'(8972);
			2906: out = 24'(-720);
			2907: out = 24'(1528);
			2908: out = 24'(-3100);
			2909: out = 24'(-14008);
			2910: out = 24'(12148);
			2911: out = 24'(15580);
			2912: out = 24'(9908);
			2913: out = 24'(-5972);
			2914: out = 24'(3180);
			2915: out = 24'(7704);
			2916: out = 24'(4540);
			2917: out = 24'(6268);
			2918: out = 24'(3348);
			2919: out = 24'(-1204);
			2920: out = 24'(-1880);
			2921: out = 24'(-7408);
			2922: out = 24'(-496);
			2923: out = 24'(11932);
			2924: out = 24'(10568);
			2925: out = 24'(-2012);
			2926: out = 24'(-12384);
			2927: out = 24'(1580);
			2928: out = 24'(8036);
			2929: out = 24'(9840);
			2930: out = 24'(-1328);
			2931: out = 24'(12540);
			2932: out = 24'(3144);
			2933: out = 24'(-5708);
			2934: out = 24'(-19248);
			2935: out = 24'(4532);
			2936: out = 24'(12888);
			2937: out = 24'(3860);
			2938: out = 24'(-1576);
			2939: out = 24'(-13200);
			2940: out = 24'(-12160);
			2941: out = 24'(13000);
			2942: out = 24'(2444);
			2943: out = 24'(3548);
			2944: out = 24'(10220);
			2945: out = 24'(-436);
			2946: out = 24'(956);
			2947: out = 24'(3120);
			2948: out = 24'(2680);
			2949: out = 24'(-3316);
			2950: out = 24'(-13676);
			2951: out = 24'(-18924);
			2952: out = 24'(8044);
			2953: out = 24'(13616);
			2954: out = 24'(5684);
			2955: out = 24'(-15180);
			2956: out = 24'(-6904);
			2957: out = 24'(3976);
			2958: out = 24'(10844);
			2959: out = 24'(124);
			2960: out = 24'(984);
			2961: out = 24'(116);
			2962: out = 24'(-16924);
			2963: out = 24'(3372);
			2964: out = 24'(-84);
			2965: out = 24'(-6164);
			2966: out = 24'(5824);
			2967: out = 24'(16000);
			2968: out = 24'(7492);
			2969: out = 24'(-23536);
			2970: out = 24'(-22644);
			2971: out = 24'(-5276);
			2972: out = 24'(15424);
			2973: out = 24'(6744);
			2974: out = 24'(-7308);
			2975: out = 24'(-13920);
			2976: out = 24'(9888);
			2977: out = 24'(-4328);
			2978: out = 24'(-564);
			2979: out = 24'(336);
			2980: out = 24'(-4172);
			2981: out = 24'(280);
			2982: out = 24'(8524);
			2983: out = 24'(9688);
			2984: out = 24'(-892);
			2985: out = 24'(-9184);
			2986: out = 24'(-4860);
			2987: out = 24'(764);
			2988: out = 24'(7588);
			2989: out = 24'(2244);
			2990: out = 24'(1476);
			2991: out = 24'(-22760);
			2992: out = 24'(-7284);
			2993: out = 24'(8268);
			2994: out = 24'(956);
			2995: out = 24'(-27692);
			2996: out = 24'(-26796);
			2997: out = 24'(18728);
			2998: out = 24'(16852);
			2999: out = 24'(11880);
			3000: out = 24'(-10748);
			3001: out = 24'(-26468);
			3002: out = 24'(-26040);
			3003: out = 24'(-6944);
			3004: out = 24'(8408);
			3005: out = 24'(9588);
			3006: out = 24'(260);
			3007: out = 24'(-8220);
			3008: out = 24'(-8200);
			3009: out = 24'(-6880);
			3010: out = 24'(-2712);
			3011: out = 24'(-124);
			3012: out = 24'(6504);
			3013: out = 24'(-856);
			3014: out = 24'(-6860);
			3015: out = 24'(5616);
			3016: out = 24'(-1020);
			3017: out = 24'(-5764);
			3018: out = 24'(-9156);
			3019: out = 24'(-132);
			3020: out = 24'(2816);
			3021: out = 24'(1360);
			3022: out = 24'(-7236);
			3023: out = 24'(196);
			3024: out = 24'(2232);
			3025: out = 24'(-3980);
			3026: out = 24'(9016);
			3027: out = 24'(-2568);
			3028: out = 24'(-12212);
			3029: out = 24'(-13280);
			3030: out = 24'(7200);
			3031: out = 24'(12172);
			3032: out = 24'(72);
			3033: out = 24'(13036);
			3034: out = 24'(252);
			3035: out = 24'(-8880);
			3036: out = 24'(-7460);
			3037: out = 24'(-10164);
			3038: out = 24'(-7308);
			3039: out = 24'(-244);
			3040: out = 24'(12564);
			3041: out = 24'(8444);
			3042: out = 24'(2568);
			3043: out = 24'(12580);
			3044: out = 24'(-10628);
			3045: out = 24'(-11940);
			3046: out = 24'(-640);
			3047: out = 24'(11420);
			3048: out = 24'(8060);
			3049: out = 24'(-1512);
			3050: out = 24'(-9516);
			3051: out = 24'(5384);
			3052: out = 24'(14164);
			3053: out = 24'(11100);
			3054: out = 24'(5456);
			3055: out = 24'(-8940);
			3056: out = 24'(-12584);
			3057: out = 24'(2412);
			3058: out = 24'(-316);
			3059: out = 24'(3820);
			3060: out = 24'(7276);
			3061: out = 24'(11736);
			3062: out = 24'(9084);
			3063: out = 24'(4412);
			3064: out = 24'(-5588);
			3065: out = 24'(5812);
			3066: out = 24'(1880);
			3067: out = 24'(-5528);
			3068: out = 24'(-2476);
			3069: out = 24'(1300);
			3070: out = 24'(4892);
			3071: out = 24'(5748);
			3072: out = 24'(1480);
			3073: out = 24'(1316);
			3074: out = 24'(3952);
			3075: out = 24'(13356);
			3076: out = 24'(2436);
			3077: out = 24'(684);
			3078: out = 24'(15976);
			3079: out = 24'(-628);
			3080: out = 24'(-1052);
			3081: out = 24'(236);
			3082: out = 24'(2032);
			3083: out = 24'(1040);
			3084: out = 24'(592);
			3085: out = 24'(476);
			3086: out = 24'(5504);
			3087: out = 24'(11440);
			3088: out = 24'(11600);
			3089: out = 24'(-16908);
			3090: out = 24'(-5108);
			3091: out = 24'(5732);
			3092: out = 24'(12916);
			3093: out = 24'(-16768);
			3094: out = 24'(-17144);
			3095: out = 24'(-5192);
			3096: out = 24'(-7836);
			3097: out = 24'(3280);
			3098: out = 24'(6744);
			3099: out = 24'(7592);
			3100: out = 24'(1324);
			3101: out = 24'(312);
			3102: out = 24'(-424);
			3103: out = 24'(652);
			3104: out = 24'(-5480);
			3105: out = 24'(-5560);
			3106: out = 24'(1320);
			3107: out = 24'(3860);
			3108: out = 24'(4912);
			3109: out = 24'(1448);
			3110: out = 24'(-3240);
			3111: out = 24'(-3812);
			3112: out = 24'(-5464);
			3113: out = 24'(-11648);
			3114: out = 24'(7912);
			3115: out = 24'(2392);
			3116: out = 24'(-2524);
			3117: out = 24'(776);
			3118: out = 24'(2808);
			3119: out = 24'(-5416);
			3120: out = 24'(-18692);
			3121: out = 24'(4436);
			3122: out = 24'(10992);
			3123: out = 24'(11600);
			3124: out = 24'(7428);
			3125: out = 24'(-2228);
			3126: out = 24'(-6024);
			3127: out = 24'(-3792);
			3128: out = 24'(-4652);
			3129: out = 24'(308);
			3130: out = 24'(5384);
			3131: out = 24'(268);
			3132: out = 24'(8476);
			3133: out = 24'(812);
			3134: out = 24'(-10440);
			3135: out = 24'(-17344);
			3136: out = 24'(-2228);
			3137: out = 24'(9564);
			3138: out = 24'(5036);
			3139: out = 24'(-9700);
			3140: out = 24'(-10060);
			3141: out = 24'(4760);
			3142: out = 24'(9572);
			3143: out = 24'(364);
			3144: out = 24'(-8828);
			3145: out = 24'(13348);
			3146: out = 24'(-17732);
			3147: out = 24'(-14116);
			3148: out = 24'(3304);
			3149: out = 24'(11232);
			3150: out = 24'(7760);
			3151: out = 24'(-292);
			3152: out = 24'(-2468);
			3153: out = 24'(-308);
			3154: out = 24'(1148);
			3155: out = 24'(-3908);
			3156: out = 24'(2020);
			3157: out = 24'(-7828);
			3158: out = 24'(-5648);
			3159: out = 24'(5288);
			3160: out = 24'(13144);
			3161: out = 24'(-824);
			3162: out = 24'(-21500);
			3163: out = 24'(-12652);
			3164: out = 24'(-4388);
			3165: out = 24'(7060);
			3166: out = 24'(7800);
			3167: out = 24'(-92);
			3168: out = 24'(-7492);
			3169: out = 24'(-5092);
			3170: out = 24'(-912);
			3171: out = 24'(6572);
			3172: out = 24'(1396);
			3173: out = 24'(-11996);
			3174: out = 24'(-8428);
			3175: out = 24'(-228);
			3176: out = 24'(7268);
			3177: out = 24'(2148);
			3178: out = 24'(2244);
			3179: out = 24'(-3472);
			3180: out = 24'(-13184);
			3181: out = 24'(6304);
			3182: out = 24'(9300);
			3183: out = 24'(5860);
			3184: out = 24'(172);
			3185: out = 24'(1304);
			3186: out = 24'(5172);
			3187: out = 24'(10368);
			3188: out = 24'(-20300);
			3189: out = 24'(-18404);
			3190: out = 24'(-516);
			3191: out = 24'(9672);
			3192: out = 24'(15340);
			3193: out = 24'(9432);
			3194: out = 24'(1120);
			3195: out = 24'(-16012);
			3196: out = 24'(-10508);
			3197: out = 24'(2196);
			3198: out = 24'(-2856);
			3199: out = 24'(10940);
			3200: out = 24'(10216);
			3201: out = 24'(5080);
			3202: out = 24'(-8864);
			3203: out = 24'(332);
			3204: out = 24'(9356);
			3205: out = 24'(-376);
			3206: out = 24'(-5548);
			3207: out = 24'(-6232);
			3208: out = 24'(4956);
			3209: out = 24'(4876);
			3210: out = 24'(8184);
			3211: out = 24'(960);
			3212: out = 24'(-8408);
			3213: out = 24'(-15844);
			3214: out = 24'(-7856);
			3215: out = 24'(4768);
			3216: out = 24'(12392);
			3217: out = 24'(-5572);
			3218: out = 24'(-21524);
			3219: out = 24'(-1460);
			3220: out = 24'(-12448);
			3221: out = 24'(-516);
			3222: out = 24'(12032);
			3223: out = 24'(8356);
			3224: out = 24'(-2204);
			3225: out = 24'(-5584);
			3226: out = 24'(9972);
			3227: out = 24'(-2616);
			3228: out = 24'(-4916);
			3229: out = 24'(-492);
			3230: out = 24'(5960);
			3231: out = 24'(7540);
			3232: out = 24'(276);
			3233: out = 24'(-10400);
			3234: out = 24'(-13416);
			3235: out = 24'(-2400);
			3236: out = 24'(12056);
			3237: out = 24'(14232);
			3238: out = 24'(6136);
			3239: out = 24'(-7688);
			3240: out = 24'(-21260);
			3241: out = 24'(-9028);
			3242: out = 24'(-372);
			3243: out = 24'(5140);
			3244: out = 24'(10156);
			3245: out = 24'(11132);
			3246: out = 24'(3352);
			3247: out = 24'(-10712);
			3248: out = 24'(-8128);
			3249: out = 24'(208);
			3250: out = 24'(7920);
			3251: out = 24'(14900);
			3252: out = 24'(-876);
			3253: out = 24'(-8272);
			3254: out = 24'(2176);
			3255: out = 24'(1200);
			3256: out = 24'(-2184);
			3257: out = 24'(-6480);
			3258: out = 24'(12080);
			3259: out = 24'(5964);
			3260: out = 24'(-1964);
			3261: out = 24'(-12372);
			3262: out = 24'(1576);
			3263: out = 24'(9252);
			3264: out = 24'(8820);
			3265: out = 24'(-11352);
			3266: out = 24'(-10052);
			3267: out = 24'(-6624);
			3268: out = 24'(-4688);
			3269: out = 24'(1496);
			3270: out = 24'(-1932);
			3271: out = 24'(-3752);
			3272: out = 24'(10008);
			3273: out = 24'(8876);
			3274: out = 24'(3164);
			3275: out = 24'(-8420);
			3276: out = 24'(3052);
			3277: out = 24'(2360);
			3278: out = 24'(352);
			3279: out = 24'(1064);
			3280: out = 24'(-972);
			3281: out = 24'(-1568);
			3282: out = 24'(-60);
			3283: out = 24'(8568);
			3284: out = 24'(7732);
			3285: out = 24'(1492);
			3286: out = 24'(-1748);
			3287: out = 24'(-5488);
			3288: out = 24'(-1444);
			3289: out = 24'(4140);
			3290: out = 24'(2588);
			3291: out = 24'(-560);
			3292: out = 24'(-1132);
			3293: out = 24'(1708);
			3294: out = 24'(3532);
			3295: out = 24'(1168);
			3296: out = 24'(-804);
			3297: out = 24'(-1056);
			3298: out = 24'(7972);
			3299: out = 24'(7252);
			3300: out = 24'(-18280);
			3301: out = 24'(-13712);
			3302: out = 24'(-4464);
			3303: out = 24'(6120);
			3304: out = 24'(1836);
			3305: out = 24'(-7128);
			3306: out = 24'(-12688);
			3307: out = 24'(3256);
			3308: out = 24'(4);
			3309: out = 24'(1576);
			3310: out = 24'(-2304);
			3311: out = 24'(-116);
			3312: out = 24'(-13008);
			3313: out = 24'(-13832);
			3314: out = 24'(12300);
			3315: out = 24'(4004);
			3316: out = 24'(4872);
			3317: out = 24'(6072);
			3318: out = 24'(-12088);
			3319: out = 24'(-10724);
			3320: out = 24'(-3900);
			3321: out = 24'(8);
			3322: out = 24'(7924);
			3323: out = 24'(3400);
			3324: out = 24'(-7076);
			3325: out = 24'(7400);
			3326: out = 24'(-1596);
			3327: out = 24'(-6280);
			3328: out = 24'(-3776);
			3329: out = 24'(8328);
			3330: out = 24'(6604);
			3331: out = 24'(-5660);
			3332: out = 24'(-4868);
			3333: out = 24'(-10172);
			3334: out = 24'(-4200);
			3335: out = 24'(8668);
			3336: out = 24'(6656);
			3337: out = 24'(3108);
			3338: out = 24'(-564);
			3339: out = 24'(-6660);
			3340: out = 24'(-1604);
			3341: out = 24'(4156);
			3342: out = 24'(6588);
			3343: out = 24'(4776);
			3344: out = 24'(-268);
			3345: out = 24'(-5516);
			3346: out = 24'(3448);
			3347: out = 24'(-4176);
			3348: out = 24'(-5104);
			3349: out = 24'(1684);
			3350: out = 24'(3984);
			3351: out = 24'(3232);
			3352: out = 24'(1756);
			3353: out = 24'(3340);
			3354: out = 24'(4032);
			3355: out = 24'(-1364);
			3356: out = 24'(-11004);
			3357: out = 24'(-18132);
			3358: out = 24'(-4180);
			3359: out = 24'(14376);
			3360: out = 24'(-6828);
			3361: out = 24'(8368);
			3362: out = 24'(5688);
			3363: out = 24'(-6608);
			3364: out = 24'(-10772);
			3365: out = 24'(-1036);
			3366: out = 24'(9132);
			3367: out = 24'(-10816);
			3368: out = 24'(2004);
			3369: out = 24'(4668);
			3370: out = 24'(308);
			3371: out = 24'(-8432);
			3372: out = 24'(-8456);
			3373: out = 24'(-3012);
			3374: out = 24'(2700);
			3375: out = 24'(1836);
			3376: out = 24'(708);
			3377: out = 24'(2652);
			3378: out = 24'(2428);
			3379: out = 24'(2980);
			3380: out = 24'(2200);
			3381: out = 24'(7124);
			3382: out = 24'(-5452);
			3383: out = 24'(-5448);
			3384: out = 24'(7780);
			3385: out = 24'(11752);
			3386: out = 24'(8836);
			3387: out = 24'(-484);
			3388: out = 24'(12068);
			3389: out = 24'(-19392);
			3390: out = 24'(-17776);
			3391: out = 24'(6736);
			3392: out = 24'(6768);
			3393: out = 24'(2388);
			3394: out = 24'(-5448);
			3395: out = 24'(980);
			3396: out = 24'(4184);
			3397: out = 24'(6748);
			3398: out = 24'(-876);
			3399: out = 24'(-1680);
			3400: out = 24'(-10416);
			3401: out = 24'(-6664);
			3402: out = 24'(9052);
			3403: out = 24'(9340);
			3404: out = 24'(5216);
			3405: out = 24'(2076);
			3406: out = 24'(-4324);
			3407: out = 24'(3760);
			3408: out = 24'(5796);
			3409: out = 24'(-4084);
			3410: out = 24'(-9952);
			3411: out = 24'(-3392);
			3412: out = 24'(11468);
			3413: out = 24'(7052);
			3414: out = 24'(2144);
			3415: out = 24'(-5940);
			3416: out = 24'(-348);
			3417: out = 24'(-9896);
			3418: out = 24'(-2028);
			3419: out = 24'(7612);
			3420: out = 24'(6040);
			3421: out = 24'(1440);
			3422: out = 24'(-3000);
			3423: out = 24'(-4296);
			3424: out = 24'(-3848);
			3425: out = 24'(-1864);
			3426: out = 24'(1268);
			3427: out = 24'(-6616);
			3428: out = 24'(4312);
			3429: out = 24'(7696);
			3430: out = 24'(-1960);
			3431: out = 24'(-5220);
			3432: out = 24'(-4232);
			3433: out = 24'(2276);
			3434: out = 24'(-3944);
			3435: out = 24'(4316);
			3436: out = 24'(3992);
			3437: out = 24'(-6560);
			3438: out = 24'(7544);
			3439: out = 24'(6112);
			3440: out = 24'(-1796);
			3441: out = 24'(-8332);
			3442: out = 24'(-3476);
			3443: out = 24'(2556);
			3444: out = 24'(-2120);
			3445: out = 24'(10184);
			3446: out = 24'(-736);
			3447: out = 24'(-12076);
			3448: out = 24'(-2416);
			3449: out = 24'(5116);
			3450: out = 24'(7488);
			3451: out = 24'(-3336);
			3452: out = 24'(980);
			3453: out = 24'(-768);
			3454: out = 24'(740);
			3455: out = 24'(-9668);
			3456: out = 24'(4248);
			3457: out = 24'(7380);
			3458: out = 24'(5096);
			3459: out = 24'(-6824);
			3460: out = 24'(-560);
			3461: out = 24'(5360);
			3462: out = 24'(-3588);
			3463: out = 24'(-6892);
			3464: out = 24'(-3108);
			3465: out = 24'(5260);
			3466: out = 24'(4812);
			3467: out = 24'(-6620);
			3468: out = 24'(-17780);
			3469: out = 24'(-16440);
			3470: out = 24'(4488);
			3471: out = 24'(14228);
			3472: out = 24'(5148);
			3473: out = 24'(7636);
			3474: out = 24'(4260);
			3475: out = 24'(3828);
			3476: out = 24'(-7612);
			3477: out = 24'(-360);
			3478: out = 24'(884);
			3479: out = 24'(1304);
			3480: out = 24'(-4932);
			3481: out = 24'(120);
			3482: out = 24'(6716);
			3483: out = 24'(12480);
			3484: out = 24'(-492);
			3485: out = 24'(-5792);
			3486: out = 24'(316);
			3487: out = 24'(-2000);
			3488: out = 24'(6764);
			3489: out = 24'(8040);
			3490: out = 24'(988);
			3491: out = 24'(-2344);
			3492: out = 24'(1612);
			3493: out = 24'(8200);
			3494: out = 24'(-856);
			3495: out = 24'(-2432);
			3496: out = 24'(-2440);
			3497: out = 24'(-2700);
			3498: out = 24'(5216);
			3499: out = 24'(5612);
			3500: out = 24'(1004);
			3501: out = 24'(-6908);
			3502: out = 24'(-1020);
			3503: out = 24'(6444);
			3504: out = 24'(4148);
			3505: out = 24'(-120);
			3506: out = 24'(-2728);
			3507: out = 24'(2576);
			3508: out = 24'(-6956);
			3509: out = 24'(4052);
			3510: out = 24'(6272);
			3511: out = 24'(1076);
			3512: out = 24'(-12272);
			3513: out = 24'(-11012);
			3514: out = 24'(-376);
			3515: out = 24'(7108);
			3516: out = 24'(3928);
			3517: out = 24'(-268);
			3518: out = 24'(964);
			3519: out = 24'(1024);
			3520: out = 24'(-124);
			3521: out = 24'(-1616);
			3522: out = 24'(1936);
			3523: out = 24'(5556);
			3524: out = 24'(6336);
			3525: out = 24'(4072);
			3526: out = 24'(-11436);
			3527: out = 24'(-12884);
			3528: out = 24'(-2952);
			3529: out = 24'(7612);
			3530: out = 24'(8156);
			3531: out = 24'(1128);
			3532: out = 24'(-11080);
			3533: out = 24'(736);
			3534: out = 24'(-3932);
			3535: out = 24'(-11488);
			3536: out = 24'(5164);
			3537: out = 24'(3212);
			3538: out = 24'(1444);
			3539: out = 24'(-4424);
			3540: out = 24'(3564);
			3541: out = 24'(1224);
			3542: out = 24'(-1348);
			3543: out = 24'(6936);
			3544: out = 24'(2348);
			3545: out = 24'(-976);
			3546: out = 24'(-4032);
			3547: out = 24'(4524);
			3548: out = 24'(-184);
			3549: out = 24'(-6908);
			3550: out = 24'(4400);
			3551: out = 24'(-368);
			3552: out = 24'(1628);
			3553: out = 24'(6276);
			3554: out = 24'(704);
			3555: out = 24'(-1596);
			3556: out = 24'(-8);
			3557: out = 24'(5284);
			3558: out = 24'(568);
			3559: out = 24'(-11112);
			3560: out = 24'(-24280);
			3561: out = 24'(-11264);
			3562: out = 24'(2660);
			3563: out = 24'(11188);
			3564: out = 24'(2480);
			3565: out = 24'(-1168);
			3566: out = 24'(-9244);
			3567: out = 24'(-12568);
			3568: out = 24'(-3844);
			3569: out = 24'(6072);
			3570: out = 24'(7532);
			3571: out = 24'(-2536);
			3572: out = 24'(-8296);
			3573: out = 24'(-8944);
			3574: out = 24'(-3524);
			3575: out = 24'(3204);
			3576: out = 24'(5068);
			3577: out = 24'(1376);
			3578: out = 24'(-8696);
			3579: out = 24'(-3260);
			3580: out = 24'(548);
			3581: out = 24'(860);
			3582: out = 24'(4768);
			3583: out = 24'(-1472);
			3584: out = 24'(-9008);
			3585: out = 24'(-4920);
			3586: out = 24'(-9912);
			3587: out = 24'(-3712);
			3588: out = 24'(3376);
			3589: out = 24'(6568);
			3590: out = 24'(-2216);
			3591: out = 24'(-8316);
			3592: out = 24'(-6772);
			3593: out = 24'(3804);
			3594: out = 24'(2440);
			3595: out = 24'(-6072);
			3596: out = 24'(-1972);
			3597: out = 24'(2996);
			3598: out = 24'(6340);
			3599: out = 24'(4956);
			3600: out = 24'(-5280);
			3601: out = 24'(-2840);
			3602: out = 24'(7564);
			3603: out = 24'(-2488);
			3604: out = 24'(100);
			3605: out = 24'(680);
			3606: out = 24'(-3136);
			3607: out = 24'(5876);
			3608: out = 24'(5052);
			3609: out = 24'(-588);
			3610: out = 24'(-22576);
			3611: out = 24'(-8732);
			3612: out = 24'(4312);
			3613: out = 24'(508);
			3614: out = 24'(4492);
			3615: out = 24'(7548);
			3616: out = 24'(8720);
			3617: out = 24'(-15528);
			3618: out = 24'(-16224);
			3619: out = 24'(-7416);
			3620: out = 24'(7180);
			3621: out = 24'(10304);
			3622: out = 24'(7392);
			3623: out = 24'(-364);
			3624: out = 24'(-16780);
			3625: out = 24'(-7452);
			3626: out = 24'(2912);
			3627: out = 24'(4220);
			3628: out = 24'(-572);
			3629: out = 24'(-400);
			3630: out = 24'(4756);
			3631: out = 24'(3920);
			3632: out = 24'(4984);
			3633: out = 24'(-964);
			3634: out = 24'(-11896);
			3635: out = 24'(5876);
			3636: out = 24'(7156);
			3637: out = 24'(1996);
			3638: out = 24'(-5280);
			3639: out = 24'(-520);
			3640: out = 24'(4956);
			3641: out = 24'(6296);
			3642: out = 24'(3144);
			3643: out = 24'(1096);
			3644: out = 24'(1108);
			3645: out = 24'(6400);
			3646: out = 24'(4368);
			3647: out = 24'(6524);
			3648: out = 24'(8984);
			3649: out = 24'(7980);
			3650: out = 24'(-2060);
			3651: out = 24'(-8548);
			3652: out = 24'(3880);
			3653: out = 24'(3972);
			3654: out = 24'(440);
			3655: out = 24'(-8680);
			3656: out = 24'(2096);
			3657: out = 24'(4772);
			3658: out = 24'(5564);
			3659: out = 24'(-1516);
			3660: out = 24'(3976);
			3661: out = 24'(5616);
			3662: out = 24'(4952);
			3663: out = 24'(-2076);
			3664: out = 24'(-2148);
			3665: out = 24'(1100);
			3666: out = 24'(4800);
			3667: out = 24'(5180);
			3668: out = 24'(3440);
			3669: out = 24'(1348);
			3670: out = 24'(948);
			3671: out = 24'(2544);
			3672: out = 24'(3112);
			3673: out = 24'(-1876);
			3674: out = 24'(3580);
			3675: out = 24'(5580);
			3676: out = 24'(4816);
			3677: out = 24'(-2908);
			3678: out = 24'(-928);
			3679: out = 24'(2620);
			3680: out = 24'(1484);
			3681: out = 24'(960);
			3682: out = 24'(-1704);
			3683: out = 24'(-1600);
			3684: out = 24'(-2112);
			3685: out = 24'(6288);
			3686: out = 24'(8880);
			3687: out = 24'(1216);
			3688: out = 24'(-8864);
			3689: out = 24'(-14712);
			3690: out = 24'(-9448);
			3691: out = 24'(4416);
			3692: out = 24'(7932);
			3693: out = 24'(3572);
			3694: out = 24'(640);
			3695: out = 24'(-7788);
			3696: out = 24'(-4400);
			3697: out = 24'(1996);
			3698: out = 24'(6700);
			3699: out = 24'(2504);
			3700: out = 24'(-2744);
			3701: out = 24'(-10640);
			3702: out = 24'(6944);
			3703: out = 24'(6056);
			3704: out = 24'(-2116);
			3705: out = 24'(-12124);
			3706: out = 24'(-104);
			3707: out = 24'(7780);
			3708: out = 24'(-632);
			3709: out = 24'(-368);
			3710: out = 24'(-4240);
			3711: out = 24'(-3572);
			3712: out = 24'(3620);
			3713: out = 24'(-384);
			3714: out = 24'(-3216);
			3715: out = 24'(384);
			3716: out = 24'(-3824);
			3717: out = 24'(-3732);
			3718: out = 24'(-1796);
			3719: out = 24'(4108);
			3720: out = 24'(3124);
			3721: out = 24'(-664);
			3722: out = 24'(-4636);
			3723: out = 24'(-5284);
			3724: out = 24'(-260);
			3725: out = 24'(2316);
			3726: out = 24'(-6064);
			3727: out = 24'(-9188);
			3728: out = 24'(-4928);
			3729: out = 24'(7000);
			3730: out = 24'(3292);
			3731: out = 24'(1676);
			3732: out = 24'(-1144);
			3733: out = 24'(-268);
			3734: out = 24'(-840);
			3735: out = 24'(-196);
			3736: out = 24'(-280);
			3737: out = 24'(-3740);
			3738: out = 24'(-4160);
			3739: out = 24'(-1372);
			3740: out = 24'(6652);
			3741: out = 24'(-1804);
			3742: out = 24'(-6816);
			3743: out = 24'(-4336);
			3744: out = 24'(-3072);
			3745: out = 24'(1748);
			3746: out = 24'(2940);
			3747: out = 24'(-1372);
			3748: out = 24'(-2044);
			3749: out = 24'(-2500);
			3750: out = 24'(-2272);
			3751: out = 24'(-3944);
			3752: out = 24'(-1580);
			3753: out = 24'(1264);
			3754: out = 24'(116);
			3755: out = 24'(1568);
			3756: out = 24'(1548);
			3757: out = 24'(2372);
			3758: out = 24'(-4340);
			3759: out = 24'(-2800);
			3760: out = 24'(-2696);
			3761: out = 24'(-8744);
			3762: out = 24'(-8020);
			3763: out = 24'(-4660);
			3764: out = 24'(1212);
			3765: out = 24'(7844);
			3766: out = 24'(7580);
			3767: out = 24'(2128);
			3768: out = 24'(-8112);
			3769: out = 24'(-3308);
			3770: out = 24'(-504);
			3771: out = 24'(-1600);
			3772: out = 24'(-4900);
			3773: out = 24'(-2376);
			3774: out = 24'(3664);
			3775: out = 24'(4248);
			3776: out = 24'(6448);
			3777: out = 24'(-580);
			3778: out = 24'(-8120);
			3779: out = 24'(-10936);
			3780: out = 24'(-2608);
			3781: out = 24'(2184);
			3782: out = 24'(-6744);
			3783: out = 24'(-476);
			3784: out = 24'(2380);
			3785: out = 24'(3840);
			3786: out = 24'(-4104);
			3787: out = 24'(-4312);
			3788: out = 24'(-2016);
			3789: out = 24'(3524);
			3790: out = 24'(1376);
			3791: out = 24'(1356);
			3792: out = 24'(1044);
			3793: out = 24'(-3696);
			3794: out = 24'(-1832);
			3795: out = 24'(-380);
			3796: out = 24'(-2872);
			3797: out = 24'(2352);
			3798: out = 24'(2696);
			3799: out = 24'(1676);
			3800: out = 24'(4328);
			3801: out = 24'(3424);
			3802: out = 24'(4624);
			3803: out = 24'(8556);
			3804: out = 24'(-4548);
			3805: out = 24'(-11856);
			3806: out = 24'(-12472);
			3807: out = 24'(1280);
			3808: out = 24'(1528);
			3809: out = 24'(3332);
			3810: out = 24'(8804);
			3811: out = 24'(-1504);
			3812: out = 24'(-5560);
			3813: out = 24'(-5668);
			3814: out = 24'(5184);
			3815: out = 24'(416);
			3816: out = 24'(-460);
			3817: out = 24'(5212);
			3818: out = 24'(824);
			3819: out = 24'(1660);
			3820: out = 24'(2512);
			3821: out = 24'(4004);
			3822: out = 24'(2844);
			3823: out = 24'(2084);
			3824: out = 24'(400);
			3825: out = 24'(4396);
			3826: out = 24'(1804);
			3827: out = 24'(-304);
			3828: out = 24'(4072);
			3829: out = 24'(3768);
			3830: out = 24'(2896);
			3831: out = 24'(368);
			3832: out = 24'(-336);
			3833: out = 24'(-1628);
			3834: out = 24'(-432);
			3835: out = 24'(6320);
			3836: out = 24'(6100);
			3837: out = 24'(3500);
			3838: out = 24'(-3812);
			3839: out = 24'(-468);
			3840: out = 24'(-4980);
			3841: out = 24'(-5268);
			3842: out = 24'(-3028);
			3843: out = 24'(6384);
			3844: out = 24'(5484);
			3845: out = 24'(-316);
			3846: out = 24'(-9752);
			3847: out = 24'(-1312);
			3848: out = 24'(7556);
			3849: out = 24'(5164);
			3850: out = 24'(-4980);
			3851: out = 24'(-5180);
			3852: out = 24'(7604);
			3853: out = 24'(2592);
			3854: out = 24'(3516);
			3855: out = 24'(-100);
			3856: out = 24'(672);
			3857: out = 24'(-296);
			3858: out = 24'(2736);
			3859: out = 24'(2052);
			3860: out = 24'(-1764);
			3861: out = 24'(-7056);
			3862: out = 24'(-4520);
			3863: out = 24'(5948);
			3864: out = 24'(5084);
			3865: out = 24'(2656);
			3866: out = 24'(1312);
			3867: out = 24'(-7428);
			3868: out = 24'(12);
			3869: out = 24'(5588);
			3870: out = 24'(4268);
			3871: out = 24'(-1888);
			3872: out = 24'(-320);
			3873: out = 24'(6248);
			3874: out = 24'(-896);
			3875: out = 24'(76);
			3876: out = 24'(-2740);
			3877: out = 24'(-11268);
			3878: out = 24'(3480);
			3879: out = 24'(8916);
			3880: out = 24'(6140);
			3881: out = 24'(-13632);
			3882: out = 24'(-5812);
			3883: out = 24'(5560);
			3884: out = 24'(5980);
			3885: out = 24'(2460);
			3886: out = 24'(-5380);
			3887: out = 24'(-8708);
			3888: out = 24'(-10072);
			3889: out = 24'(-1632);
			3890: out = 24'(3152);
			3891: out = 24'(1656);
			3892: out = 24'(192);
			3893: out = 24'(-1580);
			3894: out = 24'(-1660);
			3895: out = 24'(-24);
			3896: out = 24'(-20);
			3897: out = 24'(532);
			3898: out = 24'(2680);
			3899: out = 24'(-1876);
			3900: out = 24'(-2052);
			3901: out = 24'(-496);
			3902: out = 24'(268);
			3903: out = 24'(1020);
			3904: out = 24'(-240);
			3905: out = 24'(-3104);
			3906: out = 24'(-144);
			3907: out = 24'(1588);
			3908: out = 24'(2632);
			3909: out = 24'(1960);
			3910: out = 24'(748);
			3911: out = 24'(-1284);
			3912: out = 24'(-2404);
			3913: out = 24'(-2332);
			3914: out = 24'(-548);
			3915: out = 24'(524);
			3916: out = 24'(548);
			3917: out = 24'(-2212);
			3918: out = 24'(-3780);
			3919: out = 24'(-2936);
			3920: out = 24'(372);
			3921: out = 24'(1408);
			3922: out = 24'(212);
			3923: out = 24'(-2780);
			3924: out = 24'(-672);
			3925: out = 24'(1216);
			3926: out = 24'(1048);
			3927: out = 24'(-792);
			3928: out = 24'(-2416);
			3929: out = 24'(-2528);
			3930: out = 24'(-1768);
			3931: out = 24'(1488);
			3932: out = 24'(2772);
			3933: out = 24'(1564);
			3934: out = 24'(4064);
			3935: out = 24'(1572);
			3936: out = 24'(-2116);
			3937: out = 24'(-6544);
			3938: out = 24'(-5052);
			3939: out = 24'(-2408);
			3940: out = 24'(656);
			3941: out = 24'(-2896);
			3942: out = 24'(1760);
			3943: out = 24'(4104);
			3944: out = 24'(-3416);
			3945: out = 24'(-3720);
			3946: out = 24'(-4392);
			3947: out = 24'(-1416);
			3948: out = 24'(-9048);
			3949: out = 24'(-1908);
			3950: out = 24'(3632);
			3951: out = 24'(5340);
			3952: out = 24'(-5200);
			3953: out = 24'(-8104);
			3954: out = 24'(-2176);
			3955: out = 24'(5908);
			3956: out = 24'(3972);
			3957: out = 24'(-3484);
			3958: out = 24'(-9056);
			3959: out = 24'(-7036);
			3960: out = 24'(128);
			3961: out = 24'(5296);
			3962: out = 24'(2244);
			3963: out = 24'(-1164);
			3964: out = 24'(-4620);
			3965: out = 24'(-5940);
			3966: out = 24'(668);
			3967: out = 24'(5160);
			3968: out = 24'(4608);
			3969: out = 24'(1708);
			3970: out = 24'(-4236);
			3971: out = 24'(-5120);
			3972: out = 24'(868);
			3973: out = 24'(1452);
			3974: out = 24'(-76);
			3975: out = 24'(-2752);
			3976: out = 24'(3712);
			3977: out = 24'(3184);
			3978: out = 24'(3696);
			3979: out = 24'(3292);
			3980: out = 24'(1668);
			3981: out = 24'(216);
			3982: out = 24'(-992);
			3983: out = 24'(-14320);
			3984: out = 24'(-3524);
			3985: out = 24'(5336);
			3986: out = 24'(4260);
			3987: out = 24'(3632);
			3988: out = 24'(-1220);
			3989: out = 24'(-3880);
			3990: out = 24'(-2576);
			3991: out = 24'(1524);
			3992: out = 24'(3340);
			3993: out = 24'(340);
			3994: out = 24'(1624);
			3995: out = 24'(-208);
			3996: out = 24'(-380);
			3997: out = 24'(-1212);
			3998: out = 24'(2220);
			3999: out = 24'(2392);
			4000: out = 24'(2388);
			4001: out = 24'(-3992);
			4002: out = 24'(1364);
			4003: out = 24'(6824);
			4004: out = 24'(3860);
			4005: out = 24'(-1424);
			4006: out = 24'(-2304);
			4007: out = 24'(3732);
			4008: out = 24'(3248);
			4009: out = 24'(820);
			4010: out = 24'(-3068);
			4011: out = 24'(-1072);
			4012: out = 24'(1684);
			4013: out = 24'(3936);
			4014: out = 24'(2072);
			4015: out = 24'(1112);
			4016: out = 24'(-296);
			4017: out = 24'(844);
			4018: out = 24'(3060);
			4019: out = 24'(1220);
			4020: out = 24'(-1208);
			4021: out = 24'(-1504);
			4022: out = 24'(-3028);
			4023: out = 24'(-2404);
			4024: out = 24'(-716);
			4025: out = 24'(7004);
			4026: out = 24'(-1232);
			4027: out = 24'(-4904);
			4028: out = 24'(-4016);
			4029: out = 24'(4316);
			4030: out = 24'(3556);
			4031: out = 24'(400);
			4032: out = 24'(1664);
			4033: out = 24'(-952);
			4034: out = 24'(-820);
			4035: out = 24'(44);
			4036: out = 24'(1140);
			4037: out = 24'(72);
			4038: out = 24'(-932);
			4039: out = 24'(680);
			4040: out = 24'(2680);
			4041: out = 24'(4120);
			4042: out = 24'(1536);
			4043: out = 24'(372);
			4044: out = 24'(-7940);
			4045: out = 24'(-8560);
			4046: out = 24'(6128);
			4047: out = 24'(5364);
			4048: out = 24'(3996);
			4049: out = 24'(-652);
			4050: out = 24'(-6368);
			4051: out = 24'(-4364);
			4052: out = 24'(772);
			4053: out = 24'(-528);
			4054: out = 24'(5092);
			4055: out = 24'(1420);
			4056: out = 24'(-3540);
			4057: out = 24'(-1648);
			4058: out = 24'(920);
			4059: out = 24'(2232);
			4060: out = 24'(1380);
			4061: out = 24'(-2568);
			4062: out = 24'(-1060);
			4063: out = 24'(2500);
			4064: out = 24'(-6856);
			4065: out = 24'(-3140);
			4066: out = 24'(1488);
			4067: out = 24'(4288);
			4068: out = 24'(1960);
			4069: out = 24'(-252);
			4070: out = 24'(-1264);
			4071: out = 24'(-5332);
			4072: out = 24'(60);
			4073: out = 24'(3396);
			4074: out = 24'(1768);
			4075: out = 24'(612);
			4076: out = 24'(1108);
			4077: out = 24'(2428);
			4078: out = 24'(-3860);
			4079: out = 24'(-2644);
			4080: out = 24'(-2372);
			4081: out = 24'(-2540);
			4082: out = 24'(468);
			4083: out = 24'(1776);
			4084: out = 24'(1544);
			4085: out = 24'(412);
			4086: out = 24'(128);
			4087: out = 24'(-1364);
			4088: out = 24'(-5320);
			4089: out = 24'(-296);
			4090: out = 24'(1364);
			4091: out = 24'(1692);
			4092: out = 24'(-4832);
			4093: out = 24'(-1148);
			4094: out = 24'(348);
			4095: out = 24'(440);
			4096: out = 24'(-4948);
			4097: out = 24'(-2552);
			4098: out = 24'(708);
			4099: out = 24'(-1632);
			4100: out = 24'(-2692);
			4101: out = 24'(-268);
			4102: out = 24'(5452);
			4103: out = 24'(-876);
			4104: out = 24'(-3944);
			4105: out = 24'(-4900);
			4106: out = 24'(2604);
			4107: out = 24'(768);
			4108: out = 24'(1168);
			4109: out = 24'(1920);
			4110: out = 24'(-684);
			4111: out = 24'(-1932);
			4112: out = 24'(-2560);
			4113: out = 24'(-3088);
			4114: out = 24'(-1780);
			4115: out = 24'(640);
			4116: out = 24'(2484);
			4117: out = 24'(-5444);
			4118: out = 24'(-5684);
			4119: out = 24'(-2388);
			4120: out = 24'(-432);
			4121: out = 24'(4220);
			4122: out = 24'(2432);
			4123: out = 24'(-2312);
			4124: out = 24'(-2316);
			4125: out = 24'(-1352);
			4126: out = 24'(-432);
			4127: out = 24'(-2152);
			4128: out = 24'(124);
			4129: out = 24'(1684);
			4130: out = 24'(2156);
			4131: out = 24'(2908);
			4132: out = 24'(-1276);
			4133: out = 24'(-4088);
			4134: out = 24'(-1060);
			4135: out = 24'(2912);
			4136: out = 24'(5468);
			4137: out = 24'(4208);
			4138: out = 24'(6036);
			4139: out = 24'(2036);
			4140: out = 24'(-1056);
			4141: out = 24'(-4164);
			4142: out = 24'(1124);
			4143: out = 24'(1776);
			4144: out = 24'(232);
			4145: out = 24'(844);
			4146: out = 24'(2096);
			4147: out = 24'(2700);
			4148: out = 24'(648);
			4149: out = 24'(504);
			4150: out = 24'(-1364);
			4151: out = 24'(-2588);
			4152: out = 24'(-44);
			4153: out = 24'(1500);
			4154: out = 24'(1608);
			4155: out = 24'(-2484);
			4156: out = 24'(3132);
			4157: out = 24'(2240);
			4158: out = 24'(292);
			4159: out = 24'(-1892);
			4160: out = 24'(3208);
			4161: out = 24'(4660);
			4162: out = 24'(-504);
			4163: out = 24'(1476);
			4164: out = 24'(1464);
			4165: out = 24'(1700);
			4166: out = 24'(2136);
			4167: out = 24'(452);
			4168: out = 24'(-892);
			4169: out = 24'(-1092);
			4170: out = 24'(1424);
			4171: out = 24'(1764);
			4172: out = 24'(1500);
			4173: out = 24'(988);
			4174: out = 24'(1780);
			4175: out = 24'(1208);
			4176: out = 24'(676);
			4177: out = 24'(-8040);
			4178: out = 24'(-6108);
			4179: out = 24'(652);
			4180: out = 24'(5344);
			4181: out = 24'(3836);
			4182: out = 24'(1208);
			4183: out = 24'(-832);
			4184: out = 24'(532);
			4185: out = 24'(-4692);
			4186: out = 24'(-9024);
			4187: out = 24'(1936);
			4188: out = 24'(2652);
			4189: out = 24'(4980);
			4190: out = 24'(3744);
			4191: out = 24'(2284);
			4192: out = 24'(-3108);
			4193: out = 24'(-5208);
			4194: out = 24'(-688);
			4195: out = 24'(1372);
			4196: out = 24'(-216);
			4197: out = 24'(-5112);
			4198: out = 24'(-744);
			4199: out = 24'(1276);
			4200: out = 24'(1984);
			4201: out = 24'(-4832);
			4202: out = 24'(420);
			4203: out = 24'(2216);
			4204: out = 24'(2076);
			4205: out = 24'(-3100);
			4206: out = 24'(-1888);
			4207: out = 24'(-256);
			4208: out = 24'(-1500);
			4209: out = 24'(-2528);
			4210: out = 24'(-752);
			4211: out = 24'(2812);
			4212: out = 24'(-3352);
			4213: out = 24'(-3128);
			4214: out = 24'(-1168);
			4215: out = 24'(892);
			4216: out = 24'(612);
			4217: out = 24'(-1512);
			4218: out = 24'(-2988);
			4219: out = 24'(-1464);
			4220: out = 24'(908);
			4221: out = 24'(176);
			4222: out = 24'(-3756);
			4223: out = 24'(-4452);
			4224: out = 24'(-1168);
			4225: out = 24'(2296);
			4226: out = 24'(3376);
			4227: out = 24'(-1968);
			4228: out = 24'(-4208);
			4229: out = 24'(856);
			4230: out = 24'(2428);
			4231: out = 24'(-1404);
			4232: out = 24'(-7876);
			4233: out = 24'(-1352);
			4234: out = 24'(1888);
			4235: out = 24'(3020);
			4236: out = 24'(-1220);
			4237: out = 24'(-2768);
			4238: out = 24'(-2348);
			4239: out = 24'(588);
			4240: out = 24'(112);
			4241: out = 24'(-520);
			4242: out = 24'(-188);
			4243: out = 24'(3568);
			4244: out = 24'(1648);
			4245: out = 24'(-436);
			4246: out = 24'(-2616);
			4247: out = 24'(984);
			4248: out = 24'(1780);
			4249: out = 24'(1688);
			4250: out = 24'(-220);
			4251: out = 24'(920);
			4252: out = 24'(2356);
			4253: out = 24'(2804);
			4254: out = 24'(-4996);
			4255: out = 24'(-4972);
			4256: out = 24'(-2412);
			4257: out = 24'(2536);
			4258: out = 24'(48);
			4259: out = 24'(-84);
			4260: out = 24'(420);
			4261: out = 24'(4588);
			4262: out = 24'(640);
			4263: out = 24'(-1408);
			4264: out = 24'(868);
			4265: out = 24'(-4588);
			4266: out = 24'(-3872);
			4267: out = 24'(-1020);
			4268: out = 24'(24);
			4269: out = 24'(2700);
			4270: out = 24'(3528);
			4271: out = 24'(2060);
			4272: out = 24'(1184);
			4273: out = 24'(-2736);
			4274: out = 24'(-6044);
			4275: out = 24'(-1940);
			4276: out = 24'(-2732);
			4277: out = 24'(-1312);
			4278: out = 24'(832);
			4279: out = 24'(2128);
			4280: out = 24'(444);
			4281: out = 24'(-2036);
			4282: out = 24'(-1944);
			4283: out = 24'(-888);
			4284: out = 24'(708);
			4285: out = 24'(904);
			4286: out = 24'(2728);
			4287: out = 24'(680);
			4288: out = 24'(-416);
			4289: out = 24'(3224);
			4290: out = 24'(1668);
			4291: out = 24'(-80);
			4292: out = 24'(-2284);
			4293: out = 24'(3012);
			4294: out = 24'(3064);
			4295: out = 24'(1300);
			4296: out = 24'(-3184);
			4297: out = 24'(280);
			4298: out = 24'(2420);
			4299: out = 24'(2336);
			4300: out = 24'(-3188);
			4301: out = 24'(-3484);
			4302: out = 24'(-1760);
			4303: out = 24'(-1808);
			4304: out = 24'(1596);
			4305: out = 24'(1772);
			4306: out = 24'(-476);
			4307: out = 24'(2544);
			4308: out = 24'(220);
			4309: out = 24'(-1984);
			4310: out = 24'(-3512);
			4311: out = 24'(288);
			4312: out = 24'(1140);
			4313: out = 24'(-548);
			4314: out = 24'(-1504);
			4315: out = 24'(556);
			4316: out = 24'(2536);
			4317: out = 24'(-888);
			4318: out = 24'(2020);
			4319: out = 24'(1172);
			4320: out = 24'(-776);
			4321: out = 24'(-9676);
			4322: out = 24'(-5788);
			4323: out = 24'(1372);
			4324: out = 24'(4400);
			4325: out = 24'(3760);
			4326: out = 24'(-36);
			4327: out = 24'(-2604);
			4328: out = 24'(-1476);
			4329: out = 24'(764);
			4330: out = 24'(1504);
			4331: out = 24'(808);
			4332: out = 24'(-1632);
			4333: out = 24'(-608);
			4334: out = 24'(1036);
			4335: out = 24'(-5308);
			4336: out = 24'(-5724);
			4337: out = 24'(-3496);
			4338: out = 24'(1276);
			4339: out = 24'(2208);
			4340: out = 24'(2428);
			4341: out = 24'(1448);
			4342: out = 24'(-2356);
			4343: out = 24'(-876);
			4344: out = 24'(-496);
			4345: out = 24'(-3460);
			4346: out = 24'(-2352);
			4347: out = 24'(-1332);
			4348: out = 24'(988);
			4349: out = 24'(1168);
			4350: out = 24'(2872);
			4351: out = 24'(2200);
			4352: out = 24'(76);
			4353: out = 24'(-748);
			4354: out = 24'(-1756);
			4355: out = 24'(-2240);
			4356: out = 24'(128);
			4357: out = 24'(-1116);
			4358: out = 24'(-1512);
			4359: out = 24'(-476);
			4360: out = 24'(104);
			4361: out = 24'(244);
			4362: out = 24'(-76);
			4363: out = 24'(364);
			4364: out = 24'(-40);
			4365: out = 24'(80);
			4366: out = 24'(236);
			4367: out = 24'(24);
			4368: out = 24'(-524);
			4369: out = 24'(-836);
			4370: out = 24'(1084);
			4371: out = 24'(-464);
			4372: out = 24'(-864);
			4373: out = 24'(188);
			4374: out = 24'(716);
			4375: out = 24'(508);
			4376: out = 24'(256);
			4377: out = 24'(4124);
			4378: out = 24'(-1072);
			4379: out = 24'(-2672);
			4380: out = 24'(-584);
			4381: out = 24'(-420);
			4382: out = 24'(716);
			4383: out = 24'(552);
			4384: out = 24'(-760);
			4385: out = 24'(240);
			4386: out = 24'(-620);
			4387: out = 24'(-4096);
			4388: out = 24'(2892);
			4389: out = 24'(-544);
			4390: out = 24'(-3580);
			4391: out = 24'(-616);
			4392: out = 24'(1552);
			4393: out = 24'(2872);
			4394: out = 24'(1104);
			4395: out = 24'(2952);
			4396: out = 24'(-1408);
			4397: out = 24'(-3768);
			4398: out = 24'(252);
			4399: out = 24'(1176);
			4400: out = 24'(2556);
			4401: out = 24'(2544);
			4402: out = 24'(1480);
			4403: out = 24'(392);
			4404: out = 24'(-908);
			4405: out = 24'(-5508);
			4406: out = 24'(364);
			4407: out = 24'(1892);
			4408: out = 24'(836);
			4409: out = 24'(-932);
			4410: out = 24'(120);
			4411: out = 24'(1420);
			4412: out = 24'(980);
			4413: out = 24'(-848);
			4414: out = 24'(-684);
			4415: out = 24'(1496);
			4416: out = 24'(-288);
			4417: out = 24'(-420);
			4418: out = 24'(-1224);
			4419: out = 24'(896);
			4420: out = 24'(-680);
			4421: out = 24'(2040);
			4422: out = 24'(3484);
			4423: out = 24'(-932);
			4424: out = 24'(-4348);
			4425: out = 24'(-4800);
			4426: out = 24'(-1852);
			4427: out = 24'(684);
			4428: out = 24'(1144);
			4429: out = 24'(652);
			4430: out = 24'(-3868);
			4431: out = 24'(936);
			4432: out = 24'(2628);
			4433: out = 24'(-1224);
			4434: out = 24'(-3980);
			4435: out = 24'(-2672);
			4436: out = 24'(1644);
			4437: out = 24'(1344);
			4438: out = 24'(-424);
			4439: out = 24'(-2704);
			4440: out = 24'(-1060);
			4441: out = 24'(-512);
			4442: out = 24'(1116);
			4443: out = 24'(1308);
			4444: out = 24'(1076);
			4445: out = 24'(-288);
			4446: out = 24'(-244);
			4447: out = 24'(1616);
			4448: out = 24'(-1652);
			4449: out = 24'(-492);
			4450: out = 24'(1732);
			4451: out = 24'(224);
			4452: out = 24'(92);
			4453: out = 24'(348);
			4454: out = 24'(2888);
			4455: out = 24'(-708);
			4456: out = 24'(-1976);
			4457: out = 24'(-2672);
			4458: out = 24'(2264);
			4459: out = 24'(-804);
			4460: out = 24'(-352);
			4461: out = 24'(1836);
			4462: out = 24'(4204);
			4463: out = 24'(-816);
			4464: out = 24'(-5704);
			4465: out = 24'(2052);
			4466: out = 24'(224);
			4467: out = 24'(-948);
			4468: out = 24'(-3776);
			4469: out = 24'(2208);
			4470: out = 24'(1828);
			4471: out = 24'(196);
			4472: out = 24'(-1304);
			4473: out = 24'(-748);
			4474: out = 24'(276);
			4475: out = 24'(712);
			4476: out = 24'(248);
			4477: out = 24'(-644);
			4478: out = 24'(-1072);
			4479: out = 24'(-856);
			4480: out = 24'(368);
			4481: out = 24'(916);
			4482: out = 24'(560);
			4483: out = 24'(-2844);
			4484: out = 24'(-1516);
			4485: out = 24'(284);
			4486: out = 24'(-4740);
			4487: out = 24'(-332);
			4488: out = 24'(-976);
			4489: out = 24'(-4332);
			4490: out = 24'(636);
			4491: out = 24'(2448);
			4492: out = 24'(2484);
			4493: out = 24'(-2600);
			4494: out = 24'(152);
			4495: out = 24'(676);
			4496: out = 24'(-196);
			4497: out = 24'(-5368);
			4498: out = 24'(-3492);
			4499: out = 24'(512);
			4500: out = 24'(1688);
			4501: out = 24'(2504);
			4502: out = 24'(148);
			4503: out = 24'(-2172);
			4504: out = 24'(-88);
			4505: out = 24'(1344);
			4506: out = 24'(1308);
			4507: out = 24'(-808);
			4508: out = 24'(-84);
			4509: out = 24'(784);
			4510: out = 24'(1384);
			4511: out = 24'(164);
			4512: out = 24'(-2904);
			4513: out = 24'(-4084);
			4514: out = 24'(1904);
			4515: out = 24'(-3496);
			4516: out = 24'(-1340);
			4517: out = 24'(2560);
			4518: out = 24'(-1236);
			4519: out = 24'(-1012);
			4520: out = 24'(-248);
			4521: out = 24'(2164);
			4522: out = 24'(-2600);
			4523: out = 24'(-4640);
			4524: out = 24'(-3524);
			4525: out = 24'(2176);
			4526: out = 24'(2992);
			4527: out = 24'(1048);
			4528: out = 24'(-2900);
			4529: out = 24'(-2728);
			4530: out = 24'(-2260);
			4531: out = 24'(-1060);
			4532: out = 24'(2316);
			4533: out = 24'(1140);
			4534: out = 24'(-1060);
			4535: out = 24'(-3740);
			4536: out = 24'(-1968);
			4537: out = 24'(-1452);
			4538: out = 24'(-1656);
			4539: out = 24'(-2876);
			4540: out = 24'(-392);
			4541: out = 24'(1656);
			4542: out = 24'(1952);
			4543: out = 24'(880);
			4544: out = 24'(-440);
			4545: out = 24'(-1360);
			4546: out = 24'(-764);
			4547: out = 24'(-1812);
			4548: out = 24'(-1576);
			4549: out = 24'(-24);
			4550: out = 24'(1760);
			4551: out = 24'(1872);
			4552: out = 24'(1272);
			4553: out = 24'(1788);
			4554: out = 24'(1172);
			4555: out = 24'(-568);
			4556: out = 24'(-3664);
			4557: out = 24'(-232);
			4558: out = 24'(1448);
			4559: out = 24'(2496);
			4560: out = 24'(952);
			4561: out = 24'(2088);
			4562: out = 24'(1476);
			4563: out = 24'(492);
			4564: out = 24'(-1824);
			4565: out = 24'(-388);
			4566: out = 24'(1564);
			4567: out = 24'(1656);
			4568: out = 24'(604);
			4569: out = 24'(-556);
			4570: out = 24'(-820);
			4571: out = 24'(-912);
			4572: out = 24'(-220);
			4573: out = 24'(636);
			4574: out = 24'(680);
			4575: out = 24'(684);
			4576: out = 24'(-704);
			4577: out = 24'(-1508);
			4578: out = 24'(188);
			4579: out = 24'(1804);
			4580: out = 24'(1776);
			4581: out = 24'(1472);
			4582: out = 24'(-2584);
			4583: out = 24'(-1340);
			4584: out = 24'(3108);
			4585: out = 24'(1404);
			4586: out = 24'(652);
			4587: out = 24'(-908);
			4588: out = 24'(-732);
			4589: out = 24'(-16);
			4590: out = 24'(752);
			4591: out = 24'(416);
			4592: out = 24'(-272);
			4593: out = 24'(-348);
			4594: out = 24'(-252);
			4595: out = 24'(-1276);
			4596: out = 24'(-96);
			4597: out = 24'(800);
			4598: out = 24'(1536);
			4599: out = 24'(-1956);
			4600: out = 24'(-320);
			4601: out = 24'(1236);
			4602: out = 24'(1296);
			4603: out = 24'(400);
			4604: out = 24'(-248);
			4605: out = 24'(-144);
			4606: out = 24'(-1888);
			4607: out = 24'(156);
			4608: out = 24'(1184);
			4609: out = 24'(-336);
			4610: out = 24'(1032);
			4611: out = 24'(984);
			4612: out = 24'(628);
			4613: out = 24'(276);
			4614: out = 24'(-236);
			4615: out = 24'(-664);
			4616: out = 24'(-384);
			4617: out = 24'(-720);
			4618: out = 24'(628);
			4619: out = 24'(2004);
			4620: out = 24'(812);
			4621: out = 24'(136);
			4622: out = 24'(-432);
			4623: out = 24'(420);
			4624: out = 24'(500);
			4625: out = 24'(880);
			4626: out = 24'(100);
			4627: out = 24'(2004);
			4628: out = 24'(-2180);
			4629: out = 24'(-2964);
			4630: out = 24'(228);
			4631: out = 24'(1680);
			4632: out = 24'(-136);
			4633: out = 24'(-3152);
			4634: out = 24'(1896);
			4635: out = 24'(-1232);
			4636: out = 24'(-2188);
			4637: out = 24'(-1732);
			4638: out = 24'(-224);
			4639: out = 24'(-480);
			4640: out = 24'(-824);
			4641: out = 24'(1440);
			4642: out = 24'(464);
			4643: out = 24'(220);
			4644: out = 24'(336);
			4645: out = 24'(-736);
			4646: out = 24'(-1568);
			4647: out = 24'(-1540);
			4648: out = 24'(16);
			4649: out = 24'(708);
			4650: out = 24'(572);
			4651: out = 24'(-384);
			4652: out = 24'(-860);
			4653: out = 24'(-732);
			4654: out = 24'(184);
			4655: out = 24'(932);
			4656: out = 24'(1176);
			4657: out = 24'(220);
			4658: out = 24'(-1168);
			4659: out = 24'(-1264);
			4660: out = 24'(-1060);
			4661: out = 24'(-596);
			4662: out = 24'(-120);
			4663: out = 24'(760);
			4664: out = 24'(1208);
			4665: out = 24'(1104);
			4666: out = 24'(728);
			4667: out = 24'(-596);
			4668: out = 24'(-940);
			4669: out = 24'(1940);
			4670: out = 24'(-632);
			4671: out = 24'(-1500);
			4672: out = 24'(-880);
			4673: out = 24'(-532);
			4674: out = 24'(264);
			4675: out = 24'(876);
			4676: out = 24'(2024);
			4677: out = 24'(-728);
			4678: out = 24'(-2412);
			4679: out = 24'(-2408);
			4680: out = 24'(508);
			4681: out = 24'(984);
			4682: out = 24'(24);
			4683: out = 24'(-1288);
			4684: out = 24'(-1484);
			4685: out = 24'(-696);
			4686: out = 24'(-28);
			4687: out = 24'(-144);
			4688: out = 24'(-748);
			4689: out = 24'(-948);
			4690: out = 24'(-492);
			4691: out = 24'(460);
			4692: out = 24'(252);
			4693: out = 24'(-920);
			4694: out = 24'(-3184);
			4695: out = 24'(-1520);
			4696: out = 24'(1684);
			4697: out = 24'(2920);
			4698: out = 24'(1264);
			4699: out = 24'(-2488);
			4700: out = 24'(-4956);
			4701: out = 24'(-480);
			4702: out = 24'(2056);
			4703: out = 24'(1852);
			4704: out = 24'(-2424);
			4705: out = 24'(-1904);
			4706: out = 24'(-2640);
			4707: out = 24'(-1920);
			4708: out = 24'(2628);
			4709: out = 24'(2488);
			4710: out = 24'(824);
			4711: out = 24'(-912);
			4712: out = 24'(-1068);
			4713: out = 24'(-248);
			4714: out = 24'(672);
			4715: out = 24'(440);
			4716: out = 24'(56);
			4717: out = 24'(-172);
			4718: out = 24'(616);
			4719: out = 24'(-176);
			4720: out = 24'(-28);
			4721: out = 24'(-16);
			4722: out = 24'(1216);
			4723: out = 24'(-704);
			4724: out = 24'(-1284);
			4725: out = 24'(260);
			4726: out = 24'(320);
			4727: out = 24'(-200);
			4728: out = 24'(-1464);
			4729: out = 24'(52);
			4730: out = 24'(-1572);
			4731: out = 24'(-680);
			4732: out = 24'(1556);
			4733: out = 24'(940);
			4734: out = 24'(228);
			4735: out = 24'(-524);
			4736: out = 24'(-1788);
			4737: out = 24'(-908);
			4738: out = 24'(-1360);
			4739: out = 24'(-3020);
			4740: out = 24'(-500);
			4741: out = 24'(1200);
			4742: out = 24'(2004);
			4743: out = 24'(1204);
			4744: out = 24'(-908);
			4745: out = 24'(-2676);
			4746: out = 24'(-3216);
			4747: out = 24'(1332);
			4748: out = 24'(1372);
			4749: out = 24'(-368);
			4750: out = 24'(-1112);
			4751: out = 24'(-1208);
			4752: out = 24'(-20);
			4753: out = 24'(916);
			4754: out = 24'(284);
			4755: out = 24'(-736);
			4756: out = 24'(-1048);
			4757: out = 24'(1780);
			4758: out = 24'(-1100);
			4759: out = 24'(-1744);
			4760: out = 24'(-500);
			4761: out = 24'(1148);
			4762: out = 24'(736);
			4763: out = 24'(264);
			4764: out = 24'(2240);
			4765: out = 24'(-484);
			4766: out = 24'(-1504);
			4767: out = 24'(-1376);
			4768: out = 24'(1404);
			4769: out = 24'(864);
			4770: out = 24'(-332);
			4771: out = 24'(-264);
			4772: out = 24'(-1688);
			4773: out = 24'(-1508);
			4774: out = 24'(-548);
			4775: out = 24'(2212);
			4776: out = 24'(1116);
			4777: out = 24'(300);
			4778: out = 24'(2120);
			4779: out = 24'(-1044);
			4780: out = 24'(-1416);
			4781: out = 24'(-476);
			4782: out = 24'(-3484);
			4783: out = 24'(-1592);
			4784: out = 24'(716);
			4785: out = 24'(2028);
			4786: out = 24'(340);
			4787: out = 24'(-616);
			4788: out = 24'(-564);
			4789: out = 24'(-552);
			4790: out = 24'(76);
			4791: out = 24'(220);
			4792: out = 24'(-184);
			4793: out = 24'(232);
			4794: out = 24'(-28);
			4795: out = 24'(-628);
			4796: out = 24'(-1540);
			4797: out = 24'(-432);
			4798: out = 24'(1176);
			4799: out = 24'(1512);
			4800: out = 24'(652);
			4801: out = 24'(-856);
			4802: out = 24'(-1876);
			4803: out = 24'(-1976);
			4804: out = 24'(256);
			4805: out = 24'(1096);
			4806: out = 24'(-744);
			4807: out = 24'(-760);
			4808: out = 24'(-1548);
			4809: out = 24'(-1100);
			4810: out = 24'(444);
			4811: out = 24'(1716);
			4812: out = 24'(436);
			4813: out = 24'(-3040);
			4814: out = 24'(-612);
			4815: out = 24'(-688);
			4816: out = 24'(-988);
			4817: out = 24'(2276);
			4818: out = 24'(400);
			4819: out = 24'(184);
			4820: out = 24'(1076);
			4821: out = 24'(1384);
			4822: out = 24'(252);
			4823: out = 24'(-640);
			4824: out = 24'(624);
			4825: out = 24'(1028);
			4826: out = 24'(612);
			4827: out = 24'(-432);
			4828: out = 24'(-3104);
			4829: out = 24'(-2040);
			4830: out = 24'(640);
			4831: out = 24'(2364);
			4832: out = 24'(756);
			4833: out = 24'(-1420);
			4834: out = 24'(-2760);
			4835: out = 24'(440);
			4836: out = 24'(0);
			4837: out = 24'(-1208);
			4838: out = 24'(764);
			4839: out = 24'(-1332);
			4840: out = 24'(-1932);
			4841: out = 24'(-1768);
			4842: out = 24'(212);
			4843: out = 24'(548);
			4844: out = 24'(96);
			4845: out = 24'(164);
			4846: out = 24'(-1392);
			4847: out = 24'(-828);
			4848: out = 24'(1256);
			4849: out = 24'(-168);
			4850: out = 24'(-280);
			4851: out = 24'(-48);
			4852: out = 24'(1828);
			4853: out = 24'(-856);
			4854: out = 24'(-820);
			4855: out = 24'(1368);
			4856: out = 24'(-496);
			4857: out = 24'(1372);
			4858: out = 24'(1636);
			4859: out = 24'(-244);
			4860: out = 24'(-2088);
			4861: out = 24'(-1876);
			4862: out = 24'(380);
			4863: out = 24'(-384);
			4864: out = 24'(336);
			4865: out = 24'(252);
			4866: out = 24'(472);
			4867: out = 24'(-132);
			4868: out = 24'(-4);
			4869: out = 24'(32);
			4870: out = 24'(-88);
			4871: out = 24'(-984);
			4872: out = 24'(-868);
			4873: out = 24'(648);
			4874: out = 24'(588);
			4875: out = 24'(408);
			4876: out = 24'(-68);
			4877: out = 24'(1180);
			4878: out = 24'(564);
			4879: out = 24'(-140);
			4880: out = 24'(-1564);
			4881: out = 24'(140);
			4882: out = 24'(-8);
			4883: out = 24'(-904);
			4884: out = 24'(300);
			4885: out = 24'(108);
			4886: out = 24'(-56);
			4887: out = 24'(340);
			4888: out = 24'(-228);
			4889: out = 24'(208);
			4890: out = 24'(800);
			4891: out = 24'(856);
			4892: out = 24'(252);
			4893: out = 24'(-492);
			4894: out = 24'(-1112);
			4895: out = 24'(-180);
			4896: out = 24'(284);
			4897: out = 24'(408);
			4898: out = 24'(176);
			4899: out = 24'(548);
			4900: out = 24'(204);
			4901: out = 24'(-1424);
			4902: out = 24'(436);
			4903: out = 24'(312);
			4904: out = 24'(-436);
			4905: out = 24'(104);
			4906: out = 24'(-872);
			4907: out = 24'(-1116);
			4908: out = 24'(-1096);
			4909: out = 24'(644);
			4910: out = 24'(496);
			4911: out = 24'(-192);
			4912: out = 24'(-1332);
			4913: out = 24'(108);
			4914: out = 24'(648);
			4915: out = 24'(-208);
			4916: out = 24'(-740);
			4917: out = 24'(-96);
			4918: out = 24'(1072);
			4919: out = 24'(-1224);
			4920: out = 24'(120);
			4921: out = 24'(336);
			4922: out = 24'(452);
			4923: out = 24'(308);
			4924: out = 24'(764);
			4925: out = 24'(400);
			4926: out = 24'(-1016);
			4927: out = 24'(-868);
			4928: out = 24'(472);
			4929: out = 24'(1656);
			4930: out = 24'(-100);
			4931: out = 24'(-1024);
			4932: out = 24'(-844);
			4933: out = 24'(-1568);
			4934: out = 24'(1076);
			4935: out = 24'(1436);
			4936: out = 24'(724);
			4937: out = 24'(-3128);
			4938: out = 24'(-2112);
			4939: out = 24'(340);
			4940: out = 24'(1760);
			4941: out = 24'(-1520);
			4942: out = 24'(-2580);
			4943: out = 24'(-276);
			4944: out = 24'(624);
			4945: out = 24'(-260);
			4946: out = 24'(-2344);
			4947: out = 24'(-1192);
			4948: out = 24'(-804);
			4949: out = 24'(672);
			4950: out = 24'(576);
			4951: out = 24'(992);
			4952: out = 24'(-1340);
			4953: out = 24'(-2524);
			4954: out = 24'(-1956);
			4955: out = 24'(464);
			4956: out = 24'(1372);
			4957: out = 24'(696);
			4958: out = 24'(-1336);
			4959: out = 24'(-872);
			4960: out = 24'(372);
			4961: out = 24'(460);
			4962: out = 24'(408);
			4963: out = 24'(-476);
			4964: out = 24'(-980);
			4965: out = 24'(400);
			4966: out = 24'(-240);
			4967: out = 24'(-1512);
			4968: out = 24'(-2524);
			4969: out = 24'(-2592);
			4970: out = 24'(-1312);
			4971: out = 24'(360);
			4972: out = 24'(1240);
			4973: out = 24'(1520);
			4974: out = 24'(1000);
			4975: out = 24'(344);
			4976: out = 24'(-1268);
			4977: out = 24'(-1304);
			4978: out = 24'(32);
			4979: out = 24'(-1188);
			4980: out = 24'(408);
			4981: out = 24'(1140);
			4982: out = 24'(932);
			4983: out = 24'(-1188);
			4984: out = 24'(-1284);
			4985: out = 24'(124);
			4986: out = 24'(708);
			4987: out = 24'(584);
			4988: out = 24'(-188);
			4989: out = 24'(-176);
			4990: out = 24'(-2284);
			4991: out = 24'(-1884);
			4992: out = 24'(-384);
			4993: out = 24'(0);
			default: out = 0;
		endcase
	end
endmodule
