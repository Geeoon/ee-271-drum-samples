module closed_hihat_lookup(index, out);
	input logic unsigned [10:0] index;
	output logic signed [15:0] out;
	always_comb begin
		case(index)
			0: out = 16'(0);
			1: out = 16'(58);
			2: out = 16'(136);
			3: out = 16'(297);
			4: out = 16'(1307);
			5: out = 16'(-7945);
			6: out = 16'(11531);
			7: out = 16'(-32233);
			8: out = 16'(2660);
			9: out = 16'(18764);
			10: out = 16'(25030);
			11: out = 16'(-6370);
			12: out = 16'(10383);
			13: out = 16'(26300);
			14: out = 16'(-30392);
			15: out = 16'(28421);
			16: out = 16'(-21128);
			17: out = 16'(-21331);
			18: out = 16'(-19978);
			19: out = 16'(-32767);
			20: out = 16'(-21633);
			21: out = 16'(7570);
			22: out = 16'(-22613);
			23: out = 16'(26716);
			24: out = 16'(-29169);
			25: out = 16'(18385);
			26: out = 16'(-5193);
			27: out = 16'(-29787);
			28: out = 16'(-16740);
			29: out = 16'(4696);
			30: out = 16'(-2524);
			31: out = 16'(-21225);
			32: out = 16'(-19514);
			33: out = 16'(-2883);
			34: out = 16'(-24819);
			35: out = 16'(-25456);
			36: out = 16'(-757);
			37: out = 16'(-23698);
			38: out = 16'(27094);
			39: out = 16'(-24229);
			40: out = 16'(12825);
			41: out = 16'(17303);
			42: out = 16'(-22368);
			43: out = 16'(5157);
			44: out = 16'(31981);
			45: out = 16'(-17461);
			46: out = 16'(30359);
			47: out = 16'(-13277);
			48: out = 16'(29788);
			49: out = 16'(26357);
			50: out = 16'(4856);
			51: out = 16'(30656);
			52: out = 16'(8766);
			53: out = 16'(14752);
			54: out = 16'(-19310);
			55: out = 16'(-20949);
			56: out = 16'(-25892);
			57: out = 16'(20486);
			58: out = 16'(22830);
			59: out = 16'(-4983);
			60: out = 16'(1735);
			61: out = 16'(25648);
			62: out = 16'(-24023);
			63: out = 16'(-30199);
			64: out = 16'(-30566);
			65: out = 16'(-20486);
			66: out = 16'(32444);
			67: out = 16'(13230);
			68: out = 16'(4507);
			69: out = 16'(6085);
			70: out = 16'(-28064);
			71: out = 16'(-15251);
			72: out = 16'(-18181);
			73: out = 16'(9407);
			74: out = 16'(-10846);
			75: out = 16'(-25394);
			76: out = 16'(5104);
			77: out = 16'(1985);
			78: out = 16'(28628);
			79: out = 16'(-4314);
			80: out = 16'(-5934);
			81: out = 16'(-16181);
			82: out = 16'(16992);
			83: out = 16'(-17622);
			84: out = 16'(16512);
			85: out = 16'(14227);
			86: out = 16'(-7928);
			87: out = 16'(13063);
			88: out = 16'(-10250);
			89: out = 16'(-8411);
			90: out = 16'(15400);
			91: out = 16'(7418);
			92: out = 16'(-21302);
			93: out = 16'(-623);
			94: out = 16'(-23777);
			95: out = 16'(20332);
			96: out = 16'(-15717);
			97: out = 16'(-6198);
			98: out = 16'(5307);
			99: out = 16'(11831);
			100: out = 16'(-14907);
			101: out = 16'(-27780);
			102: out = 16'(-6313);
			103: out = 16'(264);
			104: out = 16'(29519);
			105: out = 16'(-26033);
			106: out = 16'(8942);
			107: out = 16'(-7338);
			108: out = 16'(3709);
			109: out = 16'(-4412);
			110: out = 16'(-1628);
			111: out = 16'(-23719);
			112: out = 16'(2710);
			113: out = 16'(17824);
			114: out = 16'(-3526);
			115: out = 16'(25091);
			116: out = 16'(20024);
			117: out = 16'(21219);
			118: out = 16'(-2060);
			119: out = 16'(-28281);
			120: out = 16'(8733);
			121: out = 16'(12005);
			122: out = 16'(-12917);
			123: out = 16'(-25264);
			124: out = 16'(-7991);
			125: out = 16'(-20898);
			126: out = 16'(2844);
			127: out = 16'(10660);
			128: out = 16'(-29522);
			129: out = 16'(20245);
			130: out = 16'(-26682);
			131: out = 16'(3174);
			132: out = 16'(-7976);
			133: out = 16'(-6230);
			134: out = 16'(-13470);
			135: out = 16'(495);
			136: out = 16'(-6032);
			137: out = 16'(4094);
			138: out = 16'(-3744);
			139: out = 16'(12077);
			140: out = 16'(-8647);
			141: out = 16'(4890);
			142: out = 16'(13640);
			143: out = 16'(17079);
			144: out = 16'(331);
			145: out = 16'(-4560);
			146: out = 16'(17999);
			147: out = 16'(-7671);
			148: out = 16'(18);
			149: out = 16'(-21929);
			150: out = 16'(-17755);
			151: out = 16'(-23343);
			152: out = 16'(23453);
			153: out = 16'(19537);
			154: out = 16'(11578);
			155: out = 16'(611);
			156: out = 16'(8556);
			157: out = 16'(1718);
			158: out = 16'(-22761);
			159: out = 16'(8110);
			160: out = 16'(-982);
			161: out = 16'(-8186);
			162: out = 16'(1469);
			163: out = 16'(-11320);
			164: out = 16'(-23581);
			165: out = 16'(9692);
			166: out = 16'(-10762);
			167: out = 16'(13935);
			168: out = 16'(-18389);
			169: out = 16'(1353);
			170: out = 16'(13761);
			171: out = 16'(-2321);
			172: out = 16'(-9321);
			173: out = 16'(7118);
			174: out = 16'(19165);
			175: out = 16'(-19665);
			176: out = 16'(18910);
			177: out = 16'(-17847);
			178: out = 16'(13725);
			179: out = 16'(12699);
			180: out = 16'(4944);
			181: out = 16'(-28435);
			182: out = 16'(-9466);
			183: out = 16'(3564);
			184: out = 16'(14413);
			185: out = 16'(-22364);
			186: out = 16'(14259);
			187: out = 16'(12463);
			188: out = 16'(20148);
			189: out = 16'(-13534);
			190: out = 16'(-13370);
			191: out = 16'(15641);
			192: out = 16'(16850);
			193: out = 16'(18247);
			194: out = 16'(-15997);
			195: out = 16'(-15860);
			196: out = 16'(-9148);
			197: out = 16'(14979);
			198: out = 16'(-7923);
			199: out = 16'(18090);
			200: out = 16'(10569);
			201: out = 16'(-5949);
			202: out = 16'(-10949);
			203: out = 16'(13609);
			204: out = 16'(1400);
			205: out = 16'(-1543);
			206: out = 16'(166);
			207: out = 16'(9358);
			208: out = 16'(-26106);
			209: out = 16'(14183);
			210: out = 16'(233);
			211: out = 16'(1282);
			212: out = 16'(-20664);
			213: out = 16'(9110);
			214: out = 16'(-16093);
			215: out = 16'(17848);
			216: out = 16'(-14584);
			217: out = 16'(3647);
			218: out = 16'(-8493);
			219: out = 16'(-7461);
			220: out = 16'(7102);
			221: out = 16'(-2831);
			222: out = 16'(12055);
			223: out = 16'(-772);
			224: out = 16'(5311);
			225: out = 16'(-3370);
			226: out = 16'(-538);
			227: out = 16'(-19063);
			228: out = 16'(11876);
			229: out = 16'(-14857);
			230: out = 16'(-2086);
			231: out = 16'(-7150);
			232: out = 16'(15626);
			233: out = 16'(-2161);
			234: out = 16'(-13669);
			235: out = 16'(14538);
			236: out = 16'(-19628);
			237: out = 16'(11908);
			238: out = 16'(-4087);
			239: out = 16'(-8428);
			240: out = 16'(-78);
			241: out = 16'(291);
			242: out = 16'(3856);
			243: out = 16'(3487);
			244: out = 16'(-5809);
			245: out = 16'(-7462);
			246: out = 16'(10593);
			247: out = 16'(10347);
			248: out = 16'(1636);
			249: out = 16'(-12425);
			250: out = 16'(17711);
			251: out = 16'(-591);
			252: out = 16'(-11126);
			253: out = 16'(-10699);
			254: out = 16'(-370);
			255: out = 16'(-9759);
			256: out = 16'(-17276);
			257: out = 16'(7835);
			258: out = 16'(8501);
			259: out = 16'(-7818);
			260: out = 16'(-4769);
			261: out = 16'(10754);
			262: out = 16'(-13031);
			263: out = 16'(-3277);
			264: out = 16'(4601);
			265: out = 16'(223);
			266: out = 16'(5356);
			267: out = 16'(5947);
			268: out = 16'(9005);
			269: out = 16'(-16948);
			270: out = 16'(41);
			271: out = 16'(-6585);
			272: out = 16'(-9521);
			273: out = 16'(3658);
			274: out = 16'(16616);
			275: out = 16'(12427);
			276: out = 16'(21885);
			277: out = 16'(7812);
			278: out = 16'(-9350);
			279: out = 16'(8948);
			280: out = 16'(-9319);
			281: out = 16'(8475);
			282: out = 16'(15457);
			283: out = 16'(-12288);
			284: out = 16'(4077);
			285: out = 16'(-12805);
			286: out = 16'(-12472);
			287: out = 16'(3135);
			288: out = 16'(-4139);
			289: out = 16'(-30596);
			290: out = 16'(-4450);
			291: out = 16'(-23782);
			292: out = 16'(7297);
			293: out = 16'(5528);
			294: out = 16'(7811);
			295: out = 16'(4353);
			296: out = 16'(-13603);
			297: out = 16'(9119);
			298: out = 16'(-12752);
			299: out = 16'(-3826);
			300: out = 16'(-9639);
			301: out = 16'(6325);
			302: out = 16'(-6527);
			303: out = 16'(7604);
			304: out = 16'(-5032);
			305: out = 16'(-3687);
			306: out = 16'(6999);
			307: out = 16'(2477);
			308: out = 16'(-2771);
			309: out = 16'(-8846);
			310: out = 16'(16536);
			311: out = 16'(3661);
			312: out = 16'(2717);
			313: out = 16'(15681);
			314: out = 16'(-1925);
			315: out = 16'(-3828);
			316: out = 16'(-6092);
			317: out = 16'(-14919);
			318: out = 16'(-3520);
			319: out = 16'(-18318);
			320: out = 16'(-18702);
			321: out = 16'(-16696);
			322: out = 16'(-4890);
			323: out = 16'(8201);
			324: out = 16'(2033);
			325: out = 16'(8878);
			326: out = 16'(7785);
			327: out = 16'(2438);
			328: out = 16'(8454);
			329: out = 16'(4787);
			330: out = 16'(-14251);
			331: out = 16'(879);
			332: out = 16'(1356);
			333: out = 16'(6074);
			334: out = 16'(1530);
			335: out = 16'(8817);
			336: out = 16'(-1360);
			337: out = 16'(-2271);
			338: out = 16'(-8288);
			339: out = 16'(5502);
			340: out = 16'(1857);
			341: out = 16'(4712);
			342: out = 16'(-21681);
			343: out = 16'(-320);
			344: out = 16'(5516);
			345: out = 16'(-1015);
			346: out = 16'(-1776);
			347: out = 16'(10015);
			348: out = 16'(-3062);
			349: out = 16'(14206);
			350: out = 16'(-2999);
			351: out = 16'(-9229);
			352: out = 16'(3899);
			353: out = 16'(10332);
			354: out = 16'(-318);
			355: out = 16'(-5848);
			356: out = 16'(-4598);
			357: out = 16'(2642);
			358: out = 16'(3870);
			359: out = 16'(3045);
			360: out = 16'(138);
			361: out = 16'(-209);
			362: out = 16'(1739);
			363: out = 16'(-9018);
			364: out = 16'(7469);
			365: out = 16'(7072);
			366: out = 16'(152);
			367: out = 16'(3087);
			368: out = 16'(-870);
			369: out = 16'(-535);
			370: out = 16'(7723);
			371: out = 16'(-7015);
			372: out = 16'(9954);
			373: out = 16'(3519);
			374: out = 16'(-7208);
			375: out = 16'(10820);
			376: out = 16'(-656);
			377: out = 16'(8992);
			378: out = 16'(-8841);
			379: out = 16'(-7603);
			380: out = 16'(-6535);
			381: out = 16'(7074);
			382: out = 16'(426);
			383: out = 16'(-1598);
			384: out = 16'(-7801);
			385: out = 16'(5378);
			386: out = 16'(-426);
			387: out = 16'(-3920);
			388: out = 16'(-1465);
			389: out = 16'(-8207);
			390: out = 16'(5974);
			391: out = 16'(1640);
			392: out = 16'(-3834);
			393: out = 16'(8751);
			394: out = 16'(-491);
			395: out = 16'(8485);
			396: out = 16'(-9235);
			397: out = 16'(-1400);
			398: out = 16'(12383);
			399: out = 16'(-12372);
			400: out = 16'(4896);
			401: out = 16'(-2911);
			402: out = 16'(-3303);
			403: out = 16'(1555);
			404: out = 16'(-8915);
			405: out = 16'(-5356);
			406: out = 16'(3264);
			407: out = 16'(12531);
			408: out = 16'(5618);
			409: out = 16'(-3237);
			410: out = 16'(2206);
			411: out = 16'(-1496);
			412: out = 16'(4325);
			413: out = 16'(-7661);
			414: out = 16'(4849);
			415: out = 16'(-14606);
			416: out = 16'(5858);
			417: out = 16'(3655);
			418: out = 16'(-8441);
			419: out = 16'(-16430);
			420: out = 16'(-7591);
			421: out = 16'(-3247);
			422: out = 16'(6752);
			423: out = 16'(-3579);
			424: out = 16'(1064);
			425: out = 16'(594);
			426: out = 16'(-384);
			427: out = 16'(2906);
			428: out = 16'(-969);
			429: out = 16'(-2982);
			430: out = 16'(-10685);
			431: out = 16'(6372);
			432: out = 16'(3510);
			433: out = 16'(8688);
			434: out = 16'(1985);
			435: out = 16'(-348);
			436: out = 16'(4290);
			437: out = 16'(9152);
			438: out = 16'(-1433);
			439: out = 16'(-2304);
			440: out = 16'(-5447);
			441: out = 16'(338);
			442: out = 16'(-1705);
			443: out = 16'(8416);
			444: out = 16'(3346);
			445: out = 16'(-216);
			446: out = 16'(-368);
			447: out = 16'(-2913);
			448: out = 16'(501);
			449: out = 16'(2416);
			450: out = 16'(-1112);
			451: out = 16'(-19576);
			452: out = 16'(9768);
			453: out = 16'(-8517);
			454: out = 16'(-2475);
			455: out = 16'(1206);
			456: out = 16'(-53);
			457: out = 16'(388);
			458: out = 16'(6749);
			459: out = 16'(2931);
			460: out = 16'(3246);
			461: out = 16'(8885);
			462: out = 16'(-3450);
			463: out = 16'(410);
			464: out = 16'(-31);
			465: out = 16'(130);
			466: out = 16'(4506);
			467: out = 16'(-16685);
			468: out = 16'(-2629);
			469: out = 16'(6364);
			470: out = 16'(3274);
			471: out = 16'(-2428);
			472: out = 16'(-6684);
			473: out = 16'(1701);
			474: out = 16'(4350);
			475: out = 16'(4097);
			476: out = 16'(6745);
			477: out = 16'(-2693);
			478: out = 16'(3451);
			479: out = 16'(565);
			480: out = 16'(1888);
			481: out = 16'(5935);
			482: out = 16'(4593);
			483: out = 16'(3951);
			484: out = 16'(1304);
			485: out = 16'(-3788);
			486: out = 16'(5333);
			487: out = 16'(5650);
			488: out = 16'(3326);
			489: out = 16'(-578);
			490: out = 16'(2711);
			491: out = 16'(375);
			492: out = 16'(-4118);
			493: out = 16'(-3001);
			494: out = 16'(221);
			495: out = 16'(-7564);
			496: out = 16'(8118);
			497: out = 16'(4734);
			498: out = 16'(-1876);
			499: out = 16'(-588);
			500: out = 16'(-2437);
			501: out = 16'(6066);
			502: out = 16'(-13372);
			503: out = 16'(1015);
			504: out = 16'(-4910);
			505: out = 16'(2057);
			506: out = 16'(-1120);
			507: out = 16'(1728);
			508: out = 16'(-5878);
			509: out = 16'(253);
			510: out = 16'(-8260);
			511: out = 16'(-4039);
			512: out = 16'(728);
			513: out = 16'(-3528);
			514: out = 16'(4996);
			515: out = 16'(-1632);
			516: out = 16'(-4902);
			517: out = 16'(7394);
			518: out = 16'(-5609);
			519: out = 16'(6594);
			520: out = 16'(632);
			521: out = 16'(-2397);
			522: out = 16'(866);
			523: out = 16'(1194);
			524: out = 16'(1740);
			525: out = 16'(1901);
			526: out = 16'(-2420);
			527: out = 16'(1746);
			528: out = 16'(-1733);
			529: out = 16'(3952);
			530: out = 16'(5147);
			531: out = 16'(4959);
			532: out = 16'(-1336);
			533: out = 16'(1596);
			534: out = 16'(-311);
			535: out = 16'(3521);
			536: out = 16'(-1738);
			537: out = 16'(-5766);
			538: out = 16'(-781);
			539: out = 16'(2813);
			540: out = 16'(7846);
			541: out = 16'(-2094);
			542: out = 16'(-3892);
			543: out = 16'(3653);
			544: out = 16'(3306);
			545: out = 16'(-3382);
			546: out = 16'(-307);
			547: out = 16'(111);
			548: out = 16'(4832);
			549: out = 16'(2121);
			550: out = 16'(-5269);
			551: out = 16'(1754);
			552: out = 16'(-1861);
			553: out = 16'(-5320);
			554: out = 16'(6641);
			555: out = 16'(-3239);
			556: out = 16'(-1218);
			557: out = 16'(5401);
			558: out = 16'(1318);
			559: out = 16'(-2176);
			560: out = 16'(-1527);
			561: out = 16'(-6861);
			562: out = 16'(-5782);
			563: out = 16'(1292);
			564: out = 16'(-6638);
			565: out = 16'(2551);
			566: out = 16'(-2480);
			567: out = 16'(2517);
			568: out = 16'(581);
			569: out = 16'(3229);
			570: out = 16'(-1766);
			571: out = 16'(6403);
			572: out = 16'(506);
			573: out = 16'(-6999);
			574: out = 16'(-2512);
			575: out = 16'(1875);
			576: out = 16'(-8854);
			577: out = 16'(-5812);
			578: out = 16'(-3424);
			579: out = 16'(3300);
			580: out = 16'(2528);
			581: out = 16'(1075);
			582: out = 16'(6547);
			583: out = 16'(6585);
			584: out = 16'(6623);
			585: out = 16'(1980);
			586: out = 16'(-3040);
			587: out = 16'(-3135);
			588: out = 16'(3509);
			589: out = 16'(673);
			590: out = 16'(-3018);
			591: out = 16'(-4775);
			592: out = 16'(141);
			593: out = 16'(-879);
			594: out = 16'(5082);
			595: out = 16'(-3092);
			596: out = 16'(-3592);
			597: out = 16'(5100);
			598: out = 16'(1959);
			599: out = 16'(-765);
			600: out = 16'(-2874);
			601: out = 16'(4555);
			602: out = 16'(461);
			603: out = 16'(-4552);
			604: out = 16'(2975);
			605: out = 16'(-3855);
			606: out = 16'(4695);
			607: out = 16'(1697);
			608: out = 16'(-2312);
			609: out = 16'(252);
			610: out = 16'(51);
			611: out = 16'(3967);
			612: out = 16'(1156);
			613: out = 16'(-2002);
			614: out = 16'(-115);
			615: out = 16'(1815);
			616: out = 16'(1015);
			617: out = 16'(-1162);
			618: out = 16'(-9384);
			619: out = 16'(5832);
			620: out = 16'(-324);
			621: out = 16'(-5981);
			622: out = 16'(5119);
			623: out = 16'(4857);
			624: out = 16'(-2684);
			625: out = 16'(2531);
			626: out = 16'(-1588);
			627: out = 16'(87);
			628: out = 16'(3774);
			629: out = 16'(1086);
			630: out = 16'(-5810);
			631: out = 16'(-3738);
			632: out = 16'(4321);
			633: out = 16'(3716);
			634: out = 16'(2936);
			635: out = 16'(-3802);
			636: out = 16'(-2144);
			637: out = 16'(370);
			638: out = 16'(547);
			639: out = 16'(-4094);
			640: out = 16'(-3623);
			641: out = 16'(-5092);
			642: out = 16'(608);
			643: out = 16'(-2862);
			644: out = 16'(2597);
			645: out = 16'(602);
			646: out = 16'(-1456);
			647: out = 16'(2237);
			648: out = 16'(1292);
			649: out = 16'(-3245);
			650: out = 16'(-725);
			651: out = 16'(1006);
			652: out = 16'(-408);
			653: out = 16'(1696);
			654: out = 16'(1590);
			655: out = 16'(195);
			656: out = 16'(-847);
			657: out = 16'(4);
			658: out = 16'(-1911);
			659: out = 16'(2524);
			660: out = 16'(-1228);
			661: out = 16'(-3538);
			662: out = 16'(-4014);
			663: out = 16'(3530);
			664: out = 16'(3323);
			665: out = 16'(1463);
			666: out = 16'(-2538);
			667: out = 16'(857);
			668: out = 16'(651);
			669: out = 16'(720);
			670: out = 16'(-3938);
			671: out = 16'(-4474);
			672: out = 16'(5561);
			673: out = 16'(453);
			674: out = 16'(-4908);
			675: out = 16'(-1210);
			676: out = 16'(-3610);
			677: out = 16'(4563);
			678: out = 16'(37);
			679: out = 16'(-4201);
			680: out = 16'(3016);
			681: out = 16'(1128);
			682: out = 16'(1374);
			683: out = 16'(-63);
			684: out = 16'(1546);
			685: out = 16'(6246);
			686: out = 16'(-5259);
			687: out = 16'(139);
			688: out = 16'(-1163);
			689: out = 16'(-4479);
			690: out = 16'(4395);
			691: out = 16'(-1759);
			692: out = 16'(-1458);
			693: out = 16'(2997);
			694: out = 16'(3139);
			695: out = 16'(735);
			696: out = 16'(-634);
			697: out = 16'(-2941);
			698: out = 16'(2028);
			699: out = 16'(-3637);
			700: out = 16'(-1770);
			701: out = 16'(2599);
			702: out = 16'(3352);
			703: out = 16'(1676);
			704: out = 16'(-213);
			705: out = 16'(-1436);
			706: out = 16'(-5427);
			707: out = 16'(-6592);
			708: out = 16'(3599);
			709: out = 16'(207);
			710: out = 16'(-1014);
			711: out = 16'(763);
			712: out = 16'(171);
			713: out = 16'(-1622);
			714: out = 16'(-1567);
			715: out = 16'(1299);
			716: out = 16'(2201);
			717: out = 16'(1788);
			718: out = 16'(1060);
			719: out = 16'(-659);
			720: out = 16'(-5292);
			721: out = 16'(-5064);
			722: out = 16'(-2943);
			723: out = 16'(626);
			724: out = 16'(2414);
			725: out = 16'(3849);
			726: out = 16'(1215);
			727: out = 16'(-775);
			728: out = 16'(2477);
			729: out = 16'(1135);
			730: out = 16'(-470);
			731: out = 16'(2642);
			732: out = 16'(2009);
			733: out = 16'(786);
			734: out = 16'(3222);
			735: out = 16'(-3040);
			736: out = 16'(2555);
			737: out = 16'(670);
			738: out = 16'(2011);
			739: out = 16'(-1726);
			740: out = 16'(246);
			741: out = 16'(-21);
			742: out = 16'(1873);
			743: out = 16'(3856);
			744: out = 16'(2472);
			745: out = 16'(-1043);
			746: out = 16'(-223);
			747: out = 16'(1897);
			748: out = 16'(-1821);
			749: out = 16'(-6699);
			750: out = 16'(-2687);
			751: out = 16'(2102);
			752: out = 16'(-2050);
			753: out = 16'(1626);
			754: out = 16'(-255);
			755: out = 16'(704);
			756: out = 16'(558);
			757: out = 16'(-3053);
			758: out = 16'(18);
			759: out = 16'(-1865);
			760: out = 16'(3141);
			761: out = 16'(-2657);
			762: out = 16'(2015);
			763: out = 16'(3541);
			764: out = 16'(-3146);
			765: out = 16'(1819);
			766: out = 16'(-1397);
			767: out = 16'(-619);
			768: out = 16'(370);
			769: out = 16'(609);
			770: out = 16'(-263);
			771: out = 16'(148);
			772: out = 16'(2900);
			773: out = 16'(3229);
			774: out = 16'(-1959);
			775: out = 16'(331);
			776: out = 16'(-1370);
			777: out = 16'(1228);
			778: out = 16'(-1366);
			779: out = 16'(-631);
			780: out = 16'(-4673);
			781: out = 16'(1857);
			782: out = 16'(-1163);
			783: out = 16'(2119);
			784: out = 16'(-557);
			785: out = 16'(-2515);
			786: out = 16'(-2207);
			787: out = 16'(826);
			788: out = 16'(-617);
			789: out = 16'(505);
			790: out = 16'(3286);
			791: out = 16'(-1097);
			792: out = 16'(-1873);
			793: out = 16'(349);
			794: out = 16'(1817);
			795: out = 16'(-3296);
			796: out = 16'(43);
			797: out = 16'(-5075);
			798: out = 16'(3835);
			799: out = 16'(-2627);
			800: out = 16'(2554);
			801: out = 16'(2339);
			802: out = 16'(1239);
			803: out = 16'(-2102);
			804: out = 16'(3098);
			805: out = 16'(-3112);
			806: out = 16'(-551);
			807: out = 16'(-1229);
			808: out = 16'(69);
			809: out = 16'(3014);
			810: out = 16'(-5315);
			811: out = 16'(2539);
			812: out = 16'(-2032);
			813: out = 16'(-219);
			814: out = 16'(-546);
			815: out = 16'(-491);
			816: out = 16'(2205);
			817: out = 16'(-1172);
			818: out = 16'(2502);
			819: out = 16'(763);
			820: out = 16'(-243);
			821: out = 16'(1933);
			822: out = 16'(-361);
			823: out = 16'(-283);
			824: out = 16'(-201);
			825: out = 16'(-4570);
			826: out = 16'(459);
			827: out = 16'(1);
			828: out = 16'(-3252);
			829: out = 16'(1218);
			830: out = 16'(-975);
			831: out = 16'(-1769);
			832: out = 16'(-944);
			833: out = 16'(-1217);
			834: out = 16'(1664);
			835: out = 16'(-401);
			836: out = 16'(-67);
			837: out = 16'(-1276);
			838: out = 16'(439);
			839: out = 16'(-2751);
			840: out = 16'(-1707);
			841: out = 16'(-2693);
			842: out = 16'(501);
			843: out = 16'(-2114);
			844: out = 16'(177);
			845: out = 16'(550);
			846: out = 16'(1945);
			847: out = 16'(3017);
			848: out = 16'(1692);
			849: out = 16'(1046);
			850: out = 16'(-2604);
			851: out = 16'(1304);
			852: out = 16'(1449);
			853: out = 16'(2867);
			854: out = 16'(-87);
			855: out = 16'(1510);
			856: out = 16'(-962);
			857: out = 16'(1078);
			858: out = 16'(-1058);
			859: out = 16'(998);
			860: out = 16'(-449);
			861: out = 16'(-530);
			862: out = 16'(-604);
			863: out = 16'(245);
			864: out = 16'(1062);
			865: out = 16'(-140);
			866: out = 16'(-777);
			867: out = 16'(-4445);
			868: out = 16'(1287);
			869: out = 16'(-1903);
			870: out = 16'(-1233);
			871: out = 16'(-123);
			872: out = 16'(1691);
			873: out = 16'(403);
			874: out = 16'(-610);
			875: out = 16'(251);
			876: out = 16'(1037);
			877: out = 16'(-1739);
			878: out = 16'(-3068);
			879: out = 16'(982);
			880: out = 16'(-31);
			881: out = 16'(1584);
			882: out = 16'(-738);
			883: out = 16'(-2770);
			884: out = 16'(1291);
			885: out = 16'(891);
			886: out = 16'(587);
			887: out = 16'(-46);
			888: out = 16'(407);
			889: out = 16'(-2);
			890: out = 16'(-6070);
			891: out = 16'(620);
			892: out = 16'(-961);
			893: out = 16'(-2074);
			894: out = 16'(1267);
			895: out = 16'(137);
			896: out = 16'(-2252);
			897: out = 16'(844);
			898: out = 16'(-1693);
			899: out = 16'(-493);
			900: out = 16'(-1320);
			901: out = 16'(25);
			902: out = 16'(1263);
			903: out = 16'(1078);
			904: out = 16'(2180);
			905: out = 16'(1795);
			906: out = 16'(-4195);
			907: out = 16'(-143);
			908: out = 16'(1246);
			909: out = 16'(1789);
			910: out = 16'(1239);
			911: out = 16'(277);
			912: out = 16'(2246);
			913: out = 16'(970);
			914: out = 16'(524);
			915: out = 16'(994);
			916: out = 16'(-537);
			917: out = 16'(860);
			918: out = 16'(778);
			919: out = 16'(1204);
			920: out = 16'(371);
			921: out = 16'(-528);
			922: out = 16'(-2216);
			923: out = 16'(1983);
			924: out = 16'(-1100);
			925: out = 16'(-686);
			926: out = 16'(-529);
			927: out = 16'(-158);
			928: out = 16'(905);
			929: out = 16'(-956);
			930: out = 16'(781);
			931: out = 16'(-65);
			932: out = 16'(-1232);
			933: out = 16'(-286);
			934: out = 16'(-70);
			935: out = 16'(1663);
			936: out = 16'(-768);
			937: out = 16'(-511);
			938: out = 16'(-395);
			939: out = 16'(387);
			940: out = 16'(-674);
			941: out = 16'(303);
			942: out = 16'(-2028);
			943: out = 16'(-1225);
			944: out = 16'(1612);
			945: out = 16'(-652);
			946: out = 16'(595);
			947: out = 16'(-504);
			948: out = 16'(261);
			949: out = 16'(-718);
			950: out = 16'(1082);
			951: out = 16'(-1137);
			952: out = 16'(382);
			953: out = 16'(-1390);
			954: out = 16'(-115);
			955: out = 16'(628);
			956: out = 16'(100);
			957: out = 16'(1018);
			958: out = 16'(-84);
			959: out = 16'(1525);
			960: out = 16'(-1245);
			961: out = 16'(1371);
			962: out = 16'(1889);
			963: out = 16'(1901);
			964: out = 16'(168);
			965: out = 16'(-441);
			966: out = 16'(1271);
			967: out = 16'(3);
			968: out = 16'(-80);
			969: out = 16'(-685);
			970: out = 16'(1535);
			971: out = 16'(1495);
			972: out = 16'(-2518);
			973: out = 16'(48);
			974: out = 16'(-5);
			975: out = 16'(-513);
			976: out = 16'(-60);
			977: out = 16'(658);
			978: out = 16'(-601);
			979: out = 16'(137);
			980: out = 16'(93);
			981: out = 16'(-168);
			982: out = 16'(-604);
			983: out = 16'(693);
			984: out = 16'(-529);
			985: out = 16'(164);
			986: out = 16'(-854);
			987: out = 16'(-2262);
			988: out = 16'(-1300);
			989: out = 16'(993);
			990: out = 16'(32);
			991: out = 16'(-1155);
			992: out = 16'(1152);
			993: out = 16'(217);
			994: out = 16'(928);
			995: out = 16'(417);
			996: out = 16'(-881);
			997: out = 16'(-305);
			998: out = 16'(835);
			999: out = 16'(-95);
			1000: out = 16'(597);
			1001: out = 16'(965);
			1002: out = 16'(812);
			1003: out = 16'(421);
			1004: out = 16'(-74);
			1005: out = 16'(-302);
			1006: out = 16'(-179);
			1007: out = 16'(-1004);
			1008: out = 16'(416);
			1009: out = 16'(285);
			1010: out = 16'(670);
			1011: out = 16'(-1985);
			1012: out = 16'(999);
			1013: out = 16'(193);
			1014: out = 16'(-885);
			1015: out = 16'(345);
			1016: out = 16'(-1714);
			1017: out = 16'(490);
			1018: out = 16'(15);
			1019: out = 16'(277);
			1020: out = 16'(-593);
			1021: out = 16'(386);
			1022: out = 16'(-1330);
			1023: out = 16'(-1208);
			1024: out = 16'(-1237);
			1025: out = 16'(-673);
			1026: out = 16'(-986);
			1027: out = 16'(292);
			1028: out = 16'(-640);
			1029: out = 16'(621);
			1030: out = 16'(-108);
			1031: out = 16'(-579);
			1032: out = 16'(31);
			1033: out = 16'(-319);
			1034: out = 16'(1367);
			1035: out = 16'(-264);
			1036: out = 16'(58);
			1037: out = 16'(162);
			1038: out = 16'(-11);
			1039: out = 16'(783);
			1040: out = 16'(802);
			1041: out = 16'(366);
			1042: out = 16'(-223);
			1043: out = 16'(375);
			1044: out = 16'(169);
			1045: out = 16'(1336);
			1046: out = 16'(133);
			1047: out = 16'(663);
			1048: out = 16'(-777);
			1049: out = 16'(-54);
			1050: out = 16'(496);
			1051: out = 16'(519);
			1052: out = 16'(-375);
			1053: out = 16'(-838);
			1054: out = 16'(153);
			1055: out = 16'(227);
			1056: out = 16'(-292);
			1057: out = 16'(-1052);
			1058: out = 16'(-1969);
			1059: out = 16'(-305);
			1060: out = 16'(28);
			1061: out = 16'(412);
			1062: out = 16'(445);
			1063: out = 16'(589);
			1064: out = 16'(-603);
			1065: out = 16'(105);
			1066: out = 16'(217);
			1067: out = 16'(6);
			1068: out = 16'(296);
			1069: out = 16'(-683);
			1070: out = 16'(111);
			1071: out = 16'(177);
			1072: out = 16'(-104);
			1073: out = 16'(-571);
			1074: out = 16'(-796);
			1075: out = 16'(-797);
			1076: out = 16'(399);
			1077: out = 16'(55);
			1078: out = 16'(285);
			1079: out = 16'(634);
			1080: out = 16'(-194);
			1081: out = 16'(1100);
			1082: out = 16'(-369);
			1083: out = 16'(-408);
			1084: out = 16'(-1431);
			1085: out = 16'(607);
			1086: out = 16'(-124);
			1087: out = 16'(247);
			1088: out = 16'(19);
			1089: out = 16'(32);
			1090: out = 16'(26);
			1091: out = 16'(-10);
			1092: out = 16'(-131);
			1093: out = 16'(-216);
			1094: out = 16'(64);
			1095: out = 16'(-146);
			1096: out = 16'(-190);
			1097: out = 16'(723);
			1098: out = 16'(388);
			1099: out = 16'(-352);
			1100: out = 16'(639);
			1101: out = 16'(-227);
			1102: out = 16'(209);
			1103: out = 16'(245);
			1104: out = 16'(-72);
			1105: out = 16'(-170);
			1106: out = 16'(-1087);
			1107: out = 16'(286);
			1108: out = 16'(657);
			1109: out = 16'(411);
			1110: out = 16'(-265);
			1111: out = 16'(269);
			1112: out = 16'(-413);
			1113: out = 16'(23);
			1114: out = 16'(-494);
			1115: out = 16'(-88);
			1116: out = 16'(-1426);
			1117: out = 16'(-944);
			1118: out = 16'(-326);
			1119: out = 16'(62);
			1120: out = 16'(92);
			1121: out = 16'(-379);
			1122: out = 16'(-244);
			1123: out = 16'(621);
			1124: out = 16'(-49);
			1125: out = 16'(422);
			1126: out = 16'(-22);
			1127: out = 16'(-21);
			1128: out = 16'(-726);
			1129: out = 16'(-335);
			1130: out = 16'(-62);
			1131: out = 16'(-881);
			1132: out = 16'(-725);
			1133: out = 16'(579);
			1134: out = 16'(-492);
			1135: out = 16'(-98);
			1136: out = 16'(-110);
			1137: out = 16'(-394);
			1138: out = 16'(318);
			1139: out = 16'(-916);
			1140: out = 16'(238);
			1141: out = 16'(-456);
			1142: out = 16'(151);
			1143: out = 16'(-55);
			1144: out = 16'(-176);
			1145: out = 16'(444);
			1146: out = 16'(777);
			1147: out = 16'(-183);
			1148: out = 16'(-68);
			1149: out = 16'(-24);
			1150: out = 16'(-80);
			1151: out = 16'(-62);
			1152: out = 16'(296);
			1153: out = 16'(157);
			1154: out = 16'(-96);
			1155: out = 16'(203);
			1156: out = 16'(125);
			1157: out = 16'(-545);
			1158: out = 16'(-34);
			1159: out = 16'(-547);
			1160: out = 16'(-206);
			1161: out = 16'(84);
			1162: out = 16'(4);
			1163: out = 16'(-215);
			1164: out = 16'(294);
			1165: out = 16'(-265);
			1166: out = 16'(302);
			1167: out = 16'(-235);
			1168: out = 16'(-220);
			1169: out = 16'(506);
			1170: out = 16'(127);
			1171: out = 16'(-371);
			1172: out = 16'(-187);
			1173: out = 16'(63);
			1174: out = 16'(421);
			1175: out = 16'(-1239);
			1176: out = 16'(-606);
			1177: out = 16'(657);
			1178: out = 16'(-267);
			1179: out = 16'(14);
			1180: out = 16'(-7);
			1181: out = 16'(-321);
			1182: out = 16'(-366);
			1183: out = 16'(389);
			1184: out = 16'(-447);
			1185: out = 16'(-125);
			1186: out = 16'(-227);
			1187: out = 16'(343);
			1188: out = 16'(-5);
			1189: out = 16'(-262);
			1190: out = 16'(-125);
			1191: out = 16'(560);
			1192: out = 16'(351);
			1193: out = 16'(-422);
			1194: out = 16'(279);
			1195: out = 16'(-354);
			1196: out = 16'(179);
			1197: out = 16'(-141);
			1198: out = 16'(-46);
			1199: out = 16'(-385);
			1200: out = 16'(163);
			1201: out = 16'(64);
			1202: out = 16'(-387);
			1203: out = 16'(109);
			1204: out = 16'(-247);
			1205: out = 16'(269);
			1206: out = 16'(156);
			1207: out = 16'(-776);
			1208: out = 16'(189);
			1209: out = 16'(0);
			1210: out = 16'(-483);
			1211: out = 16'(24);
			1212: out = 16'(314);
			1213: out = 16'(457);
			1214: out = 16'(-124);
			1215: out = 16'(-522);
			1216: out = 16'(84);
			1217: out = 16'(-1);
			1218: out = 16'(-217);
			1219: out = 16'(-17);
			1220: out = 16'(-391);
			1221: out = 16'(75);
			1222: out = 16'(-57);
			1223: out = 16'(63);
			1224: out = 16'(71);
			1225: out = 16'(51);
			1226: out = 16'(-109);
			1227: out = 16'(-274);
			1228: out = 16'(-333);
			1229: out = 16'(-185);
			1230: out = 16'(30);
			1231: out = 16'(191);
			1232: out = 16'(118);
			1233: out = 16'(-211);
			1234: out = 16'(181);
			1235: out = 16'(440);
			1236: out = 16'(156);
			1237: out = 16'(-201);
			1238: out = 16'(-335);
			1239: out = 16'(343);
			1240: out = 16'(93);
			1241: out = 16'(-245);
			1242: out = 16'(-631);
			1243: out = 16'(310);
			1244: out = 16'(-317);
			1245: out = 16'(102);
			1246: out = 16'(-321);
			1247: out = 16'(-47);
			1248: out = 16'(-96);
			default: out = 0;
		endcase
	end
endmodule
