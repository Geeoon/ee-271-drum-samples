module snare_lookup(index, out);
	input logic unsigned [13:0] index;
	output logic signed [15:0] out;
	always_comb begin
		case(index)
			0: out = 16'(18770);
			1: out = 16'(17990);
			2: out = 16'(23670);
			3: out = 16'(0);
			4: out = 16'(16727);
			5: out = 16'(17750);
			6: out = 16'(28006);
			7: out = 16'(8308);
			8: out = 16'(16);
			9: out = 16'(0);
			10: out = 16'(1);
			11: out = 16'(1);
			12: out = 16'(-21435);
			13: out = 16'(0);
			14: out = 16'(22666);
			15: out = 16'(1);
			16: out = 16'(2);
			17: out = 16'(16);
			18: out = 16'(24932);
			19: out = 16'(24948);
			20: out = 16'(23562);
			21: out = 16'(0);
			22: out = 16'(0);
			23: out = 16'(0);
			24: out = 16'(13);
			25: out = 16'(-69);
			26: out = 16'(-42);
			27: out = 16'(-191);
			28: out = 16'(-52);
			29: out = 16'(-982);
			30: out = 16'(-2614);
			31: out = 16'(1647);
			32: out = 16'(7171);
			33: out = 16'(6374);
			34: out = 16'(423);
			35: out = 16'(-674);
			36: out = 16'(2183);
			37: out = 16'(4318);
			38: out = 16'(3315);
			39: out = 16'(-4073);
			40: out = 16'(-5407);
			41: out = 16'(910);
			42: out = 16'(6971);
			43: out = 16'(1914);
			44: out = 16'(-9265);
			45: out = 16'(-5867);
			46: out = 16'(8736);
			47: out = 16'(9994);
			48: out = 16'(1518);
			49: out = 16'(-9887);
			50: out = 16'(-7403);
			51: out = 16'(2245);
			52: out = 16'(6871);
			53: out = 16'(8592);
			54: out = 16'(3647);
			55: out = 16'(-616);
			56: out = 16'(-4366);
			57: out = 16'(1649);
			58: out = 16'(13958);
			59: out = 16'(8119);
			60: out = 16'(-10684);
			61: out = 16'(-10784);
			62: out = 16'(-850);
			63: out = 16'(-433);
			64: out = 16'(-5174);
			65: out = 16'(-13997);
			66: out = 16'(-11329);
			67: out = 16'(5613);
			68: out = 16'(19084);
			69: out = 16'(16067);
			70: out = 16'(976);
			71: out = 16'(-10516);
			72: out = 16'(-8681);
			73: out = 16'(1746);
			74: out = 16'(12581);
			75: out = 16'(9883);
			76: out = 16'(-7718);
			77: out = 16'(-6940);
			78: out = 16'(5753);
			79: out = 16'(-1122);
			80: out = 16'(-11558);
			81: out = 16'(-16993);
			82: out = 16'(-8225);
			83: out = 16'(6572);
			84: out = 16'(22781);
			85: out = 16'(7882);
			86: out = 16'(-7089);
			87: out = 16'(-3909);
			88: out = 16'(1547);
			89: out = 16'(9372);
			90: out = 16'(1096);
			91: out = 16'(1684);
			92: out = 16'(1475);
			93: out = 16'(1186);
			94: out = 16'(-1940);
			95: out = 16'(-1972);
			96: out = 16'(-11965);
			97: out = 16'(-17898);
			98: out = 16'(-13735);
			99: out = 16'(237);
			100: out = 16'(8095);
			101: out = 16'(-4700);
			102: out = 16'(-11835);
			103: out = 16'(-3718);
			104: out = 16'(12069);
			105: out = 16'(8266);
			106: out = 16'(-3364);
			107: out = 16'(-13760);
			108: out = 16'(-5930);
			109: out = 16'(1311);
			110: out = 16'(14555);
			111: out = 16'(32248);
			112: out = 16'(21052);
			113: out = 16'(-13644);
			114: out = 16'(-31710);
			115: out = 16'(-29625);
			116: out = 16'(-14769);
			117: out = 16'(25182);
			118: out = 16'(31201);
			119: out = 16'(31299);
			120: out = 16'(30798);
			121: out = 16'(31185);
			122: out = 16'(30856);
			123: out = 16'(30389);
			124: out = 16'(21219);
			125: out = 16'(29782);
			126: out = 16'(31191);
			127: out = 16'(30781);
			128: out = 16'(30918);
			129: out = 16'(30749);
			130: out = 16'(30851);
			131: out = 16'(30464);
			132: out = 16'(28162);
			133: out = 16'(30814);
			134: out = 16'(30790);
			135: out = 16'(30714);
			136: out = 16'(30695);
			137: out = 16'(30718);
			138: out = 16'(30564);
			139: out = 16'(30568);
			140: out = 16'(30600);
			141: out = 16'(30553);
			142: out = 16'(30505);
			143: out = 16'(30581);
			144: out = 16'(30557);
			145: out = 16'(30473);
			146: out = 16'(30486);
			147: out = 16'(30473);
			148: out = 16'(30421);
			149: out = 16'(30375);
			150: out = 16'(30321);
			151: out = 16'(30303);
			152: out = 16'(30364);
			153: out = 16'(30372);
			154: out = 16'(30293);
			155: out = 16'(30228);
			156: out = 16'(30222);
			157: out = 16'(30193);
			158: out = 16'(30189);
			159: out = 16'(30131);
			160: out = 16'(30118);
			161: out = 16'(30079);
			162: out = 16'(30117);
			163: out = 16'(30102);
			164: out = 16'(30066);
			165: out = 16'(30030);
			166: out = 16'(30008);
			167: out = 16'(29941);
			168: out = 16'(29918);
			169: out = 16'(29992);
			170: out = 16'(29011);
			171: out = 16'(24247);
			172: out = 16'(26620);
			173: out = 16'(30279);
			174: out = 16'(19896);
			175: out = 16'(8215);
			176: out = 16'(9283);
			177: out = 16'(17558);
			178: out = 16'(20280);
			179: out = 16'(4734);
			180: out = 16'(-7249);
			181: out = 16'(-3920);
			182: out = 16'(10895);
			183: out = 16'(10817);
			184: out = 16'(-7541);
			185: out = 16'(-11217);
			186: out = 16'(-4488);
			187: out = 16'(-2575);
			188: out = 16'(-14923);
			189: out = 16'(-19108);
			190: out = 16'(-15315);
			191: out = 16'(-15552);
			192: out = 16'(-25236);
			193: out = 16'(-26917);
			194: out = 16'(-27661);
			195: out = 16'(-31200);
			196: out = 16'(-31114);
			197: out = 16'(-31375);
			198: out = 16'(-31019);
			199: out = 16'(-31314);
			200: out = 16'(-30870);
			201: out = 16'(-31465);
			202: out = 16'(-28465);
			203: out = 16'(-26068);
			204: out = 16'(-26714);
			205: out = 16'(-26946);
			206: out = 16'(-30527);
			207: out = 16'(-31046);
			208: out = 16'(-30997);
			209: out = 16'(-31029);
			210: out = 16'(-30884);
			211: out = 16'(-30958);
			212: out = 16'(-30693);
			213: out = 16'(-31033);
			214: out = 16'(-30682);
			215: out = 16'(-31080);
			216: out = 16'(-30399);
			217: out = 16'(-31163);
			218: out = 16'(-22490);
			219: out = 16'(-21108);
			220: out = 16'(-30972);
			221: out = 16'(-30445);
			222: out = 16'(-30828);
			223: out = 16'(-30489);
			224: out = 16'(-30718);
			225: out = 16'(-30436);
			226: out = 16'(-28366);
			227: out = 16'(-28519);
			228: out = 16'(-28153);
			229: out = 16'(-19376);
			230: out = 16'(-12644);
			231: out = 16'(-23726);
			232: out = 16'(-30378);
			233: out = 16'(-30941);
			234: out = 16'(-24856);
			235: out = 16'(-17396);
			236: out = 16'(-24247);
			237: out = 16'(-25690);
			238: out = 16'(-16177);
			239: out = 16'(-7334);
			240: out = 16'(-6742);
			241: out = 16'(-9245);
			242: out = 16'(-15967);
			243: out = 16'(-13501);
			244: out = 16'(-5105);
			245: out = 16'(2990);
			246: out = 16'(11316);
			247: out = 16'(7686);
			248: out = 16'(-597);
			249: out = 16'(2588);
			250: out = 16'(5101);
			251: out = 16'(2545);
			252: out = 16'(874);
			253: out = 16'(2400);
			254: out = 16'(608);
			255: out = 16'(13561);
			256: out = 16'(28876);
			257: out = 16'(19319);
			258: out = 16'(11304);
			259: out = 16'(9195);
			260: out = 16'(17035);
			261: out = 16'(28309);
			262: out = 16'(30675);
			263: out = 16'(30687);
			264: out = 16'(30894);
			265: out = 16'(23845);
			266: out = 16'(16016);
			267: out = 16'(17744);
			268: out = 16'(18741);
			269: out = 16'(17591);
			270: out = 16'(14908);
			271: out = 16'(23357);
			272: out = 16'(31049);
			273: out = 16'(30286);
			274: out = 16'(30730);
			275: out = 16'(30351);
			276: out = 16'(30672);
			277: out = 16'(29475);
			278: out = 16'(23368);
			279: out = 16'(23385);
			280: out = 16'(29874);
			281: out = 16'(30478);
			282: out = 16'(30406);
			283: out = 16'(30251);
			284: out = 16'(30366);
			285: out = 16'(29827);
			286: out = 16'(29572);
			287: out = 16'(30598);
			288: out = 16'(29949);
			289: out = 16'(30223);
			290: out = 16'(21598);
			291: out = 16'(22626);
			292: out = 16'(30543);
			293: out = 16'(28142);
			294: out = 16'(20592);
			295: out = 16'(20604);
			296: out = 16'(28273);
			297: out = 16'(29824);
			298: out = 16'(30509);
			299: out = 16'(28290);
			300: out = 16'(22155);
			301: out = 16'(16221);
			302: out = 16'(16683);
			303: out = 16'(18366);
			304: out = 16'(18665);
			305: out = 16'(27171);
			306: out = 16'(28552);
			307: out = 16'(14681);
			308: out = 16'(945);
			309: out = 16'(3919);
			310: out = 16'(18482);
			311: out = 16'(19637);
			312: out = 16'(3700);
			313: out = 16'(129);
			314: out = 16'(7575);
			315: out = 16'(7074);
			316: out = 16'(-782);
			317: out = 16'(1314);
			318: out = 16'(6350);
			319: out = 16'(13925);
			320: out = 16'(11605);
			321: out = 16'(6120);
			322: out = 16'(-1835);
			323: out = 16'(-4194);
			324: out = 16'(6661);
			325: out = 16'(20750);
			326: out = 16'(21200);
			327: out = 16'(4554);
			328: out = 16'(-5079);
			329: out = 16'(-2594);
			330: out = 16'(1771);
			331: out = 16'(-2702);
			332: out = 16'(-9182);
			333: out = 16'(-4649);
			334: out = 16'(5078);
			335: out = 16'(14312);
			336: out = 16'(9792);
			337: out = 16'(511);
			338: out = 16'(-7227);
			339: out = 16'(-502);
			340: out = 16'(7102);
			341: out = 16'(8494);
			342: out = 16'(7541);
			343: out = 16'(5455);
			344: out = 16'(-35);
			345: out = 16'(-6256);
			346: out = 16'(-9563);
			347: out = 16'(-9707);
			348: out = 16'(-13159);
			349: out = 16'(-11238);
			350: out = 16'(-652);
			351: out = 16'(3714);
			352: out = 16'(12526);
			353: out = 16'(13581);
			354: out = 16'(12742);
			355: out = 16'(2627);
			356: out = 16'(-1022);
			357: out = 16'(4851);
			358: out = 16'(12313);
			359: out = 16'(21958);
			360: out = 16'(16283);
			361: out = 16'(2735);
			362: out = 16'(-3839);
			363: out = 16'(-3405);
			364: out = 16'(-1713);
			365: out = 16'(-5138);
			366: out = 16'(-7361);
			367: out = 16'(-2006);
			368: out = 16'(-1111);
			369: out = 16'(-1365);
			370: out = 16'(4665);
			371: out = 16'(13367);
			372: out = 16'(14412);
			373: out = 16'(-489);
			374: out = 16'(-8387);
			375: out = 16'(-8400);
			376: out = 16'(-1358);
			377: out = 16'(3197);
			378: out = 16'(1539);
			379: out = 16'(-5299);
			380: out = 16'(-13815);
			381: out = 16'(-14595);
			382: out = 16'(-8642);
			383: out = 16'(-4118);
			384: out = 16'(396);
			385: out = 16'(3801);
			386: out = 16'(-3625);
			387: out = 16'(-22869);
			388: out = 16'(-32765);
			389: out = 16'(-23203);
			390: out = 16'(-7357);
			391: out = 16'(-3061);
			392: out = 16'(-14964);
			393: out = 16'(-24996);
			394: out = 16'(-22775);
			395: out = 16'(-15353);
			396: out = 16'(1723);
			397: out = 16'(-945);
			398: out = 16'(-15801);
			399: out = 16'(-25848);
			400: out = 16'(-22260);
			401: out = 16'(-14651);
			402: out = 16'(-15588);
			403: out = 16'(-24693);
			404: out = 16'(-29749);
			405: out = 16'(-31521);
			406: out = 16'(-28697);
			407: out = 16'(-23312);
			408: out = 16'(-29064);
			409: out = 16'(-27999);
			410: out = 16'(-18381);
			411: out = 16'(-16008);
			412: out = 16'(-27936);
			413: out = 16'(-29811);
			414: out = 16'(-21324);
			415: out = 16'(-23201);
			416: out = 16'(-30966);
			417: out = 16'(-29772);
			418: out = 16'(-25183);
			419: out = 16'(-25042);
			420: out = 16'(-29694);
			421: out = 16'(-30568);
			422: out = 16'(-31030);
			423: out = 16'(-19889);
			424: out = 16'(-19788);
			425: out = 16'(-31335);
			426: out = 16'(-30216);
			427: out = 16'(-31265);
			428: out = 16'(-30024);
			429: out = 16'(-29827);
			430: out = 16'(-21306);
			431: out = 16'(-20912);
			432: out = 16'(-30245);
			433: out = 16'(-30595);
			434: out = 16'(-30533);
			435: out = 16'(-26270);
			436: out = 16'(-18594);
			437: out = 16'(-25373);
			438: out = 16'(-31005);
			439: out = 16'(-30288);
			440: out = 16'(-30593);
			441: out = 16'(-30241);
			442: out = 16'(-30383);
			443: out = 16'(-30461);
			444: out = 16'(-29460);
			445: out = 16'(-18591);
			446: out = 16'(-11599);
			447: out = 16'(-25237);
			448: out = 16'(-30528);
			449: out = 16'(-30559);
			450: out = 16'(-27559);
			451: out = 16'(-28368);
			452: out = 16'(-29078);
			453: out = 16'(-21682);
			454: out = 16'(-21509);
			455: out = 16'(-27315);
			456: out = 16'(-30506);
			457: out = 16'(-30055);
			458: out = 16'(-29048);
			459: out = 16'(-18718);
			460: out = 16'(-9507);
			461: out = 16'(-20288);
			462: out = 16'(-30835);
			463: out = 16'(-29637);
			464: out = 16'(-29409);
			465: out = 16'(-15570);
			466: out = 16'(-11196);
			467: out = 16'(-24280);
			468: out = 16'(-30307);
			469: out = 16'(-29799);
			470: out = 16'(-24622);
			471: out = 16'(-17184);
			472: out = 16'(-17672);
			473: out = 16'(-23729);
			474: out = 16'(-21417);
			475: out = 16'(-6639);
			476: out = 16'(-10843);
			477: out = 16'(-27250);
			478: out = 16'(-30261);
			479: out = 16'(-25977);
			480: out = 16'(-12737);
			481: out = 16'(-593);
			482: out = 16'(628);
			483: out = 16'(-11189);
			484: out = 16'(-20699);
			485: out = 16'(-26772);
			486: out = 16'(-24662);
			487: out = 16'(-8816);
			488: out = 16'(2611);
			489: out = 16'(-3184);
			490: out = 16'(-4563);
			491: out = 16'(-2422);
			492: out = 16'(-4679);
			493: out = 16'(-5628);
			494: out = 16'(-10322);
			495: out = 16'(-9603);
			496: out = 16'(3589);
			497: out = 16'(15237);
			498: out = 16'(2736);
			499: out = 16'(-9575);
			500: out = 16'(1156);
			501: out = 16'(12401);
			502: out = 16'(7693);
			503: out = 16'(6312);
			504: out = 16'(14380);
			505: out = 16'(12172);
			506: out = 16'(4826);
			507: out = 16'(8001);
			508: out = 16'(9843);
			509: out = 16'(19542);
			510: out = 16'(20774);
			511: out = 16'(15713);
			512: out = 16'(23271);
			513: out = 16'(28646);
			514: out = 16'(30151);
			515: out = 16'(23198);
			516: out = 16'(19789);
			517: out = 16'(22485);
			518: out = 16'(21873);
			519: out = 16'(27261);
			520: out = 16'(31498);
			521: out = 16'(30492);
			522: out = 16'(27522);
			523: out = 16'(29563);
			524: out = 16'(28838);
			525: out = 16'(21481);
			526: out = 16'(20517);
			527: out = 16'(21860);
			528: out = 16'(27106);
			529: out = 16'(31432);
			530: out = 16'(30888);
			531: out = 16'(30429);
			532: out = 16'(27318);
			533: out = 16'(30708);
			534: out = 16'(30860);
			535: out = 16'(30946);
			536: out = 16'(30860);
			537: out = 16'(30935);
			538: out = 16'(30760);
			539: out = 16'(30832);
			540: out = 16'(30724);
			541: out = 16'(30766);
			542: out = 16'(30725);
			543: out = 16'(30723);
			544: out = 16'(30672);
			545: out = 16'(30677);
			546: out = 16'(30640);
			547: out = 16'(30630);
			548: out = 16'(30578);
			549: out = 16'(30530);
			550: out = 16'(30595);
			551: out = 16'(30475);
			552: out = 16'(30649);
			553: out = 16'(28738);
			554: out = 16'(21977);
			555: out = 16'(24677);
			556: out = 16'(30919);
			557: out = 16'(30069);
			558: out = 16'(30813);
			559: out = 16'(27921);
			560: out = 16'(21298);
			561: out = 16'(26613);
			562: out = 16'(30762);
			563: out = 16'(29958);
			564: out = 16'(30716);
			565: out = 16'(27736);
			566: out = 16'(26807);
			567: out = 16'(30892);
			568: out = 16'(29611);
			569: out = 16'(30895);
			570: out = 16'(26811);
			571: out = 16'(23132);
			572: out = 16'(29403);
			573: out = 16'(30000);
			574: out = 16'(30142);
			575: out = 16'(29890);
			576: out = 16'(30107);
			577: out = 16'(29856);
			578: out = 16'(30119);
			579: out = 16'(29719);
			580: out = 16'(30081);
			581: out = 16'(23172);
			582: out = 16'(18245);
			583: out = 16'(22195);
			584: out = 16'(23283);
			585: out = 16'(18859);
			586: out = 16'(18220);
			587: out = 16'(22364);
			588: out = 16'(19088);
			589: out = 16'(10336);
			590: out = 16'(9300);
			591: out = 16'(13053);
			592: out = 16'(24879);
			593: out = 16'(30231);
			594: out = 16'(28559);
			595: out = 16'(17029);
			596: out = 16'(9585);
			597: out = 16'(13548);
			598: out = 16'(25450);
			599: out = 16'(23019);
			600: out = 16'(15219);
			601: out = 16'(17327);
			602: out = 16'(20030);
			603: out = 16'(15143);
			604: out = 16'(6589);
			605: out = 16'(3564);
			606: out = 16'(11176);
			607: out = 16'(19139);
			608: out = 16'(10244);
			609: out = 16'(4297);
			610: out = 16'(6624);
			611: out = 16'(20813);
			612: out = 16'(15590);
			613: out = 16'(3310);
			614: out = 16'(6722);
			615: out = 16'(12023);
			616: out = 16'(9658);
			617: out = 16'(9719);
			618: out = 16'(13577);
			619: out = 16'(12237);
			620: out = 16'(-2812);
			621: out = 16'(-12039);
			622: out = 16'(-6172);
			623: out = 16'(1062);
			624: out = 16'(3153);
			625: out = 16'(-4572);
			626: out = 16'(-7563);
			627: out = 16'(-8346);
			628: out = 16'(-4328);
			629: out = 16'(-1768);
			630: out = 16'(-3040);
			631: out = 16'(2912);
			632: out = 16'(-491);
			633: out = 16'(-2526);
			634: out = 16'(-6321);
			635: out = 16'(-12252);
			636: out = 16'(-10437);
			637: out = 16'(-7522);
			638: out = 16'(-5366);
			639: out = 16'(-12933);
			640: out = 16'(-14276);
			641: out = 16'(-9204);
			642: out = 16'(-8485);
			643: out = 16'(-23647);
			644: out = 16'(-32257);
			645: out = 16'(-29904);
			646: out = 16'(-16051);
			647: out = 16'(-9916);
			648: out = 16'(-25517);
			649: out = 16'(-32164);
			650: out = 16'(-26059);
			651: out = 16'(-15698);
			652: out = 16'(-18036);
			653: out = 16'(-27668);
			654: out = 16'(-31813);
			655: out = 16'(-31140);
			656: out = 16'(-31525);
			657: out = 16'(-31332);
			658: out = 16'(-31199);
			659: out = 16'(-30085);
			660: out = 16'(-27097);
			661: out = 16'(-26970);
			662: out = 16'(-23963);
			663: out = 16'(-29077);
			664: out = 16'(-31682);
			665: out = 16'(-31035);
			666: out = 16'(-29862);
			667: out = 16'(-25375);
			668: out = 16'(-28460);
			669: out = 16'(-31147);
			670: out = 16'(-31133);
			671: out = 16'(-30995);
			672: out = 16'(-31135);
			673: out = 16'(-31006);
			674: out = 16'(-31047);
			675: out = 16'(-30904);
			676: out = 16'(-31009);
			677: out = 16'(-30522);
			678: out = 16'(-29572);
			679: out = 16'(-30966);
			680: out = 16'(-30867);
			681: out = 16'(-30842);
			682: out = 16'(-30752);
			683: out = 16'(-30775);
			684: out = 16'(-30717);
			685: out = 16'(-30703);
			686: out = 16'(-30780);
			687: out = 16'(-30754);
			688: out = 16'(-30641);
			689: out = 16'(-30186);
			690: out = 16'(-29039);
			691: out = 16'(-30442);
			692: out = 16'(-30504);
			693: out = 16'(-30789);
			694: out = 16'(-30325);
			695: out = 16'(-30816);
			696: out = 16'(-28026);
			697: out = 16'(-29096);
			698: out = 16'(-30828);
			699: out = 16'(-28736);
			700: out = 16'(-30064);
			701: out = 16'(-30476);
			702: out = 16'(-30345);
			703: out = 16'(-30419);
			704: out = 16'(-29917);
			705: out = 16'(-29102);
			706: out = 16'(-30361);
			707: out = 16'(-30178);
			708: out = 16'(-30281);
			709: out = 16'(-30211);
			710: out = 16'(-30167);
			711: out = 16'(-30214);
			712: out = 16'(-30152);
			713: out = 16'(-30089);
			714: out = 16'(-29958);
			715: out = 16'(-30211);
			716: out = 16'(-26486);
			717: out = 16'(-16133);
			718: out = 16'(-19293);
			719: out = 16'(-29581);
			720: out = 16'(-29834);
			721: out = 16'(-29647);
			722: out = 16'(-22110);
			723: out = 16'(-23300);
			724: out = 16'(-29799);
			725: out = 16'(-27286);
			726: out = 16'(-23433);
			727: out = 16'(-27241);
			728: out = 16'(-30651);
			729: out = 16'(-26898);
			730: out = 16'(-13264);
			731: out = 16'(-13230);
			732: out = 16'(-26047);
			733: out = 16'(-22419);
			734: out = 16'(-15980);
			735: out = 16'(-21934);
			736: out = 16'(-18019);
			737: out = 16'(-10796);
			738: out = 16'(-10135);
			739: out = 16'(-16841);
			740: out = 16'(-16674);
			741: out = 16'(-12733);
			742: out = 16'(2309);
			743: out = 16'(5104);
			744: out = 16'(-9414);
			745: out = 16'(-19955);
			746: out = 16'(-10066);
			747: out = 16'(2446);
			748: out = 16'(-278);
			749: out = 16'(3935);
			750: out = 16'(10107);
			751: out = 16'(4781);
			752: out = 16'(-208);
			753: out = 16'(2630);
			754: out = 16'(-2689);
			755: out = 16'(-2163);
			756: out = 16'(6470);
			757: out = 16'(7590);
			758: out = 16'(13230);
			759: out = 16'(14876);
			760: out = 16'(13010);
			761: out = 16'(10825);
			762: out = 16'(8347);
			763: out = 16'(9158);
			764: out = 16'(9059);
			765: out = 16'(10198);
			766: out = 16'(9836);
			767: out = 16'(19517);
			768: out = 16'(22820);
			769: out = 16'(14083);
			770: out = 16'(9377);
			771: out = 16'(15911);
			772: out = 16'(25046);
			773: out = 16'(29549);
			774: out = 16'(25567);
			775: out = 16'(17183);
			776: out = 16'(9415);
			777: out = 16'(4361);
			778: out = 16'(869);
			779: out = 16'(2617);
			780: out = 16'(18157);
			781: out = 16'(28130);
			782: out = 16'(14536);
			783: out = 16'(9542);
			784: out = 16'(23314);
			785: out = 16'(27224);
			786: out = 16'(12034);
			787: out = 16'(9681);
			788: out = 16'(18343);
			789: out = 16'(16716);
			790: out = 16'(22885);
			791: out = 16'(26361);
			792: out = 16'(21753);
			793: out = 16'(25406);
			794: out = 16'(29274);
			795: out = 16'(28915);
			796: out = 16'(22808);
			797: out = 16'(11867);
			798: out = 16'(10121);
			799: out = 16'(11844);
			800: out = 16'(18243);
			801: out = 16'(27562);
			802: out = 16'(31129);
			803: out = 16'(30746);
			804: out = 16'(31230);
			805: out = 16'(28364);
			806: out = 16'(23209);
			807: out = 16'(20968);
			808: out = 16'(19048);
			809: out = 16'(24122);
			810: out = 16'(24865);
			811: out = 16'(24258);
			812: out = 16'(31176);
			813: out = 16'(26182);
			814: out = 16'(18797);
			815: out = 16'(22267);
			816: out = 16'(28509);
			817: out = 16'(31288);
			818: out = 16'(24525);
			819: out = 16'(12979);
			820: out = 16'(15475);
			821: out = 16'(29417);
			822: out = 16'(28609);
			823: out = 16'(20517);
			824: out = 16'(23050);
			825: out = 16'(27799);
			826: out = 16'(23875);
			827: out = 16'(16605);
			828: out = 16'(21405);
			829: out = 16'(30659);
			830: out = 16'(27210);
			831: out = 16'(13217);
			832: out = 16'(6916);
			833: out = 16'(14952);
			834: out = 16'(22604);
			835: out = 16'(14798);
			836: out = 16'(2957);
			837: out = 16'(10378);
			838: out = 16'(22012);
			839: out = 16'(24843);
			840: out = 16'(20172);
			841: out = 16'(17642);
			842: out = 16'(13565);
			843: out = 16'(8687);
			844: out = 16'(17661);
			845: out = 16'(18309);
			846: out = 16'(9199);
			847: out = 16'(14745);
			848: out = 16'(26416);
			849: out = 16'(25255);
			850: out = 16'(6574);
			851: out = 16'(-4149);
			852: out = 16'(10576);
			853: out = 16'(28030);
			854: out = 16'(29450);
			855: out = 16'(19935);
			856: out = 16'(11733);
			857: out = 16'(7214);
			858: out = 16'(4296);
			859: out = 16'(1106);
			860: out = 16'(10716);
			861: out = 16'(20558);
			862: out = 16'(14810);
			863: out = 16'(13112);
			864: out = 16'(13685);
			865: out = 16'(13072);
			866: out = 16'(6458);
			867: out = 16'(-2880);
			868: out = 16'(-2396);
			869: out = 16'(2429);
			870: out = 16'(7507);
			871: out = 16'(9848);
			872: out = 16'(8098);
			873: out = 16'(2872);
			874: out = 16'(1481);
			875: out = 16'(1612);
			876: out = 16'(10050);
			877: out = 16'(6288);
			878: out = 16'(-6864);
			879: out = 16'(-12592);
			880: out = 16'(-9944);
			881: out = 16'(-6787);
			882: out = 16'(-3454);
			883: out = 16'(-8482);
			884: out = 16'(-11667);
			885: out = 16'(-8077);
			886: out = 16'(-2912);
			887: out = 16'(6857);
			888: out = 16'(17990);
			889: out = 16'(13892);
			890: out = 16'(-5567);
			891: out = 16'(-18618);
			892: out = 16'(-19215);
			893: out = 16'(-10752);
			894: out = 16'(-9707);
			895: out = 16'(-12689);
			896: out = 16'(-3966);
			897: out = 16'(-62);
			898: out = 16'(6740);
			899: out = 16'(11037);
			900: out = 16'(1129);
			901: out = 16'(-7221);
			902: out = 16'(-13158);
			903: out = 16'(-16652);
			904: out = 16'(-15400);
			905: out = 16'(-6293);
			906: out = 16'(-3816);
			907: out = 16'(-6293);
			908: out = 16'(-14431);
			909: out = 16'(-20197);
			910: out = 16'(-4894);
			911: out = 16'(11307);
			912: out = 16'(5558);
			913: out = 16'(-15578);
			914: out = 16'(-24499);
			915: out = 16'(-25079);
			916: out = 16'(-3915);
			917: out = 16'(13395);
			918: out = 16'(-2066);
			919: out = 16'(-14035);
			920: out = 16'(-12082);
			921: out = 16'(-2394);
			922: out = 16'(5564);
			923: out = 16'(-2139);
			924: out = 16'(-9438);
			925: out = 16'(-10347);
			926: out = 16'(-7754);
			927: out = 16'(1527);
			928: out = 16'(1367);
			929: out = 16'(-15873);
			930: out = 16'(-28068);
			931: out = 16'(-23528);
			932: out = 16'(-11488);
			933: out = 16'(-5919);
			934: out = 16'(-13941);
			935: out = 16'(-23482);
			936: out = 16'(-19585);
			937: out = 16'(-3180);
			938: out = 16'(1323);
			939: out = 16'(3358);
			940: out = 16'(1921);
			941: out = 16'(-12353);
			942: out = 16'(-22176);
			943: out = 16'(-27709);
			944: out = 16'(-13368);
			945: out = 16'(2319);
			946: out = 16'(-2210);
			947: out = 16'(-9224);
			948: out = 16'(-14597);
			949: out = 16'(-15791);
			950: out = 16'(-11964);
			951: out = 16'(-16410);
			952: out = 16'(-16361);
			953: out = 16'(-4427);
			954: out = 16'(2309);
			955: out = 16'(-13190);
			956: out = 16'(-23802);
			957: out = 16'(-20082);
			958: out = 16'(-11578);
			959: out = 16'(-3607);
			960: out = 16'(-335);
			961: out = 16'(-7939);
			962: out = 16'(-11614);
			963: out = 16'(-14472);
			964: out = 16'(-17204);
			965: out = 16'(-17995);
			966: out = 16'(-20182);
			967: out = 16'(-20585);
			968: out = 16'(-13480);
			969: out = 16'(-5550);
			970: out = 16'(-3991);
			971: out = 16'(-17654);
			972: out = 16'(-19297);
			973: out = 16'(-2246);
			974: out = 16'(-860);
			975: out = 16'(-14665);
			976: out = 16'(-21497);
			977: out = 16'(-14195);
			978: out = 16'(-11911);
			979: out = 16'(-17658);
			980: out = 16'(-14748);
			981: out = 16'(-8593);
			982: out = 16'(-5502);
			983: out = 16'(-13013);
			984: out = 16'(-14815);
			985: out = 16'(-10739);
			986: out = 16'(-6149);
			987: out = 16'(3241);
			988: out = 16'(-220);
			989: out = 16'(-16765);
			990: out = 16'(-28897);
			991: out = 16'(-24098);
			992: out = 16'(-17930);
			993: out = 16'(-3844);
			994: out = 16'(6116);
			995: out = 16'(-3953);
			996: out = 16'(-12572);
			997: out = 16'(-17390);
			998: out = 16'(-17687);
			999: out = 16'(-9038);
			1000: out = 16'(-8447);
			1001: out = 16'(-11402);
			1002: out = 16'(-17033);
			1003: out = 16'(-7551);
			1004: out = 16'(1906);
			1005: out = 16'(-13045);
			1006: out = 16'(-24723);
			1007: out = 16'(-18481);
			1008: out = 16'(-14169);
			1009: out = 16'(-12647);
			1010: out = 16'(-2232);
			1011: out = 16'(2622);
			1012: out = 16'(-18963);
			1013: out = 16'(-31203);
			1014: out = 16'(-25941);
			1015: out = 16'(-13359);
			1016: out = 16'(7758);
			1017: out = 16'(8388);
			1018: out = 16'(-16728);
			1019: out = 16'(-29216);
			1020: out = 16'(-27055);
			1021: out = 16'(-11120);
			1022: out = 16'(3032);
			1023: out = 16'(-4453);
			1024: out = 16'(-20767);
			1025: out = 16'(-23437);
			1026: out = 16'(-17567);
			1027: out = 16'(-8119);
			1028: out = 16'(-7164);
			1029: out = 16'(-13558);
			1030: out = 16'(-21979);
			1031: out = 16'(-18866);
			1032: out = 16'(-5336);
			1033: out = 16'(-513);
			1034: out = 16'(-6662);
			1035: out = 16'(-11133);
			1036: out = 16'(-12856);
			1037: out = 16'(-13947);
			1038: out = 16'(-8500);
			1039: out = 16'(-8590);
			1040: out = 16'(-16243);
			1041: out = 16'(-24659);
			1042: out = 16'(-21314);
			1043: out = 16'(-15672);
			1044: out = 16'(-10502);
			1045: out = 16'(-15577);
			1046: out = 16'(-21491);
			1047: out = 16'(-15474);
			1048: out = 16'(-10212);
			1049: out = 16'(-838);
			1050: out = 16'(-4442);
			1051: out = 16'(-5885);
			1052: out = 16'(-8632);
			1053: out = 16'(-4705);
			1054: out = 16'(-8951);
			1055: out = 16'(-13495);
			1056: out = 16'(-10683);
			1057: out = 16'(-6716);
			1058: out = 16'(-4423);
			1059: out = 16'(-4817);
			1060: out = 16'(-1326);
			1061: out = 16'(-2361);
			1062: out = 16'(-12020);
			1063: out = 16'(-18626);
			1064: out = 16'(-13394);
			1065: out = 16'(-8330);
			1066: out = 16'(-5965);
			1067: out = 16'(127);
			1068: out = 16'(358);
			1069: out = 16'(-12412);
			1070: out = 16'(-22311);
			1071: out = 16'(-8562);
			1072: out = 16'(15720);
			1073: out = 16'(13496);
			1074: out = 16'(-1487);
			1075: out = 16'(-6680);
			1076: out = 16'(-10751);
			1077: out = 16'(-4069);
			1078: out = 16'(3732);
			1079: out = 16'(5361);
			1080: out = 16'(6355);
			1081: out = 16'(-1735);
			1082: out = 16'(-2132);
			1083: out = 16'(-3944);
			1084: out = 16'(-10340);
			1085: out = 16'(5963);
			1086: out = 16'(17503);
			1087: out = 16'(6783);
			1088: out = 16'(-5591);
			1089: out = 16'(-2901);
			1090: out = 16'(5060);
			1091: out = 16'(2021);
			1092: out = 16'(1514);
			1093: out = 16'(6826);
			1094: out = 16'(3556);
			1095: out = 16'(529);
			1096: out = 16'(-148);
			1097: out = 16'(3328);
			1098: out = 16'(4015);
			1099: out = 16'(8764);
			1100: out = 16'(13578);
			1101: out = 16'(7266);
			1102: out = 16'(741);
			1103: out = 16'(1607);
			1104: out = 16'(6946);
			1105: out = 16'(13831);
			1106: out = 16'(10191);
			1107: out = 16'(1827);
			1108: out = 16'(5666);
			1109: out = 16'(7895);
			1110: out = 16'(15560);
			1111: out = 16'(15575);
			1112: out = 16'(1658);
			1113: out = 16'(2909);
			1114: out = 16'(5990);
			1115: out = 16'(4510);
			1116: out = 16'(5872);
			1117: out = 16'(1936);
			1118: out = 16'(-1399);
			1119: out = 16'(-554);
			1120: out = 16'(944);
			1121: out = 16'(-2461);
			1122: out = 16'(5326);
			1123: out = 16'(10109);
			1124: out = 16'(11848);
			1125: out = 16'(17424);
			1126: out = 16'(17586);
			1127: out = 16'(9240);
			1128: out = 16'(-5582);
			1129: out = 16'(-10448);
			1130: out = 16'(-5088);
			1131: out = 16'(10976);
			1132: out = 16'(11537);
			1133: out = 16'(4900);
			1134: out = 16'(12283);
			1135: out = 16'(12328);
			1136: out = 16'(3296);
			1137: out = 16'(10623);
			1138: out = 16'(11433);
			1139: out = 16'(6075);
			1140: out = 16'(6651);
			1141: out = 16'(13447);
			1142: out = 16'(11283);
			1143: out = 16'(670);
			1144: out = 16'(-4833);
			1145: out = 16'(2488);
			1146: out = 16'(12470);
			1147: out = 16'(15649);
			1148: out = 16'(9942);
			1149: out = 16'(5796);
			1150: out = 16'(-1008);
			1151: out = 16'(-1237);
			1152: out = 16'(-1483);
			1153: out = 16'(3327);
			1154: out = 16'(19716);
			1155: out = 16'(21704);
			1156: out = 16'(13056);
			1157: out = 16'(10769);
			1158: out = 16'(11226);
			1159: out = 16'(14141);
			1160: out = 16'(5425);
			1161: out = 16'(-1205);
			1162: out = 16'(106);
			1163: out = 16'(6090);
			1164: out = 16'(14555);
			1165: out = 16'(19834);
			1166: out = 16'(7254);
			1167: out = 16'(-1714);
			1168: out = 16'(-1549);
			1169: out = 16'(6279);
			1170: out = 16'(14898);
			1171: out = 16'(14321);
			1172: out = 16'(4719);
			1173: out = 16'(-4561);
			1174: out = 16'(3445);
			1175: out = 16'(16281);
			1176: out = 16'(18279);
			1177: out = 16'(3498);
			1178: out = 16'(907);
			1179: out = 16'(9676);
			1180: out = 16'(20229);
			1181: out = 16'(16975);
			1182: out = 16'(4830);
			1183: out = 16'(-2638);
			1184: out = 16'(347);
			1185: out = 16'(3935);
			1186: out = 16'(6038);
			1187: out = 16'(2917);
			1188: out = 16'(-2260);
			1189: out = 16'(1137);
			1190: out = 16'(10279);
			1191: out = 16'(22354);
			1192: out = 16'(28062);
			1193: out = 16'(24037);
			1194: out = 16'(4714);
			1195: out = 16'(-11314);
			1196: out = 16'(-12553);
			1197: out = 16'(388);
			1198: out = 16'(27322);
			1199: out = 16'(30143);
			1200: out = 16'(11723);
			1201: out = 16'(6503);
			1202: out = 16'(17115);
			1203: out = 16'(28767);
			1204: out = 16'(22485);
			1205: out = 16'(6034);
			1206: out = 16'(6616);
			1207: out = 16'(8121);
			1208: out = 16'(4322);
			1209: out = 16'(9500);
			1210: out = 16'(12768);
			1211: out = 16'(6152);
			1212: out = 16'(10961);
			1213: out = 16'(10461);
			1214: out = 16'(7110);
			1215: out = 16'(12065);
			1216: out = 16'(15485);
			1217: out = 16'(23225);
			1218: out = 16'(24333);
			1219: out = 16'(20439);
			1220: out = 16'(16964);
			1221: out = 16'(8964);
			1222: out = 16'(5137);
			1223: out = 16'(2685);
			1224: out = 16'(-3859);
			1225: out = 16'(444);
			1226: out = 16'(12405);
			1227: out = 16'(22950);
			1228: out = 16'(17968);
			1229: out = 16'(14844);
			1230: out = 16'(24021);
			1231: out = 16'(17230);
			1232: out = 16'(3734);
			1233: out = 16'(-1481);
			1234: out = 16'(7210);
			1235: out = 16'(10777);
			1236: out = 16'(11956);
			1237: out = 16'(16465);
			1238: out = 16'(14945);
			1239: out = 16'(15549);
			1240: out = 16'(15259);
			1241: out = 16'(8244);
			1242: out = 16'(-248);
			1243: out = 16'(-6589);
			1244: out = 16'(4783);
			1245: out = 16'(26546);
			1246: out = 16'(26704);
			1247: out = 16'(286);
			1248: out = 16'(-7888);
			1249: out = 16'(4478);
			1250: out = 16'(15846);
			1251: out = 16'(18037);
			1252: out = 16'(6230);
			1253: out = 16'(-2210);
			1254: out = 16'(-4969);
			1255: out = 16'(-799);
			1256: out = 16'(10208);
			1257: out = 16'(19727);
			1258: out = 16'(7264);
			1259: out = 16'(-5975);
			1260: out = 16'(2689);
			1261: out = 16'(6080);
			1262: out = 16'(8326);
			1263: out = 16'(9746);
			1264: out = 16'(2311);
			1265: out = 16'(-478);
			1266: out = 16'(3144);
			1267: out = 16'(11066);
			1268: out = 16'(13419);
			1269: out = 16'(5366);
			1270: out = 16'(-3125);
			1271: out = 16'(-6316);
			1272: out = 16'(-6346);
			1273: out = 16'(-146);
			1274: out = 16'(-1260);
			1275: out = 16'(-2226);
			1276: out = 16'(14569);
			1277: out = 16'(23890);
			1278: out = 16'(-650);
			1279: out = 16'(-22871);
			1280: out = 16'(-20218);
			1281: out = 16'(-5600);
			1282: out = 16'(10174);
			1283: out = 16'(20904);
			1284: out = 16'(11509);
			1285: out = 16'(-11001);
			1286: out = 16'(-17914);
			1287: out = 16'(-7440);
			1288: out = 16'(5037);
			1289: out = 16'(8521);
			1290: out = 16'(-1114);
			1291: out = 16'(-9525);
			1292: out = 16'(-10771);
			1293: out = 16'(-8081);
			1294: out = 16'(-112);
			1295: out = 16'(10097);
			1296: out = 16'(1221);
			1297: out = 16'(-14408);
			1298: out = 16'(-6881);
			1299: out = 16'(-5023);
			1300: out = 16'(5100);
			1301: out = 16'(3866);
			1302: out = 16'(-3675);
			1303: out = 16'(-4604);
			1304: out = 16'(-2054);
			1305: out = 16'(-4260);
			1306: out = 16'(-8985);
			1307: out = 16'(-12307);
			1308: out = 16'(-15423);
			1309: out = 16'(-9204);
			1310: out = 16'(819);
			1311: out = 16'(-2630);
			1312: out = 16'(-13533);
			1313: out = 16'(-23823);
			1314: out = 16'(-27742);
			1315: out = 16'(-17483);
			1316: out = 16'(110);
			1317: out = 16'(496);
			1318: out = 16'(-19600);
			1319: out = 16'(-26412);
			1320: out = 16'(-20329);
			1321: out = 16'(-11913);
			1322: out = 16'(4237);
			1323: out = 16'(-733);
			1324: out = 16'(-12594);
			1325: out = 16'(-20263);
			1326: out = 16'(-15998);
			1327: out = 16'(-3882);
			1328: out = 16'(-4328);
			1329: out = 16'(-14374);
			1330: out = 16'(-12232);
			1331: out = 16'(-8671);
			1332: out = 16'(-19143);
			1333: out = 16'(-25758);
			1334: out = 16'(-20688);
			1335: out = 16'(-5858);
			1336: out = 16'(-12507);
			1337: out = 16'(-29016);
			1338: out = 16'(-22468);
			1339: out = 16'(-13059);
			1340: out = 16'(-16545);
			1341: out = 16'(-20147);
			1342: out = 16'(-18169);
			1343: out = 16'(-15885);
			1344: out = 16'(-8458);
			1345: out = 16'(-12479);
			1346: out = 16'(-20147);
			1347: out = 16'(-24836);
			1348: out = 16'(-20542);
			1349: out = 16'(-10324);
			1350: out = 16'(-6972);
			1351: out = 16'(-3900);
			1352: out = 16'(-12650);
			1353: out = 16'(-24213);
			1354: out = 16'(-31378);
			1355: out = 16'(-23241);
			1356: out = 16'(-9857);
			1357: out = 16'(-17702);
			1358: out = 16'(-30200);
			1359: out = 16'(-24485);
			1360: out = 16'(-19195);
			1361: out = 16'(-20991);
			1362: out = 16'(-16306);
			1363: out = 16'(-11374);
			1364: out = 16'(-17254);
			1365: out = 16'(-25941);
			1366: out = 16'(-26695);
			1367: out = 16'(-29024);
			1368: out = 16'(-22035);
			1369: out = 16'(-9860);
			1370: out = 16'(-9751);
			1371: out = 16'(-9684);
			1372: out = 16'(-11863);
			1373: out = 16'(-21025);
			1374: out = 16'(-26317);
			1375: out = 16'(-30241);
			1376: out = 16'(-29567);
			1377: out = 16'(-30348);
			1378: out = 16'(-20900);
			1379: out = 16'(-6435);
			1380: out = 16'(-11764);
			1381: out = 16'(-22298);
			1382: out = 16'(-27487);
			1383: out = 16'(-24156);
			1384: out = 16'(-14306);
			1385: out = 16'(-4628);
			1386: out = 16'(-9432);
			1387: out = 16'(-22819);
			1388: out = 16'(-27548);
			1389: out = 16'(-25242);
			1390: out = 16'(-14902);
			1391: out = 16'(-20772);
			1392: out = 16'(-30155);
			1393: out = 16'(-29186);
			1394: out = 16'(-25299);
			1395: out = 16'(-16470);
			1396: out = 16'(-9422);
			1397: out = 16'(-9979);
			1398: out = 16'(-17094);
			1399: out = 16'(-27015);
			1400: out = 16'(-17330);
			1401: out = 16'(-12763);
			1402: out = 16'(-1850);
			1403: out = 16'(264);
			1404: out = 16'(-14370);
			1405: out = 16'(-22155);
			1406: out = 16'(-22405);
			1407: out = 16'(-15683);
			1408: out = 16'(-9558);
			1409: out = 16'(-17371);
			1410: out = 16'(-21091);
			1411: out = 16'(-15654);
			1412: out = 16'(-12521);
			1413: out = 16'(-8652);
			1414: out = 16'(-10334);
			1415: out = 16'(-17688);
			1416: out = 16'(-20146);
			1417: out = 16'(-18037);
			1418: out = 16'(-9744);
			1419: out = 16'(-12773);
			1420: out = 16'(-17904);
			1421: out = 16'(-2600);
			1422: out = 16'(-644);
			1423: out = 16'(-20534);
			1424: out = 16'(-23080);
			1425: out = 16'(-8391);
			1426: out = 16'(-7364);
			1427: out = 16'(-11008);
			1428: out = 16'(-11154);
			1429: out = 16'(-17049);
			1430: out = 16'(-7207);
			1431: out = 16'(11984);
			1432: out = 16'(1716);
			1433: out = 16'(-7176);
			1434: out = 16'(-8354);
			1435: out = 16'(9881);
			1436: out = 16'(7422);
			1437: out = 16'(-5796);
			1438: out = 16'(4340);
			1439: out = 16'(15506);
			1440: out = 16'(4015);
			1441: out = 16'(-18221);
			1442: out = 16'(-14324);
			1443: out = 16'(-1489);
			1444: out = 16'(4466);
			1445: out = 16'(-3388);
			1446: out = 16'(-3773);
			1447: out = 16'(3841);
			1448: out = 16'(14273);
			1449: out = 16'(12698);
			1450: out = 16'(467);
			1451: out = 16'(-4271);
			1452: out = 16'(-491);
			1453: out = 16'(11035);
			1454: out = 16'(7808);
			1455: out = 16'(5095);
			1456: out = 16'(13164);
			1457: out = 16'(15645);
			1458: out = 16'(3345);
			1459: out = 16'(-10196);
			1460: out = 16'(-3798);
			1461: out = 16'(9732);
			1462: out = 16'(12851);
			1463: out = 16'(16873);
			1464: out = 16'(23083);
			1465: out = 16'(14932);
			1466: out = 16'(-251);
			1467: out = 16'(-1511);
			1468: out = 16'(-522);
			1469: out = 16'(8284);
			1470: out = 16'(21524);
			1471: out = 16'(15306);
			1472: out = 16'(2247);
			1473: out = 16'(6896);
			1474: out = 16'(9523);
			1475: out = 16'(19230);
			1476: out = 16'(18325);
			1477: out = 16'(9656);
			1478: out = 16'(3329);
			1479: out = 16'(4305);
			1480: out = 16'(20098);
			1481: out = 16'(24078);
			1482: out = 16'(19198);
			1483: out = 16'(18904);
			1484: out = 16'(12196);
			1485: out = 16'(162);
			1486: out = 16'(3271);
			1487: out = 16'(5295);
			1488: out = 16'(8442);
			1489: out = 16'(15485);
			1490: out = 16'(18436);
			1491: out = 16'(17829);
			1492: out = 16'(24693);
			1493: out = 16'(30978);
			1494: out = 16'(18772);
			1495: out = 16'(6534);
			1496: out = 16'(4683);
			1497: out = 16'(16532);
			1498: out = 16'(26644);
			1499: out = 16'(21066);
			1500: out = 16'(19988);
			1501: out = 16'(25262);
			1502: out = 16'(23030);
			1503: out = 16'(5671);
			1504: out = 16'(-4137);
			1505: out = 16'(5272);
			1506: out = 16'(19953);
			1507: out = 16'(15766);
			1508: out = 16'(9094);
			1509: out = 16'(22232);
			1510: out = 16'(32069);
			1511: out = 16'(20777);
			1512: out = 16'(8892);
			1513: out = 16'(10670);
			1514: out = 16'(16139);
			1515: out = 16'(19152);
			1516: out = 16'(26070);
			1517: out = 16'(30348);
			1518: out = 16'(14818);
			1519: out = 16'(-3061);
			1520: out = 16'(-3723);
			1521: out = 16'(7473);
			1522: out = 16'(17261);
			1523: out = 16'(12588);
			1524: out = 16'(-113);
			1525: out = 16'(7848);
			1526: out = 16'(24571);
			1527: out = 16'(31704);
			1528: out = 16'(27262);
			1529: out = 16'(20292);
			1530: out = 16'(18461);
			1531: out = 16'(11591);
			1532: out = 16'(4403);
			1533: out = 16'(9982);
			1534: out = 16'(17932);
			1535: out = 16'(11108);
			1536: out = 16'(1617);
			1537: out = 16'(5016);
			1538: out = 16'(22665);
			1539: out = 16'(27730);
			1540: out = 16'(16241);
			1541: out = 16'(9546);
			1542: out = 16'(13470);
			1543: out = 16'(6318);
			1544: out = 16'(-1137);
			1545: out = 16'(10042);
			1546: out = 16'(17728);
			1547: out = 16'(9761);
			1548: out = 16'(9262);
			1549: out = 16'(8466);
			1550: out = 16'(11721);
			1551: out = 16'(19551);
			1552: out = 16'(12847);
			1553: out = 16'(2528);
			1554: out = 16'(-294);
			1555: out = 16'(12122);
			1556: out = 16'(24281);
			1557: out = 16'(26982);
			1558: out = 16'(13303);
			1559: out = 16'(8675);
			1560: out = 16'(13562);
			1561: out = 16'(13456);
			1562: out = 16'(6712);
			1563: out = 16'(-4701);
			1564: out = 16'(388);
			1565: out = 16'(14321);
			1566: out = 16'(22356);
			1567: out = 16'(13948);
			1568: out = 16'(-2087);
			1569: out = 16'(-3438);
			1570: out = 16'(3742);
			1571: out = 16'(10035);
			1572: out = 16'(11443);
			1573: out = 16'(785);
			1574: out = 16'(-3182);
			1575: out = 16'(1928);
			1576: out = 16'(17247);
			1577: out = 16'(28395);
			1578: out = 16'(13134);
			1579: out = 16'(-4928);
			1580: out = 16'(-7728);
			1581: out = 16'(1085);
			1582: out = 16'(2603);
			1583: out = 16'(6739);
			1584: out = 16'(9820);
			1585: out = 16'(2459);
			1586: out = 16'(-1317);
			1587: out = 16'(6729);
			1588: out = 16'(5599);
			1589: out = 16'(6098);
			1590: out = 16'(10958);
			1591: out = 16'(13699);
			1592: out = 16'(7905);
			1593: out = 16'(1883);
			1594: out = 16'(675);
			1595: out = 16'(6938);
			1596: out = 16'(18197);
			1597: out = 16'(15237);
			1598: out = 16'(253);
			1599: out = 16'(-4971);
			1600: out = 16'(1820);
			1601: out = 16'(5291);
			1602: out = 16'(-10131);
			1603: out = 16'(-15211);
			1604: out = 16'(-3524);
			1605: out = 16'(8603);
			1606: out = 16'(12850);
			1607: out = 16'(10530);
			1608: out = 16'(9381);
			1609: out = 16'(5521);
			1610: out = 16'(-4305);
			1611: out = 16'(-14768);
			1612: out = 16'(-13897);
			1613: out = 16'(-6687);
			1614: out = 16'(-5083);
			1615: out = 16'(-7250);
			1616: out = 16'(330);
			1617: out = 16'(7213);
			1618: out = 16'(495);
			1619: out = 16'(-6497);
			1620: out = 16'(-13190);
			1621: out = 16'(-10691);
			1622: out = 16'(-6875);
			1623: out = 16'(-8541);
			1624: out = 16'(-446);
			1625: out = 16'(219);
			1626: out = 16'(-7408);
			1627: out = 16'(-18224);
			1628: out = 16'(-22495);
			1629: out = 16'(-6679);
			1630: out = 16'(7908);
			1631: out = 16'(12706);
			1632: out = 16'(6691);
			1633: out = 16'(-10682);
			1634: out = 16'(-18379);
			1635: out = 16'(-17055);
			1636: out = 16'(-8529);
			1637: out = 16'(8476);
			1638: out = 16'(19412);
			1639: out = 16'(-1489);
			1640: out = 16'(-19118);
			1641: out = 16'(-19904);
			1642: out = 16'(-9844);
			1643: out = 16'(-104);
			1644: out = 16'(-2879);
			1645: out = 16'(-11372);
			1646: out = 16'(-11684);
			1647: out = 16'(3598);
			1648: out = 16'(-6180);
			1649: out = 16'(-11523);
			1650: out = 16'(-3991);
			1651: out = 16'(-5007);
			1652: out = 16'(4852);
			1653: out = 16'(4895);
			1654: out = 16'(-3595);
			1655: out = 16'(-7240);
			1656: out = 16'(-12973);
			1657: out = 16'(-9373);
			1658: out = 16'(-5347);
			1659: out = 16'(-7429);
			1660: out = 16'(-9442);
			1661: out = 16'(-11801);
			1662: out = 16'(-12737);
			1663: out = 16'(-5783);
			1664: out = 16'(-3340);
			1665: out = 16'(-6126);
			1666: out = 16'(-6402);
			1667: out = 16'(-8560);
			1668: out = 16'(-11512);
			1669: out = 16'(-19544);
			1670: out = 16'(-23734);
			1671: out = 16'(-12637);
			1672: out = 16'(-2701);
			1673: out = 16'(-5661);
			1674: out = 16'(-3285);
			1675: out = 16'(-102);
			1676: out = 16'(639);
			1677: out = 16'(-14006);
			1678: out = 16'(-23173);
			1679: out = 16'(-14285);
			1680: out = 16'(-13499);
			1681: out = 16'(-10848);
			1682: out = 16'(2060);
			1683: out = 16'(8197);
			1684: out = 16'(-12242);
			1685: out = 16'(-28428);
			1686: out = 16'(-21582);
			1687: out = 16'(-6352);
			1688: out = 16'(4341);
			1689: out = 16'(-5984);
			1690: out = 16'(-20364);
			1691: out = 16'(-18005);
			1692: out = 16'(-15255);
			1693: out = 16'(-4245);
			1694: out = 16'(-3818);
			1695: out = 16'(-15286);
			1696: out = 16'(-17008);
			1697: out = 16'(-15881);
			1698: out = 16'(-8239);
			1699: out = 16'(-14243);
			1700: out = 16'(-8507);
			1701: out = 16'(-2315);
			1702: out = 16'(-1989);
			1703: out = 16'(-387);
			1704: out = 16'(-11461);
			1705: out = 16'(-11173);
			1706: out = 16'(-1596);
			1707: out = 16'(5674);
			1708: out = 16'(-310);
			1709: out = 16'(-11118);
			1710: out = 16'(-17540);
			1711: out = 16'(-14935);
			1712: out = 16'(-13521);
			1713: out = 16'(-11617);
			1714: out = 16'(-14761);
			1715: out = 16'(-13796);
			1716: out = 16'(-10350);
			1717: out = 16'(-6281);
			1718: out = 16'(-19341);
			1719: out = 16'(-16787);
			1720: out = 16'(-4942);
			1721: out = 16'(-90);
			1722: out = 16'(-6602);
			1723: out = 16'(-13024);
			1724: out = 16'(-15904);
			1725: out = 16'(-19044);
			1726: out = 16'(-11825);
			1727: out = 16'(5715);
			1728: out = 16'(11704);
			1729: out = 16'(-2023);
			1730: out = 16'(-17099);
			1731: out = 16'(-15081);
			1732: out = 16'(2258);
			1733: out = 16'(7632);
			1734: out = 16'(-11509);
			1735: out = 16'(-19771);
			1736: out = 16'(-7036);
			1737: out = 16'(7330);
			1738: out = 16'(-6228);
			1739: out = 16'(-21127);
			1740: out = 16'(-9413);
			1741: out = 16'(6937);
			1742: out = 16'(7932);
			1743: out = 16'(-1236);
			1744: out = 16'(-2625);
			1745: out = 16'(-4000);
			1746: out = 16'(-8317);
			1747: out = 16'(-20563);
			1748: out = 16'(-13502);
			1749: out = 16'(1904);
			1750: out = 16'(-8362);
			1751: out = 16'(-28972);
			1752: out = 16'(-18154);
			1753: out = 16'(-5026);
			1754: out = 16'(1250);
			1755: out = 16'(6609);
			1756: out = 16'(9011);
			1757: out = 16'(-9736);
			1758: out = 16'(-22198);
			1759: out = 16'(-17741);
			1760: out = 16'(-7822);
			1761: out = 16'(10135);
			1762: out = 16'(12460);
			1763: out = 16'(-10347);
			1764: out = 16'(-21185);
			1765: out = 16'(-13244);
			1766: out = 16'(-351);
			1767: out = 16'(4346);
			1768: out = 16'(-3846);
			1769: out = 16'(-7656);
			1770: out = 16'(1387);
			1771: out = 16'(10380);
			1772: out = 16'(3692);
			1773: out = 16'(-9630);
			1774: out = 16'(-16701);
			1775: out = 16'(-10138);
			1776: out = 16'(-3121);
			1777: out = 16'(-8834);
			1778: out = 16'(-697);
			1779: out = 16'(784);
			1780: out = 16'(3162);
			1781: out = 16'(8945);
			1782: out = 16'(10223);
			1783: out = 16'(-5459);
			1784: out = 16'(-16272);
			1785: out = 16'(-16266);
			1786: out = 16'(-2285);
			1787: out = 16'(21091);
			1788: out = 16'(10981);
			1789: out = 16'(-15320);
			1790: out = 16'(-8866);
			1791: out = 16'(876);
			1792: out = 16'(1967);
			1793: out = 16'(164);
			1794: out = 16'(3707);
			1795: out = 16'(4272);
			1796: out = 16'(6030);
			1797: out = 16'(14302);
			1798: out = 16'(8647);
			1799: out = 16'(1409);
			1800: out = 16'(-5996);
			1801: out = 16'(-8531);
			1802: out = 16'(-2324);
			1803: out = 16'(14053);
			1804: out = 16'(17746);
			1805: out = 16'(-5101);
			1806: out = 16'(-9716);
			1807: out = 16'(4852);
			1808: out = 16'(10715);
			1809: out = 16'(5601);
			1810: out = 16'(-3413);
			1811: out = 16'(-6702);
			1812: out = 16'(-1947);
			1813: out = 16'(7926);
			1814: out = 16'(12024);
			1815: out = 16'(9491);
			1816: out = 16'(9717);
			1817: out = 16'(2036);
			1818: out = 16'(-174);
			1819: out = 16'(3690);
			1820: out = 16'(4253);
			1821: out = 16'(3483);
			1822: out = 16'(11665);
			1823: out = 16'(9736);
			1824: out = 16'(2352);
			1825: out = 16'(2075);
			1826: out = 16'(9424);
			1827: out = 16'(15862);
			1828: out = 16'(8141);
			1829: out = 16'(10236);
			1830: out = 16'(8303);
			1831: out = 16'(2009);
			1832: out = 16'(-3395);
			1833: out = 16'(1146);
			1834: out = 16'(5071);
			1835: out = 16'(9840);
			1836: out = 16'(12969);
			1837: out = 16'(8784);
			1838: out = 16'(-7396);
			1839: out = 16'(-10835);
			1840: out = 16'(-3219);
			1841: out = 16'(-413);
			1842: out = 16'(10254);
			1843: out = 16'(22018);
			1844: out = 16'(18733);
			1845: out = 16'(925);
			1846: out = 16'(-6616);
			1847: out = 16'(9016);
			1848: out = 16'(22745);
			1849: out = 16'(17074);
			1850: out = 16'(12362);
			1851: out = 16'(13349);
			1852: out = 16'(11689);
			1853: out = 16'(-1035);
			1854: out = 16'(-9623);
			1855: out = 16'(-4605);
			1856: out = 16'(485);
			1857: out = 16'(4970);
			1858: out = 16'(12809);
			1859: out = 16'(13125);
			1860: out = 16'(3867);
			1861: out = 16'(7577);
			1862: out = 16'(10482);
			1863: out = 16'(15521);
			1864: out = 16'(17432);
			1865: out = 16'(17430);
			1866: out = 16'(7718);
			1867: out = 16'(-5237);
			1868: out = 16'(-10602);
			1869: out = 16'(-2793);
			1870: out = 16'(17927);
			1871: out = 16'(27371);
			1872: out = 16'(10032);
			1873: out = 16'(-5352);
			1874: out = 16'(2266);
			1875: out = 16'(11844);
			1876: out = 16'(15629);
			1877: out = 16'(11735);
			1878: out = 16'(634);
			1879: out = 16'(-6966);
			1880: out = 16'(-5881);
			1881: out = 16'(-1587);
			1882: out = 16'(7454);
			1883: out = 16'(5524);
			1884: out = 16'(2996);
			1885: out = 16'(11663);
			1886: out = 16'(17670);
			1887: out = 16'(1794);
			1888: out = 16'(-11228);
			1889: out = 16'(-8809);
			1890: out = 16'(-424);
			1891: out = 16'(13128);
			1892: out = 16'(26984);
			1893: out = 16'(13324);
			1894: out = 16'(-4258);
			1895: out = 16'(-3055);
			1896: out = 16'(1396);
			1897: out = 16'(1755);
			1898: out = 16'(2082);
			1899: out = 16'(-1141);
			1900: out = 16'(-4421);
			1901: out = 16'(5218);
			1902: out = 16'(824);
			1903: out = 16'(-12824);
			1904: out = 16'(773);
			1905: out = 16'(12429);
			1906: out = 16'(12616);
			1907: out = 16'(7651);
			1908: out = 16'(788);
			1909: out = 16'(4979);
			1910: out = 16'(11097);
			1911: out = 16'(9807);
			1912: out = 16'(2973);
			1913: out = 16'(-5824);
			1914: out = 16'(-2579);
			1915: out = 16'(8873);
			1916: out = 16'(13025);
			1917: out = 16'(1713);
			1918: out = 16'(-2943);
			1919: out = 16'(510);
			1920: out = 16'(4436);
			1921: out = 16'(-1192);
			1922: out = 16'(-6346);
			1923: out = 16'(7661);
			1924: out = 16'(18119);
			1925: out = 16'(5545);
			1926: out = 16'(-9296);
			1927: out = 16'(-11663);
			1928: out = 16'(2426);
			1929: out = 16'(5958);
			1930: out = 16'(-694);
			1931: out = 16'(1312);
			1932: out = 16'(1986);
			1933: out = 16'(3858);
			1934: out = 16'(6877);
			1935: out = 16'(12543);
			1936: out = 16'(15520);
			1937: out = 16'(3697);
			1938: out = 16'(-9143);
			1939: out = 16'(-8219);
			1940: out = 16'(-5944);
			1941: out = 16'(1993);
			1942: out = 16'(6930);
			1943: out = 16'(-8759);
			1944: out = 16'(-15474);
			1945: out = 16'(1731);
			1946: out = 16'(15824);
			1947: out = 16'(9969);
			1948: out = 16'(11048);
			1949: out = 16'(15138);
			1950: out = 16'(6090);
			1951: out = 16'(-6967);
			1952: out = 16'(-15374);
			1953: out = 16'(-7590);
			1954: out = 16'(7201);
			1955: out = 16'(15517);
			1956: out = 16'(16);
			1957: out = 16'(-8349);
			1958: out = 16'(2291);
			1959: out = 16'(12793);
			1960: out = 16'(14351);
			1961: out = 16'(6464);
			1962: out = 16'(-4798);
			1963: out = 16'(-6884);
			1964: out = 16'(2332);
			1965: out = 16'(11547);
			1966: out = 16'(12839);
			1967: out = 16'(10774);
			1968: out = 16'(5183);
			1969: out = 16'(9098);
			1970: out = 16'(6402);
			1971: out = 16'(3467);
			1972: out = 16'(2014);
			1973: out = 16'(5038);
			1974: out = 16'(9371);
			1975: out = 16'(963);
			1976: out = 16'(4381);
			1977: out = 16'(15414);
			1978: out = 16'(10273);
			1979: out = 16'(-10652);
			1980: out = 16'(-15282);
			1981: out = 16'(-6902);
			1982: out = 16'(-2781);
			1983: out = 16'(-915);
			1984: out = 16'(2823);
			1985: out = 16'(-2946);
			1986: out = 16'(844);
			1987: out = 16'(5106);
			1988: out = 16'(5763);
			1989: out = 16'(-5864);
			1990: out = 16'(-9789);
			1991: out = 16'(-2967);
			1992: out = 16'(-262);
			1993: out = 16'(12979);
			1994: out = 16'(12718);
			1995: out = 16'(11699);
			1996: out = 16'(5216);
			1997: out = 16'(2020);
			1998: out = 16'(4735);
			1999: out = 16'(402);
			2000: out = 16'(217);
			2001: out = 16'(5709);
			2002: out = 16'(2683);
			2003: out = 16'(-375);
			2004: out = 16'(-4668);
			2005: out = 16'(-10348);
			2006: out = 16'(-3781);
			2007: out = 16'(-5320);
			2008: out = 16'(-8326);
			2009: out = 16'(2150);
			2010: out = 16'(3042);
			2011: out = 16'(-2536);
			2012: out = 16'(-7257);
			2013: out = 16'(-1456);
			2014: out = 16'(-875);
			2015: out = 16'(-7898);
			2016: out = 16'(3321);
			2017: out = 16'(12977);
			2018: out = 16'(5531);
			2019: out = 16'(-5288);
			2020: out = 16'(-464);
			2021: out = 16'(2840);
			2022: out = 16'(1886);
			2023: out = 16'(-12632);
			2024: out = 16'(-13599);
			2025: out = 16'(-8419);
			2026: out = 16'(-141);
			2027: out = 16'(-674);
			2028: out = 16'(-10683);
			2029: out = 16'(-10409);
			2030: out = 16'(-4862);
			2031: out = 16'(-3189);
			2032: out = 16'(-12786);
			2033: out = 16'(-4598);
			2034: out = 16'(-2258);
			2035: out = 16'(-3031);
			2036: out = 16'(7983);
			2037: out = 16'(8552);
			2038: out = 16'(-565);
			2039: out = 16'(-9186);
			2040: out = 16'(-10266);
			2041: out = 16'(-7967);
			2042: out = 16'(-12851);
			2043: out = 16'(-9769);
			2044: out = 16'(-4557);
			2045: out = 16'(-9343);
			2046: out = 16'(-10149);
			2047: out = 16'(-5201);
			2048: out = 16'(2252);
			2049: out = 16'(4176);
			2050: out = 16'(1585);
			2051: out = 16'(-4735);
			2052: out = 16'(-7970);
			2053: out = 16'(-3263);
			2054: out = 16'(-3983);
			2055: out = 16'(-4170);
			2056: out = 16'(-12228);
			2057: out = 16'(-19989);
			2058: out = 16'(-18323);
			2059: out = 16'(-14200);
			2060: out = 16'(-1070);
			2061: out = 16'(1596);
			2062: out = 16'(-3901);
			2063: out = 16'(53);
			2064: out = 16'(1759);
			2065: out = 16'(-10499);
			2066: out = 16'(-19962);
			2067: out = 16'(-13986);
			2068: out = 16'(-9468);
			2069: out = 16'(-5118);
			2070: out = 16'(-3773);
			2071: out = 16'(-641);
			2072: out = 16'(985);
			2073: out = 16'(-3078);
			2074: out = 16'(-12001);
			2075: out = 16'(-13047);
			2076: out = 16'(-12860);
			2077: out = 16'(-11225);
			2078: out = 16'(569);
			2079: out = 16'(9001);
			2080: out = 16'(-7906);
			2081: out = 16'(-14522);
			2082: out = 16'(-11473);
			2083: out = 16'(-9714);
			2084: out = 16'(-16538);
			2085: out = 16'(-13554);
			2086: out = 16'(2039);
			2087: out = 16'(-973);
			2088: out = 16'(-6847);
			2089: out = 16'(-12518);
			2090: out = 16'(-10990);
			2091: out = 16'(-5377);
			2092: out = 16'(-3882);
			2093: out = 16'(511);
			2094: out = 16'(-4643);
			2095: out = 16'(-7115);
			2096: out = 16'(-11561);
			2097: out = 16'(-7992);
			2098: out = 16'(5101);
			2099: out = 16'(-2950);
			2100: out = 16'(-10818);
			2101: out = 16'(-8929);
			2102: out = 16'(-4218);
			2103: out = 16'(-7854);
			2104: out = 16'(-16795);
			2105: out = 16'(-15472);
			2106: out = 16'(-7770);
			2107: out = 16'(-2686);
			2108: out = 16'(-6781);
			2109: out = 16'(-3898);
			2110: out = 16'(-6691);
			2111: out = 16'(-6748);
			2112: out = 16'(-10541);
			2113: out = 16'(-8412);
			2114: out = 16'(-9843);
			2115: out = 16'(-14152);
			2116: out = 16'(-15642);
			2117: out = 16'(-15640);
			2118: out = 16'(-5082);
			2119: out = 16'(-5107);
			2120: out = 16'(-8367);
			2121: out = 16'(-13304);
			2122: out = 16'(-13618);
			2123: out = 16'(-11384);
			2124: out = 16'(-3960);
			2125: out = 16'(3331);
			2126: out = 16'(-7815);
			2127: out = 16'(-16159);
			2128: out = 16'(-9723);
			2129: out = 16'(5087);
			2130: out = 16'(-2480);
			2131: out = 16'(-8643);
			2132: out = 16'(-1043);
			2133: out = 16'(-1376);
			2134: out = 16'(-13660);
			2135: out = 16'(-22069);
			2136: out = 16'(-13867);
			2137: out = 16'(-1541);
			2138: out = 16'(-1217);
			2139: out = 16'(-12512);
			2140: out = 16'(-9242);
			2141: out = 16'(-11020);
			2142: out = 16'(-12109);
			2143: out = 16'(-6501);
			2144: out = 16'(-8076);
			2145: out = 16'(-2887);
			2146: out = 16'(-4290);
			2147: out = 16'(-3022);
			2148: out = 16'(-4760);
			2149: out = 16'(-8012);
			2150: out = 16'(-17630);
			2151: out = 16'(-11545);
			2152: out = 16'(-4133);
			2153: out = 16'(-13079);
			2154: out = 16'(-10925);
			2155: out = 16'(623);
			2156: out = 16'(9146);
			2157: out = 16'(2286);
			2158: out = 16'(-2179);
			2159: out = 16'(-6959);
			2160: out = 16'(-3671);
			2161: out = 16'(-3828);
			2162: out = 16'(-10882);
			2163: out = 16'(-7892);
			2164: out = 16'(-8797);
			2165: out = 16'(4671);
			2166: out = 16'(9721);
			2167: out = 16'(1168);
			2168: out = 16'(-7086);
			2169: out = 16'(-7418);
			2170: out = 16'(-9214);
			2171: out = 16'(-6595);
			2172: out = 16'(3708);
			2173: out = 16'(-148);
			2174: out = 16'(-3826);
			2175: out = 16'(-2117);
			2176: out = 16'(9571);
			2177: out = 16'(8984);
			2178: out = 16'(4974);
			2179: out = 16'(1258);
			2180: out = 16'(-4379);
			2181: out = 16'(-10762);
			2182: out = 16'(-14752);
			2183: out = 16'(-1718);
			2184: out = 16'(13447);
			2185: out = 16'(12892);
			2186: out = 16'(940);
			2187: out = 16'(-2446);
			2188: out = 16'(-3361);
			2189: out = 16'(1860);
			2190: out = 16'(12753);
			2191: out = 16'(7986);
			2192: out = 16'(-2642);
			2193: out = 16'(-7786);
			2194: out = 16'(2546);
			2195: out = 16'(15427);
			2196: out = 16'(15937);
			2197: out = 16'(-1963);
			2198: out = 16'(-6812);
			2199: out = 16'(-6886);
			2200: out = 16'(-1705);
			2201: out = 16'(12928);
			2202: out = 16'(14706);
			2203: out = 16'(8891);
			2204: out = 16'(4148);
			2205: out = 16'(4354);
			2206: out = 16'(3830);
			2207: out = 16'(-912);
			2208: out = 16'(2239);
			2209: out = 16'(15977);
			2210: out = 16'(9403);
			2211: out = 16'(-4514);
			2212: out = 16'(-2662);
			2213: out = 16'(11525);
			2214: out = 16'(18202);
			2215: out = 16'(3092);
			2216: out = 16'(5794);
			2217: out = 16'(17787);
			2218: out = 16'(9912);
			2219: out = 16'(864);
			2220: out = 16'(3265);
			2221: out = 16'(5731);
			2222: out = 16'(4786);
			2223: out = 16'(6137);
			2224: out = 16'(7572);
			2225: out = 16'(3293);
			2226: out = 16'(5930);
			2227: out = 16'(10459);
			2228: out = 16'(5633);
			2229: out = 16'(3969);
			2230: out = 16'(14428);
			2231: out = 16'(17569);
			2232: out = 16'(11165);
			2233: out = 16'(7784);
			2234: out = 16'(10051);
			2235: out = 16'(16251);
			2236: out = 16'(14392);
			2237: out = 16'(7467);
			2238: out = 16'(3971);
			2239: out = 16'(1022);
			2240: out = 16'(2789);
			2241: out = 16'(7896);
			2242: out = 16'(8185);
			2243: out = 16'(9076);
			2244: out = 16'(8155);
			2245: out = 16'(11726);
			2246: out = 16'(8060);
			2247: out = 16'(5096);
			2248: out = 16'(794);
			2249: out = 16'(7778);
			2250: out = 16'(14120);
			2251: out = 16'(17359);
			2252: out = 16'(14619);
			2253: out = 16'(-180);
			2254: out = 16'(-4050);
			2255: out = 16'(7695);
			2256: out = 16'(21077);
			2257: out = 16'(15434);
			2258: out = 16'(3558);
			2259: out = 16'(-2918);
			2260: out = 16'(6369);
			2261: out = 16'(15374);
			2262: out = 16'(2800);
			2263: out = 16'(5088);
			2264: out = 16'(11230);
			2265: out = 16'(16487);
			2266: out = 16'(21043);
			2267: out = 16'(16131);
			2268: out = 16'(12726);
			2269: out = 16'(5836);
			2270: out = 16'(-1670);
			2271: out = 16'(-3643);
			2272: out = 16'(5679);
			2273: out = 16'(4845);
			2274: out = 16'(-3803);
			2275: out = 16'(4968);
			2276: out = 16'(16053);
			2277: out = 16'(12503);
			2278: out = 16'(7462);
			2279: out = 16'(-886);
			2280: out = 16'(3638);
			2281: out = 16'(6842);
			2282: out = 16'(13820);
			2283: out = 16'(18213);
			2284: out = 16'(9149);
			2285: out = 16'(7684);
			2286: out = 16'(8485);
			2287: out = 16'(6289);
			2288: out = 16'(-2392);
			2289: out = 16'(-7826);
			2290: out = 16'(2629);
			2291: out = 16'(20621);
			2292: out = 16'(14084);
			2293: out = 16'(-4901);
			2294: out = 16'(-6386);
			2295: out = 16'(8166);
			2296: out = 16'(13985);
			2297: out = 16'(1061);
			2298: out = 16'(-2244);
			2299: out = 16'(10182);
			2300: out = 16'(13495);
			2301: out = 16'(10251);
			2302: out = 16'(11438);
			2303: out = 16'(5919);
			2304: out = 16'(1415);
			2305: out = 16'(1221);
			2306: out = 16'(12888);
			2307: out = 16'(19975);
			2308: out = 16'(4334);
			2309: out = 16'(-9318);
			2310: out = 16'(-6672);
			2311: out = 16'(-282);
			2312: out = 16'(8994);
			2313: out = 16'(-400);
			2314: out = 16'(-7381);
			2315: out = 16'(7442);
			2316: out = 16'(9708);
			2317: out = 16'(-7363);
			2318: out = 16'(-11708);
			2319: out = 16'(-5288);
			2320: out = 16'(5681);
			2321: out = 16'(18624);
			2322: out = 16'(19676);
			2323: out = 16'(5789);
			2324: out = 16'(-685);
			2325: out = 16'(-7129);
			2326: out = 16'(-4076);
			2327: out = 16'(5093);
			2328: out = 16'(8597);
			2329: out = 16'(8338);
			2330: out = 16'(7404);
			2331: out = 16'(-918);
			2332: out = 16'(-11309);
			2333: out = 16'(-6754);
			2334: out = 16'(4662);
			2335: out = 16'(9459);
			2336: out = 16'(11311);
			2337: out = 16'(1299);
			2338: out = 16'(-10321);
			2339: out = 16'(-10357);
			2340: out = 16'(-1384);
			2341: out = 16'(14234);
			2342: out = 16'(9169);
			2343: out = 16'(-3124);
			2344: out = 16'(-1271);
			2345: out = 16'(7560);
			2346: out = 16'(10048);
			2347: out = 16'(5412);
			2348: out = 16'(-586);
			2349: out = 16'(2352);
			2350: out = 16'(-3848);
			2351: out = 16'(-7513);
			2352: out = 16'(-449);
			2353: out = 16'(-3098);
			2354: out = 16'(-10140);
			2355: out = 16'(-8474);
			2356: out = 16'(3252);
			2357: out = 16'(2411);
			2358: out = 16'(3402);
			2359: out = 16'(11836);
			2360: out = 16'(9040);
			2361: out = 16'(-8166);
			2362: out = 16'(-18813);
			2363: out = 16'(-8540);
			2364: out = 16'(8060);
			2365: out = 16'(4173);
			2366: out = 16'(-904);
			2367: out = 16'(-2246);
			2368: out = 16'(-7123);
			2369: out = 16'(-11710);
			2370: out = 16'(-11641);
			2371: out = 16'(-4980);
			2372: out = 16'(4130);
			2373: out = 16'(-336);
			2374: out = 16'(-1508);
			2375: out = 16'(-3716);
			2376: out = 16'(-9372);
			2377: out = 16'(4773);
			2378: out = 16'(15219);
			2379: out = 16'(7584);
			2380: out = 16'(-6630);
			2381: out = 16'(-12862);
			2382: out = 16'(-10678);
			2383: out = 16'(-2751);
			2384: out = 16'(-5331);
			2385: out = 16'(-15375);
			2386: out = 16'(-10567);
			2387: out = 16'(2483);
			2388: out = 16'(-1089);
			2389: out = 16'(-3989);
			2390: out = 16'(-4934);
			2391: out = 16'(1180);
			2392: out = 16'(4754);
			2393: out = 16'(-4038);
			2394: out = 16'(-1158);
			2395: out = 16'(6447);
			2396: out = 16'(6674);
			2397: out = 16'(-5790);
			2398: out = 16'(-12298);
			2399: out = 16'(-4919);
			2400: out = 16'(-2822);
			2401: out = 16'(-18434);
			2402: out = 16'(-14904);
			2403: out = 16'(-145);
			2404: out = 16'(-3751);
			2405: out = 16'(-10933);
			2406: out = 16'(-6903);
			2407: out = 16'(-14984);
			2408: out = 16'(-9550);
			2409: out = 16'(5544);
			2410: out = 16'(9479);
			2411: out = 16'(-4617);
			2412: out = 16'(-20642);
			2413: out = 16'(-18292);
			2414: out = 16'(-3759);
			2415: out = 16'(8490);
			2416: out = 16'(-4561);
			2417: out = 16'(-12793);
			2418: out = 16'(-11057);
			2419: out = 16'(-6001);
			2420: out = 16'(8676);
			2421: out = 16'(3528);
			2422: out = 16'(-7684);
			2423: out = 16'(-5059);
			2424: out = 16'(-6684);
			2425: out = 16'(-6238);
			2426: out = 16'(-7167);
			2427: out = 16'(-9147);
			2428: out = 16'(-6450);
			2429: out = 16'(-10216);
			2430: out = 16'(-11341);
			2431: out = 16'(-4319);
			2432: out = 16'(-5507);
			2433: out = 16'(-15457);
			2434: out = 16'(-6300);
			2435: out = 16'(5257);
			2436: out = 16'(-4826);
			2437: out = 16'(-9984);
			2438: out = 16'(-15276);
			2439: out = 16'(-14656);
			2440: out = 16'(-4996);
			2441: out = 16'(7028);
			2442: out = 16'(10842);
			2443: out = 16'(-8642);
			2444: out = 16'(-25989);
			2445: out = 16'(-18431);
			2446: out = 16'(256);
			2447: out = 16'(9384);
			2448: out = 16'(-3405);
			2449: out = 16'(-5358);
			2450: out = 16'(-5922);
			2451: out = 16'(-1741);
			2452: out = 16'(-901);
			2453: out = 16'(-1732);
			2454: out = 16'(6403);
			2455: out = 16'(6540);
			2456: out = 16'(-4031);
			2457: out = 16'(-9320);
			2458: out = 16'(-9063);
			2459: out = 16'(-3921);
			2460: out = 16'(-5724);
			2461: out = 16'(-8117);
			2462: out = 16'(-9856);
			2463: out = 16'(-4356);
			2464: out = 16'(-4069);
			2465: out = 16'(-5194);
			2466: out = 16'(-6729);
			2467: out = 16'(-2840);
			2468: out = 16'(829);
			2469: out = 16'(-2439);
			2470: out = 16'(-1486);
			2471: out = 16'(-4571);
			2472: out = 16'(-4565);
			2473: out = 16'(-3790);
			2474: out = 16'(-8168);
			2475: out = 16'(-10413);
			2476: out = 16'(-10570);
			2477: out = 16'(-14959);
			2478: out = 16'(-13367);
			2479: out = 16'(-7072);
			2480: out = 16'(-243);
			2481: out = 16'(-1818);
			2482: out = 16'(7239);
			2483: out = 16'(2108);
			2484: out = 16'(-3251);
			2485: out = 16'(-7622);
			2486: out = 16'(-4103);
			2487: out = 16'(2298);
			2488: out = 16'(-1322);
			2489: out = 16'(6304);
			2490: out = 16'(10120);
			2491: out = 16'(-4881);
			2492: out = 16'(-20853);
			2493: out = 16'(-20727);
			2494: out = 16'(-16092);
			2495: out = 16'(3901);
			2496: out = 16'(4430);
			2497: out = 16'(-11845);
			2498: out = 16'(-11108);
			2499: out = 16'(536);
			2500: out = 16'(9441);
			2501: out = 16'(2337);
			2502: out = 16'(4073);
			2503: out = 16'(-849);
			2504: out = 16'(-7861);
			2505: out = 16'(-8991);
			2506: out = 16'(-1302);
			2507: out = 16'(3967);
			2508: out = 16'(6224);
			2509: out = 16'(1592);
			2510: out = 16'(1523);
			2511: out = 16'(4410);
			2512: out = 16'(-5172);
			2513: out = 16'(-7286);
			2514: out = 16'(-2572);
			2515: out = 16'(1362);
			2516: out = 16'(3281);
			2517: out = 16'(-6558);
			2518: out = 16'(-8756);
			2519: out = 16'(452);
			2520: out = 16'(4021);
			2521: out = 16'(3304);
			2522: out = 16'(-2612);
			2523: out = 16'(-11170);
			2524: out = 16'(-5683);
			2525: out = 16'(13);
			2526: out = 16'(6720);
			2527: out = 16'(7400);
			2528: out = 16'(4190);
			2529: out = 16'(-1322);
			2530: out = 16'(-272);
			2531: out = 16'(9878);
			2532: out = 16'(6189);
			2533: out = 16'(-5255);
			2534: out = 16'(-6849);
			2535: out = 16'(-930);
			2536: out = 16'(2283);
			2537: out = 16'(2725);
			2538: out = 16'(7795);
			2539: out = 16'(8046);
			2540: out = 16'(8661);
			2541: out = 16'(2404);
			2542: out = 16'(-8380);
			2543: out = 16'(-1145);
			2544: out = 16'(3020);
			2545: out = 16'(7759);
			2546: out = 16'(9694);
			2547: out = 16'(8827);
			2548: out = 16'(8856);
			2549: out = 16'(2680);
			2550: out = 16'(1205);
			2551: out = 16'(6740);
			2552: out = 16'(6425);
			2553: out = 16'(3042);
			2554: out = 16'(-1913);
			2555: out = 16'(-915);
			2556: out = 16'(8220);
			2557: out = 16'(13530);
			2558: out = 16'(1384);
			2559: out = 16'(-9612);
			2560: out = 16'(-3271);
			2561: out = 16'(205);
			2562: out = 16'(3724);
			2563: out = 16'(3134);
			2564: out = 16'(3268);
			2565: out = 16'(1872);
			2566: out = 16'(11130);
			2567: out = 16'(17886);
			2568: out = 16'(6198);
			2569: out = 16'(-10496);
			2570: out = 16'(-11999);
			2571: out = 16'(-791);
			2572: out = 16'(2786);
			2573: out = 16'(13167);
			2574: out = 16'(13364);
			2575: out = 16'(2287);
			2576: out = 16'(-4075);
			2577: out = 16'(2668);
			2578: out = 16'(5207);
			2579: out = 16'(-1131);
			2580: out = 16'(2315);
			2581: out = 16'(8435);
			2582: out = 16'(14195);
			2583: out = 16'(7452);
			2584: out = 16'(-1956);
			2585: out = 16'(-965);
			2586: out = 16'(7097);
			2587: out = 16'(8657);
			2588: out = 16'(-2415);
			2589: out = 16'(-4506);
			2590: out = 16'(3336);
			2591: out = 16'(-3197);
			2592: out = 16'(4286);
			2593: out = 16'(19198);
			2594: out = 16'(11107);
			2595: out = 16'(-7059);
			2596: out = 16'(-6525);
			2597: out = 16'(5780);
			2598: out = 16'(8654);
			2599: out = 16'(11866);
			2600: out = 16'(5681);
			2601: out = 16'(-4796);
			2602: out = 16'(1422);
			2603: out = 16'(17267);
			2604: out = 16'(21060);
			2605: out = 16'(10289);
			2606: out = 16'(-4046);
			2607: out = 16'(-2742);
			2608: out = 16'(8723);
			2609: out = 16'(11110);
			2610: out = 16'(8094);
			2611: out = 16'(1699);
			2612: out = 16'(-2165);
			2613: out = 16'(938);
			2614: out = 16'(4757);
			2615: out = 16'(-7735);
			2616: out = 16'(-8121);
			2617: out = 16'(2115);
			2618: out = 16'(1887);
			2619: out = 16'(9741);
			2620: out = 16'(15900);
			2621: out = 16'(-2060);
			2622: out = 16'(-14493);
			2623: out = 16'(-2847);
			2624: out = 16'(3367);
			2625: out = 16'(6797);
			2626: out = 16'(11648);
			2627: out = 16'(9590);
			2628: out = 16'(8216);
			2629: out = 16'(5940);
			2630: out = 16'(-1806);
			2631: out = 16'(-217);
			2632: out = 16'(8196);
			2633: out = 16'(9141);
			2634: out = 16'(-6145);
			2635: out = 16'(-12826);
			2636: out = 16'(-2053);
			2637: out = 16'(4574);
			2638: out = 16'(12848);
			2639: out = 16'(6635);
			2640: out = 16'(-1534);
			2641: out = 16'(7805);
			2642: out = 16'(8723);
			2643: out = 16'(292);
			2644: out = 16'(-6082);
			2645: out = 16'(-5818);
			2646: out = 16'(-1018);
			2647: out = 16'(2492);
			2648: out = 16'(11905);
			2649: out = 16'(11064);
			2650: out = 16'(-3679);
			2651: out = 16'(-13117);
			2652: out = 16'(-2489);
			2653: out = 16'(3594);
			2654: out = 16'(5086);
			2655: out = 16'(310);
			2656: out = 16'(-5934);
			2657: out = 16'(-3741);
			2658: out = 16'(-2409);
			2659: out = 16'(8017);
			2660: out = 16'(12642);
			2661: out = 16'(7712);
			2662: out = 16'(4460);
			2663: out = 16'(-5247);
			2664: out = 16'(-11071);
			2665: out = 16'(-1015);
			2666: out = 16'(2866);
			2667: out = 16'(10514);
			2668: out = 16'(11386);
			2669: out = 16'(1750);
			2670: out = 16'(-4345);
			2671: out = 16'(-5893);
			2672: out = 16'(-3803);
			2673: out = 16'(-3881);
			2674: out = 16'(-4007);
			2675: out = 16'(-537);
			2676: out = 16'(3752);
			2677: out = 16'(10311);
			2678: out = 16'(6760);
			2679: out = 16'(10112);
			2680: out = 16'(11799);
			2681: out = 16'(-1518);
			2682: out = 16'(-6076);
			2683: out = 16'(-2317);
			2684: out = 16'(-2638);
			2685: out = 16'(-1003);
			2686: out = 16'(-586);
			2687: out = 16'(775);
			2688: out = 16'(1366);
			2689: out = 16'(-7426);
			2690: out = 16'(-12655);
			2691: out = 16'(-1143);
			2692: out = 16'(7846);
			2693: out = 16'(7815);
			2694: out = 16'(-12122);
			2695: out = 16'(-17243);
			2696: out = 16'(-1070);
			2697: out = 16'(19597);
			2698: out = 16'(22241);
			2699: out = 16'(-416);
			2700: out = 16'(-4983);
			2701: out = 16'(946);
			2702: out = 16'(2764);
			2703: out = 16'(5836);
			2704: out = 16'(5426);
			2705: out = 16'(-4406);
			2706: out = 16'(-9910);
			2707: out = 16'(-6992);
			2708: out = 16'(4566);
			2709: out = 16'(3951);
			2710: out = 16'(-11112);
			2711: out = 16'(-11410);
			2712: out = 16'(-1917);
			2713: out = 16'(6472);
			2714: out = 16'(4082);
			2715: out = 16'(-12951);
			2716: out = 16'(-3262);
			2717: out = 16'(4569);
			2718: out = 16'(8964);
			2719: out = 16'(16002);
			2720: out = 16'(12855);
			2721: out = 16'(-2134);
			2722: out = 16'(-14502);
			2723: out = 16'(-16796);
			2724: out = 16'(-3737);
			2725: out = 16'(5987);
			2726: out = 16'(-258);
			2727: out = 16'(-4816);
			2728: out = 16'(-3444);
			2729: out = 16'(8909);
			2730: out = 16'(7507);
			2731: out = 16'(-3175);
			2732: out = 16'(-757);
			2733: out = 16'(10720);
			2734: out = 16'(5574);
			2735: out = 16'(-6993);
			2736: out = 16'(-4808);
			2737: out = 16'(2313);
			2738: out = 16'(397);
			2739: out = 16'(-7303);
			2740: out = 16'(-4646);
			2741: out = 16'(-1674);
			2742: out = 16'(-2742);
			2743: out = 16'(-1174);
			2744: out = 16'(2828);
			2745: out = 16'(-5962);
			2746: out = 16'(-5762);
			2747: out = 16'(-120);
			2748: out = 16'(-3643);
			2749: out = 16'(-3781);
			2750: out = 16'(4125);
			2751: out = 16'(3530);
			2752: out = 16'(-4613);
			2753: out = 16'(-905);
			2754: out = 16'(-2581);
			2755: out = 16'(3267);
			2756: out = 16'(8965);
			2757: out = 16'(3543);
			2758: out = 16'(6155);
			2759: out = 16'(410);
			2760: out = 16'(-4053);
			2761: out = 16'(-6028);
			2762: out = 16'(-4221);
			2763: out = 16'(4932);
			2764: out = 16'(2882);
			2765: out = 16'(-3905);
			2766: out = 16'(205);
			2767: out = 16'(-485);
			2768: out = 16'(-3139);
			2769: out = 16'(2669);
			2770: out = 16'(853);
			2771: out = 16'(-7377);
			2772: out = 16'(-18772);
			2773: out = 16'(-13754);
			2774: out = 16'(2169);
			2775: out = 16'(12200);
			2776: out = 16'(-1470);
			2777: out = 16'(-16280);
			2778: out = 16'(-7111);
			2779: out = 16'(-785);
			2780: out = 16'(7507);
			2781: out = 16'(4741);
			2782: out = 16'(4009);
			2783: out = 16'(4503);
			2784: out = 16'(2899);
			2785: out = 16'(80);
			2786: out = 16'(-8387);
			2787: out = 16'(-11793);
			2788: out = 16'(-9511);
			2789: out = 16'(-5522);
			2790: out = 16'(-7500);
			2791: out = 16'(-4395);
			2792: out = 16'(-4724);
			2793: out = 16'(630);
			2794: out = 16'(-6970);
			2795: out = 16'(-10883);
			2796: out = 16'(-3408);
			2797: out = 16'(-2077);
			2798: out = 16'(7092);
			2799: out = 16'(11857);
			2800: out = 16'(1101);
			2801: out = 16'(-14186);
			2802: out = 16'(-8320);
			2803: out = 16'(1110);
			2804: out = 16'(6810);
			2805: out = 16'(-4976);
			2806: out = 16'(-11954);
			2807: out = 16'(-8651);
			2808: out = 16'(-6971);
			2809: out = 16'(8);
			2810: out = 16'(-1231);
			2811: out = 16'(-10790);
			2812: out = 16'(-3100);
			2813: out = 16'(8861);
			2814: out = 16'(-918);
			2815: out = 16'(-7674);
			2816: out = 16'(-5757);
			2817: out = 16'(6083);
			2818: out = 16'(352);
			2819: out = 16'(-6734);
			2820: out = 16'(4506);
			2821: out = 16'(12842);
			2822: out = 16'(605);
			2823: out = 16'(-15044);
			2824: out = 16'(-14518);
			2825: out = 16'(-2830);
			2826: out = 16'(-4038);
			2827: out = 16'(-10752);
			2828: out = 16'(-7484);
			2829: out = 16'(-7925);
			2830: out = 16'(-8570);
			2831: out = 16'(-3947);
			2832: out = 16'(-7593);
			2833: out = 16'(-4027);
			2834: out = 16'(7542);
			2835: out = 16'(7923);
			2836: out = 16'(-10965);
			2837: out = 16'(-20702);
			2838: out = 16'(-11492);
			2839: out = 16'(5388);
			2840: out = 16'(16490);
			2841: out = 16'(9562);
			2842: out = 16'(-846);
			2843: out = 16'(-11860);
			2844: out = 16'(-12738);
			2845: out = 16'(-5518);
			2846: out = 16'(2461);
			2847: out = 16'(11959);
			2848: out = 16'(4616);
			2849: out = 16'(-16399);
			2850: out = 16'(-21789);
			2851: out = 16'(-9372);
			2852: out = 16'(1312);
			2853: out = 16'(4674);
			2854: out = 16'(2713);
			2855: out = 16'(-4316);
			2856: out = 16'(-18183);
			2857: out = 16'(-11449);
			2858: out = 16'(-264);
			2859: out = 16'(6838);
			2860: out = 16'(10007);
			2861: out = 16'(-5635);
			2862: out = 16'(-19989);
			2863: out = 16'(-17719);
			2864: out = 16'(-432);
			2865: out = 16'(11599);
			2866: out = 16'(6880);
			2867: out = 16'(6795);
			2868: out = 16'(3829);
			2869: out = 16'(-1258);
			2870: out = 16'(-7828);
			2871: out = 16'(-13746);
			2872: out = 16'(-8285);
			2873: out = 16'(1478);
			2874: out = 16'(8603);
			2875: out = 16'(-305);
			2876: out = 16'(1324);
			2877: out = 16'(-1550);
			2878: out = 16'(5706);
			2879: out = 16'(1505);
			2880: out = 16'(-606);
			2881: out = 16'(1491);
			2882: out = 16'(4553);
			2883: out = 16'(4798);
			2884: out = 16'(-3432);
			2885: out = 16'(-10126);
			2886: out = 16'(-6847);
			2887: out = 16'(-3105);
			2888: out = 16'(-6971);
			2889: out = 16'(-9649);
			2890: out = 16'(-6076);
			2891: out = 16'(1536);
			2892: out = 16'(-2299);
			2893: out = 16'(-15837);
			2894: out = 16'(-20773);
			2895: out = 16'(-5744);
			2896: out = 16'(6000);
			2897: out = 16'(10626);
			2898: out = 16'(6406);
			2899: out = 16'(-6909);
			2900: out = 16'(-9698);
			2901: out = 16'(-6237);
			2902: out = 16'(-2251);
			2903: out = 16'(5884);
			2904: out = 16'(-145);
			2905: out = 16'(-3206);
			2906: out = 16'(5104);
			2907: out = 16'(10698);
			2908: out = 16'(5564);
			2909: out = 16'(-4246);
			2910: out = 16'(-9360);
			2911: out = 16'(-318);
			2912: out = 16'(3647);
			2913: out = 16'(-5662);
			2914: out = 16'(-6654);
			2915: out = 16'(-4881);
			2916: out = 16'(-6675);
			2917: out = 16'(-4494);
			2918: out = 16'(8339);
			2919: out = 16'(3139);
			2920: out = 16'(-6807);
			2921: out = 16'(7802);
			2922: out = 16'(14909);
			2923: out = 16'(8328);
			2924: out = 16'(-6742);
			2925: out = 16'(-9903);
			2926: out = 16'(554);
			2927: out = 16'(6596);
			2928: out = 16'(-684);
			2929: out = 16'(-8136);
			2930: out = 16'(-12834);
			2931: out = 16'(-15005);
			2932: out = 16'(-1899);
			2933: out = 16'(14302);
			2934: out = 16'(11859);
			2935: out = 16'(5560);
			2936: out = 16'(1287);
			2937: out = 16'(-9227);
			2938: out = 16'(-12118);
			2939: out = 16'(3575);
			2940: out = 16'(15406);
			2941: out = 16'(7971);
			2942: out = 16'(-2898);
			2943: out = 16'(-10527);
			2944: out = 16'(-5845);
			2945: out = 16'(7813);
			2946: out = 16'(11339);
			2947: out = 16'(4088);
			2948: out = 16'(6321);
			2949: out = 16'(2401);
			2950: out = 16'(-4527);
			2951: out = 16'(-5092);
			2952: out = 16'(8217);
			2953: out = 16'(16654);
			2954: out = 16'(10649);
			2955: out = 16'(-9584);
			2956: out = 16'(-11143);
			2957: out = 16'(2199);
			2958: out = 16'(18240);
			2959: out = 16'(16280);
			2960: out = 16'(872);
			2961: out = 16'(-6462);
			2962: out = 16'(-6237);
			2963: out = 16'(4674);
			2964: out = 16'(11785);
			2965: out = 16'(7064);
			2966: out = 16'(-7637);
			2967: out = 16'(-12811);
			2968: out = 16'(-1901);
			2969: out = 16'(16752);
			2970: out = 16'(14807);
			2971: out = 16'(3737);
			2972: out = 16'(-2311);
			2973: out = 16'(10701);
			2974: out = 16'(14052);
			2975: out = 16'(4390);
			2976: out = 16'(-471);
			2977: out = 16'(5088);
			2978: out = 16'(1751);
			2979: out = 16'(-3661);
			2980: out = 16'(800);
			2981: out = 16'(1186);
			2982: out = 16'(471);
			2983: out = 16'(-1937);
			2984: out = 16'(2500);
			2985: out = 16'(11347);
			2986: out = 16'(24477);
			2987: out = 16'(9979);
			2988: out = 16'(-6597);
			2989: out = 16'(-6337);
			2990: out = 16'(2108);
			2991: out = 16'(13180);
			2992: out = 16'(11929);
			2993: out = 16'(10443);
			2994: out = 16'(10997);
			2995: out = 16'(5157);
			2996: out = 16'(-10365);
			2997: out = 16'(-15963);
			2998: out = 16'(67);
			2999: out = 16'(8726);
			3000: out = 16'(2863);
			3001: out = 16'(8275);
			3002: out = 16'(7530);
			3003: out = 16'(-2273);
			3004: out = 16'(-2745);
			3005: out = 16'(-1028);
			3006: out = 16'(6700);
			3007: out = 16'(13248);
			3008: out = 16'(10889);
			3009: out = 16'(3149);
			3010: out = 16'(-1177);
			3011: out = 16'(9147);
			3012: out = 16'(19673);
			3013: out = 16'(13246);
			3014: out = 16'(-963);
			3015: out = 16'(-5065);
			3016: out = 16'(-7392);
			3017: out = 16'(-6842);
			3018: out = 16'(-4394);
			3019: out = 16'(1346);
			3020: out = 16'(9268);
			3021: out = 16'(15022);
			3022: out = 16'(13678);
			3023: out = 16'(2000);
			3024: out = 16'(-215);
			3025: out = 16'(8496);
			3026: out = 16'(18709);
			3027: out = 16'(12430);
			3028: out = 16'(-5079);
			3029: out = 16'(-11823);
			3030: out = 16'(-5626);
			3031: out = 16'(5024);
			3032: out = 16'(12451);
			3033: out = 16'(-3104);
			3034: out = 16'(-7694);
			3035: out = 16'(7330);
			3036: out = 16'(23236);
			3037: out = 16'(13395);
			3038: out = 16'(-450);
			3039: out = 16'(-4772);
			3040: out = 16'(124);
			3041: out = 16'(7437);
			3042: out = 16'(9861);
			3043: out = 16'(8364);
			3044: out = 16'(1223);
			3045: out = 16'(-4263);
			3046: out = 16'(132);
			3047: out = 16'(8714);
			3048: out = 16'(1647);
			3049: out = 16'(-17671);
			3050: out = 16'(-17118);
			3051: out = 16'(-1506);
			3052: out = 16'(10603);
			3053: out = 16'(15688);
			3054: out = 16'(12572);
			3055: out = 16'(5401);
			3056: out = 16'(-621);
			3057: out = 16'(-8042);
			3058: out = 16'(-10091);
			3059: out = 16'(-4023);
			3060: out = 16'(10899);
			3061: out = 16'(14650);
			3062: out = 16'(8295);
			3063: out = 16'(11731);
			3064: out = 16'(12101);
			3065: out = 16'(7729);
			3066: out = 16'(-4558);
			3067: out = 16'(-9979);
			3068: out = 16'(-8003);
			3069: out = 16'(4343);
			3070: out = 16'(9932);
			3071: out = 16'(1675);
			3072: out = 16'(-183);
			3073: out = 16'(1674);
			3074: out = 16'(-3333);
			3075: out = 16'(-4650);
			3076: out = 16'(-2325);
			3077: out = 16'(2529);
			3078: out = 16'(6273);
			3079: out = 16'(5518);
			3080: out = 16'(-1664);
			3081: out = 16'(-1840);
			3082: out = 16'(1888);
			3083: out = 16'(-3364);
			3084: out = 16'(-1322);
			3085: out = 16'(4396);
			3086: out = 16'(-1238);
			3087: out = 16'(-4552);
			3088: out = 16'(-581);
			3089: out = 16'(3084);
			3090: out = 16'(7836);
			3091: out = 16'(4937);
			3092: out = 16'(-6103);
			3093: out = 16'(-5619);
			3094: out = 16'(-4197);
			3095: out = 16'(3056);
			3096: out = 16'(7657);
			3097: out = 16'(1556);
			3098: out = 16'(7138);
			3099: out = 16'(12474);
			3100: out = 16'(7361);
			3101: out = 16'(-9267);
			3102: out = 16'(-19597);
			3103: out = 16'(-18830);
			3104: out = 16'(-4285);
			3105: out = 16'(11759);
			3106: out = 16'(6809);
			3107: out = 16'(3344);
			3108: out = 16'(8175);
			3109: out = 16'(5702);
			3110: out = 16'(167);
			3111: out = 16'(-5731);
			3112: out = 16'(1824);
			3113: out = 16'(13127);
			3114: out = 16'(10770);
			3115: out = 16'(-5128);
			3116: out = 16'(-14907);
			3117: out = 16'(-10286);
			3118: out = 16'(-8836);
			3119: out = 16'(-4716);
			3120: out = 16'(-455);
			3121: out = 16'(-2819);
			3122: out = 16'(2057);
			3123: out = 16'(9455);
			3124: out = 16'(11993);
			3125: out = 16'(6504);
			3126: out = 16'(-8721);
			3127: out = 16'(-16581);
			3128: out = 16'(-11674);
			3129: out = 16'(-1835);
			3130: out = 16'(-259);
			3131: out = 16'(-2500);
			3132: out = 16'(1627);
			3133: out = 16'(4699);
			3134: out = 16'(6491);
			3135: out = 16'(4835);
			3136: out = 16'(-4730);
			3137: out = 16'(-11389);
			3138: out = 16'(-3485);
			3139: out = 16'(-993);
			3140: out = 16'(-8705);
			3141: out = 16'(-12208);
			3142: out = 16'(-13444);
			3143: out = 16'(1541);
			3144: out = 16'(10542);
			3145: out = 16'(1510);
			3146: out = 16'(5523);
			3147: out = 16'(8834);
			3148: out = 16'(2401);
			3149: out = 16'(-11075);
			3150: out = 16'(-18069);
			3151: out = 16'(-12825);
			3152: out = 16'(-10119);
			3153: out = 16'(-656);
			3154: out = 16'(11346);
			3155: out = 16'(3990);
			3156: out = 16'(-2458);
			3157: out = 16'(-1848);
			3158: out = 16'(2006);
			3159: out = 16'(162);
			3160: out = 16'(-11612);
			3161: out = 16'(-18550);
			3162: out = 16'(-11052);
			3163: out = 16'(2221);
			3164: out = 16'(6754);
			3165: out = 16'(-5835);
			3166: out = 16'(-14533);
			3167: out = 16'(-6494);
			3168: out = 16'(10661);
			3169: out = 16'(10127);
			3170: out = 16'(-5359);
			3171: out = 16'(-19816);
			3172: out = 16'(-14867);
			3173: out = 16'(-3211);
			3174: out = 16'(3803);
			3175: out = 16'(8438);
			3176: out = 16'(-2477);
			3177: out = 16'(-11852);
			3178: out = 16'(-11545);
			3179: out = 16'(-9750);
			3180: out = 16'(3656);
			3181: out = 16'(12783);
			3182: out = 16'(1119);
			3183: out = 16'(-7374);
			3184: out = 16'(-7357);
			3185: out = 16'(-3584);
			3186: out = 16'(-3107);
			3187: out = 16'(-8929);
			3188: out = 16'(-17651);
			3189: out = 16'(-6739);
			3190: out = 16'(1187);
			3191: out = 16'(-711);
			3192: out = 16'(9754);
			3193: out = 16'(9531);
			3194: out = 16'(-5404);
			3195: out = 16'(-9749);
			3196: out = 16'(-10021);
			3197: out = 16'(-9138);
			3198: out = 16'(-8615);
			3199: out = 16'(4695);
			3200: out = 16'(10170);
			3201: out = 16'(-5256);
			3202: out = 16'(-11810);
			3203: out = 16'(-4609);
			3204: out = 16'(9465);
			3205: out = 16'(13371);
			3206: out = 16'(-3964);
			3207: out = 16'(-11757);
			3208: out = 16'(-8069);
			3209: out = 16'(-3737);
			3210: out = 16'(5356);
			3211: out = 16'(2113);
			3212: out = 16'(-12784);
			3213: out = 16'(-11425);
			3214: out = 16'(-4434);
			3215: out = 16'(2555);
			3216: out = 16'(770);
			3217: out = 16'(-7552);
			3218: out = 16'(-13004);
			3219: out = 16'(-8619);
			3220: out = 16'(-3258);
			3221: out = 16'(-523);
			3222: out = 16'(-8394);
			3223: out = 16'(-12308);
			3224: out = 16'(3204);
			3225: out = 16'(4628);
			3226: out = 16'(862);
			3227: out = 16'(-821);
			3228: out = 16'(-5143);
			3229: out = 16'(-8854);
			3230: out = 16'(-4151);
			3231: out = 16'(-2277);
			3232: out = 16'(-1934);
			3233: out = 16'(9505);
			3234: out = 16'(397);
			3235: out = 16'(-6402);
			3236: out = 16'(-2117);
			3237: out = 16'(2197);
			3238: out = 16'(2479);
			3239: out = 16'(-6132);
			3240: out = 16'(-751);
			3241: out = 16'(6881);
			3242: out = 16'(1548);
			3243: out = 16'(-11242);
			3244: out = 16'(-7530);
			3245: out = 16'(-253);
			3246: out = 16'(2968);
			3247: out = 16'(-1494);
			3248: out = 16'(-3167);
			3249: out = 16'(3155);
			3250: out = 16'(6045);
			3251: out = 16'(-1675);
			3252: out = 16'(-9928);
			3253: out = 16'(-9668);
			3254: out = 16'(-809);
			3255: out = 16'(-677);
			3256: out = 16'(-3360);
			3257: out = 16'(4642);
			3258: out = 16'(12168);
			3259: out = 16'(7520);
			3260: out = 16'(1910);
			3261: out = 16'(-5831);
			3262: out = 16'(-1081);
			3263: out = 16'(-605);
			3264: out = 16'(4368);
			3265: out = 16'(9135);
			3266: out = 16'(3267);
			3267: out = 16'(1825);
			3268: out = 16'(2747);
			3269: out = 16'(-5527);
			3270: out = 16'(-7222);
			3271: out = 16'(-170);
			3272: out = 16'(1893);
			3273: out = 16'(-3477);
			3274: out = 16'(-9251);
			3275: out = 16'(2907);
			3276: out = 16'(3140);
			3277: out = 16'(-11428);
			3278: out = 16'(-5823);
			3279: out = 16'(8495);
			3280: out = 16'(4027);
			3281: out = 16'(-498);
			3282: out = 16'(10023);
			3283: out = 16'(9895);
			3284: out = 16'(-6838);
			3285: out = 16'(-14417);
			3286: out = 16'(-12551);
			3287: out = 16'(-2847);
			3288: out = 16'(14326);
			3289: out = 16'(10399);
			3290: out = 16'(-3845);
			3291: out = 16'(771);
			3292: out = 16'(12206);
			3293: out = 16'(17260);
			3294: out = 16'(3295);
			3295: out = 16'(-15202);
			3296: out = 16'(-10076);
			3297: out = 16'(8170);
			3298: out = 16'(14350);
			3299: out = 16'(3056);
			3300: out = 16'(-7260);
			3301: out = 16'(-3354);
			3302: out = 16'(10570);
			3303: out = 16'(12801);
			3304: out = 16'(10626);
			3305: out = 16'(5748);
			3306: out = 16'(-1333);
			3307: out = 16'(-4571);
			3308: out = 16'(-5391);
			3309: out = 16'(7454);
			3310: out = 16'(6254);
			3311: out = 16'(-5669);
			3312: out = 16'(-602);
			3313: out = 16'(8496);
			3314: out = 16'(12330);
			3315: out = 16'(7991);
			3316: out = 16'(-2188);
			3317: out = 16'(503);
			3318: out = 16'(5022);
			3319: out = 16'(9394);
			3320: out = 16'(-2346);
			3321: out = 16'(-10196);
			3322: out = 16'(-1978);
			3323: out = 16'(4882);
			3324: out = 16'(12531);
			3325: out = 16'(13511);
			3326: out = 16'(1813);
			3327: out = 16'(-5886);
			3328: out = 16'(-8609);
			3329: out = 16'(2197);
			3330: out = 16'(13409);
			3331: out = 16'(10058);
			3332: out = 16'(4845);
			3333: out = 16'(-671);
			3334: out = 16'(-4694);
			3335: out = 16'(-15294);
			3336: out = 16'(-16043);
			3337: out = 16'(5965);
			3338: out = 16'(20756);
			3339: out = 16'(13693);
			3340: out = 16'(-795);
			3341: out = 16'(-6171);
			3342: out = 16'(4367);
			3343: out = 16'(14171);
			3344: out = 16'(15005);
			3345: out = 16'(6742);
			3346: out = 16'(975);
			3347: out = 16'(-4485);
			3348: out = 16'(2101);
			3349: out = 16'(4499);
			3350: out = 16'(515);
			3351: out = 16'(-2634);
			3352: out = 16'(435);
			3353: out = 16'(-1180);
			3354: out = 16'(3003);
			3355: out = 16'(12267);
			3356: out = 16'(5231);
			3357: out = 16'(-1061);
			3358: out = 16'(-5143);
			3359: out = 16'(-3808);
			3360: out = 16'(4263);
			3361: out = 16'(21378);
			3362: out = 16'(16510);
			3363: out = 16'(-2821);
			3364: out = 16'(-11712);
			3365: out = 16'(-2137);
			3366: out = 16'(8478);
			3367: out = 16'(11521);
			3368: out = 16'(-2164);
			3369: out = 16'(-5396);
			3370: out = 16'(3512);
			3371: out = 16'(8841);
			3372: out = 16'(9053);
			3373: out = 16'(4206);
			3374: out = 16'(-2741);
			3375: out = 16'(-5037);
			3376: out = 16'(-7588);
			3377: out = 16'(-6255);
			3378: out = 16'(897);
			3379: out = 16'(5397);
			3380: out = 16'(9684);
			3381: out = 16'(-3299);
			3382: out = 16'(-6884);
			3383: out = 16'(-3932);
			3384: out = 16'(8236);
			3385: out = 16'(18793);
			3386: out = 16'(14556);
			3387: out = 16'(453);
			3388: out = 16'(-9038);
			3389: out = 16'(-3749);
			3390: out = 16'(-3001);
			3391: out = 16'(4192);
			3392: out = 16'(6674);
			3393: out = 16'(1487);
			3394: out = 16'(-1897);
			3395: out = 16'(4279);
			3396: out = 16'(-3396);
			3397: out = 16'(-8700);
			3398: out = 16'(-1022);
			3399: out = 16'(4661);
			3400: out = 16'(-354);
			3401: out = 16'(-6147);
			3402: out = 16'(-6724);
			3403: out = 16'(-8216);
			3404: out = 16'(3924);
			3405: out = 16'(8736);
			3406: out = 16'(5190);
			3407: out = 16'(5897);
			3408: out = 16'(3500);
			3409: out = 16'(-161);
			3410: out = 16'(2700);
			3411: out = 16'(928);
			3412: out = 16'(-186);
			3413: out = 16'(8437);
			3414: out = 16'(11512);
			3415: out = 16'(-3229);
			3416: out = 16'(-14617);
			3417: out = 16'(-7941);
			3418: out = 16'(8823);
			3419: out = 16'(11500);
			3420: out = 16'(-1649);
			3421: out = 16'(-7813);
			3422: out = 16'(-724);
			3423: out = 16'(5376);
			3424: out = 16'(1532);
			3425: out = 16'(-3940);
			3426: out = 16'(1983);
			3427: out = 16'(6890);
			3428: out = 16'(3985);
			3429: out = 16'(-4340);
			3430: out = 16'(-9582);
			3431: out = 16'(-10578);
			3432: out = 16'(-15463);
			3433: out = 16'(-3366);
			3434: out = 16'(8452);
			3435: out = 16'(7061);
			3436: out = 16'(1549);
			3437: out = 16'(2784);
			3438: out = 16'(5605);
			3439: out = 16'(2984);
			3440: out = 16'(-2635);
			3441: out = 16'(-8453);
			3442: out = 16'(-5229);
			3443: out = 16'(-780);
			3444: out = 16'(3460);
			3445: out = 16'(2571);
			3446: out = 16'(-1319);
			3447: out = 16'(4129);
			3448: out = 16'(8452);
			3449: out = 16'(5609);
			3450: out = 16'(-7277);
			3451: out = 16'(-7045);
			3452: out = 16'(-6787);
			3453: out = 16'(5472);
			3454: out = 16'(4877);
			3455: out = 16'(-5283);
			3456: out = 16'(-2815);
			3457: out = 16'(6656);
			3458: out = 16'(12358);
			3459: out = 16'(2984);
			3460: out = 16'(-10314);
			3461: out = 16'(-10161);
			3462: out = 16'(-3833);
			3463: out = 16'(12221);
			3464: out = 16'(12774);
			3465: out = 16'(-4633);
			3466: out = 16'(-10100);
			3467: out = 16'(-4513);
			3468: out = 16'(-1418);
			3469: out = 16'(-1585);
			3470: out = 16'(-2769);
			3471: out = 16'(-7162);
			3472: out = 16'(-6818);
			3473: out = 16'(-11347);
			3474: out = 16'(2240);
			3475: out = 16'(4334);
			3476: out = 16'(-7011);
			3477: out = 16'(-725);
			3478: out = 16'(13926);
			3479: out = 16'(6705);
			3480: out = 16'(-10556);
			3481: out = 16'(-9486);
			3482: out = 16'(-3274);
			3483: out = 16'(-3251);
			3484: out = 16'(1056);
			3485: out = 16'(3708);
			3486: out = 16'(-2049);
			3487: out = 16'(-9731);
			3488: out = 16'(-5992);
			3489: out = 16'(4906);
			3490: out = 16'(7228);
			3491: out = 16'(6038);
			3492: out = 16'(-6513);
			3493: out = 16'(-11487);
			3494: out = 16'(-6939);
			3495: out = 16'(2816);
			3496: out = 16'(1154);
			3497: out = 16'(-7373);
			3498: out = 16'(2423);
			3499: out = 16'(6665);
			3500: out = 16'(1731);
			3501: out = 16'(6923);
			3502: out = 16'(3995);
			3503: out = 16'(-123);
			3504: out = 16'(-7169);
			3505: out = 16'(-11054);
			3506: out = 16'(-3501);
			3507: out = 16'(8000);
			3508: out = 16'(3064);
			3509: out = 16'(-15037);
			3510: out = 16'(-17073);
			3511: out = 16'(-1849);
			3512: out = 16'(8924);
			3513: out = 16'(7519);
			3514: out = 16'(3410);
			3515: out = 16'(1040);
			3516: out = 16'(-936);
			3517: out = 16'(-9104);
			3518: out = 16'(-1853);
			3519: out = 16'(11824);
			3520: out = 16'(1885);
			3521: out = 16'(-13382);
			3522: out = 16'(-10470);
			3523: out = 16'(720);
			3524: out = 16'(-2000);
			3525: out = 16'(-8831);
			3526: out = 16'(-1544);
			3527: out = 16'(3844);
			3528: out = 16'(10294);
			3529: out = 16'(8222);
			3530: out = 16'(-3239);
			3531: out = 16'(-16919);
			3532: out = 16'(-20069);
			3533: out = 16'(-6513);
			3534: out = 16'(9834);
			3535: out = 16'(17450);
			3536: out = 16'(684);
			3537: out = 16'(-11795);
			3538: out = 16'(-5247);
			3539: out = 16'(5732);
			3540: out = 16'(14427);
			3541: out = 16'(2684);
			3542: out = 16'(-6158);
			3543: out = 16'(-1157);
			3544: out = 16'(2892);
			3545: out = 16'(-235);
			3546: out = 16'(-8063);
			3547: out = 16'(-5493);
			3548: out = 16'(3846);
			3549: out = 16'(3046);
			3550: out = 16'(-1291);
			3551: out = 16'(-3552);
			3552: out = 16'(-497);
			3553: out = 16'(-1926);
			3554: out = 16'(-1685);
			3555: out = 16'(-1170);
			3556: out = 16'(-7742);
			3557: out = 16'(-9176);
			3558: out = 16'(265);
			3559: out = 16'(4719);
			3560: out = 16'(131);
			3561: out = 16'(-3439);
			3562: out = 16'(-11141);
			3563: out = 16'(-15266);
			3564: out = 16'(-3077);
			3565: out = 16'(-2292);
			3566: out = 16'(-1461);
			3567: out = 16'(6137);
			3568: out = 16'(2074);
			3569: out = 16'(3062);
			3570: out = 16'(5597);
			3571: out = 16'(8197);
			3572: out = 16'(3086);
			3573: out = 16'(-6375);
			3574: out = 16'(-3024);
			3575: out = 16'(-612);
			3576: out = 16'(-258);
			3577: out = 16'(-6876);
			3578: out = 16'(-7463);
			3579: out = 16'(-513);
			3580: out = 16'(-806);
			3581: out = 16'(-13059);
			3582: out = 16'(-11448);
			3583: out = 16'(2399);
			3584: out = 16'(6660);
			3585: out = 16'(-1802);
			3586: out = 16'(-6364);
			3587: out = 16'(-9860);
			3588: out = 16'(-4599);
			3589: out = 16'(10877);
			3590: out = 16'(16401);
			3591: out = 16'(2207);
			3592: out = 16'(-11319);
			3593: out = 16'(-11795);
			3594: out = 16'(-1493);
			3595: out = 16'(8023);
			3596: out = 16'(2201);
			3597: out = 16'(-1765);
			3598: out = 16'(4473);
			3599: out = 16'(-1508);
			3600: out = 16'(-10208);
			3601: out = 16'(-12037);
			3602: out = 16'(-9166);
			3603: out = 16'(7575);
			3604: out = 16'(19575);
			3605: out = 16'(5167);
			3606: out = 16'(-12144);
			3607: out = 16'(-10893);
			3608: out = 16'(-333);
			3609: out = 16'(8901);
			3610: out = 16'(452);
			3611: out = 16'(-4284);
			3612: out = 16'(105);
			3613: out = 16'(4794);
			3614: out = 16'(8603);
			3615: out = 16'(-808);
			3616: out = 16'(-9941);
			3617: out = 16'(-3745);
			3618: out = 16'(728);
			3619: out = 16'(4613);
			3620: out = 16'(3286);
			3621: out = 16'(-2050);
			3622: out = 16'(-184);
			3623: out = 16'(-6849);
			3624: out = 16'(-10188);
			3625: out = 16'(-6715);
			3626: out = 16'(541);
			3627: out = 16'(6339);
			3628: out = 16'(-260);
			3629: out = 16'(-1689);
			3630: out = 16'(-2419);
			3631: out = 16'(2310);
			3632: out = 16'(11334);
			3633: out = 16'(12278);
			3634: out = 16'(2636);
			3635: out = 16'(-7945);
			3636: out = 16'(-2326);
			3637: out = 16'(1244);
			3638: out = 16'(7247);
			3639: out = 16'(2684);
			3640: out = 16'(-1712);
			3641: out = 16'(-1997);
			3642: out = 16'(-3312);
			3643: out = 16'(7720);
			3644: out = 16'(11495);
			3645: out = 16'(-890);
			3646: out = 16'(-10490);
			3647: out = 16'(-7257);
			3648: out = 16'(-6542);
			3649: out = 16'(-4529);
			3650: out = 16'(811);
			3651: out = 16'(-3049);
			3652: out = 16'(-1518);
			3653: out = 16'(3747);
			3654: out = 16'(-1042);
			3655: out = 16'(-6004);
			3656: out = 16'(-9201);
			3657: out = 16'(-4900);
			3658: out = 16'(1740);
			3659: out = 16'(6682);
			3660: out = 16'(5759);
			3661: out = 16'(392);
			3662: out = 16'(722);
			3663: out = 16'(2616);
			3664: out = 16'(-1452);
			3665: out = 16'(-2378);
			3666: out = 16'(-43);
			3667: out = 16'(570);
			3668: out = 16'(2380);
			3669: out = 16'(4317);
			3670: out = 16'(-6767);
			3671: out = 16'(-10469);
			3672: out = 16'(-689);
			3673: out = 16'(6745);
			3674: out = 16'(7758);
			3675: out = 16'(6077);
			3676: out = 16'(3928);
			3677: out = 16'(-4249);
			3678: out = 16'(-9461);
			3679: out = 16'(-6502);
			3680: out = 16'(-582);
			3681: out = 16'(2485);
			3682: out = 16'(10902);
			3683: out = 16'(6808);
			3684: out = 16'(-3403);
			3685: out = 16'(-9719);
			3686: out = 16'(-12110);
			3687: out = 16'(3895);
			3688: out = 16'(15161);
			3689: out = 16'(7014);
			3690: out = 16'(2575);
			3691: out = 16'(6380);
			3692: out = 16'(-1398);
			3693: out = 16'(-13534);
			3694: out = 16'(-19040);
			3695: out = 16'(-10914);
			3696: out = 16'(10468);
			3697: out = 16'(18931);
			3698: out = 16'(4341);
			3699: out = 16'(-4508);
			3700: out = 16'(-1388);
			3701: out = 16'(8354);
			3702: out = 16'(17665);
			3703: out = 16'(6764);
			3704: out = 16'(-4435);
			3705: out = 16'(-4905);
			3706: out = 16'(-2849);
			3707: out = 16'(-5614);
			3708: out = 16'(-4296);
			3709: out = 16'(-54);
			3710: out = 16'(4490);
			3711: out = 16'(7556);
			3712: out = 16'(8362);
			3713: out = 16'(-286);
			3714: out = 16'(-4257);
			3715: out = 16'(5730);
			3716: out = 16'(3147);
			3717: out = 16'(4198);
			3718: out = 16'(2886);
			3719: out = 16'(5367);
			3720: out = 16'(4432);
			3721: out = 16'(1672);
			3722: out = 16'(5066);
			3723: out = 16'(2545);
			3724: out = 16'(-2432);
			3725: out = 16'(-8076);
			3726: out = 16'(-11896);
			3727: out = 16'(592);
			3728: out = 16'(13922);
			3729: out = 16'(3761);
			3730: out = 16'(-9248);
			3731: out = 16'(-7151);
			3732: out = 16'(11558);
			3733: out = 16'(14781);
			3734: out = 16'(-3540);
			3735: out = 16'(-2867);
			3736: out = 16'(3165);
			3737: out = 16'(2717);
			3738: out = 16'(4479);
			3739: out = 16'(7199);
			3740: out = 16'(3599);
			3741: out = 16'(-614);
			3742: out = 16'(-7193);
			3743: out = 16'(-14707);
			3744: out = 16'(-740);
			3745: out = 16'(8705);
			3746: out = 16'(3142);
			3747: out = 16'(1817);
			3748: out = 16'(8936);
			3749: out = 16'(6638);
			3750: out = 16'(3515);
			3751: out = 16'(3124);
			3752: out = 16'(693);
			3753: out = 16'(1252);
			3754: out = 16'(-8118);
			3755: out = 16'(-6650);
			3756: out = 16'(6179);
			3757: out = 16'(10377);
			3758: out = 16'(8503);
			3759: out = 16'(-1950);
			3760: out = 16'(-8425);
			3761: out = 16'(-2675);
			3762: out = 16'(4239);
			3763: out = 16'(12845);
			3764: out = 16'(14117);
			3765: out = 16'(4274);
			3766: out = 16'(1040);
			3767: out = 16'(4015);
			3768: out = 16'(-1376);
			3769: out = 16'(-537);
			3770: out = 16'(-5827);
			3771: out = 16'(-6123);
			3772: out = 16'(6597);
			3773: out = 16'(13395);
			3774: out = 16'(5721);
			3775: out = 16'(-3523);
			3776: out = 16'(-5458);
			3777: out = 16'(9579);
			3778: out = 16'(13233);
			3779: out = 16'(3519);
			3780: out = 16'(-1768);
			3781: out = 16'(-256);
			3782: out = 16'(-2036);
			3783: out = 16'(-8527);
			3784: out = 16'(-8767);
			3785: out = 16'(2945);
			3786: out = 16'(11701);
			3787: out = 16'(4515);
			3788: out = 16'(2588);
			3789: out = 16'(3494);
			3790: out = 16'(4342);
			3791: out = 16'(-2590);
			3792: out = 16'(-12771);
			3793: out = 16'(-8798);
			3794: out = 16'(-809);
			3795: out = 16'(5250);
			3796: out = 16'(11214);
			3797: out = 16'(3184);
			3798: out = 16'(5702);
			3799: out = 16'(11583);
			3800: out = 16'(10290);
			3801: out = 16'(-2106);
			3802: out = 16'(-12613);
			3803: out = 16'(-10344);
			3804: out = 16'(-359);
			3805: out = 16'(12914);
			3806: out = 16'(10224);
			3807: out = 16'(-2956);
			3808: out = 16'(446);
			3809: out = 16'(10860);
			3810: out = 16'(13908);
			3811: out = 16'(-1324);
			3812: out = 16'(-5560);
			3813: out = 16'(-692);
			3814: out = 16'(7808);
			3815: out = 16'(13155);
			3816: out = 16'(8490);
			3817: out = 16'(3419);
			3818: out = 16'(2423);
			3819: out = 16'(-1163);
			3820: out = 16'(-5647);
			3821: out = 16'(-4626);
			3822: out = 16'(-4274);
			3823: out = 16'(-7767);
			3824: out = 16'(-3670);
			3825: out = 16'(5992);
			3826: out = 16'(-1968);
			3827: out = 16'(-17426);
			3828: out = 16'(-14522);
			3829: out = 16'(-7907);
			3830: out = 16'(-3007);
			3831: out = 16'(14276);
			3832: out = 16'(14405);
			3833: out = 16'(-6926);
			3834: out = 16'(-18418);
			3835: out = 16'(-8604);
			3836: out = 16'(3123);
			3837: out = 16'(17916);
			3838: out = 16'(15661);
			3839: out = 16'(58);
			3840: out = 16'(-7464);
			3841: out = 16'(-2545);
			3842: out = 16'(7391);
			3843: out = 16'(1276);
			3844: out = 16'(-6426);
			3845: out = 16'(2303);
			3846: out = 16'(-771);
			3847: out = 16'(-9423);
			3848: out = 16'(-3388);
			3849: out = 16'(-1222);
			3850: out = 16'(3866);
			3851: out = 16'(10221);
			3852: out = 16'(8848);
			3853: out = 16'(-2647);
			3854: out = 16'(-8268);
			3855: out = 16'(-3208);
			3856: out = 16'(12486);
			3857: out = 16'(11555);
			3858: out = 16'(-1537);
			3859: out = 16'(-6696);
			3860: out = 16'(299);
			3861: out = 16'(6427);
			3862: out = 16'(967);
			3863: out = 16'(-16416);
			3864: out = 16'(-14177);
			3865: out = 16'(-1515);
			3866: out = 16'(5995);
			3867: out = 16'(7889);
			3868: out = 16'(2690);
			3869: out = 16'(6966);
			3870: out = 16'(6194);
			3871: out = 16'(-1110);
			3872: out = 16'(-9190);
			3873: out = 16'(-13450);
			3874: out = 16'(-6456);
			3875: out = 16'(3763);
			3876: out = 16'(6426);
			3877: out = 16'(3432);
			3878: out = 16'(-6340);
			3879: out = 16'(-1108);
			3880: out = 16'(632);
			3881: out = 16'(2854);
			3882: out = 16'(5610);
			3883: out = 16'(13243);
			3884: out = 16'(12286);
			3885: out = 16'(-3267);
			3886: out = 16'(-13915);
			3887: out = 16'(-12080);
			3888: out = 16'(-2404);
			3889: out = 16'(535);
			3890: out = 16'(-6147);
			3891: out = 16'(-7158);
			3892: out = 16'(-259);
			3893: out = 16'(-2183);
			3894: out = 16'(-5185);
			3895: out = 16'(-2196);
			3896: out = 16'(3991);
			3897: out = 16'(3192);
			3898: out = 16'(-8456);
			3899: out = 16'(-11406);
			3900: out = 16'(-5970);
			3901: out = 16'(7178);
			3902: out = 16'(11484);
			3903: out = 16'(-3556);
			3904: out = 16'(-6677);
			3905: out = 16'(-199);
			3906: out = 16'(347);
			3907: out = 16'(2308);
			3908: out = 16'(-5342);
			3909: out = 16'(-9941);
			3910: out = 16'(443);
			3911: out = 16'(1131);
			3912: out = 16'(-2128);
			3913: out = 16'(3539);
			3914: out = 16'(5832);
			3915: out = 16'(4531);
			3916: out = 16'(-4355);
			3917: out = 16'(-15173);
			3918: out = 16'(-6793);
			3919: out = 16'(4278);
			3920: out = 16'(3975);
			3921: out = 16'(-3973);
			3922: out = 16'(-3249);
			3923: out = 16'(-168);
			3924: out = 16'(-502);
			3925: out = 16'(-3473);
			3926: out = 16'(-9211);
			3927: out = 16'(-1794);
			3928: out = 16'(1597);
			3929: out = 16'(2230);
			3930: out = 16'(1371);
			3931: out = 16'(-2303);
			3932: out = 16'(-909);
			3933: out = 16'(1844);
			3934: out = 16'(-7956);
			3935: out = 16'(-6850);
			3936: out = 16'(-945);
			3937: out = 16'(2323);
			3938: out = 16'(7762);
			3939: out = 16'(7209);
			3940: out = 16'(2333);
			3941: out = 16'(-7073);
			3942: out = 16'(-15099);
			3943: out = 16'(-11233);
			3944: out = 16'(-5834);
			3945: out = 16'(3620);
			3946: out = 16'(8610);
			3947: out = 16'(-7337);
			3948: out = 16'(-16005);
			3949: out = 16'(-14735);
			3950: out = 16'(-2516);
			3951: out = 16'(15054);
			3952: out = 16'(19352);
			3953: out = 16'(-2167);
			3954: out = 16'(-22791);
			3955: out = 16'(-19536);
			3956: out = 16'(-6496);
			3957: out = 16'(14100);
			3958: out = 16'(12653);
			3959: out = 16'(-5451);
			3960: out = 16'(-3973);
			3961: out = 16'(7469);
			3962: out = 16'(6758);
			3963: out = 16'(-255);
			3964: out = 16'(-6964);
			3965: out = 16'(-3797);
			3966: out = 16'(-1977);
			3967: out = 16'(13);
			3968: out = 16'(-484);
			3969: out = 16'(-6889);
			3970: out = 16'(-11981);
			3971: out = 16'(-7110);
			3972: out = 16'(1300);
			3973: out = 16'(4321);
			3974: out = 16'(-1919);
			3975: out = 16'(-4658);
			3976: out = 16'(2160);
			3977: out = 16'(-887);
			3978: out = 16'(-7372);
			3979: out = 16'(-4840);
			3980: out = 16'(-2250);
			3981: out = 16'(3482);
			3982: out = 16'(8044);
			3983: out = 16'(5037);
			3984: out = 16'(-4792);
			3985: out = 16'(-9866);
			3986: out = 16'(-9867);
			3987: out = 16'(-7522);
			3988: out = 16'(1716);
			3989: out = 16'(11837);
			3990: out = 16'(7793);
			3991: out = 16'(3047);
			3992: out = 16'(2095);
			3993: out = 16'(-3379);
			3994: out = 16'(-7188);
			3995: out = 16'(-12832);
			3996: out = 16'(-5767);
			3997: out = 16'(4984);
			3998: out = 16'(3388);
			3999: out = 16'(1661);
			4000: out = 16'(1190);
			4001: out = 16'(10800);
			4002: out = 16'(13545);
			4003: out = 16'(6511);
			4004: out = 16'(-5922);
			4005: out = 16'(-8119);
			4006: out = 16'(-7411);
			4007: out = 16'(-6966);
			4008: out = 16'(-625);
			4009: out = 16'(-2157);
			4010: out = 16'(-307);
			4011: out = 16'(5232);
			4012: out = 16'(6051);
			4013: out = 16'(-3466);
			4014: out = 16'(3755);
			4015: out = 16'(8428);
			4016: out = 16'(2244);
			4017: out = 16'(-6559);
			4018: out = 16'(-9798);
			4019: out = 16'(-2693);
			4020: out = 16'(11318);
			4021: out = 16'(16180);
			4022: out = 16'(811);
			4023: out = 16'(-11183);
			4024: out = 16'(-6974);
			4025: out = 16'(1391);
			4026: out = 16'(9021);
			4027: out = 16'(3332);
			4028: out = 16'(-6496);
			4029: out = 16'(140);
			4030: out = 16'(11671);
			4031: out = 16'(7206);
			4032: out = 16'(-4080);
			4033: out = 16'(-9454);
			4034: out = 16'(4305);
			4035: out = 16'(2576);
			4036: out = 16'(-4000);
			4037: out = 16'(3902);
			4038: out = 16'(10879);
			4039: out = 16'(-778);
			4040: out = 16'(-14713);
			4041: out = 16'(-5605);
			4042: out = 16'(4217);
			4043: out = 16'(4153);
			4044: out = 16'(2313);
			4045: out = 16'(-1173);
			4046: out = 16'(-10388);
			4047: out = 16'(-10226);
			4048: out = 16'(1532);
			4049: out = 16'(9762);
			4050: out = 16'(14595);
			4051: out = 16'(8729);
			4052: out = 16'(-6203);
			4053: out = 16'(-8509);
			4054: out = 16'(-2421);
			4055: out = 16'(4327);
			4056: out = 16'(11053);
			4057: out = 16'(7346);
			4058: out = 16'(-2619);
			4059: out = 16'(699);
			4060: out = 16'(4560);
			4061: out = 16'(1684);
			4062: out = 16'(4654);
			4063: out = 16'(5934);
			4064: out = 16'(-1398);
			4065: out = 16'(2804);
			4066: out = 16'(86);
			4067: out = 16'(-3921);
			4068: out = 16'(4297);
			4069: out = 16'(12989);
			4070: out = 16'(5340);
			4071: out = 16'(-3779);
			4072: out = 16'(2198);
			4073: out = 16'(5552);
			4074: out = 16'(9043);
			4075: out = 16'(8021);
			4076: out = 16'(7050);
			4077: out = 16'(1993);
			4078: out = 16'(-6032);
			4079: out = 16'(-9336);
			4080: out = 16'(-184);
			4081: out = 16'(9804);
			4082: out = 16'(-1);
			4083: out = 16'(-9385);
			4084: out = 16'(-4682);
			4085: out = 16'(-2010);
			4086: out = 16'(5472);
			4087: out = 16'(2355);
			4088: out = 16'(-2685);
			4089: out = 16'(-1092);
			4090: out = 16'(-358);
			4091: out = 16'(6856);
			4092: out = 16'(629);
			4093: out = 16'(3550);
			4094: out = 16'(5584);
			4095: out = 16'(8000);
			4096: out = 16'(4551);
			4097: out = 16'(-5311);
			4098: out = 16'(-256);
			4099: out = 16'(6299);
			4100: out = 16'(4592);
			4101: out = 16'(-3218);
			4102: out = 16'(-1842);
			4103: out = 16'(7454);
			4104: out = 16'(7361);
			4105: out = 16'(-4614);
			4106: out = 16'(-3930);
			4107: out = 16'(388);
			4108: out = 16'(-5536);
			4109: out = 16'(-2710);
			4110: out = 16'(6425);
			4111: out = 16'(3105);
			4112: out = 16'(-3722);
			4113: out = 16'(-2048);
			4114: out = 16'(-2313);
			4115: out = 16'(-4425);
			4116: out = 16'(-4066);
			4117: out = 16'(5736);
			4118: out = 16'(4498);
			4119: out = 16'(2535);
			4120: out = 16'(8879);
			4121: out = 16'(6455);
			4122: out = 16'(-1681);
			4123: out = 16'(-10606);
			4124: out = 16'(-7085);
			4125: out = 16'(2269);
			4126: out = 16'(11429);
			4127: out = 16'(12556);
			4128: out = 16'(5467);
			4129: out = 16'(2934);
			4130: out = 16'(-585);
			4131: out = 16'(-869);
			4132: out = 16'(419);
			4133: out = 16'(6763);
			4134: out = 16'(11508);
			4135: out = 16'(5059);
			4136: out = 16'(-178);
			4137: out = 16'(1852);
			4138: out = 16'(-853);
			4139: out = 16'(-5804);
			4140: out = 16'(-8101);
			4141: out = 16'(-4983);
			4142: out = 16'(1083);
			4143: out = 16'(9892);
			4144: out = 16'(2900);
			4145: out = 16'(-9521);
			4146: out = 16'(-14862);
			4147: out = 16'(-12992);
			4148: out = 16'(-7688);
			4149: out = 16'(9575);
			4150: out = 16'(20813);
			4151: out = 16'(-2947);
			4152: out = 16'(-12509);
			4153: out = 16'(-1459);
			4154: out = 16'(10106);
			4155: out = 16'(12084);
			4156: out = 16'(1643);
			4157: out = 16'(-3596);
			4158: out = 16'(774);
			4159: out = 16'(3213);
			4160: out = 16'(3063);
			4161: out = 16'(-7868);
			4162: out = 16'(-8639);
			4163: out = 16'(2956);
			4164: out = 16'(1914);
			4165: out = 16'(3127);
			4166: out = 16'(3043);
			4167: out = 16'(550);
			4168: out = 16'(-178);
			4169: out = 16'(1436);
			4170: out = 16'(1156);
			4171: out = 16'(-6547);
			4172: out = 16'(-448);
			4173: out = 16'(10964);
			4174: out = 16'(4338);
			4175: out = 16'(-9352);
			4176: out = 16'(-11147);
			4177: out = 16'(1394);
			4178: out = 16'(13469);
			4179: out = 16'(2396);
			4180: out = 16'(-9766);
			4181: out = 16'(-7061);
			4182: out = 16'(2295);
			4183: out = 16'(3508);
			4184: out = 16'(-243);
			4185: out = 16'(-4518);
			4186: out = 16'(244);
			4187: out = 16'(8988);
			4188: out = 16'(9471);
			4189: out = 16'(8330);
			4190: out = 16'(-3792);
			4191: out = 16'(-7081);
			4192: out = 16'(-7627);
			4193: out = 16'(-2774);
			4194: out = 16'(7994);
			4195: out = 16'(9454);
			4196: out = 16'(-4957);
			4197: out = 16'(-9486);
			4198: out = 16'(-7424);
			4199: out = 16'(-7205);
			4200: out = 16'(2886);
			4201: out = 16'(3703);
			4202: out = 16'(-3472);
			4203: out = 16'(-3014);
			4204: out = 16'(5423);
			4205: out = 16'(-2051);
			4206: out = 16'(-8227);
			4207: out = 16'(-344);
			4208: out = 16'(4375);
			4209: out = 16'(6058);
			4210: out = 16'(-4677);
			4211: out = 16'(-1644);
			4212: out = 16'(7131);
			4213: out = 16'(7385);
			4214: out = 16'(2451);
			4215: out = 16'(-6132);
			4216: out = 16'(-15223);
			4217: out = 16'(-15048);
			4218: out = 16'(-4734);
			4219: out = 16'(728);
			4220: out = 16'(5981);
			4221: out = 16'(12563);
			4222: out = 16'(1205);
			4223: out = 16'(-10123);
			4224: out = 16'(-5344);
			4225: out = 16'(-1908);
			4226: out = 16'(5280);
			4227: out = 16'(8924);
			4228: out = 16'(1158);
			4229: out = 16'(-10911);
			4230: out = 16'(-11307);
			4231: out = 16'(4533);
			4232: out = 16'(8567);
			4233: out = 16'(7560);
			4234: out = 16'(1737);
			4235: out = 16'(-2098);
			4236: out = 16'(-932);
			4237: out = 16'(-2345);
			4238: out = 16'(5542);
			4239: out = 16'(8821);
			4240: out = 16'(5476);
			4241: out = 16'(-4290);
			4242: out = 16'(-9341);
			4243: out = 16'(-8010);
			4244: out = 16'(1317);
			4245: out = 16'(842);
			4246: out = 16'(-8937);
			4247: out = 16'(502);
			4248: out = 16'(3454);
			4249: out = 16'(-3923);
			4250: out = 16'(-7000);
			4251: out = 16'(-3362);
			4252: out = 16'(5924);
			4253: out = 16'(7751);
			4254: out = 16'(4175);
			4255: out = 16'(-6559);
			4256: out = 16'(-13283);
			4257: out = 16'(-10063);
			4258: out = 16'(-4354);
			4259: out = 16'(3172);
			4260: out = 16'(-944);
			4261: out = 16'(1683);
			4262: out = 16'(9815);
			4263: out = 16'(3950);
			4264: out = 16'(-708);
			4265: out = 16'(-422);
			4266: out = 16'(-3120);
			4267: out = 16'(-5638);
			4268: out = 16'(-5018);
			4269: out = 16'(-4056);
			4270: out = 16'(-2940);
			4271: out = 16'(-813);
			4272: out = 16'(-3577);
			4273: out = 16'(1586);
			4274: out = 16'(806);
			4275: out = 16'(-8322);
			4276: out = 16'(-3821);
			4277: out = 16'(9057);
			4278: out = 16'(6352);
			4279: out = 16'(-10642);
			4280: out = 16'(-14715);
			4281: out = 16'(-4939);
			4282: out = 16'(4285);
			4283: out = 16'(17086);
			4284: out = 16'(9750);
			4285: out = 16'(1226);
			4286: out = 16'(-256);
			4287: out = 16'(-741);
			4288: out = 16'(2711);
			4289: out = 16'(-3090);
			4290: out = 16'(-7224);
			4291: out = 16'(154);
			4292: out = 16'(9399);
			4293: out = 16'(535);
			4294: out = 16'(-7317);
			4295: out = 16'(-4151);
			4296: out = 16'(-238);
			4297: out = 16'(5354);
			4298: out = 16'(3576);
			4299: out = 16'(-3916);
			4300: out = 16'(-2521);
			4301: out = 16'(843);
			4302: out = 16'(914);
			4303: out = 16'(-855);
			4304: out = 16'(445);
			4305: out = 16'(4343);
			4306: out = 16'(-1319);
			4307: out = 16'(-6860);
			4308: out = 16'(-5855);
			4309: out = 16'(-1285);
			4310: out = 16'(-5589);
			4311: out = 16'(-11377);
			4312: out = 16'(-11273);
			4313: out = 16'(-4323);
			4314: out = 16'(1466);
			4315: out = 16'(5126);
			4316: out = 16'(5215);
			4317: out = 16'(1846);
			4318: out = 16'(804);
			4319: out = 16'(-2048);
			4320: out = 16'(-6098);
			4321: out = 16'(-1127);
			4322: out = 16'(4466);
			4323: out = 16'(4450);
			4324: out = 16'(928);
			4325: out = 16'(4872);
			4326: out = 16'(11216);
			4327: out = 16'(2137);
			4328: out = 16'(-12997);
			4329: out = 16'(-15151);
			4330: out = 16'(-10718);
			4331: out = 16'(-4966);
			4332: out = 16'(6398);
			4333: out = 16'(1208);
			4334: out = 16'(-9240);
			4335: out = 16'(-6124);
			4336: out = 16'(-1234);
			4337: out = 16'(7333);
			4338: out = 16'(13665);
			4339: out = 16'(8960);
			4340: out = 16'(-3608);
			4341: out = 16'(-10005);
			4342: out = 16'(-5488);
			4343: out = 16'(1081);
			4344: out = 16'(4100);
			4345: out = 16'(582);
			4346: out = 16'(-2189);
			4347: out = 16'(303);
			4348: out = 16'(-3634);
			4349: out = 16'(-11298);
			4350: out = 16'(1589);
			4351: out = 16'(6978);
			4352: out = 16'(685);
			4353: out = 16'(5422);
			4354: out = 16'(6942);
			4355: out = 16'(-6381);
			4356: out = 16'(-10080);
			4357: out = 16'(-4834);
			4358: out = 16'(3175);
			4359: out = 16'(5635);
			4360: out = 16'(9219);
			4361: out = 16'(5584);
			4362: out = 16'(3148);
			4363: out = 16'(5248);
			4364: out = 16'(8081);
			4365: out = 16'(7722);
			4366: out = 16'(-2583);
			4367: out = 16'(-11415);
			4368: out = 16'(-9073);
			4369: out = 16'(2577);
			4370: out = 16'(-2942);
			4371: out = 16'(-11270);
			4372: out = 16'(-6588);
			4373: out = 16'(-513);
			4374: out = 16'(7347);
			4375: out = 16'(13428);
			4376: out = 16'(9405);
			4377: out = 16'(-915);
			4378: out = 16'(-9605);
			4379: out = 16'(-5888);
			4380: out = 16'(2825);
			4381: out = 16'(12151);
			4382: out = 16'(5846);
			4383: out = 16'(1113);
			4384: out = 16'(7374);
			4385: out = 16'(10209);
			4386: out = 16'(-169);
			4387: out = 16'(-7723);
			4388: out = 16'(-6665);
			4389: out = 16'(1123);
			4390: out = 16'(5203);
			4391: out = 16'(2184);
			4392: out = 16'(1713);
			4393: out = 16'(2716);
			4394: out = 16'(5447);
			4395: out = 16'(-233);
			4396: out = 16'(-1419);
			4397: out = 16'(-115);
			4398: out = 16'(1216);
			4399: out = 16'(5491);
			4400: out = 16'(7321);
			4401: out = 16'(-3031);
			4402: out = 16'(-12512);
			4403: out = 16'(-11776);
			4404: out = 16'(-9836);
			4405: out = 16'(-1061);
			4406: out = 16'(4902);
			4407: out = 16'(1141);
			4408: out = 16'(-3792);
			4409: out = 16'(5717);
			4410: out = 16'(7559);
			4411: out = 16'(656);
			4412: out = 16'(-3063);
			4413: out = 16'(-2593);
			4414: out = 16'(2798);
			4415: out = 16'(4998);
			4416: out = 16'(6277);
			4417: out = 16'(2648);
			4418: out = 16'(-4452);
			4419: out = 16'(-6657);
			4420: out = 16'(1362);
			4421: out = 16'(4440);
			4422: out = 16'(1259);
			4423: out = 16'(2871);
			4424: out = 16'(3672);
			4425: out = 16'(-1968);
			4426: out = 16'(-5328);
			4427: out = 16'(-3581);
			4428: out = 16'(2770);
			4429: out = 16'(3002);
			4430: out = 16'(589);
			4431: out = 16'(1379);
			4432: out = 16'(32);
			4433: out = 16'(-896);
			4434: out = 16'(-3830);
			4435: out = 16'(2525);
			4436: out = 16'(6975);
			4437: out = 16'(1710);
			4438: out = 16'(599);
			4439: out = 16'(-645);
			4440: out = 16'(4122);
			4441: out = 16'(4273);
			4442: out = 16'(535);
			4443: out = 16'(-2388);
			4444: out = 16'(34);
			4445: out = 16'(1276);
			4446: out = 16'(-2019);
			4447: out = 16'(-262);
			4448: out = 16'(-875);
			4449: out = 16'(-1097);
			4450: out = 16'(-4496);
			4451: out = 16'(-779);
			4452: out = 16'(8989);
			4453: out = 16'(4449);
			4454: out = 16'(-3476);
			4455: out = 16'(-2443);
			4456: out = 16'(-719);
			4457: out = 16'(9584);
			4458: out = 16'(13340);
			4459: out = 16'(-2090);
			4460: out = 16'(-8337);
			4461: out = 16'(-8853);
			4462: out = 16'(2432);
			4463: out = 16'(4972);
			4464: out = 16'(-142);
			4465: out = 16'(5626);
			4466: out = 16'(13258);
			4467: out = 16'(9893);
			4468: out = 16'(-5932);
			4469: out = 16'(-15708);
			4470: out = 16'(-9676);
			4471: out = 16'(204);
			4472: out = 16'(8506);
			4473: out = 16'(11837);
			4474: out = 16'(4774);
			4475: out = 16'(-3665);
			4476: out = 16'(-170);
			4477: out = 16'(3361);
			4478: out = 16'(647);
			4479: out = 16'(-1614);
			4480: out = 16'(-5120);
			4481: out = 16'(-996);
			4482: out = 16'(3648);
			4483: out = 16'(5110);
			4484: out = 16'(1404);
			4485: out = 16'(-839);
			4486: out = 16'(-8374);
			4487: out = 16'(-9170);
			4488: out = 16'(-9065);
			4489: out = 16'(1826);
			4490: out = 16'(11631);
			4491: out = 16'(1709);
			4492: out = 16'(-2553);
			4493: out = 16'(3357);
			4494: out = 16'(8455);
			4495: out = 16'(-982);
			4496: out = 16'(-8811);
			4497: out = 16'(-4329);
			4498: out = 16'(4907);
			4499: out = 16'(4867);
			4500: out = 16'(1768);
			4501: out = 16'(-712);
			4502: out = 16'(988);
			4503: out = 16'(-2560);
			4504: out = 16'(-8636);
			4505: out = 16'(-3878);
			4506: out = 16'(5850);
			4507: out = 16'(4727);
			4508: out = 16'(337);
			4509: out = 16'(-4825);
			4510: out = 16'(-4781);
			4511: out = 16'(5843);
			4512: out = 16'(6451);
			4513: out = 16'(-2355);
			4514: out = 16'(-11074);
			4515: out = 16'(-3417);
			4516: out = 16'(10190);
			4517: out = 16'(15506);
			4518: out = 16'(7999);
			4519: out = 16'(3851);
			4520: out = 16'(523);
			4521: out = 16'(-3787);
			4522: out = 16'(-8355);
			4523: out = 16'(-12258);
			4524: out = 16'(277);
			4525: out = 16'(14610);
			4526: out = 16'(3912);
			4527: out = 16'(-7698);
			4528: out = 16'(1348);
			4529: out = 16'(6131);
			4530: out = 16'(3489);
			4531: out = 16'(-4345);
			4532: out = 16'(-3677);
			4533: out = 16'(-2979);
			4534: out = 16'(103);
			4535: out = 16'(-770);
			4536: out = 16'(3418);
			4537: out = 16'(10600);
			4538: out = 16'(11249);
			4539: out = 16'(-1824);
			4540: out = 16'(-6001);
			4541: out = 16'(-4761);
			4542: out = 16'(-1596);
			4543: out = 16'(942);
			4544: out = 16'(3224);
			4545: out = 16'(2639);
			4546: out = 16'(2591);
			4547: out = 16'(-4170);
			4548: out = 16'(-9454);
			4549: out = 16'(-1173);
			4550: out = 16'(-289);
			4551: out = 16'(4342);
			4552: out = 16'(5877);
			4553: out = 16'(5005);
			4554: out = 16'(-3586);
			4555: out = 16'(-7063);
			4556: out = 16'(-6318);
			4557: out = 16'(1815);
			4558: out = 16'(5296);
			4559: out = 16'(1495);
			4560: out = 16'(525);
			4561: out = 16'(-837);
			4562: out = 16'(-13322);
			4563: out = 16'(-15496);
			4564: out = 16'(-1320);
			4565: out = 16'(8237);
			4566: out = 16'(9868);
			4567: out = 16'(4582);
			4568: out = 16'(-342);
			4569: out = 16'(-7126);
			4570: out = 16'(489);
			4571: out = 16'(5642);
			4572: out = 16'(11775);
			4573: out = 16'(12076);
			4574: out = 16'(-1409);
			4575: out = 16'(-5539);
			4576: out = 16'(-3122);
			4577: out = 16'(1892);
			4578: out = 16'(1602);
			4579: out = 16'(-10918);
			4580: out = 16'(-5131);
			4581: out = 16'(5261);
			4582: out = 16'(5578);
			4583: out = 16'(6939);
			4584: out = 16'(7194);
			4585: out = 16'(4696);
			4586: out = 16'(-5464);
			4587: out = 16'(-13622);
			4588: out = 16'(-11433);
			4589: out = 16'(-1146);
			4590: out = 16'(-4835);
			4591: out = 16'(-4578);
			4592: out = 16'(9141);
			4593: out = 16'(6585);
			4594: out = 16'(-6435);
			4595: out = 16'(-4961);
			4596: out = 16'(-5327);
			4597: out = 16'(-1148);
			4598: out = 16'(4724);
			4599: out = 16'(7376);
			4600: out = 16'(-4340);
			4601: out = 16'(-9975);
			4602: out = 16'(-588);
			4603: out = 16'(11352);
			4604: out = 16'(12056);
			4605: out = 16'(2242);
			4606: out = 16'(-2666);
			4607: out = 16'(1412);
			4608: out = 16'(2471);
			4609: out = 16'(-6790);
			4610: out = 16'(-9604);
			4611: out = 16'(-7583);
			4612: out = 16'(-2426);
			4613: out = 16'(2783);
			4614: out = 16'(3472);
			4615: out = 16'(-1665);
			4616: out = 16'(2594);
			4617: out = 16'(5955);
			4618: out = 16'(12);
			4619: out = 16'(-11427);
			4620: out = 16'(-12847);
			4621: out = 16'(-3040);
			4622: out = 16'(7039);
			4623: out = 16'(7300);
			4624: out = 16'(-3877);
			4625: out = 16'(-9800);
			4626: out = 16'(-9976);
			4627: out = 16'(2599);
			4628: out = 16'(14591);
			4629: out = 16'(5516);
			4630: out = 16'(-4313);
			4631: out = 16'(-4483);
			4632: out = 16'(-1474);
			4633: out = 16'(3047);
			4634: out = 16'(772);
			4635: out = 16'(-5958);
			4636: out = 16'(-3397);
			4637: out = 16'(2924);
			4638: out = 16'(3952);
			4639: out = 16'(-3876);
			4640: out = 16'(-13233);
			4641: out = 16'(-10345);
			4642: out = 16'(6508);
			4643: out = 16'(10622);
			4644: out = 16'(7131);
			4645: out = 16'(3415);
			4646: out = 16'(-328);
			4647: out = 16'(-1596);
			4648: out = 16'(-8941);
			4649: out = 16'(-3535);
			4650: out = 16'(7900);
			4651: out = 16'(-2612);
			4652: out = 16'(-9199);
			4653: out = 16'(2122);
			4654: out = 16'(484);
			4655: out = 16'(-4403);
			4656: out = 16'(-6178);
			4657: out = 16'(-88);
			4658: out = 16'(1947);
			4659: out = 16'(-4115);
			4660: out = 16'(1784);
			4661: out = 16'(8726);
			4662: out = 16'(8009);
			4663: out = 16'(1671);
			4664: out = 16'(-3646);
			4665: out = 16'(-5534);
			4666: out = 16'(-6507);
			4667: out = 16'(-1602);
			4668: out = 16'(1405);
			4669: out = 16'(-1525);
			4670: out = 16'(-7139);
			4671: out = 16'(-6034);
			4672: out = 16'(10399);
			4673: out = 16'(10769);
			4674: out = 16'(-8412);
			4675: out = 16'(-11278);
			4676: out = 16'(-5176);
			4677: out = 16'(-3112);
			4678: out = 16'(81);
			4679: out = 16'(4647);
			4680: out = 16'(-1749);
			4681: out = 16'(-7598);
			4682: out = 16'(-152);
			4683: out = 16'(9820);
			4684: out = 16'(10720);
			4685: out = 16'(1515);
			4686: out = 16'(-6777);
			4687: out = 16'(577);
			4688: out = 16'(6708);
			4689: out = 16'(-4073);
			4690: out = 16'(-14004);
			4691: out = 16'(-10819);
			4692: out = 16'(-655);
			4693: out = 16'(5364);
			4694: out = 16'(1354);
			4695: out = 16'(-4010);
			4696: out = 16'(3258);
			4697: out = 16'(8556);
			4698: out = 16'(6610);
			4699: out = 16'(-1975);
			4700: out = 16'(-11623);
			4701: out = 16'(-8965);
			4702: out = 16'(-5609);
			4703: out = 16'(6840);
			4704: out = 16'(12633);
			4705: out = 16'(-553);
			4706: out = 16'(-5768);
			4707: out = 16'(2268);
			4708: out = 16'(8259);
			4709: out = 16'(6390);
			4710: out = 16'(-5328);
			4711: out = 16'(-9469);
			4712: out = 16'(-6284);
			4713: out = 16'(-2733);
			4714: out = 16'(7878);
			4715: out = 16'(3483);
			4716: out = 16'(-8418);
			4717: out = 16'(-6759);
			4718: out = 16'(745);
			4719: out = 16'(5308);
			4720: out = 16'(2443);
			4721: out = 16'(-4602);
			4722: out = 16'(-7327);
			4723: out = 16'(-9279);
			4724: out = 16'(433);
			4725: out = 16'(13423);
			4726: out = 16'(6264);
			4727: out = 16'(-7905);
			4728: out = 16'(-9348);
			4729: out = 16'(-8477);
			4730: out = 16'(-2539);
			4731: out = 16'(4289);
			4732: out = 16'(-358);
			4733: out = 16'(934);
			4734: out = 16'(8029);
			4735: out = 16'(3930);
			4736: out = 16'(-740);
			4737: out = 16'(-2389);
			4738: out = 16'(-3817);
			4739: out = 16'(4174);
			4740: out = 16'(6298);
			4741: out = 16'(5368);
			4742: out = 16'(-3327);
			4743: out = 16'(-2599);
			4744: out = 16'(6821);
			4745: out = 16'(8960);
			4746: out = 16'(-3918);
			4747: out = 16'(-8742);
			4748: out = 16'(-891);
			4749: out = 16'(4095);
			4750: out = 16'(1389);
			4751: out = 16'(-2744);
			4752: out = 16'(4835);
			4753: out = 16'(12448);
			4754: out = 16'(7114);
			4755: out = 16'(-2725);
			4756: out = 16'(-6556);
			4757: out = 16'(-2556);
			4758: out = 16'(-369);
			4759: out = 16'(-5820);
			4760: out = 16'(-4006);
			4761: out = 16'(3618);
			4762: out = 16'(4642);
			4763: out = 16'(1625);
			4764: out = 16'(1215);
			4765: out = 16'(689);
			4766: out = 16'(1220);
			4767: out = 16'(-2714);
			4768: out = 16'(3025);
			4769: out = 16'(1834);
			4770: out = 16'(4219);
			4771: out = 16'(7178);
			4772: out = 16'(5683);
			4773: out = 16'(-5368);
			4774: out = 16'(-9712);
			4775: out = 16'(-5763);
			4776: out = 16'(-920);
			4777: out = 16'(-2236);
			4778: out = 16'(-4425);
			4779: out = 16'(503);
			4780: out = 16'(-309);
			4781: out = 16'(-1542);
			4782: out = 16'(-66);
			4783: out = 16'(107);
			4784: out = 16'(1994);
			4785: out = 16'(13033);
			4786: out = 16'(17390);
			4787: out = 16'(917);
			4788: out = 16'(-15305);
			4789: out = 16'(-13389);
			4790: out = 16'(-5011);
			4791: out = 16'(6173);
			4792: out = 16'(12000);
			4793: out = 16'(-3550);
			4794: out = 16'(-7595);
			4795: out = 16'(4137);
			4796: out = 16'(12393);
			4797: out = 16'(3687);
			4798: out = 16'(-9106);
			4799: out = 16'(-7845);
			4800: out = 16'(-2379);
			4801: out = 16'(7880);
			4802: out = 16'(11427);
			4803: out = 16'(-577);
			4804: out = 16'(-8327);
			4805: out = 16'(949);
			4806: out = 16'(2677);
			4807: out = 16'(4573);
			4808: out = 16'(4886);
			4809: out = 16'(2849);
			4810: out = 16'(-3701);
			4811: out = 16'(-9488);
			4812: out = 16'(-508);
			4813: out = 16'(9257);
			4814: out = 16'(6806);
			4815: out = 16'(-5113);
			4816: out = 16'(-9562);
			4817: out = 16'(-6517);
			4818: out = 16'(6582);
			4819: out = 16'(15768);
			4820: out = 16'(4992);
			4821: out = 16'(-3151);
			4822: out = 16'(-2000);
			4823: out = 16'(6243);
			4824: out = 16'(1772);
			4825: out = 16'(-1716);
			4826: out = 16'(2534);
			4827: out = 16'(3593);
			4828: out = 16'(2937);
			4829: out = 16'(863);
			4830: out = 16'(-712);
			4831: out = 16'(-4796);
			4832: out = 16'(-7589);
			4833: out = 16'(-5022);
			4834: out = 16'(4855);
			4835: out = 16'(10097);
			4836: out = 16'(5929);
			4837: out = 16'(-4280);
			4838: out = 16'(-1837);
			4839: out = 16'(2275);
			4840: out = 16'(2634);
			4841: out = 16'(9600);
			4842: out = 16'(14254);
			4843: out = 16'(3212);
			4844: out = 16'(-11395);
			4845: out = 16'(-9044);
			4846: out = 16'(3781);
			4847: out = 16'(11062);
			4848: out = 16'(12);
			4849: out = 16'(-8145);
			4850: out = 16'(-2589);
			4851: out = 16'(2653);
			4852: out = 16'(4673);
			4853: out = 16'(-4128);
			4854: out = 16'(-10824);
			4855: out = 16'(-3546);
			4856: out = 16'(4592);
			4857: out = 16'(8603);
			4858: out = 16'(7903);
			4859: out = 16'(570);
			4860: out = 16'(-759);
			4861: out = 16'(-2118);
			4862: out = 16'(2419);
			4863: out = 16'(4664);
			4864: out = 16'(7204);
			4865: out = 16'(8414);
			4866: out = 16'(1063);
			4867: out = 16'(-13180);
			4868: out = 16'(-15096);
			4869: out = 16'(-3650);
			4870: out = 16'(1266);
			4871: out = 16'(518);
			4872: out = 16'(3026);
			4873: out = 16'(7833);
			4874: out = 16'(1753);
			4875: out = 16'(-6432);
			4876: out = 16'(-829);
			4877: out = 16'(10154);
			4878: out = 16'(10474);
			4879: out = 16'(1011);
			4880: out = 16'(-5785);
			4881: out = 16'(-5752);
			4882: out = 16'(-4592);
			4883: out = 16'(-3293);
			4884: out = 16'(-2180);
			4885: out = 16'(-39);
			4886: out = 16'(8492);
			4887: out = 16'(2033);
			4888: out = 16'(1984);
			4889: out = 16'(417);
			4890: out = 16'(-2221);
			4891: out = 16'(5805);
			4892: out = 16'(7542);
			4893: out = 16'(3361);
			4894: out = 16'(-7322);
			4895: out = 16'(-8496);
			4896: out = 16'(874);
			4897: out = 16'(5591);
			4898: out = 16'(2575);
			4899: out = 16'(-3416);
			4900: out = 16'(-8120);
			4901: out = 16'(206);
			4902: out = 16'(7968);
			4903: out = 16'(5288);
			4904: out = 16'(-4112);
			4905: out = 16'(-7732);
			4906: out = 16'(-2255);
			4907: out = 16'(4942);
			4908: out = 16'(11535);
			4909: out = 16'(3596);
			4910: out = 16'(-8333);
			4911: out = 16'(-11434);
			4912: out = 16'(-4232);
			4913: out = 16'(7973);
			4914: out = 16'(13580);
			4915: out = 16'(4990);
			4916: out = 16'(-6309);
			4917: out = 16'(-6216);
			4918: out = 16'(-4013);
			4919: out = 16'(2578);
			4920: out = 16'(5406);
			4921: out = 16'(-3711);
			4922: out = 16'(-11772);
			4923: out = 16'(-1747);
			4924: out = 16'(10575);
			4925: out = 16'(3576);
			4926: out = 16'(-5226);
			4927: out = 16'(-6156);
			4928: out = 16'(-579);
			4929: out = 16'(10243);
			4930: out = 16'(10125);
			4931: out = 16'(6408);
			4932: out = 16'(-56);
			4933: out = 16'(-6865);
			4934: out = 16'(-5914);
			4935: out = 16'(-3521);
			4936: out = 16'(3745);
			4937: out = 16'(6987);
			4938: out = 16'(-3643);
			4939: out = 16'(-11073);
			4940: out = 16'(-7041);
			4941: out = 16'(-528);
			4942: out = 16'(10362);
			4943: out = 16'(11018);
			4944: out = 16'(1557);
			4945: out = 16'(-9511);
			4946: out = 16'(-12003);
			4947: out = 16'(-8242);
			4948: out = 16'(-2478);
			4949: out = 16'(4570);
			4950: out = 16'(7681);
			4951: out = 16'(2777);
			4952: out = 16'(-5024);
			4953: out = 16'(-1090);
			4954: out = 16'(1863);
			4955: out = 16'(3958);
			4956: out = 16'(3296);
			4957: out = 16'(-1067);
			4958: out = 16'(-1716);
			4959: out = 16'(1360);
			4960: out = 16'(7833);
			4961: out = 16'(6224);
			4962: out = 16'(-2801);
			4963: out = 16'(-9846);
			4964: out = 16'(-2776);
			4965: out = 16'(-2492);
			4966: out = 16'(4646);
			4967: out = 16'(7017);
			4968: out = 16'(1588);
			4969: out = 16'(-2190);
			4970: out = 16'(1208);
			4971: out = 16'(717);
			4972: out = 16'(-5379);
			4973: out = 16'(-6731);
			4974: out = 16'(1471);
			4975: out = 16'(1870);
			4976: out = 16'(-3017);
			4977: out = 16'(-3969);
			4978: out = 16'(-4320);
			4979: out = 16'(-4195);
			4980: out = 16'(-4920);
			4981: out = 16'(-1229);
			4982: out = 16'(-1853);
			4983: out = 16'(-2127);
			4984: out = 16'(3894);
			4985: out = 16'(6801);
			4986: out = 16'(-2924);
			4987: out = 16'(-17360);
			4988: out = 16'(-8919);
			4989: out = 16'(3671);
			4990: out = 16'(9076);
			4991: out = 16'(11686);
			4992: out = 16'(4058);
			4993: out = 16'(-4783);
			4994: out = 16'(-2529);
			4995: out = 16'(-2749);
			4996: out = 16'(-1349);
			4997: out = 16'(-7127);
			4998: out = 16'(-7517);
			4999: out = 16'(7942);
			5000: out = 16'(11571);
			5001: out = 16'(2026);
			5002: out = 16'(-357);
			5003: out = 16'(1241);
			5004: out = 16'(-1519);
			5005: out = 16'(-9688);
			5006: out = 16'(-5898);
			5007: out = 16'(1517);
			5008: out = 16'(7857);
			5009: out = 16'(4771);
			5010: out = 16'(-9600);
			5011: out = 16'(-6378);
			5012: out = 16'(5340);
			5013: out = 16'(6744);
			5014: out = 16'(1254);
			5015: out = 16'(-3985);
			5016: out = 16'(-2808);
			5017: out = 16'(4817);
			5018: out = 16'(7783);
			5019: out = 16'(3052);
			5020: out = 16'(-4354);
			5021: out = 16'(-3631);
			5022: out = 16'(-432);
			5023: out = 16'(-2079);
			5024: out = 16'(-8464);
			5025: out = 16'(-10912);
			5026: out = 16'(-4127);
			5027: out = 16'(8421);
			5028: out = 16'(5027);
			5029: out = 16'(-6025);
			5030: out = 16'(-8572);
			5031: out = 16'(-409);
			5032: out = 16'(8354);
			5033: out = 16'(9871);
			5034: out = 16'(6709);
			5035: out = 16'(-1017);
			5036: out = 16'(-1550);
			5037: out = 16'(-2543);
			5038: out = 16'(-2425);
			5039: out = 16'(-3933);
			5040: out = 16'(-3958);
			5041: out = 16'(1531);
			5042: out = 16'(3466);
			5043: out = 16'(5609);
			5044: out = 16'(1425);
			5045: out = 16'(180);
			5046: out = 16'(-1466);
			5047: out = 16'(297);
			5048: out = 16'(1808);
			5049: out = 16'(597);
			5050: out = 16'(3374);
			5051: out = 16'(3751);
			5052: out = 16'(-4934);
			5053: out = 16'(-10851);
			5054: out = 16'(-9263);
			5055: out = 16'(-8314);
			5056: out = 16'(-2288);
			5057: out = 16'(4684);
			5058: out = 16'(4241);
			5059: out = 16'(-5954);
			5060: out = 16'(-10906);
			5061: out = 16'(-7607);
			5062: out = 16'(-1216);
			5063: out = 16'(3042);
			5064: out = 16'(3792);
			5065: out = 16'(5595);
			5066: out = 16'(-109);
			5067: out = 16'(-1656);
			5068: out = 16'(972);
			5069: out = 16'(1485);
			5070: out = 16'(-1622);
			5071: out = 16'(499);
			5072: out = 16'(-932);
			5073: out = 16'(649);
			5074: out = 16'(-5146);
			5075: out = 16'(-10218);
			5076: out = 16'(-1611);
			5077: out = 16'(3972);
			5078: out = 16'(5564);
			5079: out = 16'(235);
			5080: out = 16'(-3960);
			5081: out = 16'(-5682);
			5082: out = 16'(-2722);
			5083: out = 16'(8556);
			5084: out = 16'(8789);
			5085: out = 16'(4967);
			5086: out = 16'(-5110);
			5087: out = 16'(-4906);
			5088: out = 16'(3328);
			5089: out = 16'(8281);
			5090: out = 16'(9117);
			5091: out = 16'(64);
			5092: out = 16'(-3866);
			5093: out = 16'(-1891);
			5094: out = 16'(3070);
			5095: out = 16'(-735);
			5096: out = 16'(-2708);
			5097: out = 16'(3467);
			5098: out = 16'(3728);
			5099: out = 16'(-5456);
			5100: out = 16'(-6229);
			5101: out = 16'(-523);
			5102: out = 16'(1578);
			5103: out = 16'(4792);
			5104: out = 16'(3783);
			5105: out = 16'(-4141);
			5106: out = 16'(-8128);
			5107: out = 16'(-7250);
			5108: out = 16'(-5976);
			5109: out = 16'(-675);
			5110: out = 16'(13051);
			5111: out = 16'(8715);
			5112: out = 16'(-2127);
			5113: out = 16'(-1245);
			5114: out = 16'(6477);
			5115: out = 16'(11901);
			5116: out = 16'(4610);
			5117: out = 16'(-7655);
			5118: out = 16'(-6223);
			5119: out = 16'(645);
			5120: out = 16'(-4418);
			5121: out = 16'(-7497);
			5122: out = 16'(-5610);
			5123: out = 16'(1856);
			5124: out = 16'(5932);
			5125: out = 16'(6726);
			5126: out = 16'(5462);
			5127: out = 16'(-2301);
			5128: out = 16'(-4601);
			5129: out = 16'(-6713);
			5130: out = 16'(3746);
			5131: out = 16'(4300);
			5132: out = 16'(-1012);
			5133: out = 16'(4009);
			5134: out = 16'(7529);
			5135: out = 16'(2221);
			5136: out = 16'(-7968);
			5137: out = 16'(-6731);
			5138: out = 16'(2637);
			5139: out = 16'(8939);
			5140: out = 16'(2015);
			5141: out = 16'(-3403);
			5142: out = 16'(-6656);
			5143: out = 16'(2853);
			5144: out = 16'(7309);
			5145: out = 16'(-29);
			5146: out = 16'(-1071);
			5147: out = 16'(-491);
			5148: out = 16'(-1480);
			5149: out = 16'(2295);
			5150: out = 16'(5215);
			5151: out = 16'(-3508);
			5152: out = 16'(-2119);
			5153: out = 16'(4024);
			5154: out = 16'(7752);
			5155: out = 16'(5292);
			5156: out = 16'(-1448);
			5157: out = 16'(-898);
			5158: out = 16'(538);
			5159: out = 16'(-2640);
			5160: out = 16'(-6293);
			5161: out = 16'(-274);
			5162: out = 16'(1697);
			5163: out = 16'(-4932);
			5164: out = 16'(-4391);
			5165: out = 16'(-3291);
			5166: out = 16'(6594);
			5167: out = 16'(13431);
			5168: out = 16'(3498);
			5169: out = 16'(-1884);
			5170: out = 16'(-1059);
			5171: out = 16'(-1347);
			5172: out = 16'(4559);
			5173: out = 16'(5452);
			5174: out = 16'(4200);
			5175: out = 16'(-2274);
			5176: out = 16'(-8285);
			5177: out = 16'(-8200);
			5178: out = 16'(-8411);
			5179: out = 16'(530);
			5180: out = 16'(11337);
			5181: out = 16'(8159);
			5182: out = 16'(-3369);
			5183: out = 16'(-13392);
			5184: out = 16'(-8722);
			5185: out = 16'(2148);
			5186: out = 16'(11283);
			5187: out = 16'(14837);
			5188: out = 16'(-2046);
			5189: out = 16'(-11627);
			5190: out = 16'(-5478);
			5191: out = 16'(9388);
			5192: out = 16'(12276);
			5193: out = 16'(-3937);
			5194: out = 16'(-5982);
			5195: out = 16'(718);
			5196: out = 16'(6083);
			5197: out = 16'(8365);
			5198: out = 16'(-3666);
			5199: out = 16'(-6692);
			5200: out = 16'(3625);
			5201: out = 16'(8173);
			5202: out = 16'(5218);
			5203: out = 16'(-1136);
			5204: out = 16'(-926);
			5205: out = 16'(4096);
			5206: out = 16'(-2139);
			5207: out = 16'(-5534);
			5208: out = 16'(-77);
			5209: out = 16'(3289);
			5210: out = 16'(2291);
			5211: out = 16'(-5803);
			5212: out = 16'(-3705);
			5213: out = 16'(1493);
			5214: out = 16'(-1181);
			5215: out = 16'(-2267);
			5216: out = 16'(3304);
			5217: out = 16'(334);
			5218: out = 16'(-740);
			5219: out = 16'(1252);
			5220: out = 16'(-2006);
			5221: out = 16'(-4802);
			5222: out = 16'(-5857);
			5223: out = 16'(2591);
			5224: out = 16'(5442);
			5225: out = 16'(1692);
			5226: out = 16'(2408);
			5227: out = 16'(2818);
			5228: out = 16'(-6528);
			5229: out = 16'(-10234);
			5230: out = 16'(-3427);
			5231: out = 16'(6645);
			5232: out = 16'(13203);
			5233: out = 16'(2673);
			5234: out = 16'(-12573);
			5235: out = 16'(-7386);
			5236: out = 16'(5550);
			5237: out = 16'(12378);
			5238: out = 16'(10860);
			5239: out = 16'(1492);
			5240: out = 16'(-4246);
			5241: out = 16'(-203);
			5242: out = 16'(-910);
			5243: out = 16'(-2813);
			5244: out = 16'(-4608);
			5245: out = 16'(-8735);
			5246: out = 16'(387);
			5247: out = 16'(8152);
			5248: out = 16'(5960);
			5249: out = 16'(95);
			5250: out = 16'(85);
			5251: out = 16'(-4094);
			5252: out = 16'(-2823);
			5253: out = 16'(-2096);
			5254: out = 16'(-370);
			5255: out = 16'(3634);
			5256: out = 16'(1442);
			5257: out = 16'(3465);
			5258: out = 16'(3935);
			5259: out = 16'(280);
			5260: out = 16'(-1229);
			5261: out = 16'(-3449);
			5262: out = 16'(-1886);
			5263: out = 16'(3705);
			5264: out = 16'(-795);
			5265: out = 16'(-499);
			5266: out = 16'(7034);
			5267: out = 16'(8470);
			5268: out = 16'(-337);
			5269: out = 16'(-8926);
			5270: out = 16'(-10364);
			5271: out = 16'(-532);
			5272: out = 16'(2926);
			5273: out = 16'(2954);
			5274: out = 16'(3643);
			5275: out = 16'(3068);
			5276: out = 16'(-668);
			5277: out = 16'(-2286);
			5278: out = 16'(-40);
			5279: out = 16'(352);
			5280: out = 16'(-842);
			5281: out = 16'(324);
			5282: out = 16'(-613);
			5283: out = 16'(-3373);
			5284: out = 16'(-7212);
			5285: out = 16'(-3012);
			5286: out = 16'(4640);
			5287: out = 16'(7105);
			5288: out = 16'(2639);
			5289: out = 16'(2011);
			5290: out = 16'(2928);
			5291: out = 16'(-772);
			5292: out = 16'(-7508);
			5293: out = 16'(-15565);
			5294: out = 16'(-12057);
			5295: out = 16'(2570);
			5296: out = 16'(13702);
			5297: out = 16'(6551);
			5298: out = 16'(-2575);
			5299: out = 16'(-1613);
			5300: out = 16'(4881);
			5301: out = 16'(6907);
			5302: out = 16'(-3742);
			5303: out = 16'(-13084);
			5304: out = 16'(-9201);
			5305: out = 16'(7252);
			5306: out = 16'(11405);
			5307: out = 16'(-834);
			5308: out = 16'(1901);
			5309: out = 16'(7365);
			5310: out = 16'(7488);
			5311: out = 16'(-4092);
			5312: out = 16'(-6820);
			5313: out = 16'(-1660);
			5314: out = 16'(7730);
			5315: out = 16'(9019);
			5316: out = 16'(584);
			5317: out = 16'(-3475);
			5318: out = 16'(1784);
			5319: out = 16'(1837);
			5320: out = 16'(-2463);
			5321: out = 16'(758);
			5322: out = 16'(1542);
			5323: out = 16'(-4327);
			5324: out = 16'(-12488);
			5325: out = 16'(-6102);
			5326: out = 16'(-3769);
			5327: out = 16'(-4533);
			5328: out = 16'(-1893);
			5329: out = 16'(4926);
			5330: out = 16'(-867);
			5331: out = 16'(-5199);
			5332: out = 16'(2082);
			5333: out = 16'(8974);
			5334: out = 16'(7304);
			5335: out = 16'(673);
			5336: out = 16'(-3052);
			5337: out = 16'(-3529);
			5338: out = 16'(-3012);
			5339: out = 16'(-2517);
			5340: out = 16'(-8489);
			5341: out = 16'(-12589);
			5342: out = 16'(-168);
			5343: out = 16'(7525);
			5344: out = 16'(7289);
			5345: out = 16'(7636);
			5346: out = 16'(7125);
			5347: out = 16'(3030);
			5348: out = 16'(-8309);
			5349: out = 16'(-10948);
			5350: out = 16'(-6690);
			5351: out = 16'(-1903);
			5352: out = 16'(6587);
			5353: out = 16'(4662);
			5354: out = 16'(-2835);
			5355: out = 16'(-6271);
			5356: out = 16'(-3130);
			5357: out = 16'(12391);
			5358: out = 16'(16964);
			5359: out = 16'(716);
			5360: out = 16'(-15586);
			5361: out = 16'(-11873);
			5362: out = 16'(-5381);
			5363: out = 16'(4404);
			5364: out = 16'(3556);
			5365: out = 16'(-3979);
			5366: out = 16'(-1728);
			5367: out = 16'(8341);
			5368: out = 16'(10727);
			5369: out = 16'(3650);
			5370: out = 16'(-7572);
			5371: out = 16'(-10759);
			5372: out = 16'(-3583);
			5373: out = 16'(7112);
			5374: out = 16'(8593);
			5375: out = 16'(-2386);
			5376: out = 16'(-8903);
			5377: out = 16'(-1824);
			5378: out = 16'(4058);
			5379: out = 16'(517);
			5380: out = 16'(1196);
			5381: out = 16'(1202);
			5382: out = 16'(-4343);
			5383: out = 16'(-6391);
			5384: out = 16'(2284);
			5385: out = 16'(6129);
			5386: out = 16'(6504);
			5387: out = 16'(-6685);
			5388: out = 16'(-5510);
			5389: out = 16'(11);
			5390: out = 16'(-492);
			5391: out = 16'(7515);
			5392: out = 16'(8870);
			5393: out = 16'(-3205);
			5394: out = 16'(-13220);
			5395: out = 16'(-12820);
			5396: out = 16'(-8654);
			5397: out = 16'(2049);
			5398: out = 16'(7551);
			5399: out = 16'(2095);
			5400: out = 16'(-3968);
			5401: out = 16'(2587);
			5402: out = 16'(1532);
			5403: out = 16'(-395);
			5404: out = 16'(3951);
			5405: out = 16'(1546);
			5406: out = 16'(2556);
			5407: out = 16'(5257);
			5408: out = 16'(5664);
			5409: out = 16'(1200);
			5410: out = 16'(-8998);
			5411: out = 16'(-9134);
			5412: out = 16'(-5935);
			5413: out = 16'(-1841);
			5414: out = 16'(5858);
			5415: out = 16'(1398);
			5416: out = 16'(-5227);
			5417: out = 16'(607);
			5418: out = 16'(441);
			5419: out = 16'(1312);
			5420: out = 16'(3653);
			5421: out = 16'(-1329);
			5422: out = 16'(-9172);
			5423: out = 16'(-8893);
			5424: out = 16'(-216);
			5425: out = 16'(2896);
			5426: out = 16'(5573);
			5427: out = 16'(-1282);
			5428: out = 16'(-4855);
			5429: out = 16'(8037);
			5430: out = 16'(13064);
			5431: out = 16'(4635);
			5432: out = 16'(-4640);
			5433: out = 16'(-2282);
			5434: out = 16'(3315);
			5435: out = 16'(2467);
			5436: out = 16'(-1084);
			5437: out = 16'(1408);
			5438: out = 16'(-1804);
			5439: out = 16'(-4132);
			5440: out = 16'(205);
			5441: out = 16'(-2982);
			5442: out = 16'(-9657);
			5443: out = 16'(-8018);
			5444: out = 16'(-6314);
			5445: out = 16'(481);
			5446: out = 16'(9805);
			5447: out = 16'(11596);
			5448: out = 16'(-1582);
			5449: out = 16'(-7001);
			5450: out = 16'(-3082);
			5451: out = 16'(1833);
			5452: out = 16'(3683);
			5453: out = 16'(1680);
			5454: out = 16'(5743);
			5455: out = 16'(2276);
			5456: out = 16'(1436);
			5457: out = 16'(5696);
			5458: out = 16'(3997);
			5459: out = 16'(-8858);
			5460: out = 16'(-16063);
			5461: out = 16'(-11713);
			5462: out = 16'(-3447);
			5463: out = 16'(11386);
			5464: out = 16'(9166);
			5465: out = 16'(-5228);
			5466: out = 16'(-7176);
			5467: out = 16'(-2233);
			5468: out = 16'(2533);
			5469: out = 16'(3996);
			5470: out = 16'(7476);
			5471: out = 16'(3501);
			5472: out = 16'(-2563);
			5473: out = 16'(1590);
			5474: out = 16'(3930);
			5475: out = 16'(1804);
			5476: out = 16'(-3056);
			5477: out = 16'(-4728);
			5478: out = 16'(-873);
			5479: out = 16'(163);
			5480: out = 16'(4694);
			5481: out = 16'(4160);
			5482: out = 16'(-3101);
			5483: out = 16'(-13066);
			5484: out = 16'(-9587);
			5485: out = 16'(-1279);
			5486: out = 16'(6355);
			5487: out = 16'(9647);
			5488: out = 16'(5358);
			5489: out = 16'(535);
			5490: out = 16'(-2453);
			5491: out = 16'(-7156);
			5492: out = 16'(-6133);
			5493: out = 16'(143);
			5494: out = 16'(-1575);
			5495: out = 16'(-4900);
			5496: out = 16'(-4016);
			5497: out = 16'(6677);
			5498: out = 16'(6729);
			5499: out = 16'(2167);
			5500: out = 16'(5428);
			5501: out = 16'(7064);
			5502: out = 16'(8780);
			5503: out = 16'(654);
			5504: out = 16'(-2278);
			5505: out = 16'(-2652);
			5506: out = 16'(-2172);
			5507: out = 16'(-3605);
			5508: out = 16'(-1997);
			5509: out = 16'(-5833);
			5510: out = 16'(-7045);
			5511: out = 16'(-1846);
			5512: out = 16'(-452);
			5513: out = 16'(1741);
			5514: out = 16'(6552);
			5515: out = 16'(563);
			5516: out = 16'(-1011);
			5517: out = 16'(5178);
			5518: out = 16'(6787);
			5519: out = 16'(411);
			5520: out = 16'(-7733);
			5521: out = 16'(-9912);
			5522: out = 16'(-5200);
			5523: out = 16'(8392);
			5524: out = 16'(9256);
			5525: out = 16'(-3297);
			5526: out = 16'(-5204);
			5527: out = 16'(-1367);
			5528: out = 16'(6144);
			5529: out = 16'(6270);
			5530: out = 16'(1538);
			5531: out = 16'(-1676);
			5532: out = 16'(-2466);
			5533: out = 16'(247);
			5534: out = 16'(-295);
			5535: out = 16'(5560);
			5536: out = 16'(9249);
			5537: out = 16'(5679);
			5538: out = 16'(-2172);
			5539: out = 16'(-7593);
			5540: out = 16'(-3350);
			5541: out = 16'(1272);
			5542: out = 16'(2719);
			5543: out = 16'(1556);
			5544: out = 16'(3229);
			5545: out = 16'(6622);
			5546: out = 16'(10018);
			5547: out = 16'(5803);
			5548: out = 16'(-1006);
			5549: out = 16'(-4731);
			5550: out = 16'(-5620);
			5551: out = 16'(-8333);
			5552: out = 16'(-2214);
			5553: out = 16'(6811);
			5554: out = 16'(1868);
			5555: out = 16'(-6247);
			5556: out = 16'(-6688);
			5557: out = 16'(-1934);
			5558: out = 16'(6285);
			5559: out = 16'(5096);
			5560: out = 16'(-1091);
			5561: out = 16'(-3521);
			5562: out = 16'(-5092);
			5563: out = 16'(-2515);
			5564: out = 16'(8102);
			5565: out = 16'(5696);
			5566: out = 16'(-10298);
			5567: out = 16'(-6592);
			5568: out = 16'(-1379);
			5569: out = 16'(2023);
			5570: out = 16'(9500);
			5571: out = 16'(4370);
			5572: out = 16'(972);
			5573: out = 16'(1946);
			5574: out = 16'(2897);
			5575: out = 16'(3953);
			5576: out = 16'(-4097);
			5577: out = 16'(-5945);
			5578: out = 16'(2898);
			5579: out = 16'(1251);
			5580: out = 16'(-814);
			5581: out = 16'(7263);
			5582: out = 16'(6005);
			5583: out = 16'(-5572);
			5584: out = 16'(-14777);
			5585: out = 16'(-11118);
			5586: out = 16'(1624);
			5587: out = 16'(9244);
			5588: out = 16'(10807);
			5589: out = 16'(5176);
			5590: out = 16'(-3529);
			5591: out = 16'(-4163);
			5592: out = 16'(-537);
			5593: out = 16'(1148);
			5594: out = 16'(-61);
			5595: out = 16'(1230);
			5596: out = 16'(8444);
			5597: out = 16'(638);
			5598: out = 16'(2710);
			5599: out = 16'(8894);
			5600: out = 16'(9949);
			5601: out = 16'(2004);
			5602: out = 16'(-6694);
			5603: out = 16'(-8590);
			5604: out = 16'(-1310);
			5605: out = 16'(1748);
			5606: out = 16'(-3955);
			5607: out = 16'(-580);
			5608: out = 16'(7287);
			5609: out = 16'(2993);
			5610: out = 16'(-7856);
			5611: out = 16'(-9843);
			5612: out = 16'(-7456);
			5613: out = 16'(440);
			5614: out = 16'(15129);
			5615: out = 16'(6496);
			5616: out = 16'(-6737);
			5617: out = 16'(-8870);
			5618: out = 16'(1581);
			5619: out = 16'(13179);
			5620: out = 16'(9934);
			5621: out = 16'(2373);
			5622: out = 16'(-1900);
			5623: out = 16'(1352);
			5624: out = 16'(-811);
			5625: out = 16'(-4896);
			5626: out = 16'(-3763);
			5627: out = 16'(-822);
			5628: out = 16'(2770);
			5629: out = 16'(2345);
			5630: out = 16'(5435);
			5631: out = 16'(-153);
			5632: out = 16'(1407);
			5633: out = 16'(-1747);
			5634: out = 16'(976);
			5635: out = 16'(5061);
			5636: out = 16'(2543);
			5637: out = 16'(1263);
			5638: out = 16'(2200);
			5639: out = 16'(1556);
			5640: out = 16'(-4447);
			5641: out = 16'(-8469);
			5642: out = 16'(-6850);
			5643: out = 16'(-4672);
			5644: out = 16'(-3704);
			5645: out = 16'(1813);
			5646: out = 16'(3553);
			5647: out = 16'(-9447);
			5648: out = 16'(-17129);
			5649: out = 16'(-3742);
			5650: out = 16'(3424);
			5651: out = 16'(10936);
			5652: out = 16'(11324);
			5653: out = 16'(3671);
			5654: out = 16'(-8725);
			5655: out = 16'(-15077);
			5656: out = 16'(-4482);
			5657: out = 16'(8504);
			5658: out = 16'(14893);
			5659: out = 16'(6569);
			5660: out = 16'(-9190);
			5661: out = 16'(-10054);
			5662: out = 16'(-2821);
			5663: out = 16'(5750);
			5664: out = 16'(6503);
			5665: out = 16'(3812);
			5666: out = 16'(-36);
			5667: out = 16'(-2251);
			5668: out = 16'(1795);
			5669: out = 16'(349);
			5670: out = 16'(1564);
			5671: out = 16'(2460);
			5672: out = 16'(-594);
			5673: out = 16'(713);
			5674: out = 16'(5759);
			5675: out = 16'(8001);
			5676: out = 16'(6667);
			5677: out = 16'(1364);
			5678: out = 16'(-2816);
			5679: out = 16'(-4240);
			5680: out = 16'(-2868);
			5681: out = 16'(-6950);
			5682: out = 16'(-3886);
			5683: out = 16'(2576);
			5684: out = 16'(-217);
			5685: out = 16'(-5846);
			5686: out = 16'(-10170);
			5687: out = 16'(-8652);
			5688: out = 16'(835);
			5689: out = 16'(9317);
			5690: out = 16'(10076);
			5691: out = 16'(-4002);
			5692: out = 16'(-13570);
			5693: out = 16'(-6579);
			5694: out = 16'(4711);
			5695: out = 16'(12923);
			5696: out = 16'(8354);
			5697: out = 16'(-386);
			5698: out = 16'(-6250);
			5699: out = 16'(-10032);
			5700: out = 16'(-838);
			5701: out = 16'(8939);
			5702: out = 16'(4726);
			5703: out = 16'(2434);
			5704: out = 16'(2140);
			5705: out = 16'(-1406);
			5706: out = 16'(-7394);
			5707: out = 16'(-10151);
			5708: out = 16'(1105);
			5709: out = 16'(11373);
			5710: out = 16'(1641);
			5711: out = 16'(-4903);
			5712: out = 16'(1762);
			5713: out = 16'(3140);
			5714: out = 16'(2364);
			5715: out = 16'(-2990);
			5716: out = 16'(-4631);
			5717: out = 16'(-1540);
			5718: out = 16'(-1557);
			5719: out = 16'(2980);
			5720: out = 16'(1725);
			5721: out = 16'(1355);
			5722: out = 16'(5744);
			5723: out = 16'(6966);
			5724: out = 16'(43);
			5725: out = 16'(-8825);
			5726: out = 16'(-6397);
			5727: out = 16'(683);
			5728: out = 16'(7254);
			5729: out = 16'(8349);
			5730: out = 16'(4218);
			5731: out = 16'(1501);
			5732: out = 16'(1071);
			5733: out = 16'(-2523);
			5734: out = 16'(-3098);
			5735: out = 16'(-5556);
			5736: out = 16'(-4662);
			5737: out = 16'(-3471);
			5738: out = 16'(2914);
			5739: out = 16'(2918);
			5740: out = 16'(-4390);
			5741: out = 16'(-9155);
			5742: out = 16'(-5428);
			5743: out = 16'(-543);
			5744: out = 16'(5654);
			5745: out = 16'(7535);
			5746: out = 16'(419);
			5747: out = 16'(-5961);
			5748: out = 16'(-8753);
			5749: out = 16'(-2375);
			5750: out = 16'(-800);
			5751: out = 16'(-1468);
			5752: out = 16'(673);
			5753: out = 16'(1928);
			5754: out = 16'(412);
			5755: out = 16'(-793);
			5756: out = 16'(-3568);
			5757: out = 16'(-2720);
			5758: out = 16'(-761);
			5759: out = 16'(-1648);
			5760: out = 16'(4411);
			5761: out = 16'(7065);
			5762: out = 16'(-1556);
			5763: out = 16'(-11474);
			5764: out = 16'(-12881);
			5765: out = 16'(-789);
			5766: out = 16'(12298);
			5767: out = 16'(6444);
			5768: out = 16'(-5516);
			5769: out = 16'(-4557);
			5770: out = 16'(-4650);
			5771: out = 16'(-4721);
			5772: out = 16'(1386);
			5773: out = 16'(1014);
			5774: out = 16'(1790);
			5775: out = 16'(8002);
			5776: out = 16'(696);
			5777: out = 16'(-8292);
			5778: out = 16'(-10125);
			5779: out = 16'(-4550);
			5780: out = 16'(7321);
			5781: out = 16'(13712);
			5782: out = 16'(9289);
			5783: out = 16'(-3705);
			5784: out = 16'(-11174);
			5785: out = 16'(-11942);
			5786: out = 16'(-5109);
			5787: out = 16'(4812);
			5788: out = 16'(11460);
			5789: out = 16'(1645);
			5790: out = 16'(-7717);
			5791: out = 16'(-5645);
			5792: out = 16'(2368);
			5793: out = 16'(9579);
			5794: out = 16'(4468);
			5795: out = 16'(-11400);
			5796: out = 16'(-10143);
			5797: out = 16'(1730);
			5798: out = 16'(7084);
			5799: out = 16'(5355);
			5800: out = 16'(577);
			5801: out = 16'(-116);
			5802: out = 16'(6144);
			5803: out = 16'(7323);
			5804: out = 16'(2089);
			5805: out = 16'(-4217);
			5806: out = 16'(-3488);
			5807: out = 16'(1192);
			5808: out = 16'(5790);
			5809: out = 16'(7850);
			5810: out = 16'(1424);
			5811: out = 16'(-5989);
			5812: out = 16'(-4760);
			5813: out = 16'(666);
			5814: out = 16'(-1960);
			5815: out = 16'(-8010);
			5816: out = 16'(-6136);
			5817: out = 16'(2301);
			5818: out = 16'(-2279);
			5819: out = 16'(-2730);
			5820: out = 16'(4955);
			5821: out = 16'(5015);
			5822: out = 16'(-3959);
			5823: out = 16'(-3154);
			5824: out = 16'(-2889);
			5825: out = 16'(-1507);
			5826: out = 16'(4775);
			5827: out = 16'(6504);
			5828: out = 16'(2823);
			5829: out = 16'(-7258);
			5830: out = 16'(-1708);
			5831: out = 16'(7615);
			5832: out = 16'(9366);
			5833: out = 16'(-5195);
			5834: out = 16'(-10550);
			5835: out = 16'(-5466);
			5836: out = 16'(1126);
			5837: out = 16'(12217);
			5838: out = 16'(9563);
			5839: out = 16'(490);
			5840: out = 16'(-470);
			5841: out = 16'(-490);
			5842: out = 16'(-3968);
			5843: out = 16'(-6310);
			5844: out = 16'(-1030);
			5845: out = 16'(584);
			5846: out = 16'(-692);
			5847: out = 16'(5911);
			5848: out = 16'(2569);
			5849: out = 16'(-853);
			5850: out = 16'(-2484);
			5851: out = 16'(-4866);
			5852: out = 16'(807);
			5853: out = 16'(5325);
			5854: out = 16'(4641);
			5855: out = 16'(-2361);
			5856: out = 16'(-1045);
			5857: out = 16'(8067);
			5858: out = 16'(6628);
			5859: out = 16'(-3150);
			5860: out = 16'(-5982);
			5861: out = 16'(-972);
			5862: out = 16'(-4220);
			5863: out = 16'(-3187);
			5864: out = 16'(-2531);
			5865: out = 16'(-5077);
			5866: out = 16'(-3486);
			5867: out = 16'(5497);
			5868: out = 16'(7904);
			5869: out = 16'(-1770);
			5870: out = 16'(-2471);
			5871: out = 16'(7535);
			5872: out = 16'(10418);
			5873: out = 16'(-400);
			5874: out = 16'(-7323);
			5875: out = 16'(-3238);
			5876: out = 16'(3507);
			5877: out = 16'(3508);
			5878: out = 16'(-889);
			5879: out = 16'(-6115);
			5880: out = 16'(-4847);
			5881: out = 16'(900);
			5882: out = 16'(2328);
			5883: out = 16'(-3329);
			5884: out = 16'(-3814);
			5885: out = 16'(2114);
			5886: out = 16'(8256);
			5887: out = 16'(4590);
			5888: out = 16'(-1155);
			5889: out = 16'(3586);
			5890: out = 16'(4075);
			5891: out = 16'(538);
			5892: out = 16'(725);
			5893: out = 16'(-2491);
			5894: out = 16'(-8333);
			5895: out = 16'(-8478);
			5896: out = 16'(-699);
			5897: out = 16'(6082);
			5898: out = 16'(1514);
			5899: out = 16'(-627);
			5900: out = 16'(8673);
			5901: out = 16'(7988);
			5902: out = 16'(-3542);
			5903: out = 16'(-8144);
			5904: out = 16'(-6179);
			5905: out = 16'(1575);
			5906: out = 16'(7433);
			5907: out = 16'(3331);
			5908: out = 16'(-6079);
			5909: out = 16'(-5374);
			5910: out = 16'(2586);
			5911: out = 16'(11136);
			5912: out = 16'(1956);
			5913: out = 16'(-5498);
			5914: out = 16'(-282);
			5915: out = 16'(3934);
			5916: out = 16'(5260);
			5917: out = 16'(2413);
			5918: out = 16'(-654);
			5919: out = 16'(-3458);
			5920: out = 16'(-5529);
			5921: out = 16'(-12342);
			5922: out = 16'(-8293);
			5923: out = 16'(5026);
			5924: out = 16'(10578);
			5925: out = 16'(5234);
			5926: out = 16'(3135);
			5927: out = 16'(-3298);
			5928: out = 16'(-629);
			5929: out = 16'(4155);
			5930: out = 16'(2796);
			5931: out = 16'(7916);
			5932: out = 16'(4681);
			5933: out = 16'(-318);
			5934: out = 16'(-374);
			5935: out = 16'(1086);
			5936: out = 16'(774);
			5937: out = 16'(-6239);
			5938: out = 16'(-10034);
			5939: out = 16'(-537);
			5940: out = 16'(1970);
			5941: out = 16'(326);
			5942: out = 16'(2623);
			5943: out = 16'(3620);
			5944: out = 16'(-1621);
			5945: out = 16'(-10393);
			5946: out = 16'(-12067);
			5947: out = 16'(2382);
			5948: out = 16'(14015);
			5949: out = 16'(10759);
			5950: out = 16'(-5522);
			5951: out = 16'(-4613);
			5952: out = 16'(1158);
			5953: out = 16'(6425);
			5954: out = 16'(4455);
			5955: out = 16'(493);
			5956: out = 16'(-1373);
			5957: out = 16'(-103);
			5958: out = 16'(2878);
			5959: out = 16'(1688);
			5960: out = 16'(950);
			5961: out = 16'(1522);
			5962: out = 16'(-122);
			5963: out = 16'(-6408);
			5964: out = 16'(-7512);
			5965: out = 16'(-7785);
			5966: out = 16'(-8500);
			5967: out = 16'(703);
			5968: out = 16'(9420);
			5969: out = 16'(3924);
			5970: out = 16'(1210);
			5971: out = 16'(-880);
			5972: out = 16'(1840);
			5973: out = 16'(4203);
			5974: out = 16'(4671);
			5975: out = 16'(7635);
			5976: out = 16'(1365);
			5977: out = 16'(-1914);
			5978: out = 16'(-1839);
			5979: out = 16'(-2649);
			5980: out = 16'(-4098);
			5981: out = 16'(-5076);
			5982: out = 16'(-5794);
			5983: out = 16'(539);
			5984: out = 16'(4732);
			5985: out = 16'(2045);
			5986: out = 16'(-1595);
			5987: out = 16'(-3270);
			5988: out = 16'(2768);
			5989: out = 16'(4118);
			5990: out = 16'(3849);
			5991: out = 16'(1232);
			5992: out = 16'(1455);
			5993: out = 16'(-840);
			5994: out = 16'(-2291);
			5995: out = 16'(-26);
			5996: out = 16'(-3762);
			5997: out = 16'(-6667);
			5998: out = 16'(1591);
			5999: out = 16'(7057);
			6000: out = 16'(-2745);
			6001: out = 16'(-8152);
			6002: out = 16'(-3057);
			6003: out = 16'(2113);
			6004: out = 16'(5447);
			6005: out = 16'(6553);
			6006: out = 16'(-5917);
			6007: out = 16'(-7219);
			6008: out = 16'(-681);
			6009: out = 16'(2000);
			6010: out = 16'(6489);
			6011: out = 16'(-1639);
			6012: out = 16'(-5624);
			6013: out = 16'(2291);
			6014: out = 16'(7682);
			6015: out = 16'(6100);
			6016: out = 16'(-6181);
			6017: out = 16'(-10125);
			6018: out = 16'(-3269);
			6019: out = 16'(4104);
			6020: out = 16'(8008);
			6021: out = 16'(7986);
			6022: out = 16'(3036);
			6023: out = 16'(-2271);
			6024: out = 16'(-3123);
			6025: out = 16'(-1051);
			6026: out = 16'(5549);
			6027: out = 16'(6212);
			6028: out = 16'(-2514);
			6029: out = 16'(-2478);
			6030: out = 16'(3925);
			6031: out = 16'(1981);
			6032: out = 16'(-2340);
			6033: out = 16'(-4653);
			6034: out = 16'(-3833);
			6035: out = 16'(-7321);
			6036: out = 16'(-1365);
			6037: out = 16'(5209);
			6038: out = 16'(3112);
			6039: out = 16'(-1459);
			6040: out = 16'(-1143);
			6041: out = 16'(-1760);
			6042: out = 16'(-1527);
			6043: out = 16'(-4946);
			6044: out = 16'(-5221);
			6045: out = 16'(-2954);
			6046: out = 16'(2395);
			6047: out = 16'(6045);
			6048: out = 16'(9505);
			6049: out = 16'(4624);
			6050: out = 16'(-2363);
			6051: out = 16'(-867);
			6052: out = 16'(-989);
			6053: out = 16'(3082);
			6054: out = 16'(6144);
			6055: out = 16'(1947);
			6056: out = 16'(-5702);
			6057: out = 16'(-6524);
			6058: out = 16'(-3953);
			6059: out = 16'(-1652);
			6060: out = 16'(-3570);
			6061: out = 16'(-6234);
			6062: out = 16'(822);
			6063: out = 16'(2651);
			6064: out = 16'(4165);
			6065: out = 16'(1193);
			6066: out = 16'(3271);
			6067: out = 16'(2920);
			6068: out = 16'(1675);
			6069: out = 16'(1758);
			6070: out = 16'(2034);
			6071: out = 16'(1890);
			6072: out = 16'(-210);
			6073: out = 16'(2132);
			6074: out = 16'(1384);
			6075: out = 16'(-6132);
			6076: out = 16'(-11308);
			6077: out = 16'(-4414);
			6078: out = 16'(-1070);
			6079: out = 16'(-2885);
			6080: out = 16'(187);
			6081: out = 16'(3022);
			6082: out = 16'(-3354);
			6083: out = 16'(-7096);
			6084: out = 16'(-2893);
			6085: out = 16'(3750);
			6086: out = 16'(5249);
			6087: out = 16'(2395);
			6088: out = 16'(-179);
			6089: out = 16'(565);
			6090: out = 16'(473);
			6091: out = 16'(4675);
			6092: out = 16'(1200);
			6093: out = 16'(-3921);
			6094: out = 16'(-627);
			6095: out = 16'(4232);
			6096: out = 16'(2371);
			6097: out = 16'(412);
			6098: out = 16'(-972);
			6099: out = 16'(-1271);
			6100: out = 16'(-10485);
			6101: out = 16'(-9907);
			6102: out = 16'(3862);
			6103: out = 16'(6983);
			6104: out = 16'(-1331);
			6105: out = 16'(-949);
			6106: out = 16'(1400);
			6107: out = 16'(779);
			6108: out = 16'(-1598);
			6109: out = 16'(-1630);
			6110: out = 16'(3947);
			6111: out = 16'(20);
			6112: out = 16'(-1635);
			6113: out = 16'(-504);
			6114: out = 16'(2850);
			6115: out = 16'(4610);
			6116: out = 16'(978);
			6117: out = 16'(-2340);
			6118: out = 16'(-787);
			6119: out = 16'(-4472);
			6120: out = 16'(-5140);
			6121: out = 16'(-2278);
			6122: out = 16'(-6460);
			6123: out = 16'(-3768);
			6124: out = 16'(6661);
			6125: out = 16'(10528);
			6126: out = 16'(-1242);
			6127: out = 16'(-10027);
			6128: out = 16'(-1628);
			6129: out = 16'(5300);
			6130: out = 16'(10950);
			6131: out = 16'(3892);
			6132: out = 16'(-2922);
			6133: out = 16'(-4313);
			6134: out = 16'(-3605);
			6135: out = 16'(-288);
			6136: out = 16'(5497);
			6137: out = 16'(5678);
			6138: out = 16'(-1258);
			6139: out = 16'(-9385);
			6140: out = 16'(-8614);
			6141: out = 16'(2651);
			6142: out = 16'(8032);
			6143: out = 16'(-1640);
			6144: out = 16'(-4590);
			6145: out = 16'(-32);
			6146: out = 16'(236);
			6147: out = 16'(1047);
			6148: out = 16'(1049);
			6149: out = 16'(5070);
			6150: out = 16'(2059);
			6151: out = 16'(-3668);
			6152: out = 16'(-4273);
			6153: out = 16'(159);
			6154: out = 16'(4171);
			6155: out = 16'(-5778);
			6156: out = 16'(-8174);
			6157: out = 16'(-1109);
			6158: out = 16'(1970);
			6159: out = 16'(6954);
			6160: out = 16'(3819);
			6161: out = 16'(-1847);
			6162: out = 16'(-2228);
			6163: out = 16'(2547);
			6164: out = 16'(3286);
			6165: out = 16'(-2263);
			6166: out = 16'(-7474);
			6167: out = 16'(-810);
			6168: out = 16'(1427);
			6169: out = 16'(-4414);
			6170: out = 16'(-2066);
			6171: out = 16'(6011);
			6172: out = 16'(3649);
			6173: out = 16'(-3619);
			6174: out = 16'(-340);
			6175: out = 16'(929);
			6176: out = 16'(-5133);
			6177: out = 16'(-2894);
			6178: out = 16'(2084);
			6179: out = 16'(-2584);
			6180: out = 16'(-3975);
			6181: out = 16'(1434);
			6182: out = 16'(4347);
			6183: out = 16'(6032);
			6184: out = 16'(4544);
			6185: out = 16'(216);
			6186: out = 16'(492);
			6187: out = 16'(1243);
			6188: out = 16'(-5042);
			6189: out = 16'(-6032);
			6190: out = 16'(-1127);
			6191: out = 16'(238);
			6192: out = 16'(4206);
			6193: out = 16'(-233);
			6194: out = 16'(-3642);
			6195: out = 16'(4704);
			6196: out = 16'(9193);
			6197: out = 16'(7392);
			6198: out = 16'(-3798);
			6199: out = 16'(-7035);
			6200: out = 16'(-4595);
			6201: out = 16'(-914);
			6202: out = 16'(5420);
			6203: out = 16'(3091);
			6204: out = 16'(754);
			6205: out = 16'(818);
			6206: out = 16'(-5223);
			6207: out = 16'(-5287);
			6208: out = 16'(2316);
			6209: out = 16'(4725);
			6210: out = 16'(630);
			6211: out = 16'(-6381);
			6212: out = 16'(-3630);
			6213: out = 16'(1800);
			6214: out = 16'(6687);
			6215: out = 16'(4229);
			6216: out = 16'(3607);
			6217: out = 16'(2317);
			6218: out = 16'(593);
			6219: out = 16'(3468);
			6220: out = 16'(1443);
			6221: out = 16'(-800);
			6222: out = 16'(-3752);
			6223: out = 16'(-6186);
			6224: out = 16'(-6678);
			6225: out = 16'(845);
			6226: out = 16'(6211);
			6227: out = 16'(725);
			6228: out = 16'(-682);
			6229: out = 16'(13);
			6230: out = 16'(962);
			6231: out = 16'(641);
			6232: out = 16'(237);
			6233: out = 16'(1111);
			6234: out = 16'(3443);
			6235: out = 16'(821);
			6236: out = 16'(-2095);
			6237: out = 16'(-5265);
			6238: out = 16'(-5731);
			6239: out = 16'(-6734);
			6240: out = 16'(-3321);
			6241: out = 16'(-1028);
			6242: out = 16'(3113);
			6243: out = 16'(522);
			6244: out = 16'(-1744);
			6245: out = 16'(2863);
			6246: out = 16'(6525);
			6247: out = 16'(9569);
			6248: out = 16'(3452);
			6249: out = 16'(-5294);
			6250: out = 16'(-9668);
			6251: out = 16'(-6795);
			6252: out = 16'(-2503);
			6253: out = 16'(-2261);
			6254: out = 16'(-2738);
			6255: out = 16'(514);
			6256: out = 16'(694);
			6257: out = 16'(3888);
			6258: out = 16'(6647);
			6259: out = 16'(8316);
			6260: out = 16'(7239);
			6261: out = 16'(-126);
			6262: out = 16'(-6173);
			6263: out = 16'(-8377);
			6264: out = 16'(-8698);
			6265: out = 16'(-5182);
			6266: out = 16'(561);
			6267: out = 16'(3876);
			6268: out = 16'(2944);
			6269: out = 16'(3818);
			6270: out = 16'(10322);
			6271: out = 16'(5185);
			6272: out = 16'(-1085);
			6273: out = 16'(-5809);
			6274: out = 16'(166);
			6275: out = 16'(2596);
			6276: out = 16'(-1620);
			6277: out = 16'(947);
			6278: out = 16'(397);
			6279: out = 16'(-3244);
			6280: out = 16'(-2568);
			6281: out = 16'(-8032);
			6282: out = 16'(-5242);
			6283: out = 16'(4672);
			6284: out = 16'(7782);
			6285: out = 16'(4183);
			6286: out = 16'(832);
			6287: out = 16'(5634);
			6288: out = 16'(4978);
			6289: out = 16'(-1522);
			6290: out = 16'(-8536);
			6291: out = 16'(-4882);
			6292: out = 16'(847);
			6293: out = 16'(2454);
			6294: out = 16'(1505);
			6295: out = 16'(1097);
			6296: out = 16'(4454);
			6297: out = 16'(2974);
			6298: out = 16'(-890);
			6299: out = 16'(-1665);
			6300: out = 16'(-1583);
			6301: out = 16'(1155);
			6302: out = 16'(587);
			6303: out = 16'(-1841);
			6304: out = 16'(-6343);
			6305: out = 16'(-3079);
			6306: out = 16'(4482);
			6307: out = 16'(1572);
			6308: out = 16'(1723);
			6309: out = 16'(3565);
			6310: out = 16'(4485);
			6311: out = 16'(4398);
			6312: out = 16'(-2831);
			6313: out = 16'(-7969);
			6314: out = 16'(-3166);
			6315: out = 16'(3599);
			6316: out = 16'(5234);
			6317: out = 16'(2167);
			6318: out = 16'(419);
			6319: out = 16'(1322);
			6320: out = 16'(3413);
			6321: out = 16'(1284);
			6322: out = 16'(-3250);
			6323: out = 16'(-3447);
			6324: out = 16'(1456);
			6325: out = 16'(8590);
			6326: out = 16'(5103);
			6327: out = 16'(-1806);
			6328: out = 16'(-5174);
			6329: out = 16'(-1347);
			6330: out = 16'(6656);
			6331: out = 16'(7167);
			6332: out = 16'(-1919);
			6333: out = 16'(-6658);
			6334: out = 16'(-2748);
			6335: out = 16'(-3081);
			6336: out = 16'(3052);
			6337: out = 16'(6788);
			6338: out = 16'(1180);
			6339: out = 16'(-9045);
			6340: out = 16'(-8233);
			6341: out = 16'(-5965);
			6342: out = 16'(-4349);
			6343: out = 16'(3137);
			6344: out = 16'(2488);
			6345: out = 16'(-3471);
			6346: out = 16'(1523);
			6347: out = 16'(-604);
			6348: out = 16'(2663);
			6349: out = 16'(3492);
			6350: out = 16'(2694);
			6351: out = 16'(1721);
			6352: out = 16'(1349);
			6353: out = 16'(5601);
			6354: out = 16'(2685);
			6355: out = 16'(-5547);
			6356: out = 16'(-5545);
			6357: out = 16'(-1603);
			6358: out = 16'(160);
			6359: out = 16'(5803);
			6360: out = 16'(6032);
			6361: out = 16'(-632);
			6362: out = 16'(-6587);
			6363: out = 16'(-5100);
			6364: out = 16'(-702);
			6365: out = 16'(-3046);
			6366: out = 16'(-1216);
			6367: out = 16'(2160);
			6368: out = 16'(1818);
			6369: out = 16'(1920);
			6370: out = 16'(5387);
			6371: out = 16'(11744);
			6372: out = 16'(5921);
			6373: out = 16'(-6909);
			6374: out = 16'(-11574);
			6375: out = 16'(-5742);
			6376: out = 16'(686);
			6377: out = 16'(2819);
			6378: out = 16'(-2163);
			6379: out = 16'(-4002);
			6380: out = 16'(193);
			6381: out = 16'(3982);
			6382: out = 16'(6049);
			6383: out = 16'(2997);
			6384: out = 16'(-2970);
			6385: out = 16'(-433);
			6386: out = 16'(-169);
			6387: out = 16'(-978);
			6388: out = 16'(1890);
			6389: out = 16'(-2839);
			6390: out = 16'(-6822);
			6391: out = 16'(-2688);
			6392: out = 16'(3332);
			6393: out = 16'(4342);
			6394: out = 16'(2569);
			6395: out = 16'(3473);
			6396: out = 16'(4721);
			6397: out = 16'(4977);
			6398: out = 16'(2054);
			6399: out = 16'(-2418);
			6400: out = 16'(-4302);
			6401: out = 16'(-2666);
			6402: out = 16'(-1888);
			6403: out = 16'(-7718);
			6404: out = 16'(-4341);
			6405: out = 16'(4046);
			6406: out = 16'(4554);
			6407: out = 16'(3395);
			6408: out = 16'(1376);
			6409: out = 16'(776);
			6410: out = 16'(2905);
			6411: out = 16'(3239);
			6412: out = 16'(-4942);
			6413: out = 16'(-13135);
			6414: out = 16'(-10191);
			6415: out = 16'(1417);
			6416: out = 16'(9785);
			6417: out = 16'(6172);
			6418: out = 16'(373);
			6419: out = 16'(3165);
			6420: out = 16'(5483);
			6421: out = 16'(-123);
			6422: out = 16'(-7831);
			6423: out = 16'(-8066);
			6424: out = 16'(-989);
			6425: out = 16'(8286);
			6426: out = 16'(7311);
			6427: out = 16'(-4575);
			6428: out = 16'(-6863);
			6429: out = 16'(2375);
			6430: out = 16'(8980);
			6431: out = 16'(5127);
			6432: out = 16'(1287);
			6433: out = 16'(-1001);
			6434: out = 16'(-2819);
			6435: out = 16'(-3072);
			6436: out = 16'(840);
			6437: out = 16'(4278);
			6438: out = 16'(-3792);
			6439: out = 16'(-11756);
			6440: out = 16'(-4048);
			6441: out = 16'(2612);
			6442: out = 16'(5279);
			6443: out = 16'(2304);
			6444: out = 16'(-1432);
			6445: out = 16'(-2813);
			6446: out = 16'(40);
			6447: out = 16'(2631);
			6448: out = 16'(5782);
			6449: out = 16'(1889);
			6450: out = 16'(-3761);
			6451: out = 16'(-5813);
			6452: out = 16'(-2372);
			6453: out = 16'(3314);
			6454: out = 16'(7121);
			6455: out = 16'(-3973);
			6456: out = 16'(-6639);
			6457: out = 16'(-678);
			6458: out = 16'(4215);
			6459: out = 16'(5940);
			6460: out = 16'(1912);
			6461: out = 16'(-2434);
			6462: out = 16'(-6571);
			6463: out = 16'(-8035);
			6464: out = 16'(-9104);
			6465: out = 16'(834);
			6466: out = 16'(4409);
			6467: out = 16'(1377);
			6468: out = 16'(4883);
			6469: out = 16'(1872);
			6470: out = 16'(-1081);
			6471: out = 16'(-294);
			6472: out = 16'(466);
			6473: out = 16'(1355);
			6474: out = 16'(702);
			6475: out = 16'(4258);
			6476: out = 16'(4475);
			6477: out = 16'(122);
			6478: out = 16'(-5304);
			6479: out = 16'(-1833);
			6480: out = 16'(3370);
			6481: out = 16'(2221);
			6482: out = 16'(31);
			6483: out = 16'(1633);
			6484: out = 16'(4121);
			6485: out = 16'(1334);
			6486: out = 16'(-7759);
			6487: out = 16'(-10247);
			6488: out = 16'(-1220);
			6489: out = 16'(3586);
			6490: out = 16'(-4325);
			6491: out = 16'(-3765);
			6492: out = 16'(3679);
			6493: out = 16'(3198);
			6494: out = 16'(-3067);
			6495: out = 16'(-2945);
			6496: out = 16'(617);
			6497: out = 16'(3250);
			6498: out = 16'(6900);
			6499: out = 16'(-663);
			6500: out = 16'(-4431);
			6501: out = 16'(-4347);
			6502: out = 16'(-1036);
			6503: out = 16'(2329);
			6504: out = 16'(-356);
			6505: out = 16'(1555);
			6506: out = 16'(3707);
			6507: out = 16'(1531);
			6508: out = 16'(-6889);
			6509: out = 16'(-9904);
			6510: out = 16'(-3274);
			6511: out = 16'(5084);
			6512: out = 16'(6305);
			6513: out = 16'(545);
			6514: out = 16'(1555);
			6515: out = 16'(2839);
			6516: out = 16'(447);
			6517: out = 16'(-1915);
			6518: out = 16'(-3064);
			6519: out = 16'(535);
			6520: out = 16'(4188);
			6521: out = 16'(4093);
			6522: out = 16'(550);
			6523: out = 16'(462);
			6524: out = 16'(324);
			6525: out = 16'(1950);
			6526: out = 16'(-1043);
			6527: out = 16'(-5562);
			6528: out = 16'(-5699);
			6529: out = 16'(-1130);
			6530: out = 16'(2327);
			6531: out = 16'(195);
			6532: out = 16'(-5647);
			6533: out = 16'(-4188);
			6534: out = 16'(-3552);
			6535: out = 16'(-1119);
			6536: out = 16'(981);
			6537: out = 16'(205);
			6538: out = 16'(-3169);
			6539: out = 16'(-2081);
			6540: out = 16'(267);
			6541: out = 16'(983);
			6542: out = 16'(1630);
			6543: out = 16'(-768);
			6544: out = 16'(1748);
			6545: out = 16'(5068);
			6546: out = 16'(5313);
			6547: out = 16'(1532);
			6548: out = 16'(-3041);
			6549: out = 16'(-4538);
			6550: out = 16'(-2147);
			6551: out = 16'(-4052);
			6552: out = 16'(-5134);
			6553: out = 16'(-1758);
			6554: out = 16'(1685);
			6555: out = 16'(8117);
			6556: out = 16'(4851);
			6557: out = 16'(2413);
			6558: out = 16'(-3408);
			6559: out = 16'(-2788);
			6560: out = 16'(811);
			6561: out = 16'(-154);
			6562: out = 16'(4223);
			6563: out = 16'(3060);
			6564: out = 16'(1915);
			6565: out = 16'(1194);
			6566: out = 16'(1396);
			6567: out = 16'(-5296);
			6568: out = 16'(-6374);
			6569: out = 16'(-2167);
			6570: out = 16'(-128);
			6571: out = 16'(-2635);
			6572: out = 16'(129);
			6573: out = 16'(-3065);
			6574: out = 16'(-6541);
			6575: out = 16'(-2097);
			6576: out = 16'(1251);
			6577: out = 16'(3696);
			6578: out = 16'(2617);
			6579: out = 16'(-1458);
			6580: out = 16'(-5720);
			6581: out = 16'(-5430);
			6582: out = 16'(2574);
			6583: out = 16'(7763);
			6584: out = 16'(7870);
			6585: out = 16'(-3380);
			6586: out = 16'(-11542);
			6587: out = 16'(-4623);
			6588: out = 16'(5936);
			6589: out = 16'(12628);
			6590: out = 16'(6127);
			6591: out = 16'(-2989);
			6592: out = 16'(-3949);
			6593: out = 16'(1346);
			6594: out = 16'(1061);
			6595: out = 16'(-6820);
			6596: out = 16'(-5680);
			6597: out = 16'(-3);
			6598: out = 16'(1440);
			6599: out = 16'(7135);
			6600: out = 16'(2239);
			6601: out = 16'(2473);
			6602: out = 16'(7023);
			6603: out = 16'(4785);
			6604: out = 16'(-2436);
			6605: out = 16'(-8560);
			6606: out = 16'(-6837);
			6607: out = 16'(-2508);
			6608: out = 16'(5038);
			6609: out = 16'(8888);
			6610: out = 16'(1845);
			6611: out = 16'(557);
			6612: out = 16'(839);
			6613: out = 16'(-155);
			6614: out = 16'(2630);
			6615: out = 16'(-1441);
			6616: out = 16'(-550);
			6617: out = 16'(5103);
			6618: out = 16'(6215);
			6619: out = 16'(-4289);
			6620: out = 16'(-11524);
			6621: out = 16'(-10893);
			6622: out = 16'(-1663);
			6623: out = 16'(6796);
			6624: out = 16'(7693);
			6625: out = 16'(-1946);
			6626: out = 16'(-2792);
			6627: out = 16'(405);
			6628: out = 16'(684);
			6629: out = 16'(7502);
			6630: out = 16'(6522);
			6631: out = 16'(-600);
			6632: out = 16'(-1796);
			6633: out = 16'(1989);
			6634: out = 16'(-1219);
			6635: out = 16'(-11601);
			6636: out = 16'(-10781);
			6637: out = 16'(107);
			6638: out = 16'(1283);
			6639: out = 16'(5654);
			6640: out = 16'(6813);
			6641: out = 16'(3969);
			6642: out = 16'(-265);
			6643: out = 16'(-2591);
			6644: out = 16'(241);
			6645: out = 16'(2399);
			6646: out = 16'(348);
			6647: out = 16'(-3461);
			6648: out = 16'(-2235);
			6649: out = 16'(-2631);
			6650: out = 16'(-2938);
			6651: out = 16'(3221);
			6652: out = 16'(4812);
			6653: out = 16'(504);
			6654: out = 16'(2072);
			6655: out = 16'(2270);
			6656: out = 16'(1061);
			6657: out = 16'(766);
			6658: out = 16'(-1162);
			6659: out = 16'(-5103);
			6660: out = 16'(-2284);
			6661: out = 16'(1876);
			6662: out = 16'(6622);
			6663: out = 16'(5302);
			6664: out = 16'(5309);
			6665: out = 16'(4895);
			6666: out = 16'(2663);
			6667: out = 16'(809);
			6668: out = 16'(-2291);
			6669: out = 16'(-4246);
			6670: out = 16'(-5514);
			6671: out = 16'(-1584);
			6672: out = 16'(865);
			6673: out = 16'(-631);
			6674: out = 16'(-6349);
			6675: out = 16'(-4856);
			6676: out = 16'(-172);
			6677: out = 16'(7058);
			6678: out = 16'(8128);
			6679: out = 16'(1368);
			6680: out = 16'(-2098);
			6681: out = 16'(-4460);
			6682: out = 16'(-119);
			6683: out = 16'(-1599);
			6684: out = 16'(-1220);
			6685: out = 16'(5842);
			6686: out = 16'(5004);
			6687: out = 16'(-3178);
			6688: out = 16'(-9107);
			6689: out = 16'(-10154);
			6690: out = 16'(2560);
			6691: out = 16'(10239);
			6692: out = 16'(3388);
			6693: out = 16'(-2251);
			6694: out = 16'(-227);
			6695: out = 16'(3254);
			6696: out = 16'(291);
			6697: out = 16'(-5901);
			6698: out = 16'(-3479);
			6699: out = 16'(5685);
			6700: out = 16'(8106);
			6701: out = 16'(4291);
			6702: out = 16'(1601);
			6703: out = 16'(-632);
			6704: out = 16'(875);
			6705: out = 16'(-1473);
			6706: out = 16'(-3589);
			6707: out = 16'(2700);
			6708: out = 16'(4358);
			6709: out = 16'(-4824);
			6710: out = 16'(-10079);
			6711: out = 16'(-4711);
			6712: out = 16'(2573);
			6713: out = 16'(1960);
			6714: out = 16'(1659);
			6715: out = 16'(3203);
			6716: out = 16'(-1288);
			6717: out = 16'(-4143);
			6718: out = 16'(-1475);
			6719: out = 16'(4428);
			6720: out = 16'(2951);
			6721: out = 16'(-4197);
			6722: out = 16'(-7998);
			6723: out = 16'(-2027);
			6724: out = 16'(8376);
			6725: out = 16'(4956);
			6726: out = 16'(-335);
			6727: out = 16'(1134);
			6728: out = 16'(1666);
			6729: out = 16'(904);
			6730: out = 16'(630);
			6731: out = 16'(2962);
			6732: out = 16'(5504);
			6733: out = 16'(-955);
			6734: out = 16'(-7483);
			6735: out = 16'(-6654);
			6736: out = 16'(-3651);
			6737: out = 16'(2892);
			6738: out = 16'(1923);
			6739: out = 16'(-2781);
			6740: out = 16'(1434);
			6741: out = 16'(5630);
			6742: out = 16'(1224);
			6743: out = 16'(-8743);
			6744: out = 16'(-10966);
			6745: out = 16'(-1759);
			6746: out = 16'(5910);
			6747: out = 16'(5670);
			6748: out = 16'(4008);
			6749: out = 16'(4012);
			6750: out = 16'(1627);
			6751: out = 16'(1402);
			6752: out = 16'(-1206);
			6753: out = 16'(-5703);
			6754: out = 16'(-8032);
			6755: out = 16'(591);
			6756: out = 16'(6383);
			6757: out = 16'(559);
			6758: out = 16'(-247);
			6759: out = 16'(2845);
			6760: out = 16'(5445);
			6761: out = 16'(1126);
			6762: out = 16'(-614);
			6763: out = 16'(1596);
			6764: out = 16'(3854);
			6765: out = 16'(2004);
			6766: out = 16'(-2236);
			6767: out = 16'(-864);
			6768: out = 16'(591);
			6769: out = 16'(83);
			6770: out = 16'(-1503);
			6771: out = 16'(-2521);
			6772: out = 16'(-4253);
			6773: out = 16'(-2368);
			6774: out = 16'(-359);
			6775: out = 16'(-996);
			6776: out = 16'(-1291);
			6777: out = 16'(-2624);
			6778: out = 16'(-7296);
			6779: out = 16'(-4284);
			6780: out = 16'(6455);
			6781: out = 16'(10783);
			6782: out = 16'(-2016);
			6783: out = 16'(-13530);
			6784: out = 16'(-8926);
			6785: out = 16'(1110);
			6786: out = 16'(9566);
			6787: out = 16'(6804);
			6788: out = 16'(-3059);
			6789: out = 16'(-4105);
			6790: out = 16'(2417);
			6791: out = 16'(2561);
			6792: out = 16'(-1048);
			6793: out = 16'(-6635);
			6794: out = 16'(-3779);
			6795: out = 16'(4565);
			6796: out = 16'(2631);
			6797: out = 16'(2703);
			6798: out = 16'(3032);
			6799: out = 16'(3841);
			6800: out = 16'(2701);
			6801: out = 16'(-1072);
			6802: out = 16'(-8769);
			6803: out = 16'(-6830);
			6804: out = 16'(-4120);
			6805: out = 16'(-3894);
			6806: out = 16'(6003);
			6807: out = 16'(8996);
			6808: out = 16'(-856);
			6809: out = 16'(-2638);
			6810: out = 16'(-2518);
			6811: out = 16'(1077);
			6812: out = 16'(2891);
			6813: out = 16'(4032);
			6814: out = 16'(4473);
			6815: out = 16'(110);
			6816: out = 16'(2992);
			6817: out = 16'(3803);
			6818: out = 16'(-519);
			6819: out = 16'(-3824);
			6820: out = 16'(-2373);
			6821: out = 16'(-2778);
			6822: out = 16'(887);
			6823: out = 16'(2627);
			6824: out = 16'(359);
			6825: out = 16'(-1320);
			6826: out = 16'(696);
			6827: out = 16'(5354);
			6828: out = 16'(3877);
			6829: out = 16'(-3399);
			6830: out = 16'(-3415);
			6831: out = 16'(-1647);
			6832: out = 16'(-3842);
			6833: out = 16'(-2332);
			6834: out = 16'(3238);
			6835: out = 16'(-969);
			6836: out = 16'(-7916);
			6837: out = 16'(-4547);
			6838: out = 16'(846);
			6839: out = 16'(3945);
			6840: out = 16'(2471);
			6841: out = 16'(-5303);
			6842: out = 16'(-5379);
			6843: out = 16'(-1693);
			6844: out = 16'(8654);
			6845: out = 16'(9226);
			6846: out = 16'(-236);
			6847: out = 16'(-4123);
			6848: out = 16'(-2359);
			6849: out = 16'(-794);
			6850: out = 16'(-891);
			6851: out = 16'(-2496);
			6852: out = 16'(-3144);
			6853: out = 16'(4427);
			6854: out = 16'(7668);
			6855: out = 16'(-1780);
			6856: out = 16'(-9715);
			6857: out = 16'(-7067);
			6858: out = 16'(2031);
			6859: out = 16'(4642);
			6860: out = 16'(7676);
			6861: out = 16'(4692);
			6862: out = 16'(-2290);
			6863: out = 16'(-7461);
			6864: out = 16'(-7770);
			6865: out = 16'(390);
			6866: out = 16'(4677);
			6867: out = 16'(2574);
			6868: out = 16'(2140);
			6869: out = 16'(3754);
			6870: out = 16'(2778);
			6871: out = 16'(3513);
			6872: out = 16'(1198);
			6873: out = 16'(-1031);
			6874: out = 16'(-7648);
			6875: out = 16'(-6707);
			6876: out = 16'(-2450);
			6877: out = 16'(1108);
			6878: out = 16'(1700);
			6879: out = 16'(-2827);
			6880: out = 16'(-1861);
			6881: out = 16'(4867);
			6882: out = 16'(4193);
			6883: out = 16'(-3512);
			6884: out = 16'(-8855);
			6885: out = 16'(-7146);
			6886: out = 16'(965);
			6887: out = 16'(11009);
			6888: out = 16'(8436);
			6889: out = 16'(-931);
			6890: out = 16'(-4996);
			6891: out = 16'(-4822);
			6892: out = 16'(-1785);
			6893: out = 16'(3431);
			6894: out = 16'(5930);
			6895: out = 16'(257);
			6896: out = 16'(253);
			6897: out = 16'(-197);
			6898: out = 16'(-1592);
			6899: out = 16'(1015);
			6900: out = 16'(-2884);
			6901: out = 16'(1242);
			6902: out = 16'(5666);
			6903: out = 16'(63);
			6904: out = 16'(-659);
			6905: out = 16'(814);
			6906: out = 16'(-1100);
			6907: out = 16'(-4592);
			6908: out = 16'(-6465);
			6909: out = 16'(954);
			6910: out = 16'(4064);
			6911: out = 16'(1467);
			6912: out = 16'(-344);
			6913: out = 16'(-167);
			6914: out = 16'(-139);
			6915: out = 16'(-5569);
			6916: out = 16'(-3899);
			6917: out = 16'(2520);
			6918: out = 16'(4164);
			6919: out = 16'(4496);
			6920: out = 16'(4131);
			6921: out = 16'(1825);
			6922: out = 16'(-4570);
			6923: out = 16'(-7605);
			6924: out = 16'(-974);
			6925: out = 16'(2146);
			6926: out = 16'(4173);
			6927: out = 16'(3357);
			6928: out = 16'(-2097);
			6929: out = 16'(-5787);
			6930: out = 16'(-4022);
			6931: out = 16'(3436);
			6932: out = 16'(1618);
			6933: out = 16'(-3230);
			6934: out = 16'(-3);
			6935: out = 16'(1055);
			6936: out = 16'(3164);
			6937: out = 16'(4866);
			6938: out = 16'(3011);
			6939: out = 16'(3912);
			6940: out = 16'(-462);
			6941: out = 16'(-3501);
			6942: out = 16'(-2560);
			6943: out = 16'(-1658);
			6944: out = 16'(2318);
			6945: out = 16'(1988);
			6946: out = 16'(-2122);
			6947: out = 16'(-2889);
			6948: out = 16'(-1358);
			6949: out = 16'(-466);
			6950: out = 16'(2560);
			6951: out = 16'(2432);
			6952: out = 16'(1079);
			6953: out = 16'(1495);
			6954: out = 16'(-3919);
			6955: out = 16'(-7339);
			6956: out = 16'(-1066);
			6957: out = 16'(3458);
			6958: out = 16'(-236);
			6959: out = 16'(1864);
			6960: out = 16'(3188);
			6961: out = 16'(1101);
			6962: out = 16'(45);
			6963: out = 16'(-1398);
			6964: out = 16'(-573);
			6965: out = 16'(-174);
			6966: out = 16'(4561);
			6967: out = 16'(6661);
			6968: out = 16'(-1581);
			6969: out = 16'(-9334);
			6970: out = 16'(-6150);
			6971: out = 16'(591);
			6972: out = 16'(4805);
			6973: out = 16'(1824);
			6974: out = 16'(3852);
			6975: out = 16'(1371);
			6976: out = 16'(-4800);
			6977: out = 16'(-407);
			6978: out = 16'(6818);
			6979: out = 16'(4468);
			6980: out = 16'(-6504);
			6981: out = 16'(-10202);
			6982: out = 16'(-4774);
			6983: out = 16'(2459);
			6984: out = 16'(9968);
			6985: out = 16'(2046);
			6986: out = 16'(-6781);
			6987: out = 16'(-726);
			6988: out = 16'(6310);
			6989: out = 16'(7603);
			6990: out = 16'(2244);
			6991: out = 16'(-2399);
			6992: out = 16'(-337);
			6993: out = 16'(569);
			6994: out = 16'(-508);
			6995: out = 16'(-978);
			6996: out = 16'(853);
			6997: out = 16'(5233);
			6998: out = 16'(3817);
			6999: out = 16'(-6320);
			7000: out = 16'(-7688);
			7001: out = 16'(-1119);
			7002: out = 16'(3114);
			7003: out = 16'(1210);
			7004: out = 16'(2006);
			7005: out = 16'(4067);
			7006: out = 16'(-842);
			7007: out = 16'(-4146);
			7008: out = 16'(-472);
			7009: out = 16'(5290);
			7010: out = 16'(6068);
			7011: out = 16'(-3841);
			7012: out = 16'(-6182);
			7013: out = 16'(-2467);
			7014: out = 16'(-1888);
			7015: out = 16'(1363);
			7016: out = 16'(1871);
			7017: out = 16'(-2544);
			7018: out = 16'(-5681);
			7019: out = 16'(214);
			7020: out = 16'(4399);
			7021: out = 16'(3062);
			7022: out = 16'(2670);
			7023: out = 16'(1686);
			7024: out = 16'(-1488);
			7025: out = 16'(-203);
			7026: out = 16'(-810);
			7027: out = 16'(-864);
			7028: out = 16'(2848);
			7029: out = 16'(2954);
			7030: out = 16'(354);
			7031: out = 16'(-1737);
			7032: out = 16'(-1985);
			7033: out = 16'(638);
			7034: out = 16'(469);
			7035: out = 16'(-3723);
			7036: out = 16'(-2201);
			7037: out = 16'(821);
			7038: out = 16'(5660);
			7039: out = 16'(897);
			7040: out = 16'(-784);
			7041: out = 16'(3407);
			7042: out = 16'(1775);
			7043: out = 16'(-3377);
			7044: out = 16'(-583);
			7045: out = 16'(2219);
			7046: out = 16'(-272);
			7047: out = 16'(-5508);
			7048: out = 16'(-4230);
			7049: out = 16'(-2785);
			7050: out = 16'(-2330);
			7051: out = 16'(1457);
			7052: out = 16'(1031);
			7053: out = 16'(-304);
			7054: out = 16'(-37);
			7055: out = 16'(1544);
			7056: out = 16'(444);
			7057: out = 16'(-1851);
			7058: out = 16'(-368);
			7059: out = 16'(1879);
			7060: out = 16'(4106);
			7061: out = 16'(1420);
			7062: out = 16'(-2399);
			7063: out = 16'(92);
			7064: out = 16'(5852);
			7065: out = 16'(3701);
			7066: out = 16'(-2566);
			7067: out = 16'(517);
			7068: out = 16'(863);
			7069: out = 16'(-1806);
			7070: out = 16'(-3948);
			7071: out = 16'(-5010);
			7072: out = 16'(1149);
			7073: out = 16'(3242);
			7074: out = 16'(-2164);
			7075: out = 16'(292);
			7076: out = 16'(1395);
			7077: out = 16'(2795);
			7078: out = 16'(4851);
			7079: out = 16'(1959);
			7080: out = 16'(-1801);
			7081: out = 16'(-7301);
			7082: out = 16'(-4768);
			7083: out = 16'(-386);
			7084: out = 16'(4241);
			7085: out = 16'(3531);
			7086: out = 16'(1856);
			7087: out = 16'(3901);
			7088: out = 16'(-88);
			7089: out = 16'(-6295);
			7090: out = 16'(-7349);
			7091: out = 16'(-1807);
			7092: out = 16'(2823);
			7093: out = 16'(3587);
			7094: out = 16'(5020);
			7095: out = 16'(4898);
			7096: out = 16'(-1037);
			7097: out = 16'(-5861);
			7098: out = 16'(-4087);
			7099: out = 16'(-1245);
			7100: out = 16'(-1526);
			7101: out = 16'(-1062);
			7102: out = 16'(3620);
			7103: out = 16'(4920);
			7104: out = 16'(-2134);
			7105: out = 16'(-3106);
			7106: out = 16'(-42);
			7107: out = 16'(1004);
			7108: out = 16'(1379);
			7109: out = 16'(1119);
			7110: out = 16'(-116);
			7111: out = 16'(-2477);
			7112: out = 16'(-4034);
			7113: out = 16'(-934);
			7114: out = 16'(1282);
			7115: out = 16'(-498);
			7116: out = 16'(2212);
			7117: out = 16'(6872);
			7118: out = 16'(2916);
			7119: out = 16'(-4122);
			7120: out = 16'(-7904);
			7121: out = 16'(-1030);
			7122: out = 16'(6932);
			7123: out = 16'(5896);
			7124: out = 16'(765);
			7125: out = 16'(-1501);
			7126: out = 16'(-1623);
			7127: out = 16'(-4112);
			7128: out = 16'(-3482);
			7129: out = 16'(2961);
			7130: out = 16'(6914);
			7131: out = 16'(-1430);
			7132: out = 16'(-10114);
			7133: out = 16'(-5048);
			7134: out = 16'(2461);
			7135: out = 16'(5587);
			7136: out = 16'(2412);
			7137: out = 16'(-4887);
			7138: out = 16'(-7162);
			7139: out = 16'(-145);
			7140: out = 16'(7762);
			7141: out = 16'(6818);
			7142: out = 16'(-557);
			7143: out = 16'(-3536);
			7144: out = 16'(1680);
			7145: out = 16'(3549);
			7146: out = 16'(4302);
			7147: out = 16'(2418);
			7148: out = 16'(1258);
			7149: out = 16'(390);
			7150: out = 16'(-870);
			7151: out = 16'(-2063);
			7152: out = 16'(-2241);
			7153: out = 16'(-1501);
			7154: out = 16'(-3517);
			7155: out = 16'(-1435);
			7156: out = 16'(414);
			7157: out = 16'(1844);
			7158: out = 16'(-1748);
			7159: out = 16'(-5947);
			7160: out = 16'(-5557);
			7161: out = 16'(142);
			7162: out = 16'(6162);
			7163: out = 16'(3416);
			7164: out = 16'(79);
			7165: out = 16'(-1147);
			7166: out = 16'(1240);
			7167: out = 16'(4092);
			7168: out = 16'(329);
			7169: out = 16'(116);
			7170: out = 16'(3460);
			7171: out = 16'(4298);
			7172: out = 16'(-4165);
			7173: out = 16'(-10627);
			7174: out = 16'(-4288);
			7175: out = 16'(3518);
			7176: out = 16'(1861);
			7177: out = 16'(-5614);
			7178: out = 16'(-3857);
			7179: out = 16'(1084);
			7180: out = 16'(3504);
			7181: out = 16'(6739);
			7182: out = 16'(3215);
			7183: out = 16'(-2450);
			7184: out = 16'(-6513);
			7185: out = 16'(-2411);
			7186: out = 16'(5404);
			7187: out = 16'(6722);
			7188: out = 16'(632);
			7189: out = 16'(-6050);
			7190: out = 16'(-3337);
			7191: out = 16'(5265);
			7192: out = 16'(4831);
			7193: out = 16'(106);
			7194: out = 16'(-4429);
			7195: out = 16'(-2244);
			7196: out = 16'(538);
			7197: out = 16'(-2662);
			7198: out = 16'(42);
			7199: out = 16'(3978);
			7200: out = 16'(3357);
			7201: out = 16'(-3124);
			7202: out = 16'(-4830);
			7203: out = 16'(-2186);
			7204: out = 16'(1006);
			7205: out = 16'(328);
			7206: out = 16'(-1946);
			7207: out = 16'(-89);
			7208: out = 16'(1944);
			7209: out = 16'(-2412);
			7210: out = 16'(-3305);
			7211: out = 16'(-1628);
			7212: out = 16'(3377);
			7213: out = 16'(6988);
			7214: out = 16'(2424);
			7215: out = 16'(-3069);
			7216: out = 16'(-5732);
			7217: out = 16'(594);
			7218: out = 16'(2065);
			7219: out = 16'(-228);
			7220: out = 16'(-1472);
			7221: out = 16'(2672);
			7222: out = 16'(6669);
			7223: out = 16'(1862);
			7224: out = 16'(925);
			7225: out = 16'(911);
			7226: out = 16'(883);
			7227: out = 16'(-237);
			7228: out = 16'(-2768);
			7229: out = 16'(-934);
			7230: out = 16'(3076);
			7231: out = 16'(2503);
			7232: out = 16'(-575);
			7233: out = 16'(1281);
			7234: out = 16'(3452);
			7235: out = 16'(-518);
			7236: out = 16'(-6971);
			7237: out = 16'(-6057);
			7238: out = 16'(-2267);
			7239: out = 16'(-1908);
			7240: out = 16'(1033);
			7241: out = 16'(716);
			7242: out = 16'(-4477);
			7243: out = 16'(-5539);
			7244: out = 16'(-1553);
			7245: out = 16'(2615);
			7246: out = 16'(1977);
			7247: out = 16'(1363);
			7248: out = 16'(-3692);
			7249: out = 16'(-6247);
			7250: out = 16'(-4334);
			7251: out = 16'(-118);
			7252: out = 16'(3086);
			7253: out = 16'(55);
			7254: out = 16'(753);
			7255: out = 16'(1308);
			7256: out = 16'(-561);
			7257: out = 16'(418);
			7258: out = 16'(1975);
			7259: out = 16'(334);
			7260: out = 16'(820);
			7261: out = 16'(-2491);
			7262: out = 16'(-2214);
			7263: out = 16'(-169);
			7264: out = 16'(-1373);
			7265: out = 16'(2693);
			7266: out = 16'(3018);
			7267: out = 16'(-4125);
			7268: out = 16'(-5327);
			7269: out = 16'(-283);
			7270: out = 16'(-1318);
			7271: out = 16'(420);
			7272: out = 16'(3962);
			7273: out = 16'(1977);
			7274: out = 16'(-6028);
			7275: out = 16'(-5930);
			7276: out = 16'(3558);
			7277: out = 16'(7297);
			7278: out = 16'(3466);
			7279: out = 16'(-1934);
			7280: out = 16'(-1119);
			7281: out = 16'(893);
			7282: out = 16'(-1500);
			7283: out = 16'(-4215);
			7284: out = 16'(-5429);
			7285: out = 16'(-402);
			7286: out = 16'(5780);
			7287: out = 16'(6845);
			7288: out = 16'(-500);
			7289: out = 16'(-2587);
			7290: out = 16'(1763);
			7291: out = 16'(4433);
			7292: out = 16'(4956);
			7293: out = 16'(465);
			7294: out = 16'(-5198);
			7295: out = 16'(-7576);
			7296: out = 16'(-3564);
			7297: out = 16'(-4301);
			7298: out = 16'(-1730);
			7299: out = 16'(3611);
			7300: out = 16'(5435);
			7301: out = 16'(3256);
			7302: out = 16'(-1301);
			7303: out = 16'(-4552);
			7304: out = 16'(-638);
			7305: out = 16'(4572);
			7306: out = 16'(3269);
			7307: out = 16'(-1238);
			7308: out = 16'(-192);
			7309: out = 16'(369);
			7310: out = 16'(-2039);
			7311: out = 16'(461);
			7312: out = 16'(-2618);
			7313: out = 16'(-2647);
			7314: out = 16'(1124);
			7315: out = 16'(2218);
			7316: out = 16'(3392);
			7317: out = 16'(4803);
			7318: out = 16'(3339);
			7319: out = 16'(2619);
			7320: out = 16'(482);
			7321: out = 16'(-816);
			7322: out = 16'(-2877);
			7323: out = 16'(-3904);
			7324: out = 16'(1632);
			7325: out = 16'(1810);
			7326: out = 16'(-46);
			7327: out = 16'(2920);
			7328: out = 16'(3066);
			7329: out = 16'(-1367);
			7330: out = 16'(-6843);
			7331: out = 16'(-8645);
			7332: out = 16'(-3045);
			7333: out = 16'(169);
			7334: out = 16'(6079);
			7335: out = 16'(4855);
			7336: out = 16'(1023);
			7337: out = 16'(633);
			7338: out = 16'(-242);
			7339: out = 16'(2233);
			7340: out = 16'(3456);
			7341: out = 16'(3061);
			7342: out = 16'(-720);
			7343: out = 16'(-616);
			7344: out = 16'(1944);
			7345: out = 16'(999);
			7346: out = 16'(593);
			7347: out = 16'(-848);
			7348: out = 16'(-2875);
			7349: out = 16'(-4256);
			7350: out = 16'(2303);
			7351: out = 16'(1105);
			7352: out = 16'(-3937);
			7353: out = 16'(-705);
			7354: out = 16'(3132);
			7355: out = 16'(3207);
			7356: out = 16'(-3260);
			7357: out = 16'(-518);
			7358: out = 16'(2872);
			7359: out = 16'(5806);
			7360: out = 16'(4431);
			7361: out = 16'(670);
			7362: out = 16'(-3955);
			7363: out = 16'(-5837);
			7364: out = 16'(-8108);
			7365: out = 16'(-2496);
			7366: out = 16'(5953);
			7367: out = 16'(-446);
			7368: out = 16'(-8715);
			7369: out = 16'(-3432);
			7370: out = 16'(761);
			7371: out = 16'(4365);
			7372: out = 16'(6755);
			7373: out = 16'(4834);
			7374: out = 16'(-1606);
			7375: out = 16'(-6449);
			7376: out = 16'(-5925);
			7377: out = 16'(-2829);
			7378: out = 16'(3622);
			7379: out = 16'(7022);
			7380: out = 16'(4695);
			7381: out = 16'(1344);
			7382: out = 16'(464);
			7383: out = 16'(2683);
			7384: out = 16'(4577);
			7385: out = 16'(1125);
			7386: out = 16'(-3747);
			7387: out = 16'(-2922);
			7388: out = 16'(2615);
			7389: out = 16'(2021);
			7390: out = 16'(-4889);
			7391: out = 16'(-4931);
			7392: out = 16'(-371);
			7393: out = 16'(631);
			7394: out = 16'(-570);
			7395: out = 16'(2760);
			7396: out = 16'(-1837);
			7397: out = 16'(-1906);
			7398: out = 16'(2429);
			7399: out = 16'(7317);
			7400: out = 16'(2743);
			7401: out = 16'(-6090);
			7402: out = 16'(-7729);
			7403: out = 16'(-1120);
			7404: out = 16'(4223);
			7405: out = 16'(-18);
			7406: out = 16'(-4801);
			7407: out = 16'(-2737);
			7408: out = 16'(40);
			7409: out = 16'(2658);
			7410: out = 16'(5387);
			7411: out = 16'(2520);
			7412: out = 16'(-395);
			7413: out = 16'(-3670);
			7414: out = 16'(-4049);
			7415: out = 16'(724);
			7416: out = 16'(2749);
			7417: out = 16'(4912);
			7418: out = 16'(7512);
			7419: out = 16'(1900);
			7420: out = 16'(-2955);
			7421: out = 16'(-5971);
			7422: out = 16'(-2393);
			7423: out = 16'(3352);
			7424: out = 16'(2939);
			7425: out = 16'(-155);
			7426: out = 16'(261);
			7427: out = 16'(-3996);
			7428: out = 16'(-4101);
			7429: out = 16'(1922);
			7430: out = 16'(-289);
			7431: out = 16'(1331);
			7432: out = 16'(5358);
			7433: out = 16'(4294);
			7434: out = 16'(-5542);
			7435: out = 16'(-9361);
			7436: out = 16'(-4952);
			7437: out = 16'(2776);
			7438: out = 16'(6852);
			7439: out = 16'(4146);
			7440: out = 16'(-2904);
			7441: out = 16'(-4219);
			7442: out = 16'(-4012);
			7443: out = 16'(-1254);
			7444: out = 16'(6696);
			7445: out = 16'(7761);
			7446: out = 16'(-2237);
			7447: out = 16'(-5666);
			7448: out = 16'(-4035);
			7449: out = 16'(-546);
			7450: out = 16'(3852);
			7451: out = 16'(817);
			7452: out = 16'(-934);
			7453: out = 16'(1835);
			7454: out = 16'(7906);
			7455: out = 16'(5699);
			7456: out = 16'(-955);
			7457: out = 16'(-3496);
			7458: out = 16'(-66);
			7459: out = 16'(3200);
			7460: out = 16'(4493);
			7461: out = 16'(2321);
			7462: out = 16'(822);
			7463: out = 16'(-905);
			7464: out = 16'(-3752);
			7465: out = 16'(-7575);
			7466: out = 16'(-4716);
			7467: out = 16'(1291);
			7468: out = 16'(-742);
			7469: out = 16'(-4719);
			7470: out = 16'(828);
			7471: out = 16'(3731);
			7472: out = 16'(1932);
			7473: out = 16'(-1586);
			7474: out = 16'(-1055);
			7475: out = 16'(-3358);
			7476: out = 16'(-4391);
			7477: out = 16'(2326);
			7478: out = 16'(6131);
			7479: out = 16'(1689);
			7480: out = 16'(-499);
			7481: out = 16'(1437);
			7482: out = 16'(2590);
			7483: out = 16'(-1240);
			7484: out = 16'(-7854);
			7485: out = 16'(-6607);
			7486: out = 16'(-1873);
			7487: out = 16'(4327);
			7488: out = 16'(3499);
			7489: out = 16'(-925);
			7490: out = 16'(-3490);
			7491: out = 16'(-921);
			7492: out = 16'(6078);
			7493: out = 16'(6347);
			7494: out = 16'(106);
			7495: out = 16'(-4427);
			7496: out = 16'(-2715);
			7497: out = 16'(3025);
			7498: out = 16'(3081);
			7499: out = 16'(-2391);
			7500: out = 16'(-1666);
			7501: out = 16'(2494);
			7502: out = 16'(479);
			7503: out = 16'(-785);
			7504: out = 16'(-189);
			7505: out = 16'(1169);
			7506: out = 16'(4790);
			7507: out = 16'(1365);
			7508: out = 16'(-257);
			7509: out = 16'(-261);
			7510: out = 16'(-1198);
			7511: out = 16'(2214);
			7512: out = 16'(182);
			7513: out = 16'(-329);
			7514: out = 16'(423);
			7515: out = 16'(-1793);
			7516: out = 16'(-1934);
			7517: out = 16'(-1744);
			7518: out = 16'(-1014);
			7519: out = 16'(2286);
			7520: out = 16'(556);
			7521: out = 16'(-995);
			7522: out = 16'(1357);
			7523: out = 16'(2674);
			7524: out = 16'(1329);
			7525: out = 16'(-3298);
			7526: out = 16'(-5028);
			7527: out = 16'(-3125);
			7528: out = 16'(809);
			7529: out = 16'(4316);
			7530: out = 16'(1452);
			7531: out = 16'(-2220);
			7532: out = 16'(-557);
			7533: out = 16'(1133);
			7534: out = 16'(-3648);
			7535: out = 16'(-5320);
			7536: out = 16'(-1274);
			7537: out = 16'(-486);
			7538: out = 16'(1696);
			7539: out = 16'(-383);
			7540: out = 16'(-3919);
			7541: out = 16'(206);
			7542: out = 16'(5315);
			7543: out = 16'(3740);
			7544: out = 16'(-981);
			7545: out = 16'(-3252);
			7546: out = 16'(-1410);
			7547: out = 16'(5855);
			7548: out = 16'(4628);
			7549: out = 16'(-2705);
			7550: out = 16'(-6453);
			7551: out = 16'(-2011);
			7552: out = 16'(5507);
			7553: out = 16'(4745);
			7554: out = 16'(-2825);
			7555: out = 16'(-1707);
			7556: out = 16'(1612);
			7557: out = 16'(2342);
			7558: out = 16'(1727);
			7559: out = 16'(17);
			7560: out = 16'(-3313);
			7561: out = 16'(-5568);
			7562: out = 16'(-6361);
			7563: out = 16'(199);
			7564: out = 16'(6770);
			7565: out = 16'(2144);
			7566: out = 16'(-6000);
			7567: out = 16'(-1231);
			7568: out = 16'(2329);
			7569: out = 16'(725);
			7570: out = 16'(405);
			7571: out = 16'(-265);
			7572: out = 16'(-3351);
			7573: out = 16'(-1763);
			7574: out = 16'(-279);
			7575: out = 16'(-3159);
			7576: out = 16'(1969);
			7577: out = 16'(2901);
			7578: out = 16'(3537);
			7579: out = 16'(384);
			7580: out = 16'(-4170);
			7581: out = 16'(348);
			7582: out = 16'(5776);
			7583: out = 16'(6414);
			7584: out = 16'(1276);
			7585: out = 16'(-5206);
			7586: out = 16'(-4486);
			7587: out = 16'(-2833);
			7588: out = 16'(-562);
			7589: out = 16'(1793);
			7590: out = 16'(2826);
			7591: out = 16'(-2151);
			7592: out = 16'(-3213);
			7593: out = 16'(2914);
			7594: out = 16'(1838);
			7595: out = 16'(3466);
			7596: out = 16'(4204);
			7597: out = 16'(5237);
			7598: out = 16'(1359);
			7599: out = 16'(-3544);
			7600: out = 16'(-4756);
			7601: out = 16'(-985);
			7602: out = 16'(2384);
			7603: out = 16'(-1131);
			7604: out = 16'(-3777);
			7605: out = 16'(-1039);
			7606: out = 16'(1172);
			7607: out = 16'(1246);
			7608: out = 16'(-743);
			7609: out = 16'(1743);
			7610: out = 16'(2432);
			7611: out = 16'(2779);
			7612: out = 16'(781);
			7613: out = 16'(-2548);
			7614: out = 16'(-4623);
			7615: out = 16'(-3720);
			7616: out = 16'(381);
			7617: out = 16'(-1021);
			7618: out = 16'(-3014);
			7619: out = 16'(15);
			7620: out = 16'(2991);
			7621: out = 16'(3479);
			7622: out = 16'(-1452);
			7623: out = 16'(-3713);
			7624: out = 16'(-1033);
			7625: out = 16'(2052);
			7626: out = 16'(1318);
			7627: out = 16'(-103);
			7628: out = 16'(2218);
			7629: out = 16'(2031);
			7630: out = 16'(-392);
			7631: out = 16'(1284);
			7632: out = 16'(377);
			7633: out = 16'(-1700);
			7634: out = 16'(-2163);
			7635: out = 16'(1189);
			7636: out = 16'(3507);
			7637: out = 16'(-2111);
			7638: out = 16'(-3622);
			7639: out = 16'(-1690);
			7640: out = 16'(-533);
			7641: out = 16'(1734);
			7642: out = 16'(948);
			7643: out = 16'(-2696);
			7644: out = 16'(-2856);
			7645: out = 16'(989);
			7646: out = 16'(-1460);
			7647: out = 16'(-4528);
			7648: out = 16'(-2902);
			7649: out = 16'(736);
			7650: out = 16'(271);
			7651: out = 16'(-311);
			7652: out = 16'(2167);
			7653: out = 16'(5976);
			7654: out = 16'(2970);
			7655: out = 16'(-5282);
			7656: out = 16'(-9783);
			7657: out = 16'(-4887);
			7658: out = 16'(3087);
			7659: out = 16'(1534);
			7660: out = 16'(-1447);
			7661: out = 16'(951);
			7662: out = 16'(4062);
			7663: out = 16'(6106);
			7664: out = 16'(-970);
			7665: out = 16'(-4750);
			7666: out = 16'(-937);
			7667: out = 16'(3004);
			7668: out = 16'(4249);
			7669: out = 16'(4473);
			7670: out = 16'(3762);
			7671: out = 16'(-349);
			7672: out = 16'(-7121);
			7673: out = 16'(-8905);
			7674: out = 16'(-4691);
			7675: out = 16'(-359);
			7676: out = 16'(2781);
			7677: out = 16'(2498);
			7678: out = 16'(-1890);
			7679: out = 16'(-2225);
			7680: out = 16'(3182);
			7681: out = 16'(6879);
			7682: out = 16'(6139);
			7683: out = 16'(-1928);
			7684: out = 16'(-4825);
			7685: out = 16'(-1443);
			7686: out = 16'(-1106);
			7687: out = 16'(2872);
			7688: out = 16'(4126);
			7689: out = 16'(960);
			7690: out = 16'(-1219);
			7691: out = 16'(-482);
			7692: out = 16'(495);
			7693: out = 16'(-1370);
			7694: out = 16'(-418);
			7695: out = 16'(1380);
			7696: out = 16'(4371);
			7697: out = 16'(6677);
			7698: out = 16'(1121);
			7699: out = 16'(-3492);
			7700: out = 16'(-4134);
			7701: out = 16'(-2905);
			7702: out = 16'(-815);
			7703: out = 16'(1960);
			7704: out = 16'(3488);
			7705: out = 16'(-302);
			7706: out = 16'(-5252);
			7707: out = 16'(-2796);
			7708: out = 16'(-28);
			7709: out = 16'(3824);
			7710: out = 16'(1015);
			7711: out = 16'(-2448);
			7712: out = 16'(-2410);
			7713: out = 16'(517);
			7714: out = 16'(3401);
			7715: out = 16'(5544);
			7716: out = 16'(1677);
			7717: out = 16'(-3120);
			7718: out = 16'(-1966);
			7719: out = 16'(-1088);
			7720: out = 16'(435);
			7721: out = 16'(2458);
			7722: out = 16'(1840);
			7723: out = 16'(-120);
			7724: out = 16'(-3010);
			7725: out = 16'(-2075);
			7726: out = 16'(-2270);
			7727: out = 16'(-2573);
			7728: out = 16'(599);
			7729: out = 16'(4886);
			7730: out = 16'(2355);
			7731: out = 16'(-634);
			7732: out = 16'(-986);
			7733: out = 16'(2596);
			7734: out = 16'(3620);
			7735: out = 16'(679);
			7736: out = 16'(2079);
			7737: out = 16'(1266);
			7738: out = 16'(-1842);
			7739: out = 16'(-3827);
			7740: out = 16'(-1095);
			7741: out = 16'(99);
			7742: out = 16'(-352);
			7743: out = 16'(-573);
			7744: out = 16'(-2040);
			7745: out = 16'(-6851);
			7746: out = 16'(-4428);
			7747: out = 16'(990);
			7748: out = 16'(2938);
			7749: out = 16'(1476);
			7750: out = 16'(1507);
			7751: out = 16'(1767);
			7752: out = 16'(-1358);
			7753: out = 16'(754);
			7754: out = 16'(-1412);
			7755: out = 16'(3064);
			7756: out = 16'(5926);
			7757: out = 16'(3247);
			7758: out = 16'(2165);
			7759: out = 16'(908);
			7760: out = 16'(-164);
			7761: out = 16'(-1275);
			7762: out = 16'(-4781);
			7763: out = 16'(-3393);
			7764: out = 16'(2344);
			7765: out = 16'(2205);
			7766: out = 16'(-2353);
			7767: out = 16'(-1038);
			7768: out = 16'(178);
			7769: out = 16'(793);
			7770: out = 16'(900);
			7771: out = 16'(306);
			7772: out = 16'(2211);
			7773: out = 16'(1883);
			7774: out = 16'(1771);
			7775: out = 16'(-1393);
			7776: out = 16'(-4436);
			7777: out = 16'(-3578);
			7778: out = 16'(-1850);
			7779: out = 16'(664);
			7780: out = 16'(2648);
			7781: out = 16'(2471);
			7782: out = 16'(1681);
			7783: out = 16'(-1477);
			7784: out = 16'(931);
			7785: out = 16'(2879);
			7786: out = 16'(-590);
			7787: out = 16'(692);
			7788: out = 16'(3050);
			7789: out = 16'(-1321);
			7790: out = 16'(-4673);
			7791: out = 16'(-1512);
			7792: out = 16'(1225);
			7793: out = 16'(-55);
			7794: out = 16'(-5297);
			7795: out = 16'(-4595);
			7796: out = 16'(190);
			7797: out = 16'(2194);
			7798: out = 16'(2477);
			7799: out = 16'(-2671);
			7800: out = 16'(-6875);
			7801: out = 16'(-417);
			7802: out = 16'(3572);
			7803: out = 16'(4217);
			7804: out = 16'(1651);
			7805: out = 16'(-4381);
			7806: out = 16'(-1447);
			7807: out = 16'(166);
			7808: out = 16'(2284);
			7809: out = 16'(4878);
			7810: out = 16'(3287);
			7811: out = 16'(1076);
			7812: out = 16'(-3366);
			7813: out = 16'(-6731);
			7814: out = 16'(-5575);
			7815: out = 16'(-1162);
			7816: out = 16'(4610);
			7817: out = 16'(6122);
			7818: out = 16'(3351);
			7819: out = 16'(-1133);
			7820: out = 16'(-2694);
			7821: out = 16'(-89);
			7822: out = 16'(2888);
			7823: out = 16'(2891);
			7824: out = 16'(-1946);
			7825: out = 16'(-469);
			7826: out = 16'(3946);
			7827: out = 16'(5670);
			7828: out = 16'(-893);
			7829: out = 16'(-4063);
			7830: out = 16'(-4014);
			7831: out = 16'(-1271);
			7832: out = 16'(-1240);
			7833: out = 16'(260);
			7834: out = 16'(-24);
			7835: out = 16'(-1246);
			7836: out = 16'(68);
			7837: out = 16'(3828);
			7838: out = 16'(7776);
			7839: out = 16'(2335);
			7840: out = 16'(-3641);
			7841: out = 16'(-4615);
			7842: out = 16'(-815);
			7843: out = 16'(615);
			7844: out = 16'(-4579);
			7845: out = 16'(-1903);
			7846: out = 16'(3680);
			7847: out = 16'(3135);
			7848: out = 16'(-1695);
			7849: out = 16'(-3374);
			7850: out = 16'(72);
			7851: out = 16'(1047);
			7852: out = 16'(2831);
			7853: out = 16'(5310);
			7854: out = 16'(820);
			7855: out = 16'(-7153);
			7856: out = 16'(-9117);
			7857: out = 16'(-6802);
			7858: out = 16'(-640);
			7859: out = 16'(6109);
			7860: out = 16'(229);
			7861: out = 16'(-3478);
			7862: out = 16'(1295);
			7863: out = 16'(6339);
			7864: out = 16'(4528);
			7865: out = 16'(-3754);
			7866: out = 16'(-5403);
			7867: out = 16'(-1746);
			7868: out = 16'(4597);
			7869: out = 16'(7297);
			7870: out = 16'(-1102);
			7871: out = 16'(-5333);
			7872: out = 16'(-1743);
			7873: out = 16'(-237);
			7874: out = 16'(3268);
			7875: out = 16'(2088);
			7876: out = 16'(-236);
			7877: out = 16'(-1060);
			7878: out = 16'(-756);
			7879: out = 16'(-915);
			7880: out = 16'(-631);
			7881: out = 16'(-1102);
			7882: out = 16'(2397);
			7883: out = 16'(2024);
			7884: out = 16'(-142);
			7885: out = 16'(494);
			7886: out = 16'(-398);
			7887: out = 16'(-3435);
			7888: out = 16'(-5752);
			7889: out = 16'(-3481);
			7890: out = 16'(3816);
			7891: out = 16'(5107);
			7892: out = 16'(726);
			7893: out = 16'(-1397);
			7894: out = 16'(-1173);
			7895: out = 16'(2517);
			7896: out = 16'(5770);
			7897: out = 16'(4552);
			7898: out = 16'(-707);
			7899: out = 16'(-3704);
			7900: out = 16'(-1523);
			7901: out = 16'(-1083);
			7902: out = 16'(-963);
			7903: out = 16'(-1563);
			7904: out = 16'(404);
			7905: out = 16'(2146);
			7906: out = 16'(-183);
			7907: out = 16'(-2155);
			7908: out = 16'(-1073);
			7909: out = 16'(205);
			7910: out = 16'(-1903);
			7911: out = 16'(1410);
			7912: out = 16'(186);
			7913: out = 16'(-548);
			7914: out = 16'(547);
			7915: out = 16'(412);
			7916: out = 16'(442);
			7917: out = 16'(-465);
			7918: out = 16'(866);
			7919: out = 16'(4150);
			7920: out = 16'(5044);
			7921: out = 16'(648);
			7922: out = 16'(-4668);
			7923: out = 16'(-5350);
			7924: out = 16'(210);
			7925: out = 16'(3146);
			7926: out = 16'(1054);
			7927: out = 16'(-3446);
			7928: out = 16'(-2589);
			7929: out = 16'(784);
			7930: out = 16'(3187);
			7931: out = 16'(-2697);
			7932: out = 16'(-3367);
			7933: out = 16'(446);
			7934: out = 16'(3030);
			7935: out = 16'(4094);
			7936: out = 16'(492);
			7937: out = 16'(-245);
			7938: out = 16'(-586);
			7939: out = 16'(-1048);
			7940: out = 16'(496);
			7941: out = 16'(365);
			7942: out = 16'(2614);
			7943: out = 16'(3449);
			7944: out = 16'(1283);
			7945: out = 16'(-754);
			7946: out = 16'(-1913);
			7947: out = 16'(331);
			7948: out = 16'(3077);
			7949: out = 16'(1222);
			7950: out = 16'(-3377);
			7951: out = 16'(-1838);
			7952: out = 16'(-1116);
			7953: out = 16'(-1044);
			7954: out = 16'(-3640);
			7955: out = 16'(-1883);
			7956: out = 16'(416);
			7957: out = 16'(-508);
			7958: out = 16'(2493);
			7959: out = 16'(2337);
			7960: out = 16'(904);
			7961: out = 16'(-3533);
			7962: out = 16'(-2328);
			7963: out = 16'(-2720);
			7964: out = 16'(414);
			7965: out = 16'(2188);
			7966: out = 16'(-270);
			7967: out = 16'(-3330);
			7968: out = 16'(-242);
			7969: out = 16'(3626);
			7970: out = 16'(1000);
			7971: out = 16'(-3634);
			7972: out = 16'(-3103);
			7973: out = 16'(2577);
			7974: out = 16'(-833);
			7975: out = 16'(-1566);
			7976: out = 16'(4160);
			7977: out = 16'(2839);
			7978: out = 16'(-2656);
			7979: out = 16'(-1400);
			7980: out = 16'(128);
			7981: out = 16'(-658);
			7982: out = 16'(-1988);
			7983: out = 16'(-1288);
			7984: out = 16'(-1110);
			7985: out = 16'(670);
			7986: out = 16'(1250);
			7987: out = 16'(-2857);
			7988: out = 16'(-1411);
			7989: out = 16'(-118);
			7990: out = 16'(1093);
			7991: out = 16'(4772);
			7992: out = 16'(2578);
			7993: out = 16'(-411);
			7994: out = 16'(-1810);
			7995: out = 16'(-1122);
			7996: out = 16'(46);
			7997: out = 16'(-261);
			7998: out = 16'(724);
			7999: out = 16'(2294);
			8000: out = 16'(1931);
			8001: out = 16'(1237);
			8002: out = 16'(-1417);
			8003: out = 16'(-3387);
			8004: out = 16'(-6255);
			8005: out = 16'(-3928);
			8006: out = 16'(3168);
			8007: out = 16'(5757);
			8008: out = 16'(23);
			8009: out = 16'(-2440);
			8010: out = 16'(163);
			8011: out = 16'(1758);
			8012: out = 16'(901);
			8013: out = 16'(-1293);
			8014: out = 16'(-4485);
			8015: out = 16'(-3062);
			8016: out = 16'(2595);
			8017: out = 16'(3241);
			8018: out = 16'(398);
			8019: out = 16'(-2671);
			8020: out = 16'(-190);
			8021: out = 16'(5586);
			8022: out = 16'(5971);
			8023: out = 16'(573);
			8024: out = 16'(-5799);
			8025: out = 16'(-5084);
			8026: out = 16'(-3335);
			8027: out = 16'(1377);
			8028: out = 16'(4181);
			8029: out = 16'(90);
			8030: out = 16'(-5865);
			8031: out = 16'(-3693);
			8032: out = 16'(-170);
			8033: out = 16'(1661);
			8034: out = 16'(4007);
			8035: out = 16'(1399);
			8036: out = 16'(-3059);
			8037: out = 16'(-1799);
			8038: out = 16'(-973);
			8039: out = 16'(-1050);
			8040: out = 16'(215);
			8041: out = 16'(-807);
			8042: out = 16'(1212);
			8043: out = 16'(2477);
			8044: out = 16'(1829);
			8045: out = 16'(628);
			8046: out = 16'(1749);
			8047: out = 16'(-562);
			8048: out = 16'(-2783);
			8049: out = 16'(-1954);
			8050: out = 16'(-2279);
			8051: out = 16'(3880);
			8052: out = 16'(7133);
			8053: out = 16'(1004);
			8054: out = 16'(-3886);
			8055: out = 16'(-4328);
			8056: out = 16'(-284);
			8057: out = 16'(5492);
			8058: out = 16'(4577);
			8059: out = 16'(-1669);
			8060: out = 16'(-5983);
			8061: out = 16'(-4092);
			8062: out = 16'(3571);
			8063: out = 16'(5907);
			8064: out = 16'(1733);
			8065: out = 16'(-3753);
			8066: out = 16'(-2638);
			8067: out = 16'(-3717);
			8068: out = 16'(-2346);
			8069: out = 16'(1321);
			8070: out = 16'(2535);
			8071: out = 16'(3555);
			8072: out = 16'(1337);
			8073: out = 16'(-2611);
			8074: out = 16'(-1535);
			8075: out = 16'(2596);
			8076: out = 16'(3215);
			8077: out = 16'(1549);
			8078: out = 16'(-2706);
			8079: out = 16'(-4668);
			8080: out = 16'(-810);
			8081: out = 16'(2700);
			8082: out = 16'(2918);
			8083: out = 16'(1346);
			8084: out = 16'(1165);
			8085: out = 16'(1289);
			8086: out = 16'(530);
			8087: out = 16'(-1146);
			8088: out = 16'(-3631);
			8089: out = 16'(-2572);
			8090: out = 16'(3507);
			8091: out = 16'(2626);
			8092: out = 16'(-2210);
			8093: out = 16'(-1242);
			8094: out = 16'(3285);
			8095: out = 16'(6063);
			8096: out = 16'(1321);
			8097: out = 16'(-3171);
			8098: out = 16'(-1975);
			8099: out = 16'(846);
			8100: out = 16'(2824);
			8101: out = 16'(599);
			8102: out = 16'(-2163);
			8103: out = 16'(-955);
			8104: out = 16'(2357);
			8105: out = 16'(1595);
			8106: out = 16'(2271);
			8107: out = 16'(2492);
			8108: out = 16'(1898);
			8109: out = 16'(-1584);
			8110: out = 16'(-3345);
			8111: out = 16'(-2828);
			8112: out = 16'(-3602);
			8113: out = 16'(-4959);
			8114: out = 16'(381);
			8115: out = 16'(1852);
			8116: out = 16'(204);
			8117: out = 16'(-332);
			8118: out = 16'(3811);
			8119: out = 16'(4730);
			8120: out = 16'(-2040);
			8121: out = 16'(-5934);
			8122: out = 16'(-3648);
			8123: out = 16'(-1019);
			8124: out = 16'(-553);
			8125: out = 16'(593);
			8126: out = 16'(-164);
			8127: out = 16'(-1687);
			8128: out = 16'(128);
			8129: out = 16'(-519);
			8130: out = 16'(-2209);
			8131: out = 16'(1751);
			8132: out = 16'(4583);
			8133: out = 16'(3262);
			8134: out = 16'(-570);
			8135: out = 16'(-1961);
			8136: out = 16'(256);
			8137: out = 16'(1037);
			8138: out = 16'(-976);
			8139: out = 16'(-2223);
			8140: out = 16'(-1769);
			8141: out = 16'(-633);
			8142: out = 16'(2970);
			8143: out = 16'(3544);
			8144: out = 16'(-4458);
			8145: out = 16'(-7139);
			8146: out = 16'(-1051);
			8147: out = 16'(4500);
			8148: out = 16'(4598);
			8149: out = 16'(1295);
			8150: out = 16'(-489);
			8151: out = 16'(-93);
			8152: out = 16'(3185);
			8153: out = 16'(3400);
			8154: out = 16'(562);
			8155: out = 16'(-97);
			8156: out = 16'(-781);
			8157: out = 16'(-572);
			8158: out = 16'(167);
			8159: out = 16'(1264);
			8160: out = 16'(2227);
			8161: out = 16'(-168);
			8162: out = 16'(-2873);
			8163: out = 16'(-2068);
			8164: out = 16'(-2291);
			8165: out = 16'(-1326);
			8166: out = 16'(865);
			8167: out = 16'(1342);
			8168: out = 16'(-863);
			8169: out = 16'(1018);
			8170: out = 16'(3062);
			8171: out = 16'(-619);
			8172: out = 16'(-3281);
			8173: out = 16'(-2273);
			8174: out = 16'(355);
			8175: out = 16'(574);
			8176: out = 16'(722);
			8177: out = 16'(2028);
			8178: out = 16'(1348);
			8179: out = 16'(478);
			8180: out = 16'(-2125);
			8181: out = 16'(-2116);
			8182: out = 16'(3065);
			8183: out = 16'(3351);
			8184: out = 16'(-918);
			8185: out = 16'(-1885);
			8186: out = 16'(-315);
			8187: out = 16'(357);
			8188: out = 16'(2062);
			8189: out = 16'(4243);
			8190: out = 16'(1216);
			8191: out = 16'(-3124);
			8192: out = 16'(-3395);
			8193: out = 16'(-4382);
			8194: out = 16'(1485);
			8195: out = 16'(7141);
			8196: out = 16'(2490);
			8197: out = 16'(-2413);
			8198: out = 16'(-1000);
			8199: out = 16'(1756);
			8200: out = 16'(3043);
			8201: out = 16'(324);
			8202: out = 16'(471);
			8203: out = 16'(1743);
			8204: out = 16'(1869);
			8205: out = 16'(3226);
			8206: out = 16'(2675);
			8207: out = 16'(-1480);
			8208: out = 16'(-5444);
			8209: out = 16'(-5674);
			8210: out = 16'(-1647);
			8211: out = 16'(3149);
			8212: out = 16'(-1072);
			8213: out = 16'(-5453);
			8214: out = 16'(-2545);
			8215: out = 16'(1732);
			8216: out = 16'(1513);
			8217: out = 16'(304);
			8218: out = 16'(-3);
			8219: out = 16'(-3895);
			8220: out = 16'(-3500);
			8221: out = 16'(-352);
			8222: out = 16'(3100);
			8223: out = 16'(4524);
			8224: out = 16'(-80);
			8225: out = 16'(-5304);
			8226: out = 16'(-5320);
			8227: out = 16'(299);
			8228: out = 16'(3220);
			8229: out = 16'(-2990);
			8230: out = 16'(-1746);
			8231: out = 16'(3268);
			8232: out = 16'(2803);
			8233: out = 16'(990);
			8234: out = 16'(-134);
			8235: out = 16'(39);
			8236: out = 16'(1055);
			8237: out = 16'(312);
			8238: out = 16'(-2494);
			8239: out = 16'(-1849);
			8240: out = 16'(3147);
			8241: out = 16'(5216);
			8242: out = 16'(554);
			8243: out = 16'(-5349);
			8244: out = 16'(-3156);
			8245: out = 16'(1709);
			8246: out = 16'(3879);
			8247: out = 16'(-152);
			8248: out = 16'(-3323);
			8249: out = 16'(-1091);
			8250: out = 16'(-1768);
			8251: out = 16'(1311);
			8252: out = 16'(4566);
			8253: out = 16'(-333);
			8254: out = 16'(-2117);
			8255: out = 16'(-622);
			8256: out = 16'(-448);
			8257: out = 16'(-3160);
			8258: out = 16'(-3146);
			8259: out = 16'(-1026);
			8260: out = 16'(2824);
			8261: out = 16'(6757);
			8262: out = 16'(4729);
			8263: out = 16'(-2259);
			8264: out = 16'(-4528);
			8265: out = 16'(-1531);
			8266: out = 16'(304);
			8267: out = 16'(2230);
			8268: out = 16'(3701);
			8269: out = 16'(1358);
			8270: out = 16'(-3812);
			8271: out = 16'(-3314);
			8272: out = 16'(1102);
			8273: out = 16'(2545);
			8274: out = 16'(2472);
			8275: out = 16'(-2285);
			8276: out = 16'(-6100);
			8277: out = 16'(-2134);
			8278: out = 16'(2054);
			8279: out = 16'(3399);
			8280: out = 16'(-1034);
			8281: out = 16'(-1562);
			8282: out = 16'(1846);
			8283: out = 16'(1057);
			8284: out = 16'(133);
			8285: out = 16'(714);
			8286: out = 16'(-559);
			8287: out = 16'(-1212);
			8288: out = 16'(-309);
			8289: out = 16'(34);
			8290: out = 16'(457);
			8291: out = 16'(-2521);
			8292: out = 16'(-2048);
			8293: out = 16'(2445);
			8294: out = 16'(1449);
			8295: out = 16'(-544);
			8296: out = 16'(1406);
			8297: out = 16'(1013);
			8298: out = 16'(-5628);
			8299: out = 16'(-8053);
			8300: out = 16'(-3081);
			8301: out = 16'(691);
			8302: out = 16'(5385);
			8303: out = 16'(5188);
			8304: out = 16'(-622);
			8305: out = 16'(-3035);
			8306: out = 16'(-1187);
			8307: out = 16'(3877);
			8308: out = 16'(5612);
			8309: out = 16'(2217);
			8310: out = 16'(-1129);
			8311: out = 16'(-650);
			8312: out = 16'(-188);
			8313: out = 16'(-486);
			8314: out = 16'(-3335);
			8315: out = 16'(-2931);
			8316: out = 16'(-460);
			8317: out = 16'(756);
			8318: out = 16'(2247);
			8319: out = 16'(1528);
			8320: out = 16'(-2153);
			8321: out = 16'(-1750);
			8322: out = 16'(356);
			8323: out = 16'(-2862);
			8324: out = 16'(-2891);
			8325: out = 16'(-1247);
			8326: out = 16'(-73);
			8327: out = 16'(3236);
			8328: out = 16'(2905);
			8329: out = 16'(2604);
			8330: out = 16'(1383);
			8331: out = 16'(-1024);
			8332: out = 16'(-3526);
			8333: out = 16'(-2115);
			8334: out = 16'(399);
			8335: out = 16'(1519);
			8336: out = 16'(2885);
			8337: out = 16'(706);
			8338: out = 16'(1822);
			8339: out = 16'(1831);
			8340: out = 16'(-1221);
			8341: out = 16'(-604);
			8342: out = 16'(665);
			8343: out = 16'(1946);
			8344: out = 16'(2498);
			8345: out = 16'(468);
			8346: out = 16'(-1051);
			8347: out = 16'(-1185);
			8348: out = 16'(-1990);
			8349: out = 16'(-2040);
			8350: out = 16'(-2383);
			8351: out = 16'(-1952);
			8352: out = 16'(-2588);
			8353: out = 16'(-2533);
			8354: out = 16'(1663);
			8355: out = 16'(3821);
			8356: out = 16'(1399);
			8357: out = 16'(-1633);
			8358: out = 16'(-1362);
			8359: out = 16'(-224);
			8360: out = 16'(319);
			8361: out = 16'(835);
			8362: out = 16'(2286);
			8363: out = 16'(691);
			8364: out = 16'(344);
			8365: out = 16'(-541);
			8366: out = 16'(-975);
			8367: out = 16'(-1247);
			8368: out = 16'(-1541);
			8369: out = 16'(-246);
			8370: out = 16'(1248);
			8371: out = 16'(3453);
			8372: out = 16'(361);
			8373: out = 16'(-1961);
			8374: out = 16'(-3523);
			8375: out = 16'(-1511);
			8376: out = 16'(1508);
			8377: out = 16'(3169);
			8378: out = 16'(1483);
			8379: out = 16'(734);
			8380: out = 16'(1786);
			8381: out = 16'(1143);
			8382: out = 16'(-983);
			8383: out = 16'(-1243);
			8384: out = 16'(-2487);
			8385: out = 16'(-2994);
			8386: out = 16'(-252);
			8387: out = 16'(3529);
			8388: out = 16'(820);
			8389: out = 16'(-1697);
			8390: out = 16'(-719);
			8391: out = 16'(-585);
			8392: out = 16'(-3110);
			8393: out = 16'(-4494);
			8394: out = 16'(2141);
			8395: out = 16'(1120);
			8396: out = 16'(653);
			8397: out = 16'(5055);
			8398: out = 16'(3531);
			8399: out = 16'(-500);
			8400: out = 16'(-4645);
			8401: out = 16'(-2184);
			8402: out = 16'(3925);
			8403: out = 16'(4987);
			8404: out = 16'(181);
			8405: out = 16'(-3413);
			8406: out = 16'(-3475);
			8407: out = 16'(-1406);
			8408: out = 16'(205);
			8409: out = 16'(-281);
			8410: out = 16'(-1057);
			8411: out = 16'(-40);
			8412: out = 16'(-1043);
			8413: out = 16'(-339);
			8414: out = 16'(871);
			8415: out = 16'(1853);
			8416: out = 16'(2543);
			8417: out = 16'(-1191);
			8418: out = 16'(-1524);
			8419: out = 16'(-791);
			8420: out = 16'(1573);
			8421: out = 16'(662);
			8422: out = 16'(-1361);
			8423: out = 16'(1487);
			8424: out = 16'(-67);
			8425: out = 16'(1341);
			8426: out = 16'(2126);
			8427: out = 16'(1390);
			8428: out = 16'(-127);
			8429: out = 16'(81);
			8430: out = 16'(-1510);
			8431: out = 16'(463);
			8432: out = 16'(2219);
			8433: out = 16'(875);
			8434: out = 16'(-511);
			8435: out = 16'(-1752);
			8436: out = 16'(-607);
			8437: out = 16'(-849);
			8438: out = 16'(714);
			8439: out = 16'(2241);
			8440: out = 16'(-1849);
			8441: out = 16'(-3467);
			8442: out = 16'(-367);
			8443: out = 16'(4029);
			8444: out = 16'(-857);
			8445: out = 16'(-4893);
			8446: out = 16'(-170);
			8447: out = 16'(3906);
			8448: out = 16'(3260);
			8449: out = 16'(792);
			8450: out = 16'(-606);
			8451: out = 16'(-162);
			8452: out = 16'(-1186);
			8453: out = 16'(-3784);
			8454: out = 16'(-154);
			8455: out = 16'(2855);
			8456: out = 16'(127);
			8457: out = 16'(-2176);
			8458: out = 16'(-1571);
			8459: out = 16'(-635);
			8460: out = 16'(-220);
			8461: out = 16'(965);
			8462: out = 16'(1639);
			8463: out = 16'(1809);
			8464: out = 16'(2213);
			8465: out = 16'(-686);
			8466: out = 16'(-2595);
			8467: out = 16'(-2499);
			8468: out = 16'(-1457);
			8469: out = 16'(1788);
			8470: out = 16'(2603);
			8471: out = 16'(1900);
			8472: out = 16'(2384);
			8473: out = 16'(2192);
			8474: out = 16'(-2833);
			8475: out = 16'(-4102);
			8476: out = 16'(-4853);
			8477: out = 16'(635);
			8478: out = 16'(5981);
			8479: out = 16'(3566);
			8480: out = 16'(-2585);
			8481: out = 16'(-1817);
			8482: out = 16'(-3);
			8483: out = 16'(1518);
			8484: out = 16'(1897);
			8485: out = 16'(-448);
			8486: out = 16'(-1749);
			8487: out = 16'(-1115);
			8488: out = 16'(-1282);
			8489: out = 16'(-1895);
			8490: out = 16'(589);
			8491: out = 16'(444);
			8492: out = 16'(807);
			8493: out = 16'(2373);
			8494: out = 16'(3096);
			8495: out = 16'(-313);
			8496: out = 16'(-2226);
			8497: out = 16'(-1260);
			8498: out = 16'(521);
			8499: out = 16'(1936);
			8500: out = 16'(231);
			8501: out = 16'(-3041);
			8502: out = 16'(540);
			8503: out = 16'(2167);
			8504: out = 16'(680);
			8505: out = 16'(-2129);
			8506: out = 16'(-1152);
			8507: out = 16'(-334);
			8508: out = 16'(272);
			8509: out = 16'(2628);
			8510: out = 16'(4004);
			8511: out = 16'(1327);
			8512: out = 16'(-2963);
			8513: out = 16'(-310);
			8514: out = 16'(1475);
			8515: out = 16'(878);
			8516: out = 16'(-2029);
			8517: out = 16'(-3786);
			8518: out = 16'(-1287);
			8519: out = 16'(1092);
			8520: out = 16'(1);
			8521: out = 16'(-997);
			8522: out = 16'(608);
			8523: out = 16'(579);
			8524: out = 16'(334);
			8525: out = 16'(465);
			8526: out = 16'(2645);
			8527: out = 16'(1037);
			8528: out = 16'(-2801);
			8529: out = 16'(-276);
			8530: out = 16'(1823);
			8531: out = 16'(1673);
			8532: out = 16'(-226);
			8533: out = 16'(-2902);
			8534: out = 16'(-3723);
			8535: out = 16'(-4315);
			8536: out = 16'(378);
			8537: out = 16'(4789);
			8538: out = 16'(2696);
			8539: out = 16'(-2333);
			8540: out = 16'(-4834);
			8541: out = 16'(-3380);
			8542: out = 16'(-243);
			8543: out = 16'(4558);
			8544: out = 16'(2248);
			8545: out = 16'(-3211);
			8546: out = 16'(-1469);
			8547: out = 16'(700);
			8548: out = 16'(2255);
			8549: out = 16'(1750);
			8550: out = 16'(-2950);
			8551: out = 16'(-1247);
			8552: out = 16'(3694);
			8553: out = 16'(3520);
			8554: out = 16'(-381);
			8555: out = 16'(-4192);
			8556: out = 16'(-1768);
			8557: out = 16'(3097);
			8558: out = 16'(2277);
			8559: out = 16'(-1736);
			8560: out = 16'(-3069);
			8561: out = 16'(-693);
			8562: out = 16'(2440);
			8563: out = 16'(3188);
			8564: out = 16'(610);
			8565: out = 16'(7);
			8566: out = 16'(-86);
			8567: out = 16'(38);
			8568: out = 16'(608);
			8569: out = 16'(-2850);
			8570: out = 16'(-2655);
			8571: out = 16'(959);
			8572: out = 16'(2370);
			8573: out = 16'(237);
			8574: out = 16'(-2049);
			8575: out = 16'(-104);
			8576: out = 16'(4602);
			8577: out = 16'(1875);
			8578: out = 16'(-4213);
			8579: out = 16'(-4321);
			8580: out = 16'(-2348);
			8581: out = 16'(2114);
			8582: out = 16'(3528);
			8583: out = 16'(1092);
			8584: out = 16'(908);
			8585: out = 16'(3226);
			8586: out = 16'(718);
			8587: out = 16'(-3809);
			8588: out = 16'(-7114);
			8589: out = 16'(-2888);
			8590: out = 16'(1025);
			8591: out = 16'(654);
			8592: out = 16'(2909);
			8593: out = 16'(2753);
			8594: out = 16'(648);
			8595: out = 16'(-2903);
			8596: out = 16'(-2028);
			8597: out = 16'(-1863);
			8598: out = 16'(-278);
			8599: out = 16'(3828);
			8600: out = 16'(3941);
			8601: out = 16'(531);
			8602: out = 16'(-899);
			8603: out = 16'(-364);
			8604: out = 16'(2069);
			8605: out = 16'(409);
			8606: out = 16'(-1676);
			8607: out = 16'(-282);
			8608: out = 16'(-146);
			8609: out = 16'(-410);
			8610: out = 16'(2087);
			8611: out = 16'(1887);
			8612: out = 16'(-2574);
			8613: out = 16'(-4961);
			8614: out = 16'(-1260);
			8615: out = 16'(2459);
			8616: out = 16'(479);
			8617: out = 16'(-378);
			8618: out = 16'(-1158);
			8619: out = 16'(-1299);
			8620: out = 16'(-707);
			8621: out = 16'(-848);
			8622: out = 16'(629);
			8623: out = 16'(-72);
			8624: out = 16'(285);
			8625: out = 16'(-468);
			8626: out = 16'(-634);
			8627: out = 16'(1197);
			8628: out = 16'(1498);
			8629: out = 16'(3182);
			8630: out = 16'(1628);
			8631: out = 16'(-3949);
			8632: out = 16'(-4253);
			8633: out = 16'(1562);
			8634: out = 16'(3554);
			8635: out = 16'(-90);
			8636: out = 16'(-6268);
			8637: out = 16'(-2438);
			8638: out = 16'(2491);
			8639: out = 16'(4566);
			8640: out = 16'(2287);
			8641: out = 16'(1567);
			8642: out = 16'(1788);
			8643: out = 16'(581);
			8644: out = 16'(415);
			8645: out = 16'(-865);
			8646: out = 16'(-687);
			8647: out = 16'(-798);
			8648: out = 16'(-448);
			8649: out = 16'(-1803);
			8650: out = 16'(-122);
			8651: out = 16'(-612);
			8652: out = 16'(-1148);
			8653: out = 16'(-419);
			8654: out = 16'(67);
			8655: out = 16'(-1834);
			8656: out = 16'(-2141);
			8657: out = 16'(1641);
			8658: out = 16'(1946);
			8659: out = 16'(3595);
			8660: out = 16'(2323);
			8661: out = 16'(1016);
			8662: out = 16'(-135);
			8663: out = 16'(-1544);
			8664: out = 16'(-3316);
			8665: out = 16'(-2468);
			8666: out = 16'(1809);
			8667: out = 16'(862);
			8668: out = 16'(-403);
			8669: out = 16'(2062);
			8670: out = 16'(1268);
			8671: out = 16'(-1472);
			8672: out = 16'(-2778);
			8673: out = 16'(-4154);
			8674: out = 16'(-531);
			8675: out = 16'(3401);
			8676: out = 16'(4349);
			8677: out = 16'(-597);
			8678: out = 16'(-3551);
			8679: out = 16'(-1693);
			8680: out = 16'(936);
			8681: out = 16'(1422);
			8682: out = 16'(-789);
			8683: out = 16'(-1287);
			8684: out = 16'(971);
			8685: out = 16'(3340);
			8686: out = 16'(39);
			8687: out = 16'(-963);
			8688: out = 16'(-1926);
			8689: out = 16'(840);
			8690: out = 16'(723);
			8691: out = 16'(44);
			8692: out = 16'(1446);
			8693: out = 16'(2104);
			8694: out = 16'(-594);
			8695: out = 16'(-3974);
			8696: out = 16'(-3258);
			8697: out = 16'(329);
			8698: out = 16'(1426);
			8699: out = 16'(1488);
			8700: out = 16'(2821);
			8701: out = 16'(2220);
			8702: out = 16'(-1296);
			8703: out = 16'(-4379);
			8704: out = 16'(-3519);
			8705: out = 16'(-4339);
			8706: out = 16'(-2506);
			8707: out = 16'(2587);
			8708: out = 16'(2602);
			8709: out = 16'(-568);
			8710: out = 16'(-533);
			8711: out = 16'(174);
			8712: out = 16'(1638);
			8713: out = 16'(5);
			8714: out = 16'(-1421);
			8715: out = 16'(-948);
			8716: out = 16'(-608);
			8717: out = 16'(863);
			8718: out = 16'(2233);
			8719: out = 16'(281);
			8720: out = 16'(-4816);
			8721: out = 16'(-3880);
			8722: out = 16'(-1327);
			8723: out = 16'(1011);
			8724: out = 16'(4151);
			8725: out = 16'(1152);
			8726: out = 16'(-628);
			8727: out = 16'(1662);
			8728: out = 16'(2425);
			8729: out = 16'(2258);
			8730: out = 16'(168);
			8731: out = 16'(-3322);
			8732: out = 16'(-1516);
			8733: out = 16'(-1909);
			8734: out = 16'(-1374);
			8735: out = 16'(1860);
			8736: out = 16'(1860);
			8737: out = 16'(-66);
			8738: out = 16'(59);
			8739: out = 16'(3023);
			8740: out = 16'(145);
			8741: out = 16'(-4723);
			8742: out = 16'(-2601);
			8743: out = 16'(2195);
			8744: out = 16'(1872);
			8745: out = 16'(1532);
			8746: out = 16'(2439);
			8747: out = 16'(1569);
			8748: out = 16'(-2012);
			8749: out = 16'(-6298);
			8750: out = 16'(-4932);
			8751: out = 16'(1493);
			8752: out = 16'(3844);
			8753: out = 16'(-452);
			8754: out = 16'(-1609);
			8755: out = 16'(-1055);
			8756: out = 16'(1251);
			8757: out = 16'(5581);
			8758: out = 16'(2939);
			8759: out = 16'(-1599);
			8760: out = 16'(-3443);
			8761: out = 16'(-2035);
			8762: out = 16'(-1510);
			8763: out = 16'(456);
			8764: out = 16'(1225);
			8765: out = 16'(788);
			8766: out = 16'(1094);
			8767: out = 16'(1457);
			8768: out = 16'(1365);
			8769: out = 16'(-142);
			8770: out = 16'(-139);
			8771: out = 16'(302);
			8772: out = 16'(2304);
			8773: out = 16'(2423);
			8774: out = 16'(1532);
			8775: out = 16'(-313);
			8776: out = 16'(-469);
			8777: out = 16'(-1891);
			8778: out = 16'(-3396);
			8779: out = 16'(-1920);
			8780: out = 16'(-432);
			8781: out = 16'(1);
			8782: out = 16'(1838);
			8783: out = 16'(213);
			8784: out = 16'(-2553);
			8785: out = 16'(-1723);
			8786: out = 16'(-1347);
			8787: out = 16'(1188);
			8788: out = 16'(1434);
			8789: out = 16'(1189);
			8790: out = 16'(996);
			8791: out = 16'(2240);
			8792: out = 16'(1569);
			8793: out = 16'(-2476);
			8794: out = 16'(-3771);
			8795: out = 16'(-1876);
			8796: out = 16'(2314);
			8797: out = 16'(2950);
			8798: out = 16'(-431);
			8799: out = 16'(-2001);
			8800: out = 16'(-1259);
			8801: out = 16'(-349);
			8802: out = 16'(1150);
			8803: out = 16'(1519);
			8804: out = 16'(-168);
			8805: out = 16'(-5);
			8806: out = 16'(89);
			8807: out = 16'(-1099);
			8808: out = 16'(-2646);
			8809: out = 16'(-5760);
			8810: out = 16'(-1065);
			8811: out = 16'(3566);
			8812: out = 16'(3389);
			8813: out = 16'(2197);
			8814: out = 16'(1331);
			8815: out = 16'(-940);
			8816: out = 16'(-2110);
			8817: out = 16'(-2829);
			8818: out = 16'(-3016);
			8819: out = 16'(-628);
			8820: out = 16'(1125);
			8821: out = 16'(2616);
			8822: out = 16'(2572);
			8823: out = 16'(838);
			8824: out = 16'(958);
			8825: out = 16'(2158);
			8826: out = 16'(1490);
			8827: out = 16'(-521);
			8828: out = 16'(-2297);
			8829: out = 16'(199);
			8830: out = 16'(3762);
			8831: out = 16'(2987);
			8832: out = 16'(-3511);
			8833: out = 16'(-3412);
			8834: out = 16'(173);
			8835: out = 16'(2313);
			8836: out = 16'(256);
			8837: out = 16'(-1580);
			8838: out = 16'(1508);
			8839: out = 16'(3164);
			8840: out = 16'(1913);
			8841: out = 16'(440);
			8842: out = 16'(70);
			8843: out = 16'(399);
			8844: out = 16'(-797);
			8845: out = 16'(-1057);
			8846: out = 16'(-46);
			8847: out = 16'(465);
			8848: out = 16'(-2230);
			8849: out = 16'(-1055);
			8850: out = 16'(276);
			8851: out = 16'(-1774);
			8852: out = 16'(-1171);
			8853: out = 16'(583);
			8854: out = 16'(1254);
			8855: out = 16'(2010);
			8856: out = 16'(2144);
			8857: out = 16'(-550);
			8858: out = 16'(-2423);
			8859: out = 16'(-2643);
			8860: out = 16'(-597);
			8861: out = 16'(1115);
			8862: out = 16'(1047);
			8863: out = 16'(1675);
			8864: out = 16'(2122);
			8865: out = 16'(1010);
			8866: out = 16'(-1635);
			8867: out = 16'(-2683);
			8868: out = 16'(-824);
			8869: out = 16'(-1549);
			8870: out = 16'(-552);
			8871: out = 16'(2779);
			8872: out = 16'(2549);
			8873: out = 16'(-4079);
			8874: out = 16'(-7217);
			8875: out = 16'(-4285);
			8876: out = 16'(-459);
			8877: out = 16'(5213);
			8878: out = 16'(4897);
			8879: out = 16'(-1559);
			8880: out = 16'(-6055);
			8881: out = 16'(-4152);
			8882: out = 16'(-454);
			8883: out = 16'(2345);
			8884: out = 16'(4067);
			8885: out = 16'(1670);
			8886: out = 16'(-4455);
			8887: out = 16'(-5679);
			8888: out = 16'(-2471);
			8889: out = 16'(2666);
			8890: out = 16'(6213);
			8891: out = 16'(2773);
			8892: out = 16'(-1131);
			8893: out = 16'(-3626);
			8894: out = 16'(-331);
			8895: out = 16'(3890);
			8896: out = 16'(3618);
			8897: out = 16'(1332);
			8898: out = 16'(-1275);
			8899: out = 16'(-2678);
			8900: out = 16'(-944);
			8901: out = 16'(2646);
			8902: out = 16'(2266);
			8903: out = 16'(-645);
			8904: out = 16'(529);
			8905: out = 16'(442);
			8906: out = 16'(-1397);
			8907: out = 16'(-2174);
			8908: out = 16'(-3856);
			8909: out = 16'(646);
			8910: out = 16'(4490);
			8911: out = 16'(2592);
			8912: out = 16'(-1120);
			8913: out = 16'(-1104);
			8914: out = 16'(663);
			8915: out = 16'(1724);
			8916: out = 16'(869);
			8917: out = 16'(1536);
			8918: out = 16'(-578);
			8919: out = 16'(-1069);
			8920: out = 16'(396);
			8921: out = 16'(-343);
			8922: out = 16'(-1344);
			8923: out = 16'(297);
			8924: out = 16'(243);
			8925: out = 16'(395);
			8926: out = 16'(1589);
			8927: out = 16'(2227);
			8928: out = 16'(1445);
			8929: out = 16'(-191);
			8930: out = 16'(-999);
			8931: out = 16'(-220);
			8932: out = 16'(-1667);
			8933: out = 16'(-1767);
			8934: out = 16'(-2128);
			8935: out = 16'(-2738);
			8936: out = 16'(1943);
			8937: out = 16'(4481);
			8938: out = 16'(848);
			8939: out = 16'(-2370);
			8940: out = 16'(-1106);
			8941: out = 16'(467);
			8942: out = 16'(2351);
			8943: out = 16'(2463);
			8944: out = 16'(569);
			8945: out = 16'(-103);
			8946: out = 16'(307);
			8947: out = 16'(-66);
			8948: out = 16'(-594);
			8949: out = 16'(-3030);
			8950: out = 16'(-2606);
			8951: out = 16'(820);
			8952: out = 16'(2551);
			8953: out = 16'(-1588);
			8954: out = 16'(-3809);
			8955: out = 16'(-1624);
			8956: out = 16'(796);
			8957: out = 16'(2187);
			8958: out = 16'(2387);
			8959: out = 16'(360);
			8960: out = 16'(-2725);
			8961: out = 16'(-814);
			8962: out = 16'(886);
			8963: out = 16'(-65);
			8964: out = 16'(-1909);
			8965: out = 16'(-3382);
			8966: out = 16'(259);
			8967: out = 16'(4523);
			8968: out = 16'(2991);
			8969: out = 16'(795);
			8970: out = 16'(-223);
			8971: out = 16'(1167);
			8972: out = 16'(-418);
			8973: out = 16'(-1698);
			8974: out = 16'(-824);
			8975: out = 16'(2280);
			8976: out = 16'(2899);
			8977: out = 16'(-833);
			8978: out = 16'(-1314);
			8979: out = 16'(-496);
			8980: out = 16'(-905);
			8981: out = 16'(538);
			8982: out = 16'(1363);
			8983: out = 16'(-1662);
			8984: out = 16'(-748);
			8985: out = 16'(-214);
			8986: out = 16'(926);
			8987: out = 16'(3287);
			8988: out = 16'(1651);
			8989: out = 16'(-1577);
			8990: out = 16'(-1665);
			8991: out = 16'(-896);
			8992: out = 16'(-2102);
			8993: out = 16'(-5109);
			8994: out = 16'(-732);
			8995: out = 16'(2184);
			8996: out = 16'(2684);
			8997: out = 16'(2207);
			8998: out = 16'(1975);
			8999: out = 16'(1742);
			9000: out = 16'(265);
			9001: out = 16'(-1289);
			9002: out = 16'(-2037);
			9003: out = 16'(-324);
			9004: out = 16'(2190);
			9005: out = 16'(1025);
			9006: out = 16'(-2818);
			9007: out = 16'(-2166);
			9008: out = 16'(1882);
			9009: out = 16'(2941);
			9010: out = 16'(-2121);
			9011: out = 16'(-4937);
			9012: out = 16'(-2789);
			9013: out = 16'(-1254);
			9014: out = 16'(1942);
			9015: out = 16'(2715);
			9016: out = 16'(-46);
			9017: out = 16'(-1958);
			9018: out = 16'(107);
			9019: out = 16'(522);
			9020: out = 16'(1417);
			9021: out = 16'(1769);
			9022: out = 16'(396);
			9023: out = 16'(379);
			9024: out = 16'(904);
			9025: out = 16'(754);
			9026: out = 16'(810);
			9027: out = 16'(173);
			9028: out = 16'(1311);
			9029: out = 16'(-308);
			9030: out = 16'(-1792);
			9031: out = 16'(-628);
			9032: out = 16'(607);
			9033: out = 16'(-2102);
			9034: out = 16'(-2685);
			9035: out = 16'(378);
			9036: out = 16'(-574);
			9037: out = 16'(196);
			9038: out = 16'(2967);
			9039: out = 16'(815);
			9040: out = 16'(-4645);
			9041: out = 16'(-4672);
			9042: out = 16'(-1423);
			9043: out = 16'(2257);
			9044: out = 16'(3519);
			9045: out = 16'(-575);
			9046: out = 16'(-5503);
			9047: out = 16'(-2022);
			9048: out = 16'(3312);
			9049: out = 16'(3633);
			9050: out = 16'(2051);
			9051: out = 16'(1351);
			9052: out = 16'(1082);
			9053: out = 16'(497);
			9054: out = 16'(-1984);
			9055: out = 16'(-2642);
			9056: out = 16'(597);
			9057: out = 16'(-243);
			9058: out = 16'(-974);
			9059: out = 16'(-537);
			9060: out = 16'(-960);
			9061: out = 16'(865);
			9062: out = 16'(1011);
			9063: out = 16'(-1137);
			9064: out = 16'(-767);
			9065: out = 16'(293);
			9066: out = 16'(2164);
			9067: out = 16'(1928);
			9068: out = 16'(675);
			9069: out = 16'(503);
			9070: out = 16'(-415);
			9071: out = 16'(-3166);
			9072: out = 16'(-2036);
			9073: out = 16'(-316);
			9074: out = 16'(1167);
			9075: out = 16'(1817);
			9076: out = 16'(-792);
			9077: out = 16'(-3418);
			9078: out = 16'(-2087);
			9079: out = 16'(2215);
			9080: out = 16'(3448);
			9081: out = 16'(1013);
			9082: out = 16'(-1131);
			9083: out = 16'(-354);
			9084: out = 16'(2357);
			9085: out = 16'(-873);
			9086: out = 16'(-1714);
			9087: out = 16'(-470);
			9088: out = 16'(-266);
			9089: out = 16'(689);
			9090: out = 16'(3046);
			9091: out = 16'(991);
			9092: out = 16'(-1929);
			9093: out = 16'(-2959);
			9094: out = 16'(-233);
			9095: out = 16'(3542);
			9096: out = 16'(862);
			9097: out = 16'(-2446);
			9098: out = 16'(-563);
			9099: out = 16'(1054);
			9100: out = 16'(-1347);
			9101: out = 16'(-5200);
			9102: out = 16'(-3028);
			9103: out = 16'(-121);
			9104: out = 16'(79);
			9105: out = 16'(3652);
			9106: out = 16'(4363);
			9107: out = 16'(-324);
			9108: out = 16'(-4597);
			9109: out = 16'(-3330);
			9110: out = 16'(256);
			9111: out = 16'(859);
			9112: out = 16'(-70);
			9113: out = 16'(1445);
			9114: out = 16'(-825);
			9115: out = 16'(-1323);
			9116: out = 16'(597);
			9117: out = 16'(1552);
			9118: out = 16'(2903);
			9119: out = 16'(1846);
			9120: out = 16'(-2237);
			9121: out = 16'(-3886);
			9122: out = 16'(-2078);
			9123: out = 16'(1001);
			9124: out = 16'(4557);
			9125: out = 16'(2962);
			9126: out = 16'(-1318);
			9127: out = 16'(-2237);
			9128: out = 16'(-675);
			9129: out = 16'(1029);
			9130: out = 16'(-2249);
			9131: out = 16'(-569);
			9132: out = 16'(2322);
			9133: out = 16'(2091);
			9134: out = 16'(-782);
			9135: out = 16'(-1207);
			9136: out = 16'(1658);
			9137: out = 16'(2119);
			9138: out = 16'(1059);
			9139: out = 16'(-474);
			9140: out = 16'(-971);
			9141: out = 16'(-190);
			9142: out = 16'(-491);
			9143: out = 16'(-881);
			9144: out = 16'(897);
			9145: out = 16'(2519);
			9146: out = 16'(-124);
			9147: out = 16'(-3652);
			9148: out = 16'(-2710);
			9149: out = 16'(-354);
			9150: out = 16'(1877);
			9151: out = 16'(-310);
			9152: out = 16'(-251);
			9153: out = 16'(634);
			9154: out = 16'(-283);
			9155: out = 16'(-3202);
			9156: out = 16'(-493);
			9157: out = 16'(1696);
			9158: out = 16'(-221);
			9159: out = 16'(656);
			9160: out = 16'(1171);
			9161: out = 16'(-257);
			9162: out = 16'(1142);
			9163: out = 16'(1850);
			9164: out = 16'(508);
			9165: out = 16'(-2002);
			9166: out = 16'(-1649);
			9167: out = 16'(-73);
			9168: out = 16'(-231);
			9169: out = 16'(-348);
			9170: out = 16'(189);
			9171: out = 16'(1725);
			9172: out = 16'(-393);
			9173: out = 16'(1133);
			9174: out = 16'(3141);
			9175: out = 16'(1964);
			9176: out = 16'(-1459);
			9177: out = 16'(-2325);
			9178: out = 16'(-1878);
			9179: out = 16'(-1400);
			9180: out = 16'(76);
			9181: out = 16'(-1200);
			9182: out = 16'(-1189);
			9183: out = 16'(2095);
			9184: out = 16'(3782);
			9185: out = 16'(1100);
			9186: out = 16'(-3233);
			9187: out = 16'(-2928);
			9188: out = 16'(1526);
			9189: out = 16'(4710);
			9190: out = 16'(1449);
			9191: out = 16'(-1871);
			9192: out = 16'(-684);
			9193: out = 16'(2904);
			9194: out = 16'(1950);
			9195: out = 16'(-972);
			9196: out = 16'(-1837);
			9197: out = 16'(78);
			9198: out = 16'(604);
			9199: out = 16'(1369);
			9200: out = 16'(936);
			9201: out = 16'(186);
			9202: out = 16'(-3630);
			9203: out = 16'(-3606);
			9204: out = 16'(-616);
			9205: out = 16'(-947);
			9206: out = 16'(1039);
			9207: out = 16'(3024);
			9208: out = 16'(473);
			9209: out = 16'(-2612);
			9210: out = 16'(-2799);
			9211: out = 16'(-1827);
			9212: out = 16'(2234);
			9213: out = 16'(3207);
			9214: out = 16'(1942);
			9215: out = 16'(-1410);
			9216: out = 16'(-1388);
			9217: out = 16'(-513);
			9218: out = 16'(427);
			9219: out = 16'(494);
			9220: out = 16'(-830);
			9221: out = 16'(696);
			9222: out = 16'(697);
			9223: out = 16'(2639);
			9224: out = 16'(2222);
			9225: out = 16'(1511);
			9226: out = 16'(340);
			9227: out = 16'(-555);
			9228: out = 16'(844);
			9229: out = 16'(1117);
			9230: out = 16'(38);
			9231: out = 16'(-1343);
			9232: out = 16'(-2075);
			9233: out = 16'(-1296);
			9234: out = 16'(-750);
			9235: out = 16'(-3136);
			9236: out = 16'(-3696);
			9237: out = 16'(-2784);
			9238: out = 16'(-1578);
			9239: out = 16'(2082);
			9240: out = 16'(4944);
			9241: out = 16'(2723);
			9242: out = 16'(-2469);
			9243: out = 16'(-4303);
			9244: out = 16'(-1478);
			9245: out = 16'(1907);
			9246: out = 16'(2459);
			9247: out = 16'(2741);
			9248: out = 16'(1318);
			9249: out = 16'(-2943);
			9250: out = 16'(-4606);
			9251: out = 16'(-2710);
			9252: out = 16'(875);
			9253: out = 16'(2713);
			9254: out = 16'(2254);
			9255: out = 16'(-775);
			9256: out = 16'(-2598);
			9257: out = 16'(-1964);
			9258: out = 16'(976);
			9259: out = 16'(4341);
			9260: out = 16'(4229);
			9261: out = 16'(790);
			9262: out = 16'(-1616);
			9263: out = 16'(-795);
			9264: out = 16'(-1368);
			9265: out = 16'(-2265);
			9266: out = 16'(-1663);
			9267: out = 16'(221);
			9268: out = 16'(663);
			9269: out = 16'(2242);
			9270: out = 16'(2998);
			9271: out = 16'(2647);
			9272: out = 16'(1117);
			9273: out = 16'(-172);
			9274: out = 16'(-1212);
			9275: out = 16'(-1308);
			9276: out = 16'(-1309);
			9277: out = 16'(-1105);
			9278: out = 16'(-675);
			9279: out = 16'(131);
			9280: out = 16'(668);
			9281: out = 16'(463);
			9282: out = 16'(-1295);
			9283: out = 16'(-2314);
			9284: out = 16'(-1296);
			9285: out = 16'(244);
			9286: out = 16'(2801);
			9287: out = 16'(1757);
			9288: out = 16'(-538);
			9289: out = 16'(-2229);
			9290: out = 16'(-906);
			9291: out = 16'(1603);
			9292: out = 16'(-332);
			9293: out = 16'(287);
			9294: out = 16'(790);
			9295: out = 16'(720);
			9296: out = 16'(2479);
			9297: out = 16'(3094);
			9298: out = 16'(1505);
			9299: out = 16'(-781);
			9300: out = 16'(-3111);
			9301: out = 16'(-2050);
			9302: out = 16'(-1355);
			9303: out = 16'(-1619);
			9304: out = 16'(-757);
			9305: out = 16'(-4);
			9306: out = 16'(-10);
			9307: out = 16'(1176);
			9308: out = 16'(2427);
			9309: out = 16'(638);
			9310: out = 16'(-2039);
			9311: out = 16'(-1667);
			9312: out = 16'(-1598);
			9313: out = 16'(-751);
			9314: out = 16'(742);
			9315: out = 16'(1738);
			9316: out = 16'(1798);
			9317: out = 16'(1917);
			9318: out = 16'(543);
			9319: out = 16'(374);
			9320: out = 16'(914);
			9321: out = 16'(452);
			9322: out = 16'(-456);
			9323: out = 16'(-210);
			9324: out = 16'(2288);
			9325: out = 16'(1154);
			9326: out = 16'(-1784);
			9327: out = 16'(-2615);
			9328: out = 16'(-970);
			9329: out = 16'(697);
			9330: out = 16'(741);
			9331: out = 16'(549);
			9332: out = 16'(-1090);
			9333: out = 16'(-1116);
			9334: out = 16'(478);
			9335: out = 16'(1297);
			9336: out = 16'(-2541);
			9337: out = 16'(-2511);
			9338: out = 16'(-395);
			9339: out = 16'(1717);
			9340: out = 16'(1289);
			9341: out = 16'(331);
			9342: out = 16'(1281);
			9343: out = 16'(1216);
			9344: out = 16'(571);
			9345: out = 16'(-2579);
			9346: out = 16'(-2776);
			9347: out = 16'(-1781);
			9348: out = 16'(533);
			9349: out = 16'(2867);
			9350: out = 16'(1211);
			9351: out = 16'(453);
			9352: out = 16'(438);
			9353: out = 16'(389);
			9354: out = 16'(-1441);
			9355: out = 16'(-1448);
			9356: out = 16'(904);
			9357: out = 16'(267);
			9358: out = 16'(509);
			9359: out = 16'(1614);
			9360: out = 16'(1287);
			9361: out = 16'(-121);
			9362: out = 16'(-1749);
			9363: out = 16'(-1051);
			9364: out = 16'(-1688);
			9365: out = 16'(-1908);
			9366: out = 16'(118);
			9367: out = 16'(1494);
			9368: out = 16'(22);
			9369: out = 16'(-1323);
			9370: out = 16'(-1698);
			9371: out = 16'(-322);
			9372: out = 16'(-678);
			9373: out = 16'(-786);
			9374: out = 16'(2292);
			9375: out = 16'(1190);
			9376: out = 16'(263);
			9377: out = 16'(1786);
			9378: out = 16'(1346);
			9379: out = 16'(-2435);
			9380: out = 16'(-3420);
			9381: out = 16'(-2182);
			9382: out = 16'(498);
			9383: out = 16'(127);
			9384: out = 16'(-778);
			9385: out = 16'(-117);
			9386: out = 16'(769);
			9387: out = 16'(2873);
			9388: out = 16'(2613);
			9389: out = 16'(-185);
			9390: out = 16'(-3795);
			9391: out = 16'(-2011);
			9392: out = 16'(-1915);
			9393: out = 16'(-1180);
			9394: out = 16'(2830);
			9395: out = 16'(3163);
			9396: out = 16'(-633);
			9397: out = 16'(-1734);
			9398: out = 16'(430);
			9399: out = 16'(2369);
			9400: out = 16'(833);
			9401: out = 16'(-1746);
			9402: out = 16'(-2208);
			9403: out = 16'(-1407);
			9404: out = 16'(1266);
			9405: out = 16'(2654);
			9406: out = 16'(-954);
			9407: out = 16'(-5464);
			9408: out = 16'(-3038);
			9409: out = 16'(2051);
			9410: out = 16'(3125);
			9411: out = 16'(2538);
			9412: out = 16'(-7);
			9413: out = 16'(-2003);
			9414: out = 16'(-222);
			9415: out = 16'(184);
			9416: out = 16'(2274);
			9417: out = 16'(1823);
			9418: out = 16'(-430);
			9419: out = 16'(-570);
			9420: out = 16'(-595);
			9421: out = 16'(95);
			9422: out = 16'(-345);
			9423: out = 16'(-1639);
			9424: out = 16'(713);
			9425: out = 16'(721);
			9426: out = 16'(445);
			9427: out = 16'(-261);
			9428: out = 16'(-503);
			9429: out = 16'(682);
			9430: out = 16'(2555);
			9431: out = 16'(2160);
			9432: out = 16'(223);
			9433: out = 16'(-527);
			9434: out = 16'(-255);
			9435: out = 16'(481);
			9436: out = 16'(-990);
			9437: out = 16'(-1405);
			9438: out = 16'(-1322);
			9439: out = 16'(-148);
			9440: out = 16'(-1219);
			9441: out = 16'(-704);
			9442: out = 16'(-2021);
			9443: out = 16'(-1651);
			9444: out = 16'(704);
			9445: out = 16'(2294);
			9446: out = 16'(2511);
			9447: out = 16'(-355);
			9448: out = 16'(-361);
			9449: out = 16'(-587);
			9450: out = 16'(-40);
			9451: out = 16'(469);
			9452: out = 16'(-118);
			9453: out = 16'(1587);
			9454: out = 16'(2392);
			9455: out = 16'(-1065);
			9456: out = 16'(-3197);
			9457: out = 16'(-3074);
			9458: out = 16'(-1688);
			9459: out = 16'(1326);
			9460: out = 16'(2399);
			9461: out = 16'(219);
			9462: out = 16'(-689);
			9463: out = 16'(-1259);
			9464: out = 16'(233);
			9465: out = 16'(1521);
			9466: out = 16'(-1272);
			9467: out = 16'(-1357);
			9468: out = 16'(1260);
			9469: out = 16'(1053);
			9470: out = 16'(-2044);
			9471: out = 16'(-2323);
			9472: out = 16'(-949);
			9473: out = 16'(-159);
			9474: out = 16'(2050);
			9475: out = 16'(637);
			9476: out = 16'(-1987);
			9477: out = 16'(-373);
			9478: out = 16'(2338);
			9479: out = 16'(3386);
			9480: out = 16'(-146);
			9481: out = 16'(348);
			9482: out = 16'(2271);
			9483: out = 16'(2128);
			9484: out = 16'(-2348);
			9485: out = 16'(-3352);
			9486: out = 16'(-1179);
			9487: out = 16'(-236);
			9488: out = 16'(234);
			9489: out = 16'(562);
			9490: out = 16'(1290);
			9491: out = 16'(-105);
			9492: out = 16'(-798);
			9493: out = 16'(-209);
			9494: out = 16'(285);
			9495: out = 16'(1143);
			9496: out = 16'(665);
			9497: out = 16'(-746);
			9498: out = 16'(-1393);
			9499: out = 16'(-1921);
			9500: out = 16'(-1727);
			9501: out = 16'(1974);
			9502: out = 16'(3449);
			9503: out = 16'(-1004);
			9504: out = 16'(-3560);
			9505: out = 16'(-1709);
			9506: out = 16'(515);
			9507: out = 16'(3795);
			9508: out = 16'(2770);
			9509: out = 16'(-491);
			9510: out = 16'(-707);
			9511: out = 16'(-599);
			9512: out = 16'(757);
			9513: out = 16'(-17);
			9514: out = 16'(-1139);
			9515: out = 16'(615);
			9516: out = 16'(973);
			9517: out = 16'(134);
			9518: out = 16'(-1218);
			9519: out = 16'(-2425);
			9520: out = 16'(-1732);
			9521: out = 16'(-306);
			9522: out = 16'(-240);
			9523: out = 16'(1356);
			9524: out = 16'(1082);
			9525: out = 16'(-237);
			9526: out = 16'(-2463);
			9527: out = 16'(-3441);
			9528: out = 16'(772);
			9529: out = 16'(3011);
			9530: out = 16'(2327);
			9531: out = 16'(1166);
			9532: out = 16'(589);
			9533: out = 16'(-815);
			9534: out = 16'(-2107);
			9535: out = 16'(-1580);
			9536: out = 16'(-683);
			9537: out = 16'(-805);
			9538: out = 16'(1216);
			9539: out = 16'(611);
			9540: out = 16'(-614);
			9541: out = 16'(1932);
			9542: out = 16'(2255);
			9543: out = 16'(1168);
			9544: out = 16'(-76);
			9545: out = 16'(13);
			9546: out = 16'(-898);
			9547: out = 16'(-1280);
			9548: out = 16'(1844);
			9549: out = 16'(2146);
			9550: out = 16'(-45);
			9551: out = 16'(92);
			9552: out = 16'(-419);
			9553: out = 16'(351);
			9554: out = 16'(698);
			9555: out = 16'(-710);
			9556: out = 16'(243);
			9557: out = 16'(2375);
			9558: out = 16'(573);
			9559: out = 16'(-3189);
			9560: out = 16'(-4558);
			9561: out = 16'(-699);
			9562: out = 16'(1071);
			9563: out = 16'(-520);
			9564: out = 16'(1387);
			9565: out = 16'(2669);
			9566: out = 16'(407);
			9567: out = 16'(-4407);
			9568: out = 16'(-4732);
			9569: out = 16'(-1409);
			9570: out = 16'(1522);
			9571: out = 16'(3146);
			9572: out = 16'(2441);
			9573: out = 16'(-604);
			9574: out = 16'(-3817);
			9575: out = 16'(-2143);
			9576: out = 16'(240);
			9577: out = 16'(3468);
			9578: out = 16'(2009);
			9579: out = 16'(-2113);
			9580: out = 16'(-2473);
			9581: out = 16'(322);
			9582: out = 16'(3853);
			9583: out = 16'(1981);
			9584: out = 16'(-876);
			9585: out = 16'(107);
			9586: out = 16'(1122);
			9587: out = 16'(1169);
			9588: out = 16'(1632);
			9589: out = 16'(-183);
			9590: out = 16'(-2036);
			9591: out = 16'(-3983);
			9592: out = 16'(-2704);
			9593: out = 16'(1556);
			9594: out = 16'(1821);
			9595: out = 16'(-1327);
			9596: out = 16'(-397);
			9597: out = 16'(315);
			9598: out = 16'(-1490);
			9599: out = 16'(-656);
			9600: out = 16'(498);
			9601: out = 16'(1780);
			9602: out = 16'(1261);
			9603: out = 16'(-884);
			9604: out = 16'(-1349);
			9605: out = 16'(-165);
			9606: out = 16'(947);
			9607: out = 16'(130);
			9608: out = 16'(-572);
			9609: out = 16'(-70);
			9610: out = 16'(1998);
			9611: out = 16'(3929);
			9612: out = 16'(1782);
			9613: out = 16'(-2082);
			9614: out = 16'(-3020);
			9615: out = 16'(-1100);
			9616: out = 16'(729);
			9617: out = 16'(2414);
			9618: out = 16'(1005);
			9619: out = 16'(-318);
			9620: out = 16'(561);
			9621: out = 16'(-144);
			9622: out = 16'(-2440);
			9623: out = 16'(-2856);
			9624: out = 16'(-2417);
			9625: out = 16'(499);
			9626: out = 16'(2550);
			9627: out = 16'(2459);
			9628: out = 16'(-7);
			9629: out = 16'(-1008);
			9630: out = 16'(-1656);
			9631: out = 16'(796);
			9632: out = 16'(2814);
			9633: out = 16'(1191);
			9634: out = 16'(-2004);
			9635: out = 16'(-1900);
			9636: out = 16'(166);
			9637: out = 16'(1356);
			9638: out = 16'(-1017);
			9639: out = 16'(-2661);
			9640: out = 16'(-539);
			9641: out = 16'(1248);
			9642: out = 16'(2347);
			9643: out = 16'(1242);
			9644: out = 16'(-2014);
			9645: out = 16'(-1914);
			9646: out = 16'(341);
			9647: out = 16'(1823);
			9648: out = 16'(884);
			9649: out = 16'(-1010);
			9650: out = 16'(128);
			9651: out = 16'(931);
			9652: out = 16'(-1014);
			9653: out = 16'(-1126);
			9654: out = 16'(178);
			9655: out = 16'(381);
			9656: out = 16'(-763);
			9657: out = 16'(-215);
			9658: out = 16'(1030);
			9659: out = 16'(719);
			9660: out = 16'(-216);
			9661: out = 16'(-3185);
			9662: out = 16'(-4360);
			9663: out = 16'(364);
			9664: out = 16'(4232);
			9665: out = 16'(2808);
			9666: out = 16'(-1176);
			9667: out = 16'(-2419);
			9668: out = 16'(650);
			9669: out = 16'(3373);
			9670: out = 16'(1770);
			9671: out = 16'(36);
			9672: out = 16'(1035);
			9673: out = 16'(2172);
			9674: out = 16'(446);
			9675: out = 16'(-2986);
			9676: out = 16'(-2252);
			9677: out = 16'(297);
			9678: out = 16'(30);
			9679: out = 16'(-906);
			9680: out = 16'(-159);
			9681: out = 16'(616);
			9682: out = 16'(1063);
			9683: out = 16'(1187);
			9684: out = 16'(1023);
			9685: out = 16'(136);
			9686: out = 16'(665);
			9687: out = 16'(659);
			9688: out = 16'(1067);
			9689: out = 16'(699);
			9690: out = 16'(-870);
			9691: out = 16'(-522);
			9692: out = 16'(341);
			9693: out = 16'(-496);
			9694: out = 16'(-2233);
			9695: out = 16'(-2664);
			9696: out = 16'(-796);
			9697: out = 16'(791);
			9698: out = 16'(1211);
			9699: out = 16'(-1464);
			9700: out = 16'(-2143);
			9701: out = 16'(415);
			9702: out = 16'(816);
			9703: out = 16'(68);
			9704: out = 16'(193);
			9705: out = 16'(1728);
			9706: out = 16'(1306);
			9707: out = 16'(34);
			9708: out = 16'(288);
			9709: out = 16'(1106);
			9710: out = 16'(1100);
			9711: out = 16'(-1347);
			9712: out = 16'(-1466);
			9713: out = 16'(-536);
			9714: out = 16'(1485);
			9715: out = 16'(547);
			9716: out = 16'(-1652);
			9717: out = 16'(-2248);
			9718: out = 16'(226);
			9719: out = 16'(2295);
			9720: out = 16'(402);
			9721: out = 16'(-603);
			9722: out = 16'(615);
			9723: out = 16'(2071);
			9724: out = 16'(-47);
			9725: out = 16'(-2426);
			9726: out = 16'(-1448);
			9727: out = 16'(-410);
			9728: out = 16'(-1617);
			9729: out = 16'(-2124);
			9730: out = 16'(-223);
			9731: out = 16'(-413);
			9732: out = 16'(395);
			9733: out = 16'(636);
			9734: out = 16'(-398);
			9735: out = 16'(-2843);
			9736: out = 16'(-2049);
			9737: out = 16'(1388);
			9738: out = 16'(1614);
			9739: out = 16'(1900);
			9740: out = 16'(2403);
			9741: out = 16'(1309);
			9742: out = 16'(-2423);
			9743: out = 16'(-5126);
			9744: out = 16'(-4598);
			9745: out = 16'(-434);
			9746: out = 16'(2992);
			9747: out = 16'(1575);
			9748: out = 16'(-255);
			9749: out = 16'(321);
			9750: out = 16'(1370);
			9751: out = 16'(1979);
			9752: out = 16'(365);
			9753: out = 16'(1082);
			9754: out = 16'(2811);
			9755: out = 16'(1272);
			9756: out = 16'(-2009);
			9757: out = 16'(-2824);
			9758: out = 16'(-360);
			9759: out = 16'(-206);
			9760: out = 16'(-3631);
			9761: out = 16'(-2126);
			9762: out = 16'(885);
			9763: out = 16'(836);
			9764: out = 16'(1600);
			9765: out = 16'(3206);
			9766: out = 16'(1306);
			9767: out = 16'(-2440);
			9768: out = 16'(-5161);
			9769: out = 16'(-2578);
			9770: out = 16'(1330);
			9771: out = 16'(2092);
			9772: out = 16'(803);
			9773: out = 16'(-984);
			9774: out = 16'(-1772);
			9775: out = 16'(-592);
			9776: out = 16'(2009);
			9777: out = 16'(1819);
			9778: out = 16'(128);
			9779: out = 16'(-1248);
			9780: out = 16'(-2498);
			9781: out = 16'(-920);
			9782: out = 16'(307);
			9783: out = 16'(1687);
			9784: out = 16'(2673);
			9785: out = 16'(311);
			9786: out = 16'(-2338);
			9787: out = 16'(-3006);
			9788: out = 16'(-1193);
			9789: out = 16'(2842);
			9790: out = 16'(2841);
			9791: out = 16'(70);
			9792: out = 16'(-1865);
			9793: out = 16'(-249);
			9794: out = 16'(2276);
			9795: out = 16'(2254);
			9796: out = 16'(-688);
			9797: out = 16'(-769);
			9798: out = 16'(-502);
			9799: out = 16'(-503);
			9800: out = 16'(645);
			9801: out = 16'(497);
			9802: out = 16'(-1181);
			9803: out = 16'(-1536);
			9804: out = 16'(-375);
			9805: out = 16'(-303);
			9806: out = 16'(-1349);
			9807: out = 16'(222);
			9808: out = 16'(1146);
			9809: out = 16'(1863);
			9810: out = 16'(467);
			9811: out = 16'(262);
			9812: out = 16'(1361);
			9813: out = 16'(1122);
			9814: out = 16'(-957);
			9815: out = 16'(-2177);
			9816: out = 16'(-887);
			9817: out = 16'(120);
			9818: out = 16'(358);
			9819: out = 16'(640);
			9820: out = 16'(1608);
			9821: out = 16'(311);
			9822: out = 16'(-2048);
			9823: out = 16'(-2146);
			9824: out = 16'(-1348);
			9825: out = 16'(764);
			9826: out = 16'(1987);
			9827: out = 16'(-121);
			9828: out = 16'(-2121);
			9829: out = 16'(-1829);
			9830: out = 16'(653);
			9831: out = 16'(2113);
			9832: out = 16'(1372);
			9833: out = 16'(542);
			9834: out = 16'(-1896);
			9835: out = 16'(-3224);
			9836: out = 16'(-2182);
			9837: out = 16'(1081);
			9838: out = 16'(3592);
			9839: out = 16'(176);
			9840: out = 16'(-1310);
			9841: out = 16'(1251);
			9842: out = 16'(1562);
			9843: out = 16'(1229);
			9844: out = 16'(-213);
			9845: out = 16'(-580);
			9846: out = 16'(-1367);
			9847: out = 16'(-2422);
			9848: out = 16'(-122);
			9849: out = 16'(694);
			9850: out = 16'(-39);
			9851: out = 16'(580);
			9852: out = 16'(518);
			9853: out = 16'(-637);
			9854: out = 16'(-973);
			9855: out = 16'(364);
			9856: out = 16'(1591);
			9857: out = 16'(862);
			9858: out = 16'(-771);
			9859: out = 16'(-1175);
			9860: out = 16'(1631);
			9861: out = 16'(2835);
			9862: out = 16'(-784);
			9863: out = 16'(-2966);
			9864: out = 16'(-1734);
			9865: out = 16'(680);
			9866: out = 16'(1168);
			9867: out = 16'(1659);
			9868: out = 16'(1049);
			9869: out = 16'(430);
			9870: out = 16'(-130);
			9871: out = 16'(130);
			9872: out = 16'(-82);
			9873: out = 16'(-1567);
			9874: out = 16'(-1370);
			9875: out = 16'(-514);
			9876: out = 16'(298);
			9877: out = 16'(417);
			9878: out = 16'(633);
			9879: out = 16'(-323);
			9880: out = 16'(114);
			9881: out = 16'(1013);
			9882: out = 16'(696);
			9883: out = 16'(-247);
			9884: out = 16'(-205);
			9885: out = 16'(-750);
			9886: out = 16'(-1127);
			9887: out = 16'(-847);
			9888: out = 16'(-1318);
			9889: out = 16'(1174);
			9890: out = 16'(2330);
			9891: out = 16'(-475);
			9892: out = 16'(-1758);
			9893: out = 16'(-965);
			9894: out = 16'(446);
			9895: out = 16'(2449);
			9896: out = 16'(1307);
			9897: out = 16'(-1708);
			9898: out = 16'(-3341);
			9899: out = 16'(-870);
			9900: out = 16'(3030);
			9901: out = 16'(2216);
			9902: out = 16'(-76);
			9903: out = 16'(-349);
			9904: out = 16'(1080);
			9905: out = 16'(604);
			9906: out = 16'(386);
			9907: out = 16'(-469);
			9908: out = 16'(-251);
			9909: out = 16'(781);
			9910: out = 16'(1014);
			9911: out = 16'(-296);
			9912: out = 16'(-1367);
			9913: out = 16'(-261);
			9914: out = 16'(669);
			9915: out = 16'(78);
			9916: out = 16'(-755);
			9917: out = 16'(-151);
			9918: out = 16'(681);
			9919: out = 16'(911);
			9920: out = 16'(-715);
			9921: out = 16'(-2143);
			9922: out = 16'(-1948);
			9923: out = 16'(298);
			9924: out = 16'(2551);
			9925: out = 16'(1106);
			9926: out = 16'(-695);
			9927: out = 16'(-1060);
			9928: out = 16'(1297);
			9929: out = 16'(2081);
			9930: out = 16'(323);
			9931: out = 16'(-1753);
			9932: out = 16'(-1525);
			9933: out = 16'(116);
			9934: out = 16'(305);
			9935: out = 16'(-19);
			9936: out = 16'(-1466);
			9937: out = 16'(-2115);
			9938: out = 16'(-936);
			9939: out = 16'(1359);
			9940: out = 16'(2259);
			9941: out = 16'(1758);
			9942: out = 16'(31);
			9943: out = 16'(-2221);
			9944: out = 16'(-1136);
			9945: out = 16'(-244);
			9946: out = 16'(757);
			9947: out = 16'(2001);
			9948: out = 16'(455);
			9949: out = 16'(49);
			9950: out = 16'(1251);
			9951: out = 16'(810);
			9952: out = 16'(-428);
			9953: out = 16'(-2007);
			9954: out = 16'(-1937);
			9955: out = 16'(-417);
			9956: out = 16'(709);
			9957: out = 16'(1896);
			9958: out = 16'(2211);
			9959: out = 16'(1822);
			9960: out = 16'(-414);
			9961: out = 16'(-718);
			9962: out = 16'(-283);
			9963: out = 16'(779);
			9964: out = 16'(-174);
			9965: out = 16'(147);
			9966: out = 16'(1699);
			9967: out = 16'(483);
			9968: out = 16'(-2200);
			9969: out = 16'(-1286);
			9970: out = 16'(-1034);
			9971: out = 16'(-272);
			9972: out = 16'(1267);
			9973: out = 16'(633);
			9974: out = 16'(-1638);
			9975: out = 16'(-2565);
			9976: out = 16'(27);
			9977: out = 16'(1233);
			9978: out = 16'(1434);
			9979: out = 16'(1157);
			9980: out = 16'(1067);
			9981: out = 16'(-1425);
			9982: out = 16'(-2299);
			9983: out = 16'(-911);
			9984: out = 16'(1714);
			9985: out = 16'(1922);
			9986: out = 16'(-1615);
			9987: out = 16'(-3003);
			9988: out = 16'(-1018);
			9989: out = 16'(688);
			9990: out = 16'(703);
			9991: out = 16'(181);
			9992: out = 16'(21);
			9993: out = 16'(796);
			9994: out = 16'(1355);
			9995: out = 16'(-628);
			9996: out = 16'(-1809);
			9997: out = 16'(-1343);
			9998: out = 16'(1335);
			9999: out = 16'(1538);
			10000: out = 16'(1015);
			10001: out = 16'(1183);
			10002: out = 16'(1998);
			10003: out = 16'(737);
			10004: out = 16'(-1828);
			10005: out = 16'(-2846);
			10006: out = 16'(-1451);
			10007: out = 16'(436);
			10008: out = 16'(1409);
			10009: out = 16'(1000);
			10010: out = 16'(-391);
			10011: out = 16'(-720);
			10012: out = 16'(356);
			10013: out = 16'(1326);
			10014: out = 16'(-582);
			10015: out = 16'(-3322);
			10016: out = 16'(-2268);
			10017: out = 16'(375);
			10018: out = 16'(1516);
			10019: out = 16'(670);
			10020: out = 16'(-1820);
			10021: out = 16'(-1148);
			10022: out = 16'(1702);
			10023: out = 16'(2454);
			10024: out = 16'(302);
			10025: out = 16'(-3027);
			10026: out = 16'(-1386);
			10027: out = 16'(972);
			10028: out = 16'(1642);
			10029: out = 16'(1693);
			10030: out = 16'(524);
			10031: out = 16'(-646);
			10032: out = 16'(-3);
			10033: out = 16'(-935);
			10034: out = 16'(-1694);
			10035: out = 16'(-316);
			10036: out = 16'(704);
			10037: out = 16'(-869);
			10038: out = 16'(-181);
			10039: out = 16'(-167);
			10040: out = 16'(367);
			10041: out = 16'(1841);
			10042: out = 16'(38);
			10043: out = 16'(420);
			10044: out = 16'(570);
			10045: out = 16'(1913);
			10046: out = 16'(1035);
			10047: out = 16'(-193);
			10048: out = 16'(511);
			10049: out = 16'(1105);
			10050: out = 16'(132);
			10051: out = 16'(-393);
			10052: out = 16'(-95);
			10053: out = 16'(-168);
			10054: out = 16'(-1331);
			10055: out = 16'(-2560);
			10056: out = 16'(-1688);
			10057: out = 16'(-540);
			10058: out = 16'(-88);
			10059: out = 16'(700);
			10060: out = 16'(2207);
			10061: out = 16'(1036);
			10062: out = 16'(-1186);
			10063: out = 16'(-2641);
			10064: out = 16'(-2101);
			10065: out = 16'(610);
			10066: out = 16'(-348);
			10067: out = 16'(-9);
			10068: out = 16'(449);
			10069: out = 16'(-138);
			10070: out = 16'(265);
			10071: out = 16'(467);
			10072: out = 16'(1069);
			10073: out = 16'(1879);
			10074: out = 16'(198);
			10075: out = 16'(-1781);
			10076: out = 16'(-2526);
			10077: out = 16'(-1739);
			10078: out = 16'(723);
			10079: out = 16'(1131);
			10080: out = 16'(-1961);
			10081: out = 16'(-1379);
			10082: out = 16'(1208);
			10083: out = 16'(1589);
			10084: out = 16'(897);
			10085: out = 16'(317);
			10086: out = 16'(-494);
			10087: out = 16'(-958);
			10088: out = 16'(371);
			10089: out = 16'(448);
			10090: out = 16'(-668);
			10091: out = 16'(-1020);
			10092: out = 16'(699);
			10093: out = 16'(1023);
			10094: out = 16'(964);
			10095: out = 16'(2276);
			10096: out = 16'(1534);
			10097: out = 16'(-994);
			10098: out = 16'(-3471);
			10099: out = 16'(-2652);
			10100: out = 16'(-21);
			10101: out = 16'(2544);
			10102: out = 16'(1069);
			10103: out = 16'(-1915);
			10104: out = 16'(-1441);
			10105: out = 16'(31);
			10106: out = 16'(1449);
			10107: out = 16'(1346);
			10108: out = 16'(-1481);
			10109: out = 16'(-2564);
			10110: out = 16'(-1063);
			10111: out = 16'(1009);
			10112: out = 16'(1624);
			10113: out = 16'(1127);
			10114: out = 16'(289);
			10115: out = 16'(-1168);
			10116: out = 16'(59);
			10117: out = 16'(1480);
			10118: out = 16'(1485);
			10119: out = 16'(640);
			10120: out = 16'(-569);
			10121: out = 16'(-1068);
			10122: out = 16'(-1362);
			10123: out = 16'(-89);
			10124: out = 16'(468);
			10125: out = 16'(-1298);
			10126: out = 16'(-1382);
			10127: out = 16'(1176);
			10128: out = 16'(359);
			10129: out = 16'(-1931);
			10130: out = 16'(-2050);
			10131: out = 16'(-7);
			10132: out = 16'(704);
			10133: out = 16'(339);
			10134: out = 16'(587);
			10135: out = 16'(1003);
			10136: out = 16'(904);
			10137: out = 16'(491);
			10138: out = 16'(-697);
			10139: out = 16'(-1440);
			10140: out = 16'(-795);
			10141: out = 16'(-70);
			10142: out = 16'(1670);
			10143: out = 16'(2878);
			10144: out = 16'(1502);
			10145: out = 16'(-1196);
			10146: out = 16'(-2014);
			10147: out = 16'(-1520);
			10148: out = 16'(88);
			10149: out = 16'(89);
			10150: out = 16'(51);
			10151: out = 16'(712);
			10152: out = 16'(872);
			10153: out = 16'(-328);
			10154: out = 16'(-602);
			10155: out = 16'(677);
			10156: out = 16'(831);
			10157: out = 16'(-1597);
			10158: out = 16'(-1747);
			10159: out = 16'(612);
			10160: out = 16'(-113);
			10161: out = 16'(-385);
			10162: out = 16'(1221);
			10163: out = 16'(1259);
			10164: out = 16'(-1333);
			10165: out = 16'(-4941);
			10166: out = 16'(-4289);
			10167: out = 16'(317);
			10168: out = 16'(3661);
			10169: out = 16'(2522);
			10170: out = 16'(-614);
			10171: out = 16'(-1238);
			10172: out = 16'(-887);
			10173: out = 16'(1684);
			10174: out = 16'(947);
			10175: out = 16'(869);
			10176: out = 16'(1467);
			10177: out = 16'(800);
			10178: out = 16'(-41);
			10179: out = 16'(-718);
			10180: out = 16'(-1300);
			10181: out = 16'(-502);
			10182: out = 16'(-782);
			10183: out = 16'(-686);
			10184: out = 16'(-38);
			10185: out = 16'(410);
			10186: out = 16'(847);
			10187: out = 16'(-358);
			10188: out = 16'(-1835);
			10189: out = 16'(-1210);
			10190: out = 16'(377);
			10191: out = 16'(1799);
			10192: out = 16'(610);
			10193: out = 16'(304);
			10194: out = 16'(709);
			10195: out = 16'(935);
			10196: out = 16'(120);
			10197: out = 16'(-73);
			10198: out = 16'(-710);
			10199: out = 16'(-458);
			10200: out = 16'(-310);
			10201: out = 16'(151);
			10202: out = 16'(1414);
			10203: out = 16'(680);
			10204: out = 16'(-1982);
			10205: out = 16'(-3135);
			10206: out = 16'(-2160);
			10207: out = 16'(-677);
			10208: out = 16'(1616);
			10209: out = 16'(1223);
			10210: out = 16'(-252);
			10211: out = 16'(-1104);
			10212: out = 16'(-60);
			10213: out = 16'(942);
			10214: out = 16'(1122);
			10215: out = 16'(328);
			10216: out = 16'(-810);
			10217: out = 16'(-779);
			10218: out = 16'(-648);
			10219: out = 16'(833);
			10220: out = 16'(2287);
			10221: out = 16'(1302);
			10222: out = 16'(-500);
			10223: out = 16'(-1095);
			10224: out = 16'(-770);
			10225: out = 16'(639);
			10226: out = 16'(1181);
			10227: out = 16'(-252);
			10228: out = 16'(-1154);
			10229: out = 16'(-757);
			10230: out = 16'(3);
			10231: out = 16'(656);
			10232: out = 16'(641);
			10233: out = 16'(-468);
			10234: out = 16'(557);
			10235: out = 16'(1054);
			10236: out = 16'(27);
			10237: out = 16'(-1375);
			10238: out = 16'(-1967);
			10239: out = 16'(-736);
			10240: out = 16'(1115);
			10241: out = 16'(1570);
			10242: out = 16'(-457);
			10243: out = 16'(-11);
			10244: out = 16'(1618);
			10245: out = 16'(1338);
			10246: out = 16'(-1304);
			10247: out = 16'(-3438);
			10248: out = 16'(-1808);
			10249: out = 16'(1182);
			10250: out = 16'(3263);
			10251: out = 16'(1838);
			10252: out = 16'(-765);
			10253: out = 16'(-1549);
			10254: out = 16'(332);
			10255: out = 16'(1668);
			10256: out = 16'(2205);
			10257: out = 16'(438);
			10258: out = 16'(-716);
			10259: out = 16'(-938);
			10260: out = 16'(-885);
			10261: out = 16'(-541);
			10262: out = 16'(-1277);
			10263: out = 16'(-2561);
			10264: out = 16'(-1252);
			10265: out = 16'(841);
			10266: out = 16'(322);
			10267: out = 16'(547);
			10268: out = 16'(2147);
			10269: out = 16'(1688);
			10270: out = 16'(-1263);
			10271: out = 16'(-3153);
			10272: out = 16'(-2009);
			10273: out = 16'(319);
			10274: out = 16'(2798);
			10275: out = 16'(2138);
			10276: out = 16'(-1168);
			10277: out = 16'(-3170);
			10278: out = 16'(-1924);
			10279: out = 16'(1338);
			10280: out = 16'(1658);
			10281: out = 16'(642);
			10282: out = 16'(298);
			10283: out = 16'(-105);
			10284: out = 16'(-1422);
			10285: out = 16'(-1269);
			10286: out = 16'(431);
			10287: out = 16'(1449);
			10288: out = 16'(2067);
			10289: out = 16'(365);
			10290: out = 16'(-1780);
			10291: out = 16'(-1541);
			10292: out = 16'(568);
			10293: out = 16'(2205);
			10294: out = 16'(1134);
			10295: out = 16'(-909);
			10296: out = 16'(-1082);
			10297: out = 16'(238);
			10298: out = 16'(2227);
			10299: out = 16'(1404);
			10300: out = 16'(-1218);
			10301: out = 16'(-1407);
			10302: out = 16'(-656);
			10303: out = 16'(-614);
			10304: out = 16'(73);
			10305: out = 16'(416);
			10306: out = 16'(236);
			10307: out = 16'(-65);
			10308: out = 16'(758);
			10309: out = 16'(712);
			10310: out = 16'(-157);
			10311: out = 16'(1057);
			10312: out = 16'(1491);
			10313: out = 16'(1167);
			10314: out = 16'(-314);
			10315: out = 16'(-1276);
			10316: out = 16'(-996);
			10317: out = 16'(628);
			10318: out = 16'(472);
			10319: out = 16'(-1535);
			10320: out = 16'(-2133);
			10321: out = 16'(-243);
			10322: out = 16'(1324);
			10323: out = 16'(-81);
			10324: out = 16'(-1686);
			10325: out = 16'(-196);
			10326: out = 16'(925);
			10327: out = 16'(1136);
			10328: out = 16'(-1);
			10329: out = 16'(44);
			10330: out = 16'(1053);
			10331: out = 16'(568);
			10332: out = 16'(-224);
			10333: out = 16'(-1036);
			10334: out = 16'(-122);
			10335: out = 16'(57);
			10336: out = 16'(-120);
			10337: out = 16'(642);
			10338: out = 16'(-55);
			10339: out = 16'(-482);
			10340: out = 16'(143);
			10341: out = 16'(327);
			10342: out = 16'(7);
			10343: out = 16'(156);
			10344: out = 16'(131);
			10345: out = 16'(-669);
			10346: out = 16'(-879);
			10347: out = 16'(-1160);
			10348: out = 16'(-635);
			10349: out = 16'(9);
			10350: out = 16'(419);
			10351: out = 16'(-390);
			10352: out = 16'(-1045);
			10353: out = 16'(-143);
			10354: out = 16'(390);
			10355: out = 16'(659);
			10356: out = 16'(-1140);
			10357: out = 16'(-30);
			10358: out = 16'(1019);
			10359: out = 16'(359);
			10360: out = 16'(609);
			10361: out = 16'(1190);
			10362: out = 16'(-472);
			10363: out = 16'(-1292);
			10364: out = 16'(246);
			10365: out = 16'(120);
			10366: out = 16'(-560);
			10367: out = 16'(-2166);
			10368: out = 16'(-1349);
			10369: out = 16'(924);
			10370: out = 16'(2430);
			10371: out = 16'(2015);
			10372: out = 16'(-47);
			10373: out = 16'(-840);
			10374: out = 16'(-1072);
			10375: out = 16'(116);
			10376: out = 16'(544);
			10377: out = 16'(801);
			10378: out = 16'(782);
			10379: out = 16'(967);
			10380: out = 16'(-970);
			10381: out = 16'(-1765);
			10382: out = 16'(-123);
			10383: out = 16'(647);
			10384: out = 16'(-234);
			10385: out = 16'(-21);
			10386: out = 16'(487);
			10387: out = 16'(-1423);
			10388: out = 16'(-2518);
			10389: out = 16'(-1469);
			10390: out = 16'(271);
			10391: out = 16'(1601);
			10392: out = 16'(1617);
			10393: out = 16'(155);
			10394: out = 16'(-1768);
			10395: out = 16'(-1834);
			10396: out = 16'(945);
			10397: out = 16'(2472);
			10398: out = 16'(611);
			10399: out = 16'(-1811);
			10400: out = 16'(-1546);
			10401: out = 16'(102);
			10402: out = 16'(1113);
			10403: out = 16'(615);
			10404: out = 16'(1);
			10405: out = 16'(1520);
			10406: out = 16'(2215);
			10407: out = 16'(-144);
			10408: out = 16'(-1026);
			10409: out = 16'(-885);
			10410: out = 16'(868);
			10411: out = 16'(91);
			10412: out = 16'(-391);
			10413: out = 16'(1354);
			10414: out = 16'(1273);
			10415: out = 16'(-338);
			10416: out = 16'(-293);
			10417: out = 16'(-153);
			10418: out = 16'(159);
			10419: out = 16'(-1054);
			10420: out = 16'(-1280);
			10421: out = 16'(329);
			10422: out = 16'(34);
			10423: out = 16'(-1059);
			10424: out = 16'(-764);
			10425: out = 16'(-693);
			10426: out = 16'(-2413);
			10427: out = 16'(-789);
			10428: out = 16'(951);
			10429: out = 16'(486);
			10430: out = 16'(1207);
			10431: out = 16'(844);
			10432: out = 16'(-1092);
			10433: out = 16'(-1792);
			10434: out = 16'(-567);
			10435: out = 16'(1866);
			10436: out = 16'(1298);
			10437: out = 16'(-214);
			10438: out = 16'(-68);
			10439: out = 16'(942);
			10440: out = 16'(1405);
			10441: out = 16'(-265);
			10442: out = 16'(-2190);
			10443: out = 16'(-940);
			10444: out = 16'(778);
			10445: out = 16'(659);
			10446: out = 16'(-276);
			10447: out = 16'(-550);
			10448: out = 16'(20);
			10449: out = 16'(1418);
			10450: out = 16'(1773);
			10451: out = 16'(1183);
			10452: out = 16'(475);
			10453: out = 16'(170);
			10454: out = 16'(-172);
			10455: out = 16'(217);
			10456: out = 16'(-269);
			10457: out = 16'(-1147);
			10458: out = 16'(-1627);
			10459: out = 16'(-449);
			10460: out = 16'(631);
			10461: out = 16'(-564);
			10462: out = 16'(-1416);
			10463: out = 16'(634);
			10464: out = 16'(1160);
			10465: out = 16'(-76);
			10466: out = 16'(-1484);
			10467: out = 16'(-475);
			10468: out = 16'(-118);
			10469: out = 16'(-36);
			10470: out = 16'(721);
			10471: out = 16'(-152);
			10472: out = 16'(-1476);
			10473: out = 16'(-1220);
			10474: out = 16'(-109);
			10475: out = 16'(16);
			10476: out = 16'(530);
			10477: out = 16'(919);
			10478: out = 16'(1157);
			10479: out = 16'(465);
			10480: out = 16'(-272);
			10481: out = 16'(-521);
			10482: out = 16'(53);
			10483: out = 16'(698);
			10484: out = 16'(-380);
			10485: out = 16'(-613);
			10486: out = 16'(-527);
			10487: out = 16'(-427);
			10488: out = 16'(404);
			10489: out = 16'(1294);
			10490: out = 16'(-333);
			10491: out = 16'(-1588);
			10492: out = 16'(-82);
			10493: out = 16'(1585);
			10494: out = 16'(31);
			10495: out = 16'(-697);
			10496: out = 16'(542);
			10497: out = 16'(520);
			10498: out = 16'(-512);
			10499: out = 16'(276);
			10500: out = 16'(361);
			10501: out = 16'(240);
			10502: out = 16'(-171);
			10503: out = 16'(-1037);
			10504: out = 16'(489);
			10505: out = 16'(823);
			10506: out = 16'(-483);
			10507: out = 16'(-763);
			10508: out = 16'(-619);
			10509: out = 16'(-840);
			10510: out = 16'(-318);
			10511: out = 16'(17);
			10512: out = 16'(649);
			10513: out = 16'(512);
			10514: out = 16'(506);
			10515: out = 16'(-168);
			10516: out = 16'(-14);
			10517: out = 16'(-229);
			10518: out = 16'(-1177);
			10519: out = 16'(-149);
			10520: out = 16'(738);
			10521: out = 16'(305);
			10522: out = 16'(-1640);
			10523: out = 16'(-1120);
			10524: out = 16'(299);
			10525: out = 16'(936);
			10526: out = 16'(164);
			10527: out = 16'(-85);
			10528: out = 16'(-234);
			10529: out = 16'(-564);
			10530: out = 16'(630);
			10531: out = 16'(739);
			10532: out = 16'(770);
			10533: out = 16'(-745);
			10534: out = 16'(-1427);
			10535: out = 16'(-292);
			10536: out = 16'(495);
			10537: out = 16'(1034);
			10538: out = 16'(518);
			10539: out = 16'(-1530);
			10540: out = 16'(-2068);
			10541: out = 16'(-524);
			10542: out = 16'(1062);
			10543: out = 16'(1062);
			10544: out = 16'(-139);
			10545: out = 16'(-390);
			10546: out = 16'(-386);
			10547: out = 16'(-472);
			10548: out = 16'(173);
			10549: out = 16'(1143);
			10550: out = 16'(359);
			10551: out = 16'(154);
			10552: out = 16'(-127);
			10553: out = 16'(479);
			10554: out = 16'(579);
			10555: out = 16'(-716);
			10556: out = 16'(-1561);
			10557: out = 16'(-382);
			10558: out = 16'(-43);
			10559: out = 16'(-972);
			10560: out = 16'(-421);
			10561: out = 16'(357);
			10562: out = 16'(186);
			10563: out = 16'(718);
			10564: out = 16'(968);
			10565: out = 16'(-480);
			10566: out = 16'(-2219);
			10567: out = 16'(-2003);
			10568: out = 16'(294);
			10569: out = 16'(1607);
			10570: out = 16'(921);
			10571: out = 16'(286);
			10572: out = 16'(735);
			10573: out = 16'(666);
			10574: out = 16'(353);
			10575: out = 16'(-616);
			10576: out = 16'(-1130);
			10577: out = 16'(-572);
			10578: out = 16'(1145);
			10579: out = 16'(621);
			10580: out = 16'(-609);
			10581: out = 16'(-755);
			10582: out = 16'(-479);
			10583: out = 16'(-486);
			10584: out = 16'(365);
			10585: out = 16'(1752);
			10586: out = 16'(862);
			10587: out = 16'(-782);
			10588: out = 16'(-1676);
			10589: out = 16'(-367);
			10590: out = 16'(1427);
			10591: out = 16'(101);
			10592: out = 16'(-787);
			10593: out = 16'(-159);
			10594: out = 16'(-115);
			10595: out = 16'(-759);
			10596: out = 16'(-556);
			10597: out = 16'(337);
			10598: out = 16'(412);
			10599: out = 16'(152);
			10600: out = 16'(562);
			10601: out = 16'(-143);
			10602: out = 16'(-436);
			10603: out = 16'(-1263);
			10604: out = 16'(-152);
			10605: out = 16'(665);
			10606: out = 16'(317);
			10607: out = 16'(1145);
			10608: out = 16'(493);
			10609: out = 16'(-932);
			10610: out = 16'(-1147);
			10611: out = 16'(-331);
			10612: out = 16'(582);
			10613: out = 16'(404);
			10614: out = 16'(1132);
			10615: out = 16'(1384);
			10616: out = 16'(74);
			10617: out = 16'(-1474);
			10618: out = 16'(-1583);
			10619: out = 16'(-184);
			10620: out = 16'(909);
			10621: out = 16'(68);
			10622: out = 16'(-978);
			10623: out = 16'(-801);
			10624: out = 16'(-1134);
			10625: out = 16'(-1118);
			10626: out = 16'(1409);
			10627: out = 16'(889);
			10628: out = 16'(-547);
			10629: out = 16'(309);
			10630: out = 16'(1196);
			10631: out = 16'(-83);
			10632: out = 16'(-1907);
			10633: out = 16'(-1818);
			10634: out = 16'(-492);
			10635: out = 16'(1527);
			10636: out = 16'(2062);
			10637: out = 16'(-450);
			10638: out = 16'(-857);
			10639: out = 16'(8);
			10640: out = 16'(1920);
			10641: out = 16'(1777);
			10642: out = 16'(450);
			10643: out = 16'(-41);
			10644: out = 16'(669);
			10645: out = 16'(427);
			10646: out = 16'(-824);
			10647: out = 16'(-1603);
			10648: out = 16'(-544);
			10649: out = 16'(110);
			10650: out = 16'(-612);
			10651: out = 16'(36);
			10652: out = 16'(793);
			10653: out = 16'(96);
			10654: out = 16'(-1043);
			10655: out = 16'(-1658);
			10656: out = 16'(-1233);
			10657: out = 16'(-631);
			10658: out = 16'(452);
			10659: out = 16'(1782);
			10660: out = 16'(666);
			10661: out = 16'(-262);
			10662: out = 16'(362);
			10663: out = 16'(766);
			10664: out = 16'(295);
			10665: out = 16'(-1425);
			10666: out = 16'(-1341);
			10667: out = 16'(623);
			10668: out = 16'(328);
			10669: out = 16'(-109);
			10670: out = 16'(808);
			10671: out = 16'(838);
			10672: out = 16'(784);
			10673: out = 16'(-36);
			10674: out = 16'(-519);
			10675: out = 16'(-170);
			10676: out = 16'(-549);
			10677: out = 16'(554);
			10678: out = 16'(653);
			10679: out = 16'(-38);
			10680: out = 16'(-443);
			10681: out = 16'(356);
			10682: out = 16'(527);
			10683: out = 16'(756);
			10684: out = 16'(-297);
			10685: out = 16'(-772);
			10686: out = 16'(-166);
			10687: out = 16'(309);
			10688: out = 16'(761);
			10689: out = 16'(-69);
			10690: out = 16'(-855);
			10691: out = 16'(-30);
			10692: out = 16'(806);
			10693: out = 16'(600);
			10694: out = 16'(-146);
			10695: out = 16'(-875);
			10696: out = 16'(-301);
			10697: out = 16'(-391);
			10698: out = 16'(483);
			10699: out = 16'(1047);
			10700: out = 16'(-289);
			10701: out = 16'(-2399);
			10702: out = 16'(-1884);
			10703: out = 16'(-842);
			10704: out = 16'(-112);
			10705: out = 16'(1118);
			10706: out = 16'(687);
			10707: out = 16'(-442);
			10708: out = 16'(-42);
			10709: out = 16'(874);
			10710: out = 16'(509);
			10711: out = 16'(-66);
			10712: out = 16'(-454);
			10713: out = 16'(-42);
			10714: out = 16'(-753);
			10715: out = 16'(-935);
			10716: out = 16'(870);
			10717: out = 16'(1232);
			10718: out = 16'(291);
			10719: out = 16'(-685);
			10720: out = 16'(-1013);
			10721: out = 16'(-410);
			10722: out = 16'(1400);
			10723: out = 16'(1761);
			10724: out = 16'(-444);
			10725: out = 16'(-2171);
			10726: out = 16'(-943);
			10727: out = 16'(1164);
			10728: out = 16'(1363);
			10729: out = 16'(-304);
			10730: out = 16'(-664);
			10731: out = 16'(930);
			10732: out = 16'(1095);
			10733: out = 16'(99);
			10734: out = 16'(-732);
			10735: out = 16'(-128);
			10736: out = 16'(-112);
			10737: out = 16'(-653);
			10738: out = 16'(-858);
			10739: out = 16'(-115);
			10740: out = 16'(1307);
			10741: out = 16'(1129);
			10742: out = 16'(-848);
			10743: out = 16'(-1975);
			10744: out = 16'(-1503);
			10745: out = 16'(1080);
			10746: out = 16'(2523);
			10747: out = 16'(998);
			10748: out = 16'(-1531);
			10749: out = 16'(-2087);
			10750: out = 16'(-637);
			10751: out = 16'(1247);
			10752: out = 16'(1469);
			10753: out = 16'(-324);
			10754: out = 16'(-1068);
			10755: out = 16'(-477);
			10756: out = 16'(-119);
			10757: out = 16'(829);
			10758: out = 16'(141);
			10759: out = 16'(128);
			10760: out = 16'(956);
			10761: out = 16'(434);
			10762: out = 16'(-331);
			10763: out = 16'(-1301);
			10764: out = 16'(-1109);
			10765: out = 16'(212);
			10766: out = 16'(1387);
			10767: out = 16'(-64);
			10768: out = 16'(-666);
			10769: out = 16'(529);
			10770: out = 16'(710);
			10771: out = 16'(262);
			10772: out = 16'(-663);
			10773: out = 16'(-172);
			10774: out = 16'(305);
			10775: out = 16'(1268);
			10776: out = 16'(1060);
			10777: out = 16'(-172);
			10778: out = 16'(-1770);
			10779: out = 16'(-1508);
			10780: out = 16'(-385);
			10781: out = 16'(127);
			10782: out = 16'(245);
			10783: out = 16'(479);
			10784: out = 16'(111);
			10785: out = 16'(147);
			10786: out = 16'(220);
			10787: out = 16'(16);
			10788: out = 16'(-316);
			10789: out = 16'(-243);
			10790: out = 16'(367);
			10791: out = 16'(-432);
			10792: out = 16'(-1084);
			10793: out = 16'(-366);
			10794: out = 16'(593);
			10795: out = 16'(1039);
			10796: out = 16'(789);
			10797: out = 16'(622);
			10798: out = 16'(712);
			10799: out = 16'(157);
			10800: out = 16'(-722);
			10801: out = 16'(-1295);
			10802: out = 16'(-1886);
			10803: out = 16'(-1438);
			10804: out = 16'(104);
			10805: out = 16'(465);
			10806: out = 16'(416);
			10807: out = 16'(729);
			10808: out = 16'(1398);
			10809: out = 16'(1284);
			10810: out = 16'(-469);
			10811: out = 16'(-1824);
			10812: out = 16'(-1858);
			10813: out = 16'(-1042);
			10814: out = 16'(690);
			10815: out = 16'(1713);
			10816: out = 16'(666);
			10817: out = 16'(-163);
			10818: out = 16'(147);
			10819: out = 16'(370);
			10820: out = 16'(2);
			10821: out = 16'(-1013);
			10822: out = 16'(-762);
			10823: out = 16'(251);
			10824: out = 16'(1161);
			10825: out = 16'(113);
			10826: out = 16'(-881);
			10827: out = 16'(-201);
			10828: out = 16'(1174);
			10829: out = 16'(953);
			10830: out = 16'(-301);
			10831: out = 16'(-328);
			10832: out = 16'(267);
			10833: out = 16'(295);
			10834: out = 16'(-205);
			10835: out = 16'(-351);
			10836: out = 16'(-272);
			10837: out = 16'(-691);
			10838: out = 16'(-919);
			10839: out = 16'(-280);
			10840: out = 16'(-228);
			10841: out = 16'(-48);
			10842: out = 16'(554);
			10843: out = 16'(714);
			10844: out = 16'(-298);
			10845: out = 16'(-1823);
			10846: out = 16'(-1778);
			10847: out = 16'(-8);
			10848: out = 16'(1326);
			10849: out = 16'(1089);
			10850: out = 16'(124);
			10851: out = 16'(-222);
			10852: out = 16'(-270);
			10853: out = 16'(413);
			10854: out = 16'(582);
			10855: out = 16'(-460);
			10856: out = 16'(-616);
			10857: out = 16'(-157);
			10858: out = 16'(720);
			10859: out = 16'(986);
			10860: out = 16'(455);
			10861: out = 16'(63);
			10862: out = 16'(8);
			10863: out = 16'(-249);
			10864: out = 16'(-1355);
			10865: out = 16'(-1934);
			10866: out = 16'(-306);
			10867: out = 16'(781);
			10868: out = 16'(-205);
			10869: out = 16'(-718);
			10870: out = 16'(144);
			10871: out = 16'(855);
			10872: out = 16'(353);
			10873: out = 16'(-1665);
			10874: out = 16'(-1297);
			10875: out = 16'(-143);
			10876: out = 16'(523);
			10877: out = 16'(1229);
			10878: out = 16'(1210);
			10879: out = 16'(137);
			10880: out = 16'(-817);
			10881: out = 16'(-1442);
			10882: out = 16'(-1493);
			10883: out = 16'(-332);
			10884: out = 16'(215);
			10885: out = 16'(636);
			10886: out = 16'(930);
			10887: out = 16'(536);
			10888: out = 16'(-479);
			10889: out = 16'(-302);
			10890: out = 16'(473);
			10891: out = 16'(214);
			10892: out = 16'(-74);
			10893: out = 16'(247);
			10894: out = 16'(507);
			10895: out = 16'(-582);
			10896: out = 16'(-792);
			10897: out = 16'(-339);
			10898: out = 16'(560);
			10899: out = 16'(17);
			10900: out = 16'(-796);
			10901: out = 16'(-90);
			10902: out = 16'(524);
			10903: out = 16'(893);
			10904: out = 16'(428);
			10905: out = 16'(228);
			10906: out = 16'(-594);
			10907: out = 16'(-1182);
			10908: out = 16'(-712);
			10909: out = 16'(719);
			10910: out = 16'(1481);
			10911: out = 16'(43);
			10912: out = 16'(-966);
			10913: out = 16'(-375);
			10914: out = 16'(420);
			10915: out = 16'(398);
			10916: out = 16'(-1258);
			10917: out = 16'(-1439);
			10918: out = 16'(-49);
			10919: out = 16'(628);
			10920: out = 16'(654);
			10921: out = 16'(157);
			10922: out = 16'(251);
			10923: out = 16'(-71);
			10924: out = 16'(-1017);
			10925: out = 16'(-46);
			10926: out = 16'(691);
			10927: out = 16'(-63);
			10928: out = 16'(-289);
			10929: out = 16'(574);
			10930: out = 16'(311);
			10931: out = 16'(-1506);
			10932: out = 16'(-2437);
			10933: out = 16'(-1236);
			10934: out = 16'(207);
			10935: out = 16'(1079);
			10936: out = 16'(1389);
			10937: out = 16'(507);
			10938: out = 16'(-792);
			10939: out = 16'(-1270);
			10940: out = 16'(-418);
			10941: out = 16'(1012);
			10942: out = 16'(1594);
			10943: out = 16'(-228);
			10944: out = 16'(-1523);
			10945: out = 16'(-1275);
			10946: out = 16'(509);
			10947: out = 16'(1367);
			10948: out = 16'(85);
			10949: out = 16'(-440);
			10950: out = 16'(845);
			10951: out = 16'(1085);
			10952: out = 16'(-301);
			10953: out = 16'(-1889);
			10954: out = 16'(-1082);
			10955: out = 16'(198);
			10956: out = 16'(320);
			10957: out = 16'(885);
			10958: out = 16'(621);
			10959: out = 16'(-259);
			10960: out = 16'(-262);
			10961: out = 16'(-396);
			10962: out = 16'(-928);
			10963: out = 16'(-767);
			10964: out = 16'(133);
			10965: out = 16'(602);
			10966: out = 16'(183);
			10967: out = 16'(583);
			10968: out = 16'(742);
			10969: out = 16'(491);
			10970: out = 16'(139);
			10971: out = 16'(-346);
			10972: out = 16'(420);
			10973: out = 16'(855);
			10974: out = 16'(406);
			10975: out = 16'(-510);
			10976: out = 16'(-469);
			10977: out = 16'(-63);
			10978: out = 16'(-176);
			10979: out = 16'(-1291);
			10980: out = 16'(-631);
			10981: out = 16'(282);
			10982: out = 16'(521);
			10983: out = 16'(884);
			10984: out = 16'(1025);
			10985: out = 16'(349);
			10986: out = 16'(-1244);
			10987: out = 16'(-1323);
			10988: out = 16'(-189);
			10989: out = 16'(524);
			10990: out = 16'(143);
			10991: out = 16'(-467);
			10992: out = 16'(-62);
			10993: out = 16'(594);
			10994: out = 16'(213);
			10995: out = 16'(180);
			10996: out = 16'(41);
			10997: out = 16'(-155);
			10998: out = 16'(-53);
			10999: out = 16'(-381);
			11000: out = 16'(-907);
			11001: out = 16'(-489);
			11002: out = 16'(505);
			11003: out = 16'(1126);
			11004: out = 16'(816);
			11005: out = 16'(-106);
			11006: out = 16'(-394);
			11007: out = 16'(-383);
			11008: out = 16'(191);
			11009: out = 16'(1452);
			11010: out = 16'(555);
			11011: out = 16'(-801);
			11012: out = 16'(-711);
			11013: out = 16'(185);
			11014: out = 16'(731);
			11015: out = 16'(-177);
			11016: out = 16'(-1583);
			11017: out = 16'(-694);
			11018: out = 16'(785);
			11019: out = 16'(1087);
			11020: out = 16'(-706);
			11021: out = 16'(-772);
			11022: out = 16'(283);
			11023: out = 16'(791);
			11024: out = 16'(658);
			11025: out = 16'(211);
			11026: out = 16'(-129);
			11027: out = 16'(333);
			11028: out = 16'(800);
			11029: out = 16'(60);
			11030: out = 16'(-1132);
			11031: out = 16'(-1488);
			11032: out = 16'(-342);
			11033: out = 16'(-33);
			11034: out = 16'(340);
			11035: out = 16'(179);
			11036: out = 16'(455);
			11037: out = 16'(10);
			11038: out = 16'(-1221);
			11039: out = 16'(-595);
			11040: out = 16'(481);
			11041: out = 16'(1357);
			11042: out = 16'(671);
			11043: out = 16'(-32);
			11044: out = 16'(-276);
			11045: out = 16'(47);
			11046: out = 16'(142);
			11047: out = 16'(-126);
			11048: out = 16'(-7);
			11049: out = 16'(174);
			11050: out = 16'(73);
			11051: out = 16'(-457);
			11052: out = 16'(-213);
			11053: out = 16'(-466);
			11054: out = 16'(-360);
			11055: out = 16'(-359);
			11056: out = 16'(-786);
			11057: out = 16'(-308);
			11058: out = 16'(190);
			11059: out = 16'(332);
			11060: out = 16'(497);
			11061: out = 16'(448);
			11062: out = 16'(764);
			11063: out = 16'(-321);
			11064: out = 16'(-935);
			11065: out = 16'(435);
			11066: out = 16'(1043);
			11067: out = 16'(233);
			11068: out = 16'(-733);
			11069: out = 16'(-1351);
			11070: out = 16'(-99);
			11071: out = 16'(893);
			11072: out = 16'(567);
			11073: out = 16'(-112);
			11074: out = 16'(-36);
			11075: out = 16'(603);
			11076: out = 16'(532);
			11077: out = 16'(23);
			11078: out = 16'(-908);
			11079: out = 16'(-843);
			11080: out = 16'(486);
			11081: out = 16'(266);
			11082: out = 16'(-596);
			11083: out = 16'(-836);
			11084: out = 16'(-912);
			11085: out = 16'(522);
			11086: out = 16'(1731);
			11087: out = 16'(688);
			11088: out = 16'(-1537);
			11089: out = 16'(-2291);
			11090: out = 16'(-1648);
			11091: out = 16'(574);
			11092: out = 16'(2022);
			11093: out = 16'(480);
			11094: out = 16'(-602);
			11095: out = 16'(-51);
			11096: out = 16'(500);
			11097: out = 16'(271);
			11098: out = 16'(-478);
			11099: out = 16'(-457);
			11100: out = 16'(737);
			11101: out = 16'(1769);
			11102: out = 16'(573);
			11103: out = 16'(-1188);
			11104: out = 16'(-1348);
			11105: out = 16'(-465);
			11106: out = 16'(191);
			11107: out = 16'(661);
			11108: out = 16'(823);
			11109: out = 16'(-280);
			11110: out = 16'(-903);
			11111: out = 16'(-177);
			11112: out = 16'(38);
			11113: out = 16'(-5);
			11114: out = 16'(-759);
			11115: out = 16'(-723);
			11116: out = 16'(167);
			11117: out = 16'(548);
			11118: out = 16'(885);
			11119: out = 16'(-29);
			11120: out = 16'(-825);
			11121: out = 16'(-218);
			11122: out = 16'(346);
			11123: out = 16'(619);
			11124: out = 16'(730);
			11125: out = 16'(710);
			11126: out = 16'(-37);
			11127: out = 16'(-1298);
			11128: out = 16'(-1841);
			11129: out = 16'(-441);
			11130: out = 16'(728);
			11131: out = 16'(-30);
			11132: out = 16'(-711);
			11133: out = 16'(-697);
			11134: out = 16'(-231);
			11135: out = 16'(388);
			11136: out = 16'(1084);
			11137: out = 16'(1118);
			11138: out = 16'(-318);
			11139: out = 16'(-1540);
			11140: out = 16'(-1510);
			11141: out = 16'(354);
			11142: out = 16'(1261);
			11143: out = 16'(259);
			11144: out = 16'(-387);
			11145: out = 16'(-286);
			11146: out = 16'(-216);
			11147: out = 16'(991);
			11148: out = 16'(545);
			11149: out = 16'(-20);
			11150: out = 16'(-6);
			11151: out = 16'(6);
			11152: out = 16'(144);
			11153: out = 16'(-784);
			11154: out = 16'(-552);
			11155: out = 16'(733);
			11156: out = 16'(782);
			11157: out = 16'(319);
			11158: out = 16'(97);
			11159: out = 16'(91);
			11160: out = 16'(-506);
			11161: out = 16'(-761);
			11162: out = 16'(-469);
			11163: out = 16'(-72);
			11164: out = 16'(108);
			11165: out = 16'(-553);
			11166: out = 16'(-617);
			11167: out = 16'(127);
			11168: out = 16'(630);
			11169: out = 16'(764);
			11170: out = 16'(-1);
			11171: out = 16'(-1390);
			11172: out = 16'(-1857);
			11173: out = 16'(-256);
			11174: out = 16'(1222);
			11175: out = 16'(794);
			11176: out = 16'(374);
			11177: out = 16'(64);
			11178: out = 16'(233);
			11179: out = 16'(-28);
			11180: out = 16'(147);
			11181: out = 16'(66);
			11182: out = 16'(-113);
			11183: out = 16'(-92);
			11184: out = 16'(-467);
			11185: out = 16'(690);
			11186: out = 16'(1047);
			11187: out = 16'(-118);
			11188: out = 16'(-691);
			11189: out = 16'(-323);
			11190: out = 16'(383);
			11191: out = 16'(685);
			11192: out = 16'(472);
			11193: out = 16'(271);
			11194: out = 16'(-159);
			11195: out = 16'(-329);
			11196: out = 16'(-115);
			11197: out = 16'(264);
			11198: out = 16'(331);
			11199: out = 16'(-424);
			11200: out = 16'(-923);
			11201: out = 16'(-215);
			11202: out = 16'(695);
			11203: out = 16'(199);
			11204: out = 16'(-1493);
			11205: out = 16'(-1388);
			11206: out = 16'(-149);
			11207: out = 16'(634);
			11208: out = 16'(640);
			11209: out = 16'(317);
			11210: out = 16'(373);
			11211: out = 16'(-1);
			11212: out = 16'(-483);
			11213: out = 16'(-1191);
			11214: out = 16'(-1176);
			11215: out = 16'(-886);
			11216: out = 16'(-48);
			11217: out = 16'(744);
			11218: out = 16'(128);
			11219: out = 16'(-57);
			11220: out = 16'(749);
			11221: out = 16'(596);
			11222: out = 16'(87);
			11223: out = 16'(-377);
			11224: out = 16'(-73);
			11225: out = 16'(-10);
			11226: out = 16'(85);
			11227: out = 16'(411);
			11228: out = 16'(-101);
			11229: out = 16'(-1089);
			11230: out = 16'(-850);
			11231: out = 16'(229);
			11232: out = 16'(570);
			11233: out = 16'(621);
			11234: out = 16'(-141);
			11235: out = 16'(28);
			11236: out = 16'(-112);
			11237: out = 16'(-419);
			11238: out = 16'(22);
			11239: out = 16'(-208);
			11240: out = 16'(-267);
			11241: out = 16'(410);
			11242: out = 16'(-20);
			11243: out = 16'(-1093);
			11244: out = 16'(-1331);
			11245: out = 16'(-406);
			11246: out = 16'(523);
			11247: out = 16'(1026);
			11248: out = 16'(1118);
			11249: out = 16'(363);
			11250: out = 16'(-680);
			11251: out = 16'(-1510);
			11252: out = 16'(-1065);
			11253: out = 16'(-446);
			11254: out = 16'(53);
			11255: out = 16'(844);
			11256: out = 16'(257);
			11257: out = 16'(-660);
			11258: out = 16'(-232);
			11259: out = 16'(722);
			11260: out = 16'(1317);
			11261: out = 16'(224);
			11262: out = 16'(-857);
			11263: out = 16'(-823);
			11264: out = 16'(-77);
			11265: out = 16'(670);
			11266: out = 16'(308);
			11267: out = 16'(-252);
			11268: out = 16'(-509);
			11269: out = 16'(93);
			11270: out = 16'(155);
			11271: out = 16'(-214);
			11272: out = 16'(255);
			11273: out = 16'(173);
			11274: out = 16'(481);
			11275: out = 16'(545);
			11276: out = 16'(44);
			11277: out = 16'(433);
			11278: out = 16'(405);
			11279: out = 16'(-6);
			11280: out = 16'(-385);
			11281: out = 16'(-535);
			11282: out = 16'(-263);
			11283: out = 16'(-227);
			11284: out = 16'(-59);
			11285: out = 16'(-16);
			11286: out = 16'(-88);
			11287: out = 16'(-41);
			11288: out = 16'(202);
			11289: out = 16'(115);
			11290: out = 16'(-86);
			11291: out = 16'(-511);
			11292: out = 16'(220);
			11293: out = 16'(633);
			11294: out = 16'(-261);
			11295: out = 16'(-1207);
			11296: out = 16'(-686);
			11297: out = 16'(13);
			11298: out = 16'(-161);
			11299: out = 16'(-287);
			11300: out = 16'(379);
			11301: out = 16'(374);
			11302: out = 16'(-422);
			11303: out = 16'(-696);
			11304: out = 16'(-230);
			11305: out = 16'(-177);
			11306: out = 16'(295);
			11307: out = 16'(757);
			11308: out = 16'(224);
			11309: out = 16'(-722);
			11310: out = 16'(-780);
			11311: out = 16'(-14);
			11312: out = 16'(542);
			11313: out = 16'(-11);
			11314: out = 16'(81);
			11315: out = 16'(112);
			11316: out = 16'(-215);
			11317: out = 16'(15);
			11318: out = 16'(61);
			11319: out = 16'(239);
			11320: out = 16'(414);
			11321: out = 16'(-199);
			11322: out = 16'(-585);
			11323: out = 16'(-503);
			11324: out = 16'(-667);
			11325: out = 16'(-153);
			11326: out = 16'(634);
			11327: out = 16'(-161);
			11328: out = 16'(-972);
			11329: out = 16'(-563);
			11330: out = 16'(-402);
			11331: out = 16'(631);
			11332: out = 16'(1427);
			11333: out = 16'(609);
			11334: out = 16'(-702);
			11335: out = 16'(-1324);
			11336: out = 16'(-613);
			11337: out = 16'(194);
			11338: out = 16'(699);
			11339: out = 16'(295);
			11340: out = 16'(61);
			11341: out = 16'(521);
			11342: out = 16'(434);
			11343: out = 16'(-117);
			11344: out = 16'(-127);
			11345: out = 16'(-215);
			11346: out = 16'(83);
			11347: out = 16'(120);
			11348: out = 16'(246);
			11349: out = 16'(-87);
			11350: out = 16'(-212);
			11351: out = 16'(-214);
			11352: out = 16'(258);
			11353: out = 16'(600);
			11354: out = 16'(-26);
			11355: out = 16'(-735);
			11356: out = 16'(-243);
			11357: out = 16'(5);
			11358: out = 16'(-421);
			11359: out = 16'(-531);
			11360: out = 16'(-518);
			11361: out = 16'(370);
			11362: out = 16'(848);
			11363: out = 16'(811);
			11364: out = 16'(218);
			11365: out = 16'(-349);
			11366: out = 16'(-370);
			11367: out = 16'(-403);
			11368: out = 16'(-18);
			11369: out = 16'(67);
			11370: out = 16'(-574);
			11371: out = 16'(93);
			11372: out = 16'(917);
			11373: out = 16'(-68);
			11374: out = 16'(-803);
			11375: out = 16'(-566);
			11376: out = 16'(398);
			11377: out = 16'(553);
			11378: out = 16'(-196);
			11379: out = 16'(133);
			11380: out = 16'(384);
			11381: out = 16'(529);
			11382: out = 16'(561);
			11383: out = 16'(360);
			11384: out = 16'(-179);
			11385: out = 16'(-416);
			11386: out = 16'(-786);
			11387: out = 16'(-266);
			11388: out = 16'(312);
			11389: out = 16'(-229);
			11390: out = 16'(-983);
			11391: out = 16'(-678);
			11392: out = 16'(-273);
			11393: out = 16'(3);
			11394: out = 16'(631);
			11395: out = 16'(714);
			11396: out = 16'(-31);
			11397: out = 16'(-563);
			11398: out = 16'(-1133);
			11399: out = 16'(-681);
			11400: out = 16'(542);
			11401: out = 16'(1062);
			11402: out = 16'(536);
			11403: out = 16'(-260);
			11404: out = 16'(-666);
			11405: out = 16'(63);
			11406: out = 16'(847);
			11407: out = 16'(794);
			11408: out = 16'(163);
			11409: out = 16'(-455);
			11410: out = 16'(-598);
			11411: out = 16'(-575);
			11412: out = 16'(-128);
			11413: out = 16'(67);
			11414: out = 16'(-309);
			11415: out = 16'(-44);
			11416: out = 16'(69);
			11417: out = 16'(146);
			11418: out = 16'(194);
			11419: out = 16'(406);
			11420: out = 16'(789);
			11421: out = 16'(430);
			11422: out = 16'(-62);
			11423: out = 16'(-348);
			11424: out = 16'(-54);
			11425: out = 16'(347);
			11426: out = 16'(-32);
			11427: out = 16'(-434);
			11428: out = 16'(93);
			11429: out = 16'(139);
			11430: out = 16'(-407);
			11431: out = 16'(-450);
			11432: out = 16'(-496);
			11433: out = 16'(-174);
			11434: out = 16'(-222);
			11435: out = 16'(106);
			11436: out = 16'(456);
			11437: out = 16'(306);
			11438: out = 16'(283);
			11439: out = 16'(407);
			11440: out = 16'(-58);
			11441: out = 16'(-726);
			11442: out = 16'(-336);
			11443: out = 16'(219);
			11444: out = 16'(264);
			11445: out = 16'(-397);
			11446: out = 16'(-331);
			11447: out = 16'(163);
			11448: out = 16'(278);
			11449: out = 16'(204);
			11450: out = 16'(-236);
			11451: out = 16'(-278);
			11452: out = 16'(-54);
			11453: out = 16'(621);
			11454: out = 16'(547);
			11455: out = 16'(-277);
			11456: out = 16'(-798);
			11457: out = 16'(-72);
			11458: out = 16'(554);
			11459: out = 16'(395);
			11460: out = 16'(-690);
			11461: out = 16'(-523);
			11462: out = 16'(234);
			11463: out = 16'(181);
			11464: out = 16'(850);
			11465: out = 16'(1082);
			11466: out = 16'(328);
			11467: out = 16'(-928);
			11468: out = 16'(-1300);
			11469: out = 16'(-830);
			11470: out = 16'(360);
			11471: out = 16'(585);
			11472: out = 16'(-53);
			11473: out = 16'(-173);
			11474: out = 16'(136);
			11475: out = 16'(-188);
			11476: out = 16'(-354);
			11477: out = 16'(-782);
			11478: out = 16'(-535);
			11479: out = 16'(212);
			11480: out = 16'(778);
			11481: out = 16'(671);
			11482: out = 16'(-12);
			11483: out = 16'(52);
			11484: out = 16'(467);
			11485: out = 16'(457);
			11486: out = 16'(-503);
			11487: out = 16'(-1081);
			11488: out = 16'(-336);
			11489: out = 16'(438);
			11490: out = 16'(-23);
			11491: out = 16'(-568);
			11492: out = 16'(-360);
			11493: out = 16'(590);
			11494: out = 16'(856);
			11495: out = 16'(-10);
			11496: out = 16'(-251);
			11497: out = 16'(49);
			11498: out = 16'(462);
			11499: out = 16'(560);
			11500: out = 16'(362);
			11501: out = 16'(-48);
			11502: out = 16'(-562);
			11503: out = 16'(-994);
			11504: out = 16'(-753);
			11505: out = 16'(221);
			11506: out = 16'(605);
			11507: out = 16'(-346);
			11508: out = 16'(-781);
			11509: out = 16'(-108);
			11510: out = 16'(130);
			11511: out = 16'(338);
			11512: out = 16'(731);
			11513: out = 16'(690);
			11514: out = 16'(-335);
			11515: out = 16'(-882);
			11516: out = 16'(-642);
			11517: out = 16'(-24);
			11518: out = 16'(132);
			11519: out = 16'(-143);
			11520: out = 16'(-246);
			11521: out = 16'(152);
			11522: out = 16'(214);
			11523: out = 16'(-86);
			11524: out = 16'(-210);
			11525: out = 16'(-126);
			11526: out = 16'(282);
			11527: out = 16'(348);
			11528: out = 16'(-247);
			11529: out = 16'(-233);
			11530: out = 16'(-23);
			11531: out = 16'(308);
			11532: out = 16'(422);
			11533: out = 16'(-115);
			11534: out = 16'(-290);
			11535: out = 16'(-184);
			11536: out = 16'(412);
			11537: out = 16'(794);
			11538: out = 16'(327);
			11539: out = 16'(-544);
			11540: out = 16'(-836);
			11541: out = 16'(-464);
			11542: out = 16'(268);
			11543: out = 16'(607);
			11544: out = 16'(269);
			11545: out = 16'(-153);
			11546: out = 16'(-185);
			11547: out = 16'(-11);
			11548: out = 16'(-607);
			11549: out = 16'(-828);
			11550: out = 16'(-392);
			11551: out = 16'(195);
			11552: out = 16'(337);
			11553: out = 16'(540);
			11554: out = 16'(761);
			11555: out = 16'(315);
			11556: out = 16'(-367);
			11557: out = 16'(-790);
			11558: out = 16'(-643);
			11559: out = 16'(-219);
			11560: out = 16'(293);
			11561: out = 16'(482);
			11562: out = 16'(129);
			11563: out = 16'(186);
			11564: out = 16'(374);
			11565: out = 16'(485);
			11566: out = 16'(-170);
			11567: out = 16'(-603);
			11568: out = 16'(-655);
			11569: out = 16'(-133);
			11570: out = 16'(314);
			11571: out = 16'(27);
			11572: out = 16'(-493);
			11573: out = 16'(-424);
			11574: out = 16'(88);
			11575: out = 16'(278);
			11576: out = 16'(-240);
			11577: out = 16'(-731);
			11578: out = 16'(-562);
			11579: out = 16'(43);
			11580: out = 16'(331);
			11581: out = 16'(221);
			11582: out = 16'(-208);
			11583: out = 16'(-543);
			11584: out = 16'(-382);
			11585: out = 16'(-362);
			11586: out = 16'(128);
			11587: out = 16'(894);
			11588: out = 16'(523);
			11589: out = 16'(-190);
			11590: out = 16'(-538);
			11591: out = 16'(-254);
			11592: out = 16'(266);
			11593: out = 16'(-110);
			11594: out = 16'(-219);
			11595: out = 16'(13);
			11596: out = 16'(259);
			11597: out = 16'(126);
			11598: out = 16'(193);
			11599: out = 16'(165);
			11600: out = 16'(-382);
			11601: out = 16'(-718);
			11602: out = 16'(-441);
			11603: out = 16'(-156);
			11604: out = 16'(445);
			11605: out = 16'(365);
			11606: out = 16'(98);
			11607: out = 16'(-41);
			11608: out = 16'(-97);
			11609: out = 16'(140);
			11610: out = 16'(-297);
			11611: out = 16'(-602);
			11612: out = 16'(-236);
			11613: out = 16'(449);
			11614: out = 16'(429);
			11615: out = 16'(44);
			11616: out = 16'(113);
			11617: out = 16'(78);
			11618: out = 16'(-395);
			11619: out = 16'(-368);
			11620: out = 16'(-299);
			11621: out = 16'(-135);
			11622: out = 16'(-47);
			11623: out = 16'(-49);
			11624: out = 16'(-30);
			11625: out = 16'(-91);
			11626: out = 16'(399);
			11627: out = 16'(517);
			11628: out = 16'(-293);
			11629: out = 16'(-1000);
			11630: out = 16'(-810);
			11631: out = 16'(-313);
			11632: out = 16'(394);
			11633: out = 16'(545);
			11634: out = 16'(139);
			11635: out = 16'(-348);
			11636: out = 16'(-564);
			11637: out = 16'(34);
			11638: out = 16'(163);
			11639: out = 16'(483);
			11640: out = 16'(40);
			11641: out = 16'(-315);
			11642: out = 16'(-352);
			11643: out = 16'(-53);
			11644: out = 16'(402);
			11645: out = 16'(216);
			11646: out = 16'(-129);
			11647: out = 16'(183);
			11648: out = 16'(180);
			11649: out = 16'(-109);
			11650: out = 16'(-371);
			11651: out = 16'(-485);
			11652: out = 16'(-439);
			11653: out = 16'(-587);
			11654: out = 16'(-107);
			11655: out = 16'(416);
			11656: out = 16'(-47);
			11657: out = 16'(-202);
			11658: out = 16'(297);
			11659: out = 16'(56);
			11660: out = 16'(-709);
			11661: out = 16'(-1111);
			11662: out = 16'(-521);
			11663: out = 16'(-30);
			11664: out = 16'(510);
			11665: out = 16'(533);
			11666: out = 16'(-122);
			11667: out = 16'(-93);
			11668: out = 16'(-187);
			11669: out = 16'(254);
			11670: out = 16'(284);
			11671: out = 16'(19);
			11672: out = 16'(-10);
			11673: out = 16'(-180);
			11674: out = 16'(-152);
			11675: out = 16'(37);
			11676: out = 16'(-12);
			11677: out = 16'(-533);
			11678: out = 16'(-475);
			11679: out = 16'(-191);
			11680: out = 16'(-211);
			11681: out = 16'(98);
			11682: out = 16'(420);
			11683: out = 16'(-31);
			11684: out = 16'(-228);
			11685: out = 16'(34);
			11686: out = 16'(-123);
			11687: out = 16'(169);
			11688: out = 16'(-231);
			11689: out = 16'(-57);
			11690: out = 16'(180);
			11691: out = 16'(142);
			11692: out = 16'(469);
			11693: out = 16'(446);
			11694: out = 16'(36);
			11695: out = 16'(-566);
			11696: out = 16'(-562);
			11697: out = 16'(-647);
			11698: out = 16'(-62);
			11699: out = 16'(173);
			11700: out = 16'(48);
			11701: out = 16'(240);
			11702: out = 16'(280);
			11703: out = 16'(26);
			11704: out = 16'(-211);
			11705: out = 16'(60);
			11706: out = 16'(99);
			11707: out = 16'(202);
			11708: out = 16'(-101);
			11709: out = 16'(-292);
			11710: out = 16'(159);
			11711: out = 16'(631);
			11712: out = 16'(294);
			11713: out = 16'(-193);
			11714: out = 16'(48);
			11715: out = 16'(239);
			11716: out = 16'(-140);
			11717: out = 16'(-337);
			11718: out = 16'(-318);
			11719: out = 16'(-217);
			11720: out = 16'(66);
			11721: out = 16'(-163);
			11722: out = 16'(-267);
			11723: out = 16'(164);
			11724: out = 16'(553);
			11725: out = 16'(282);
			11726: out = 16'(-431);
			11727: out = 16'(-461);
			11728: out = 16'(-24);
			11729: out = 16'(203);
			11730: out = 16'(-40);
			11731: out = 16'(289);
			11732: out = 16'(665);
			11733: out = 16'(296);
			11734: out = 16'(-453);
			11735: out = 16'(-573);
			11736: out = 16'(-66);
			11737: out = 16'(611);
			11738: out = 16'(88);
			11739: out = 16'(-529);
			11740: out = 16'(-203);
			11741: out = 16'(57);
			11742: out = 16'(-417);
			11743: out = 16'(-671);
			11744: out = 16'(-299);
			default: out = 0;
		endcase
	end
endmodule
