module snare_lookup(index, out);
	input logic unsigned [13:0] index;
	output logic signed [23:0] out;
	always_comb begin
		case(index)
			0: out = 24'(75080);
			1: out = 24'(71960);
			2: out = 24'(94680);
			3: out = 24'(0);
			4: out = 24'(66908);
			5: out = 24'(71000);
			6: out = 24'(112024);
			7: out = 24'(33232);
			8: out = 24'(64);
			9: out = 24'(0);
			10: out = 24'(4);
			11: out = 24'(4);
			12: out = 24'(-85740);
			13: out = 24'(0);
			14: out = 24'(90664);
			15: out = 24'(4);
			16: out = 24'(8);
			17: out = 24'(64);
			18: out = 24'(99728);
			19: out = 24'(99792);
			20: out = 24'(94248);
			21: out = 24'(0);
			22: out = 24'(0);
			23: out = 24'(0);
			24: out = 24'(52);
			25: out = 24'(-276);
			26: out = 24'(-168);
			27: out = 24'(-764);
			28: out = 24'(-208);
			29: out = 24'(-3928);
			30: out = 24'(-10456);
			31: out = 24'(6588);
			32: out = 24'(28684);
			33: out = 24'(25496);
			34: out = 24'(1692);
			35: out = 24'(-2696);
			36: out = 24'(8732);
			37: out = 24'(17272);
			38: out = 24'(13260);
			39: out = 24'(-16292);
			40: out = 24'(-21628);
			41: out = 24'(3640);
			42: out = 24'(27884);
			43: out = 24'(7656);
			44: out = 24'(-37060);
			45: out = 24'(-23468);
			46: out = 24'(34944);
			47: out = 24'(39976);
			48: out = 24'(6072);
			49: out = 24'(-39548);
			50: out = 24'(-29612);
			51: out = 24'(8980);
			52: out = 24'(27484);
			53: out = 24'(34368);
			54: out = 24'(14588);
			55: out = 24'(-2464);
			56: out = 24'(-17464);
			57: out = 24'(6596);
			58: out = 24'(55832);
			59: out = 24'(32476);
			60: out = 24'(-42736);
			61: out = 24'(-43136);
			62: out = 24'(-3400);
			63: out = 24'(-1732);
			64: out = 24'(-20696);
			65: out = 24'(-55988);
			66: out = 24'(-45316);
			67: out = 24'(22452);
			68: out = 24'(76336);
			69: out = 24'(64268);
			70: out = 24'(3904);
			71: out = 24'(-42064);
			72: out = 24'(-34724);
			73: out = 24'(6984);
			74: out = 24'(50324);
			75: out = 24'(39532);
			76: out = 24'(-30872);
			77: out = 24'(-27760);
			78: out = 24'(23012);
			79: out = 24'(-4488);
			80: out = 24'(-46232);
			81: out = 24'(-67972);
			82: out = 24'(-32900);
			83: out = 24'(26288);
			84: out = 24'(91124);
			85: out = 24'(31528);
			86: out = 24'(-28356);
			87: out = 24'(-15636);
			88: out = 24'(6188);
			89: out = 24'(37488);
			90: out = 24'(4384);
			91: out = 24'(6736);
			92: out = 24'(5900);
			93: out = 24'(4744);
			94: out = 24'(-7760);
			95: out = 24'(-7888);
			96: out = 24'(-47860);
			97: out = 24'(-71592);
			98: out = 24'(-54940);
			99: out = 24'(948);
			100: out = 24'(32380);
			101: out = 24'(-18800);
			102: out = 24'(-47340);
			103: out = 24'(-14872);
			104: out = 24'(48276);
			105: out = 24'(33064);
			106: out = 24'(-13456);
			107: out = 24'(-55040);
			108: out = 24'(-23720);
			109: out = 24'(5244);
			110: out = 24'(58220);
			111: out = 24'(128992);
			112: out = 24'(84208);
			113: out = 24'(-54576);
			114: out = 24'(-126840);
			115: out = 24'(-118500);
			116: out = 24'(-59076);
			117: out = 24'(100728);
			118: out = 24'(124804);
			119: out = 24'(125196);
			120: out = 24'(123192);
			121: out = 24'(124740);
			122: out = 24'(123424);
			123: out = 24'(121556);
			124: out = 24'(84876);
			125: out = 24'(119128);
			126: out = 24'(124764);
			127: out = 24'(123124);
			128: out = 24'(123672);
			129: out = 24'(122996);
			130: out = 24'(123404);
			131: out = 24'(121856);
			132: out = 24'(112648);
			133: out = 24'(123256);
			134: out = 24'(123160);
			135: out = 24'(122856);
			136: out = 24'(122780);
			137: out = 24'(122872);
			138: out = 24'(122256);
			139: out = 24'(122272);
			140: out = 24'(122400);
			141: out = 24'(122212);
			142: out = 24'(122020);
			143: out = 24'(122324);
			144: out = 24'(122228);
			145: out = 24'(121892);
			146: out = 24'(121944);
			147: out = 24'(121892);
			148: out = 24'(121684);
			149: out = 24'(121500);
			150: out = 24'(121284);
			151: out = 24'(121212);
			152: out = 24'(121456);
			153: out = 24'(121488);
			154: out = 24'(121172);
			155: out = 24'(120912);
			156: out = 24'(120888);
			157: out = 24'(120772);
			158: out = 24'(120756);
			159: out = 24'(120524);
			160: out = 24'(120472);
			161: out = 24'(120316);
			162: out = 24'(120468);
			163: out = 24'(120408);
			164: out = 24'(120264);
			165: out = 24'(120120);
			166: out = 24'(120032);
			167: out = 24'(119764);
			168: out = 24'(119672);
			169: out = 24'(119968);
			170: out = 24'(116044);
			171: out = 24'(96988);
			172: out = 24'(106480);
			173: out = 24'(121116);
			174: out = 24'(79584);
			175: out = 24'(32860);
			176: out = 24'(37132);
			177: out = 24'(70232);
			178: out = 24'(81120);
			179: out = 24'(18936);
			180: out = 24'(-28996);
			181: out = 24'(-15680);
			182: out = 24'(43580);
			183: out = 24'(43268);
			184: out = 24'(-30164);
			185: out = 24'(-44868);
			186: out = 24'(-17952);
			187: out = 24'(-10300);
			188: out = 24'(-59692);
			189: out = 24'(-76432);
			190: out = 24'(-61260);
			191: out = 24'(-62208);
			192: out = 24'(-100944);
			193: out = 24'(-107668);
			194: out = 24'(-110644);
			195: out = 24'(-124800);
			196: out = 24'(-124456);
			197: out = 24'(-125500);
			198: out = 24'(-124076);
			199: out = 24'(-125256);
			200: out = 24'(-123480);
			201: out = 24'(-125860);
			202: out = 24'(-113860);
			203: out = 24'(-104272);
			204: out = 24'(-106856);
			205: out = 24'(-107784);
			206: out = 24'(-122108);
			207: out = 24'(-124184);
			208: out = 24'(-123988);
			209: out = 24'(-124116);
			210: out = 24'(-123536);
			211: out = 24'(-123832);
			212: out = 24'(-122772);
			213: out = 24'(-124132);
			214: out = 24'(-122728);
			215: out = 24'(-124320);
			216: out = 24'(-121596);
			217: out = 24'(-124652);
			218: out = 24'(-89960);
			219: out = 24'(-84432);
			220: out = 24'(-123888);
			221: out = 24'(-121780);
			222: out = 24'(-123312);
			223: out = 24'(-121956);
			224: out = 24'(-122872);
			225: out = 24'(-121744);
			226: out = 24'(-113464);
			227: out = 24'(-114076);
			228: out = 24'(-112612);
			229: out = 24'(-77504);
			230: out = 24'(-50576);
			231: out = 24'(-94904);
			232: out = 24'(-121512);
			233: out = 24'(-123764);
			234: out = 24'(-99424);
			235: out = 24'(-69584);
			236: out = 24'(-96988);
			237: out = 24'(-102760);
			238: out = 24'(-64708);
			239: out = 24'(-29336);
			240: out = 24'(-26968);
			241: out = 24'(-36980);
			242: out = 24'(-63868);
			243: out = 24'(-54004);
			244: out = 24'(-20420);
			245: out = 24'(11960);
			246: out = 24'(45264);
			247: out = 24'(30744);
			248: out = 24'(-2388);
			249: out = 24'(10352);
			250: out = 24'(20404);
			251: out = 24'(10180);
			252: out = 24'(3496);
			253: out = 24'(9600);
			254: out = 24'(2432);
			255: out = 24'(54244);
			256: out = 24'(115504);
			257: out = 24'(77276);
			258: out = 24'(45216);
			259: out = 24'(36780);
			260: out = 24'(68140);
			261: out = 24'(113236);
			262: out = 24'(122700);
			263: out = 24'(122748);
			264: out = 24'(123576);
			265: out = 24'(95380);
			266: out = 24'(64064);
			267: out = 24'(70976);
			268: out = 24'(74964);
			269: out = 24'(70364);
			270: out = 24'(59632);
			271: out = 24'(93428);
			272: out = 24'(124196);
			273: out = 24'(121144);
			274: out = 24'(122920);
			275: out = 24'(121404);
			276: out = 24'(122688);
			277: out = 24'(117900);
			278: out = 24'(93472);
			279: out = 24'(93540);
			280: out = 24'(119496);
			281: out = 24'(121912);
			282: out = 24'(121624);
			283: out = 24'(121004);
			284: out = 24'(121464);
			285: out = 24'(119308);
			286: out = 24'(118288);
			287: out = 24'(122392);
			288: out = 24'(119796);
			289: out = 24'(120892);
			290: out = 24'(86392);
			291: out = 24'(90504);
			292: out = 24'(122172);
			293: out = 24'(112568);
			294: out = 24'(82368);
			295: out = 24'(82416);
			296: out = 24'(113092);
			297: out = 24'(119296);
			298: out = 24'(122036);
			299: out = 24'(113160);
			300: out = 24'(88620);
			301: out = 24'(64884);
			302: out = 24'(66732);
			303: out = 24'(73464);
			304: out = 24'(74660);
			305: out = 24'(108684);
			306: out = 24'(114208);
			307: out = 24'(58724);
			308: out = 24'(3780);
			309: out = 24'(15676);
			310: out = 24'(73928);
			311: out = 24'(78548);
			312: out = 24'(14800);
			313: out = 24'(516);
			314: out = 24'(30300);
			315: out = 24'(28296);
			316: out = 24'(-3128);
			317: out = 24'(5256);
			318: out = 24'(25400);
			319: out = 24'(55700);
			320: out = 24'(46420);
			321: out = 24'(24480);
			322: out = 24'(-7340);
			323: out = 24'(-16776);
			324: out = 24'(26644);
			325: out = 24'(83000);
			326: out = 24'(84800);
			327: out = 24'(18216);
			328: out = 24'(-20316);
			329: out = 24'(-10376);
			330: out = 24'(7084);
			331: out = 24'(-10808);
			332: out = 24'(-36728);
			333: out = 24'(-18596);
			334: out = 24'(20312);
			335: out = 24'(57248);
			336: out = 24'(39168);
			337: out = 24'(2044);
			338: out = 24'(-28908);
			339: out = 24'(-2008);
			340: out = 24'(28408);
			341: out = 24'(33976);
			342: out = 24'(30164);
			343: out = 24'(21820);
			344: out = 24'(-140);
			345: out = 24'(-25024);
			346: out = 24'(-38252);
			347: out = 24'(-38828);
			348: out = 24'(-52636);
			349: out = 24'(-44952);
			350: out = 24'(-2608);
			351: out = 24'(14856);
			352: out = 24'(50104);
			353: out = 24'(54324);
			354: out = 24'(50968);
			355: out = 24'(10508);
			356: out = 24'(-4088);
			357: out = 24'(19404);
			358: out = 24'(49252);
			359: out = 24'(87832);
			360: out = 24'(65132);
			361: out = 24'(10940);
			362: out = 24'(-15356);
			363: out = 24'(-13620);
			364: out = 24'(-6852);
			365: out = 24'(-20552);
			366: out = 24'(-29444);
			367: out = 24'(-8024);
			368: out = 24'(-4444);
			369: out = 24'(-5460);
			370: out = 24'(18660);
			371: out = 24'(53468);
			372: out = 24'(57648);
			373: out = 24'(-1956);
			374: out = 24'(-33548);
			375: out = 24'(-33600);
			376: out = 24'(-5432);
			377: out = 24'(12788);
			378: out = 24'(6156);
			379: out = 24'(-21196);
			380: out = 24'(-55260);
			381: out = 24'(-58380);
			382: out = 24'(-34568);
			383: out = 24'(-16472);
			384: out = 24'(1584);
			385: out = 24'(15204);
			386: out = 24'(-14500);
			387: out = 24'(-91476);
			388: out = 24'(-131060);
			389: out = 24'(-92812);
			390: out = 24'(-29428);
			391: out = 24'(-12244);
			392: out = 24'(-59856);
			393: out = 24'(-99984);
			394: out = 24'(-91100);
			395: out = 24'(-61412);
			396: out = 24'(6892);
			397: out = 24'(-3780);
			398: out = 24'(-63204);
			399: out = 24'(-103392);
			400: out = 24'(-89040);
			401: out = 24'(-58604);
			402: out = 24'(-62352);
			403: out = 24'(-98772);
			404: out = 24'(-118996);
			405: out = 24'(-126084);
			406: out = 24'(-114788);
			407: out = 24'(-93248);
			408: out = 24'(-116256);
			409: out = 24'(-111996);
			410: out = 24'(-73524);
			411: out = 24'(-64032);
			412: out = 24'(-111744);
			413: out = 24'(-119244);
			414: out = 24'(-85296);
			415: out = 24'(-92804);
			416: out = 24'(-123864);
			417: out = 24'(-119088);
			418: out = 24'(-100732);
			419: out = 24'(-100168);
			420: out = 24'(-118776);
			421: out = 24'(-122272);
			422: out = 24'(-124120);
			423: out = 24'(-79556);
			424: out = 24'(-79152);
			425: out = 24'(-125340);
			426: out = 24'(-120864);
			427: out = 24'(-125060);
			428: out = 24'(-120096);
			429: out = 24'(-119308);
			430: out = 24'(-85224);
			431: out = 24'(-83648);
			432: out = 24'(-120980);
			433: out = 24'(-122380);
			434: out = 24'(-122132);
			435: out = 24'(-105080);
			436: out = 24'(-74376);
			437: out = 24'(-101492);
			438: out = 24'(-124020);
			439: out = 24'(-121152);
			440: out = 24'(-122372);
			441: out = 24'(-120964);
			442: out = 24'(-121532);
			443: out = 24'(-121844);
			444: out = 24'(-117840);
			445: out = 24'(-74364);
			446: out = 24'(-46396);
			447: out = 24'(-100948);
			448: out = 24'(-122112);
			449: out = 24'(-122236);
			450: out = 24'(-110236);
			451: out = 24'(-113472);
			452: out = 24'(-116312);
			453: out = 24'(-86728);
			454: out = 24'(-86036);
			455: out = 24'(-109260);
			456: out = 24'(-122024);
			457: out = 24'(-120220);
			458: out = 24'(-116192);
			459: out = 24'(-74872);
			460: out = 24'(-38028);
			461: out = 24'(-81152);
			462: out = 24'(-123340);
			463: out = 24'(-118548);
			464: out = 24'(-117636);
			465: out = 24'(-62280);
			466: out = 24'(-44784);
			467: out = 24'(-97120);
			468: out = 24'(-121228);
			469: out = 24'(-119196);
			470: out = 24'(-98488);
			471: out = 24'(-68736);
			472: out = 24'(-70688);
			473: out = 24'(-94916);
			474: out = 24'(-85668);
			475: out = 24'(-26556);
			476: out = 24'(-43372);
			477: out = 24'(-109000);
			478: out = 24'(-121044);
			479: out = 24'(-103908);
			480: out = 24'(-50948);
			481: out = 24'(-2372);
			482: out = 24'(2512);
			483: out = 24'(-44756);
			484: out = 24'(-82796);
			485: out = 24'(-107088);
			486: out = 24'(-98648);
			487: out = 24'(-35264);
			488: out = 24'(10444);
			489: out = 24'(-12736);
			490: out = 24'(-18252);
			491: out = 24'(-9688);
			492: out = 24'(-18716);
			493: out = 24'(-22512);
			494: out = 24'(-41288);
			495: out = 24'(-38412);
			496: out = 24'(14356);
			497: out = 24'(60948);
			498: out = 24'(10944);
			499: out = 24'(-38300);
			500: out = 24'(4624);
			501: out = 24'(49604);
			502: out = 24'(30772);
			503: out = 24'(25248);
			504: out = 24'(57520);
			505: out = 24'(48688);
			506: out = 24'(19304);
			507: out = 24'(32004);
			508: out = 24'(39372);
			509: out = 24'(78168);
			510: out = 24'(83096);
			511: out = 24'(62852);
			512: out = 24'(93084);
			513: out = 24'(114584);
			514: out = 24'(120604);
			515: out = 24'(92792);
			516: out = 24'(79156);
			517: out = 24'(89940);
			518: out = 24'(87492);
			519: out = 24'(109044);
			520: out = 24'(125992);
			521: out = 24'(121968);
			522: out = 24'(110088);
			523: out = 24'(118252);
			524: out = 24'(115352);
			525: out = 24'(85924);
			526: out = 24'(82068);
			527: out = 24'(87440);
			528: out = 24'(108424);
			529: out = 24'(125728);
			530: out = 24'(123552);
			531: out = 24'(121716);
			532: out = 24'(109272);
			533: out = 24'(122832);
			534: out = 24'(123440);
			535: out = 24'(123784);
			536: out = 24'(123440);
			537: out = 24'(123740);
			538: out = 24'(123040);
			539: out = 24'(123328);
			540: out = 24'(122896);
			541: out = 24'(123064);
			542: out = 24'(122900);
			543: out = 24'(122892);
			544: out = 24'(122688);
			545: out = 24'(122708);
			546: out = 24'(122560);
			547: out = 24'(122520);
			548: out = 24'(122312);
			549: out = 24'(122120);
			550: out = 24'(122380);
			551: out = 24'(121900);
			552: out = 24'(122596);
			553: out = 24'(114952);
			554: out = 24'(87908);
			555: out = 24'(98708);
			556: out = 24'(123676);
			557: out = 24'(120276);
			558: out = 24'(123252);
			559: out = 24'(111684);
			560: out = 24'(85192);
			561: out = 24'(106452);
			562: out = 24'(123048);
			563: out = 24'(119832);
			564: out = 24'(122864);
			565: out = 24'(110944);
			566: out = 24'(107228);
			567: out = 24'(123568);
			568: out = 24'(118444);
			569: out = 24'(123580);
			570: out = 24'(107244);
			571: out = 24'(92528);
			572: out = 24'(117612);
			573: out = 24'(120000);
			574: out = 24'(120568);
			575: out = 24'(119560);
			576: out = 24'(120428);
			577: out = 24'(119424);
			578: out = 24'(120476);
			579: out = 24'(118876);
			580: out = 24'(120324);
			581: out = 24'(92688);
			582: out = 24'(72980);
			583: out = 24'(88780);
			584: out = 24'(93132);
			585: out = 24'(75436);
			586: out = 24'(72880);
			587: out = 24'(89456);
			588: out = 24'(76352);
			589: out = 24'(41344);
			590: out = 24'(37200);
			591: out = 24'(52212);
			592: out = 24'(99516);
			593: out = 24'(120924);
			594: out = 24'(114236);
			595: out = 24'(68116);
			596: out = 24'(38340);
			597: out = 24'(54192);
			598: out = 24'(101800);
			599: out = 24'(92076);
			600: out = 24'(60876);
			601: out = 24'(69308);
			602: out = 24'(80120);
			603: out = 24'(60572);
			604: out = 24'(26356);
			605: out = 24'(14256);
			606: out = 24'(44704);
			607: out = 24'(76556);
			608: out = 24'(40976);
			609: out = 24'(17188);
			610: out = 24'(26496);
			611: out = 24'(83252);
			612: out = 24'(62360);
			613: out = 24'(13240);
			614: out = 24'(26888);
			615: out = 24'(48092);
			616: out = 24'(38632);
			617: out = 24'(38876);
			618: out = 24'(54308);
			619: out = 24'(48948);
			620: out = 24'(-11248);
			621: out = 24'(-48156);
			622: out = 24'(-24688);
			623: out = 24'(4248);
			624: out = 24'(12612);
			625: out = 24'(-18288);
			626: out = 24'(-30252);
			627: out = 24'(-33384);
			628: out = 24'(-17312);
			629: out = 24'(-7072);
			630: out = 24'(-12160);
			631: out = 24'(11648);
			632: out = 24'(-1964);
			633: out = 24'(-10104);
			634: out = 24'(-25284);
			635: out = 24'(-49008);
			636: out = 24'(-41748);
			637: out = 24'(-30088);
			638: out = 24'(-21464);
			639: out = 24'(-51732);
			640: out = 24'(-57104);
			641: out = 24'(-36816);
			642: out = 24'(-33940);
			643: out = 24'(-94588);
			644: out = 24'(-129028);
			645: out = 24'(-119616);
			646: out = 24'(-64204);
			647: out = 24'(-39664);
			648: out = 24'(-102068);
			649: out = 24'(-128656);
			650: out = 24'(-104236);
			651: out = 24'(-62792);
			652: out = 24'(-72144);
			653: out = 24'(-110672);
			654: out = 24'(-127252);
			655: out = 24'(-124560);
			656: out = 24'(-126100);
			657: out = 24'(-125328);
			658: out = 24'(-124796);
			659: out = 24'(-120340);
			660: out = 24'(-108388);
			661: out = 24'(-107880);
			662: out = 24'(-95852);
			663: out = 24'(-116308);
			664: out = 24'(-126728);
			665: out = 24'(-124140);
			666: out = 24'(-119448);
			667: out = 24'(-101500);
			668: out = 24'(-113840);
			669: out = 24'(-124588);
			670: out = 24'(-124532);
			671: out = 24'(-123980);
			672: out = 24'(-124540);
			673: out = 24'(-124024);
			674: out = 24'(-124188);
			675: out = 24'(-123616);
			676: out = 24'(-124036);
			677: out = 24'(-122088);
			678: out = 24'(-118288);
			679: out = 24'(-123864);
			680: out = 24'(-123468);
			681: out = 24'(-123368);
			682: out = 24'(-123008);
			683: out = 24'(-123100);
			684: out = 24'(-122868);
			685: out = 24'(-122812);
			686: out = 24'(-123120);
			687: out = 24'(-123016);
			688: out = 24'(-122564);
			689: out = 24'(-120744);
			690: out = 24'(-116156);
			691: out = 24'(-121768);
			692: out = 24'(-122016);
			693: out = 24'(-123156);
			694: out = 24'(-121300);
			695: out = 24'(-123264);
			696: out = 24'(-112104);
			697: out = 24'(-116384);
			698: out = 24'(-123312);
			699: out = 24'(-114944);
			700: out = 24'(-120256);
			701: out = 24'(-121904);
			702: out = 24'(-121380);
			703: out = 24'(-121676);
			704: out = 24'(-119668);
			705: out = 24'(-116408);
			706: out = 24'(-121444);
			707: out = 24'(-120712);
			708: out = 24'(-121124);
			709: out = 24'(-120844);
			710: out = 24'(-120668);
			711: out = 24'(-120856);
			712: out = 24'(-120608);
			713: out = 24'(-120356);
			714: out = 24'(-119832);
			715: out = 24'(-120844);
			716: out = 24'(-105944);
			717: out = 24'(-64532);
			718: out = 24'(-77172);
			719: out = 24'(-118324);
			720: out = 24'(-119336);
			721: out = 24'(-118588);
			722: out = 24'(-88440);
			723: out = 24'(-93200);
			724: out = 24'(-119196);
			725: out = 24'(-109144);
			726: out = 24'(-93732);
			727: out = 24'(-108964);
			728: out = 24'(-122604);
			729: out = 24'(-107592);
			730: out = 24'(-53056);
			731: out = 24'(-52920);
			732: out = 24'(-104188);
			733: out = 24'(-89676);
			734: out = 24'(-63920);
			735: out = 24'(-87736);
			736: out = 24'(-72076);
			737: out = 24'(-43184);
			738: out = 24'(-40540);
			739: out = 24'(-67364);
			740: out = 24'(-66696);
			741: out = 24'(-50932);
			742: out = 24'(9236);
			743: out = 24'(20416);
			744: out = 24'(-37656);
			745: out = 24'(-79820);
			746: out = 24'(-40264);
			747: out = 24'(9784);
			748: out = 24'(-1112);
			749: out = 24'(15740);
			750: out = 24'(40428);
			751: out = 24'(19124);
			752: out = 24'(-832);
			753: out = 24'(10520);
			754: out = 24'(-10756);
			755: out = 24'(-8652);
			756: out = 24'(25880);
			757: out = 24'(30360);
			758: out = 24'(52920);
			759: out = 24'(59504);
			760: out = 24'(52040);
			761: out = 24'(43300);
			762: out = 24'(33388);
			763: out = 24'(36632);
			764: out = 24'(36236);
			765: out = 24'(40792);
			766: out = 24'(39344);
			767: out = 24'(78068);
			768: out = 24'(91280);
			769: out = 24'(56332);
			770: out = 24'(37508);
			771: out = 24'(63644);
			772: out = 24'(100184);
			773: out = 24'(118196);
			774: out = 24'(102268);
			775: out = 24'(68732);
			776: out = 24'(37660);
			777: out = 24'(17444);
			778: out = 24'(3476);
			779: out = 24'(10468);
			780: out = 24'(72628);
			781: out = 24'(112520);
			782: out = 24'(58144);
			783: out = 24'(38168);
			784: out = 24'(93256);
			785: out = 24'(108896);
			786: out = 24'(48136);
			787: out = 24'(38724);
			788: out = 24'(73372);
			789: out = 24'(66864);
			790: out = 24'(91540);
			791: out = 24'(105444);
			792: out = 24'(87012);
			793: out = 24'(101624);
			794: out = 24'(117096);
			795: out = 24'(115660);
			796: out = 24'(91232);
			797: out = 24'(47468);
			798: out = 24'(40484);
			799: out = 24'(47376);
			800: out = 24'(72972);
			801: out = 24'(110248);
			802: out = 24'(124516);
			803: out = 24'(122984);
			804: out = 24'(124920);
			805: out = 24'(113456);
			806: out = 24'(92836);
			807: out = 24'(83872);
			808: out = 24'(76192);
			809: out = 24'(96488);
			810: out = 24'(99460);
			811: out = 24'(97032);
			812: out = 24'(124704);
			813: out = 24'(104728);
			814: out = 24'(75188);
			815: out = 24'(89068);
			816: out = 24'(114036);
			817: out = 24'(125152);
			818: out = 24'(98100);
			819: out = 24'(51916);
			820: out = 24'(61900);
			821: out = 24'(117668);
			822: out = 24'(114436);
			823: out = 24'(82068);
			824: out = 24'(92200);
			825: out = 24'(111196);
			826: out = 24'(95500);
			827: out = 24'(66420);
			828: out = 24'(85620);
			829: out = 24'(122636);
			830: out = 24'(108840);
			831: out = 24'(52868);
			832: out = 24'(27664);
			833: out = 24'(59808);
			834: out = 24'(90416);
			835: out = 24'(59192);
			836: out = 24'(11828);
			837: out = 24'(41512);
			838: out = 24'(88048);
			839: out = 24'(99372);
			840: out = 24'(80688);
			841: out = 24'(70568);
			842: out = 24'(54260);
			843: out = 24'(34748);
			844: out = 24'(70644);
			845: out = 24'(73236);
			846: out = 24'(36796);
			847: out = 24'(58980);
			848: out = 24'(105664);
			849: out = 24'(101020);
			850: out = 24'(26296);
			851: out = 24'(-16596);
			852: out = 24'(42304);
			853: out = 24'(112120);
			854: out = 24'(117800);
			855: out = 24'(79740);
			856: out = 24'(46932);
			857: out = 24'(28856);
			858: out = 24'(17184);
			859: out = 24'(4424);
			860: out = 24'(42864);
			861: out = 24'(82232);
			862: out = 24'(59240);
			863: out = 24'(52448);
			864: out = 24'(54740);
			865: out = 24'(52288);
			866: out = 24'(25832);
			867: out = 24'(-11520);
			868: out = 24'(-9584);
			869: out = 24'(9716);
			870: out = 24'(30028);
			871: out = 24'(39392);
			872: out = 24'(32392);
			873: out = 24'(11488);
			874: out = 24'(5924);
			875: out = 24'(6448);
			876: out = 24'(40200);
			877: out = 24'(25152);
			878: out = 24'(-27456);
			879: out = 24'(-50368);
			880: out = 24'(-39776);
			881: out = 24'(-27148);
			882: out = 24'(-13816);
			883: out = 24'(-33928);
			884: out = 24'(-46668);
			885: out = 24'(-32308);
			886: out = 24'(-11648);
			887: out = 24'(27428);
			888: out = 24'(71960);
			889: out = 24'(55568);
			890: out = 24'(-22268);
			891: out = 24'(-74472);
			892: out = 24'(-76860);
			893: out = 24'(-43008);
			894: out = 24'(-38828);
			895: out = 24'(-50756);
			896: out = 24'(-15864);
			897: out = 24'(-248);
			898: out = 24'(26960);
			899: out = 24'(44148);
			900: out = 24'(4516);
			901: out = 24'(-28884);
			902: out = 24'(-52632);
			903: out = 24'(-66608);
			904: out = 24'(-61600);
			905: out = 24'(-25172);
			906: out = 24'(-15264);
			907: out = 24'(-25172);
			908: out = 24'(-57724);
			909: out = 24'(-80788);
			910: out = 24'(-19576);
			911: out = 24'(45228);
			912: out = 24'(22232);
			913: out = 24'(-62312);
			914: out = 24'(-97996);
			915: out = 24'(-100316);
			916: out = 24'(-15660);
			917: out = 24'(53580);
			918: out = 24'(-8264);
			919: out = 24'(-56140);
			920: out = 24'(-48328);
			921: out = 24'(-9576);
			922: out = 24'(22256);
			923: out = 24'(-8556);
			924: out = 24'(-37752);
			925: out = 24'(-41388);
			926: out = 24'(-31016);
			927: out = 24'(6108);
			928: out = 24'(5468);
			929: out = 24'(-63492);
			930: out = 24'(-112272);
			931: out = 24'(-94112);
			932: out = 24'(-45952);
			933: out = 24'(-23676);
			934: out = 24'(-55764);
			935: out = 24'(-93928);
			936: out = 24'(-78340);
			937: out = 24'(-12720);
			938: out = 24'(5292);
			939: out = 24'(13432);
			940: out = 24'(7684);
			941: out = 24'(-49412);
			942: out = 24'(-88704);
			943: out = 24'(-110836);
			944: out = 24'(-53472);
			945: out = 24'(9276);
			946: out = 24'(-8840);
			947: out = 24'(-36896);
			948: out = 24'(-58388);
			949: out = 24'(-63164);
			950: out = 24'(-47856);
			951: out = 24'(-65640);
			952: out = 24'(-65444);
			953: out = 24'(-17708);
			954: out = 24'(9236);
			955: out = 24'(-52760);
			956: out = 24'(-95208);
			957: out = 24'(-80328);
			958: out = 24'(-46312);
			959: out = 24'(-14428);
			960: out = 24'(-1340);
			961: out = 24'(-31756);
			962: out = 24'(-46456);
			963: out = 24'(-57888);
			964: out = 24'(-68816);
			965: out = 24'(-71980);
			966: out = 24'(-80728);
			967: out = 24'(-82340);
			968: out = 24'(-53920);
			969: out = 24'(-22200);
			970: out = 24'(-15964);
			971: out = 24'(-70616);
			972: out = 24'(-77188);
			973: out = 24'(-8984);
			974: out = 24'(-3440);
			975: out = 24'(-58660);
			976: out = 24'(-85988);
			977: out = 24'(-56780);
			978: out = 24'(-47644);
			979: out = 24'(-70632);
			980: out = 24'(-58992);
			981: out = 24'(-34372);
			982: out = 24'(-22008);
			983: out = 24'(-52052);
			984: out = 24'(-59260);
			985: out = 24'(-42956);
			986: out = 24'(-24596);
			987: out = 24'(12964);
			988: out = 24'(-880);
			989: out = 24'(-67060);
			990: out = 24'(-115588);
			991: out = 24'(-96392);
			992: out = 24'(-71720);
			993: out = 24'(-15376);
			994: out = 24'(24464);
			995: out = 24'(-15812);
			996: out = 24'(-50288);
			997: out = 24'(-69560);
			998: out = 24'(-70748);
			999: out = 24'(-36152);
			1000: out = 24'(-33788);
			1001: out = 24'(-45608);
			1002: out = 24'(-68132);
			1003: out = 24'(-30204);
			1004: out = 24'(7624);
			1005: out = 24'(-52180);
			1006: out = 24'(-98892);
			1007: out = 24'(-73924);
			1008: out = 24'(-56676);
			1009: out = 24'(-50588);
			1010: out = 24'(-8928);
			1011: out = 24'(10488);
			1012: out = 24'(-75852);
			1013: out = 24'(-124812);
			1014: out = 24'(-103764);
			1015: out = 24'(-53436);
			1016: out = 24'(31032);
			1017: out = 24'(33552);
			1018: out = 24'(-66912);
			1019: out = 24'(-116864);
			1020: out = 24'(-108220);
			1021: out = 24'(-44480);
			1022: out = 24'(12128);
			1023: out = 24'(-17812);
			1024: out = 24'(-83068);
			1025: out = 24'(-93748);
			1026: out = 24'(-70268);
			1027: out = 24'(-32476);
			1028: out = 24'(-28656);
			1029: out = 24'(-54232);
			1030: out = 24'(-87916);
			1031: out = 24'(-75464);
			1032: out = 24'(-21344);
			1033: out = 24'(-2052);
			1034: out = 24'(-26648);
			1035: out = 24'(-44532);
			1036: out = 24'(-51424);
			1037: out = 24'(-55788);
			1038: out = 24'(-34000);
			1039: out = 24'(-34360);
			1040: out = 24'(-64972);
			1041: out = 24'(-98636);
			1042: out = 24'(-85256);
			1043: out = 24'(-62688);
			1044: out = 24'(-42008);
			1045: out = 24'(-62308);
			1046: out = 24'(-85964);
			1047: out = 24'(-61896);
			1048: out = 24'(-40848);
			1049: out = 24'(-3352);
			1050: out = 24'(-17768);
			1051: out = 24'(-23540);
			1052: out = 24'(-34528);
			1053: out = 24'(-18820);
			1054: out = 24'(-35804);
			1055: out = 24'(-53980);
			1056: out = 24'(-42732);
			1057: out = 24'(-26864);
			1058: out = 24'(-17692);
			1059: out = 24'(-19268);
			1060: out = 24'(-5304);
			1061: out = 24'(-9444);
			1062: out = 24'(-48080);
			1063: out = 24'(-74504);
			1064: out = 24'(-53576);
			1065: out = 24'(-33320);
			1066: out = 24'(-23860);
			1067: out = 24'(508);
			1068: out = 24'(1432);
			1069: out = 24'(-49648);
			1070: out = 24'(-89244);
			1071: out = 24'(-34248);
			1072: out = 24'(62880);
			1073: out = 24'(53984);
			1074: out = 24'(-5948);
			1075: out = 24'(-26720);
			1076: out = 24'(-43004);
			1077: out = 24'(-16276);
			1078: out = 24'(14928);
			1079: out = 24'(21444);
			1080: out = 24'(25420);
			1081: out = 24'(-6940);
			1082: out = 24'(-8528);
			1083: out = 24'(-15776);
			1084: out = 24'(-41360);
			1085: out = 24'(23852);
			1086: out = 24'(70012);
			1087: out = 24'(27132);
			1088: out = 24'(-22364);
			1089: out = 24'(-11604);
			1090: out = 24'(20240);
			1091: out = 24'(8084);
			1092: out = 24'(6056);
			1093: out = 24'(27304);
			1094: out = 24'(14224);
			1095: out = 24'(2116);
			1096: out = 24'(-592);
			1097: out = 24'(13312);
			1098: out = 24'(16060);
			1099: out = 24'(35056);
			1100: out = 24'(54312);
			1101: out = 24'(29064);
			1102: out = 24'(2964);
			1103: out = 24'(6428);
			1104: out = 24'(27784);
			1105: out = 24'(55324);
			1106: out = 24'(40764);
			1107: out = 24'(7308);
			1108: out = 24'(22664);
			1109: out = 24'(31580);
			1110: out = 24'(62240);
			1111: out = 24'(62300);
			1112: out = 24'(6632);
			1113: out = 24'(11636);
			1114: out = 24'(23960);
			1115: out = 24'(18040);
			1116: out = 24'(23488);
			1117: out = 24'(7744);
			1118: out = 24'(-5596);
			1119: out = 24'(-2216);
			1120: out = 24'(3776);
			1121: out = 24'(-9844);
			1122: out = 24'(21304);
			1123: out = 24'(40436);
			1124: out = 24'(47392);
			1125: out = 24'(69696);
			1126: out = 24'(70344);
			1127: out = 24'(36960);
			1128: out = 24'(-22328);
			1129: out = 24'(-41792);
			1130: out = 24'(-20352);
			1131: out = 24'(43904);
			1132: out = 24'(46148);
			1133: out = 24'(19600);
			1134: out = 24'(49132);
			1135: out = 24'(49312);
			1136: out = 24'(13184);
			1137: out = 24'(42492);
			1138: out = 24'(45732);
			1139: out = 24'(24300);
			1140: out = 24'(26604);
			1141: out = 24'(53788);
			1142: out = 24'(45132);
			1143: out = 24'(2680);
			1144: out = 24'(-19332);
			1145: out = 24'(9952);
			1146: out = 24'(49880);
			1147: out = 24'(62596);
			1148: out = 24'(39768);
			1149: out = 24'(23184);
			1150: out = 24'(-4032);
			1151: out = 24'(-4948);
			1152: out = 24'(-5932);
			1153: out = 24'(13308);
			1154: out = 24'(78864);
			1155: out = 24'(86816);
			1156: out = 24'(52224);
			1157: out = 24'(43076);
			1158: out = 24'(44904);
			1159: out = 24'(56564);
			1160: out = 24'(21700);
			1161: out = 24'(-4820);
			1162: out = 24'(424);
			1163: out = 24'(24360);
			1164: out = 24'(58220);
			1165: out = 24'(79336);
			1166: out = 24'(29016);
			1167: out = 24'(-6856);
			1168: out = 24'(-6196);
			1169: out = 24'(25116);
			1170: out = 24'(59592);
			1171: out = 24'(57284);
			1172: out = 24'(18876);
			1173: out = 24'(-18244);
			1174: out = 24'(13780);
			1175: out = 24'(65124);
			1176: out = 24'(73116);
			1177: out = 24'(13992);
			1178: out = 24'(3628);
			1179: out = 24'(38704);
			1180: out = 24'(80916);
			1181: out = 24'(67900);
			1182: out = 24'(19320);
			1183: out = 24'(-10552);
			1184: out = 24'(1388);
			1185: out = 24'(15740);
			1186: out = 24'(24152);
			1187: out = 24'(11668);
			1188: out = 24'(-9040);
			1189: out = 24'(4548);
			1190: out = 24'(41116);
			1191: out = 24'(89416);
			1192: out = 24'(112248);
			1193: out = 24'(96148);
			1194: out = 24'(18856);
			1195: out = 24'(-45256);
			1196: out = 24'(-50212);
			1197: out = 24'(1552);
			1198: out = 24'(109288);
			1199: out = 24'(120572);
			1200: out = 24'(46892);
			1201: out = 24'(26012);
			1202: out = 24'(68460);
			1203: out = 24'(115068);
			1204: out = 24'(89940);
			1205: out = 24'(24136);
			1206: out = 24'(26464);
			1207: out = 24'(32484);
			1208: out = 24'(17288);
			1209: out = 24'(38000);
			1210: out = 24'(51072);
			1211: out = 24'(24608);
			1212: out = 24'(43844);
			1213: out = 24'(41844);
			1214: out = 24'(28440);
			1215: out = 24'(48260);
			1216: out = 24'(61940);
			1217: out = 24'(92900);
			1218: out = 24'(97332);
			1219: out = 24'(81756);
			1220: out = 24'(67856);
			1221: out = 24'(35856);
			1222: out = 24'(20548);
			1223: out = 24'(10740);
			1224: out = 24'(-15436);
			1225: out = 24'(1776);
			1226: out = 24'(49620);
			1227: out = 24'(91800);
			1228: out = 24'(71872);
			1229: out = 24'(59376);
			1230: out = 24'(96084);
			1231: out = 24'(68920);
			1232: out = 24'(14936);
			1233: out = 24'(-5924);
			1234: out = 24'(28840);
			1235: out = 24'(43108);
			1236: out = 24'(47824);
			1237: out = 24'(65860);
			1238: out = 24'(59780);
			1239: out = 24'(62196);
			1240: out = 24'(61036);
			1241: out = 24'(32976);
			1242: out = 24'(-992);
			1243: out = 24'(-26356);
			1244: out = 24'(19132);
			1245: out = 24'(106184);
			1246: out = 24'(106816);
			1247: out = 24'(1144);
			1248: out = 24'(-31552);
			1249: out = 24'(17912);
			1250: out = 24'(63384);
			1251: out = 24'(72148);
			1252: out = 24'(24920);
			1253: out = 24'(-8840);
			1254: out = 24'(-19876);
			1255: out = 24'(-3196);
			1256: out = 24'(40832);
			1257: out = 24'(78908);
			1258: out = 24'(29056);
			1259: out = 24'(-23900);
			1260: out = 24'(10756);
			1261: out = 24'(24320);
			1262: out = 24'(33304);
			1263: out = 24'(38984);
			1264: out = 24'(9244);
			1265: out = 24'(-1912);
			1266: out = 24'(12576);
			1267: out = 24'(44264);
			1268: out = 24'(53676);
			1269: out = 24'(21464);
			1270: out = 24'(-12500);
			1271: out = 24'(-25264);
			1272: out = 24'(-25384);
			1273: out = 24'(-584);
			1274: out = 24'(-5040);
			1275: out = 24'(-8904);
			1276: out = 24'(58276);
			1277: out = 24'(95560);
			1278: out = 24'(-2600);
			1279: out = 24'(-91484);
			1280: out = 24'(-80872);
			1281: out = 24'(-22400);
			1282: out = 24'(40696);
			1283: out = 24'(83616);
			1284: out = 24'(46036);
			1285: out = 24'(-44004);
			1286: out = 24'(-71656);
			1287: out = 24'(-29760);
			1288: out = 24'(20148);
			1289: out = 24'(34084);
			1290: out = 24'(-4456);
			1291: out = 24'(-38100);
			1292: out = 24'(-43084);
			1293: out = 24'(-32324);
			1294: out = 24'(-448);
			1295: out = 24'(40388);
			1296: out = 24'(4884);
			1297: out = 24'(-57632);
			1298: out = 24'(-27524);
			1299: out = 24'(-20092);
			1300: out = 24'(20400);
			1301: out = 24'(15464);
			1302: out = 24'(-14700);
			1303: out = 24'(-18416);
			1304: out = 24'(-8216);
			1305: out = 24'(-17040);
			1306: out = 24'(-35940);
			1307: out = 24'(-49228);
			1308: out = 24'(-61692);
			1309: out = 24'(-36816);
			1310: out = 24'(3276);
			1311: out = 24'(-10520);
			1312: out = 24'(-54132);
			1313: out = 24'(-95292);
			1314: out = 24'(-110968);
			1315: out = 24'(-69932);
			1316: out = 24'(440);
			1317: out = 24'(1984);
			1318: out = 24'(-78400);
			1319: out = 24'(-105648);
			1320: out = 24'(-81316);
			1321: out = 24'(-47652);
			1322: out = 24'(16948);
			1323: out = 24'(-2932);
			1324: out = 24'(-50376);
			1325: out = 24'(-81052);
			1326: out = 24'(-63992);
			1327: out = 24'(-15528);
			1328: out = 24'(-17312);
			1329: out = 24'(-57496);
			1330: out = 24'(-48928);
			1331: out = 24'(-34684);
			1332: out = 24'(-76572);
			1333: out = 24'(-103032);
			1334: out = 24'(-82752);
			1335: out = 24'(-23432);
			1336: out = 24'(-50028);
			1337: out = 24'(-116064);
			1338: out = 24'(-89872);
			1339: out = 24'(-52236);
			1340: out = 24'(-66180);
			1341: out = 24'(-80588);
			1342: out = 24'(-72676);
			1343: out = 24'(-63540);
			1344: out = 24'(-33832);
			1345: out = 24'(-49916);
			1346: out = 24'(-80588);
			1347: out = 24'(-99344);
			1348: out = 24'(-82168);
			1349: out = 24'(-41296);
			1350: out = 24'(-27888);
			1351: out = 24'(-15600);
			1352: out = 24'(-50600);
			1353: out = 24'(-96852);
			1354: out = 24'(-125512);
			1355: out = 24'(-92964);
			1356: out = 24'(-39428);
			1357: out = 24'(-70808);
			1358: out = 24'(-120800);
			1359: out = 24'(-97940);
			1360: out = 24'(-76780);
			1361: out = 24'(-83964);
			1362: out = 24'(-65224);
			1363: out = 24'(-45496);
			1364: out = 24'(-69016);
			1365: out = 24'(-103764);
			1366: out = 24'(-106780);
			1367: out = 24'(-116096);
			1368: out = 24'(-88140);
			1369: out = 24'(-39440);
			1370: out = 24'(-39004);
			1371: out = 24'(-38736);
			1372: out = 24'(-47452);
			1373: out = 24'(-84100);
			1374: out = 24'(-105268);
			1375: out = 24'(-120964);
			1376: out = 24'(-118268);
			1377: out = 24'(-121392);
			1378: out = 24'(-83600);
			1379: out = 24'(-25740);
			1380: out = 24'(-47056);
			1381: out = 24'(-89192);
			1382: out = 24'(-109948);
			1383: out = 24'(-96624);
			1384: out = 24'(-57224);
			1385: out = 24'(-18512);
			1386: out = 24'(-37728);
			1387: out = 24'(-91276);
			1388: out = 24'(-110192);
			1389: out = 24'(-100968);
			1390: out = 24'(-59608);
			1391: out = 24'(-83088);
			1392: out = 24'(-120620);
			1393: out = 24'(-116744);
			1394: out = 24'(-101196);
			1395: out = 24'(-65880);
			1396: out = 24'(-37688);
			1397: out = 24'(-39916);
			1398: out = 24'(-68376);
			1399: out = 24'(-108060);
			1400: out = 24'(-69320);
			1401: out = 24'(-51052);
			1402: out = 24'(-7400);
			1403: out = 24'(1056);
			1404: out = 24'(-57480);
			1405: out = 24'(-88620);
			1406: out = 24'(-89620);
			1407: out = 24'(-62732);
			1408: out = 24'(-38232);
			1409: out = 24'(-69484);
			1410: out = 24'(-84364);
			1411: out = 24'(-62616);
			1412: out = 24'(-50084);
			1413: out = 24'(-34608);
			1414: out = 24'(-41336);
			1415: out = 24'(-70752);
			1416: out = 24'(-80584);
			1417: out = 24'(-72148);
			1418: out = 24'(-38976);
			1419: out = 24'(-51092);
			1420: out = 24'(-71616);
			1421: out = 24'(-10400);
			1422: out = 24'(-2576);
			1423: out = 24'(-82136);
			1424: out = 24'(-92320);
			1425: out = 24'(-33564);
			1426: out = 24'(-29456);
			1427: out = 24'(-44032);
			1428: out = 24'(-44616);
			1429: out = 24'(-68196);
			1430: out = 24'(-28828);
			1431: out = 24'(47936);
			1432: out = 24'(6864);
			1433: out = 24'(-28704);
			1434: out = 24'(-33416);
			1435: out = 24'(39524);
			1436: out = 24'(29688);
			1437: out = 24'(-23184);
			1438: out = 24'(17360);
			1439: out = 24'(62024);
			1440: out = 24'(16060);
			1441: out = 24'(-72884);
			1442: out = 24'(-57296);
			1443: out = 24'(-5956);
			1444: out = 24'(17864);
			1445: out = 24'(-13552);
			1446: out = 24'(-15092);
			1447: out = 24'(15364);
			1448: out = 24'(57092);
			1449: out = 24'(50792);
			1450: out = 24'(1868);
			1451: out = 24'(-17084);
			1452: out = 24'(-1964);
			1453: out = 24'(44140);
			1454: out = 24'(31232);
			1455: out = 24'(20380);
			1456: out = 24'(52656);
			1457: out = 24'(62580);
			1458: out = 24'(13380);
			1459: out = 24'(-40784);
			1460: out = 24'(-15192);
			1461: out = 24'(38928);
			1462: out = 24'(51404);
			1463: out = 24'(67492);
			1464: out = 24'(92332);
			1465: out = 24'(59728);
			1466: out = 24'(-1004);
			1467: out = 24'(-6044);
			1468: out = 24'(-2088);
			1469: out = 24'(33136);
			1470: out = 24'(86096);
			1471: out = 24'(61224);
			1472: out = 24'(8988);
			1473: out = 24'(27584);
			1474: out = 24'(38092);
			1475: out = 24'(76920);
			1476: out = 24'(73300);
			1477: out = 24'(38624);
			1478: out = 24'(13316);
			1479: out = 24'(17220);
			1480: out = 24'(80392);
			1481: out = 24'(96312);
			1482: out = 24'(76792);
			1483: out = 24'(75616);
			1484: out = 24'(48784);
			1485: out = 24'(648);
			1486: out = 24'(13084);
			1487: out = 24'(21180);
			1488: out = 24'(33768);
			1489: out = 24'(61940);
			1490: out = 24'(73744);
			1491: out = 24'(71316);
			1492: out = 24'(98772);
			1493: out = 24'(123912);
			1494: out = 24'(75088);
			1495: out = 24'(26136);
			1496: out = 24'(18732);
			1497: out = 24'(66128);
			1498: out = 24'(106576);
			1499: out = 24'(84264);
			1500: out = 24'(79952);
			1501: out = 24'(101048);
			1502: out = 24'(92120);
			1503: out = 24'(22684);
			1504: out = 24'(-16548);
			1505: out = 24'(21088);
			1506: out = 24'(79812);
			1507: out = 24'(63064);
			1508: out = 24'(36376);
			1509: out = 24'(88928);
			1510: out = 24'(128276);
			1511: out = 24'(83108);
			1512: out = 24'(35568);
			1513: out = 24'(42680);
			1514: out = 24'(64556);
			1515: out = 24'(76608);
			1516: out = 24'(104280);
			1517: out = 24'(121392);
			1518: out = 24'(59272);
			1519: out = 24'(-12244);
			1520: out = 24'(-14892);
			1521: out = 24'(29892);
			1522: out = 24'(69044);
			1523: out = 24'(50352);
			1524: out = 24'(-452);
			1525: out = 24'(31392);
			1526: out = 24'(98284);
			1527: out = 24'(126816);
			1528: out = 24'(109048);
			1529: out = 24'(81168);
			1530: out = 24'(73844);
			1531: out = 24'(46364);
			1532: out = 24'(17612);
			1533: out = 24'(39928);
			1534: out = 24'(71728);
			1535: out = 24'(44432);
			1536: out = 24'(6468);
			1537: out = 24'(20064);
			1538: out = 24'(90660);
			1539: out = 24'(110920);
			1540: out = 24'(64964);
			1541: out = 24'(38184);
			1542: out = 24'(53880);
			1543: out = 24'(25272);
			1544: out = 24'(-4548);
			1545: out = 24'(40168);
			1546: out = 24'(70912);
			1547: out = 24'(39044);
			1548: out = 24'(37048);
			1549: out = 24'(33864);
			1550: out = 24'(46884);
			1551: out = 24'(78204);
			1552: out = 24'(51388);
			1553: out = 24'(10112);
			1554: out = 24'(-1176);
			1555: out = 24'(48488);
			1556: out = 24'(97124);
			1557: out = 24'(107928);
			1558: out = 24'(53212);
			1559: out = 24'(34700);
			1560: out = 24'(54248);
			1561: out = 24'(53824);
			1562: out = 24'(26848);
			1563: out = 24'(-18804);
			1564: out = 24'(1552);
			1565: out = 24'(57284);
			1566: out = 24'(89424);
			1567: out = 24'(55792);
			1568: out = 24'(-8348);
			1569: out = 24'(-13752);
			1570: out = 24'(14968);
			1571: out = 24'(40140);
			1572: out = 24'(45772);
			1573: out = 24'(3140);
			1574: out = 24'(-12728);
			1575: out = 24'(7712);
			1576: out = 24'(68988);
			1577: out = 24'(113580);
			1578: out = 24'(52536);
			1579: out = 24'(-19712);
			1580: out = 24'(-30912);
			1581: out = 24'(4340);
			1582: out = 24'(10412);
			1583: out = 24'(26956);
			1584: out = 24'(39280);
			1585: out = 24'(9836);
			1586: out = 24'(-5268);
			1587: out = 24'(26916);
			1588: out = 24'(22396);
			1589: out = 24'(24392);
			1590: out = 24'(43832);
			1591: out = 24'(54796);
			1592: out = 24'(31620);
			1593: out = 24'(7532);
			1594: out = 24'(2700);
			1595: out = 24'(27752);
			1596: out = 24'(72788);
			1597: out = 24'(60948);
			1598: out = 24'(1012);
			1599: out = 24'(-19884);
			1600: out = 24'(7280);
			1601: out = 24'(21164);
			1602: out = 24'(-40524);
			1603: out = 24'(-60844);
			1604: out = 24'(-14096);
			1605: out = 24'(34412);
			1606: out = 24'(51400);
			1607: out = 24'(42120);
			1608: out = 24'(37524);
			1609: out = 24'(22084);
			1610: out = 24'(-17220);
			1611: out = 24'(-59072);
			1612: out = 24'(-55588);
			1613: out = 24'(-26748);
			1614: out = 24'(-20332);
			1615: out = 24'(-29000);
			1616: out = 24'(1320);
			1617: out = 24'(28852);
			1618: out = 24'(1980);
			1619: out = 24'(-25988);
			1620: out = 24'(-52760);
			1621: out = 24'(-42764);
			1622: out = 24'(-27500);
			1623: out = 24'(-34164);
			1624: out = 24'(-1784);
			1625: out = 24'(876);
			1626: out = 24'(-29632);
			1627: out = 24'(-72896);
			1628: out = 24'(-89980);
			1629: out = 24'(-26716);
			1630: out = 24'(31632);
			1631: out = 24'(50824);
			1632: out = 24'(26764);
			1633: out = 24'(-42728);
			1634: out = 24'(-73516);
			1635: out = 24'(-68220);
			1636: out = 24'(-34116);
			1637: out = 24'(33904);
			1638: out = 24'(77648);
			1639: out = 24'(-5956);
			1640: out = 24'(-76472);
			1641: out = 24'(-79616);
			1642: out = 24'(-39376);
			1643: out = 24'(-416);
			1644: out = 24'(-11516);
			1645: out = 24'(-45488);
			1646: out = 24'(-46736);
			1647: out = 24'(14392);
			1648: out = 24'(-24720);
			1649: out = 24'(-46092);
			1650: out = 24'(-15964);
			1651: out = 24'(-20028);
			1652: out = 24'(19408);
			1653: out = 24'(19580);
			1654: out = 24'(-14380);
			1655: out = 24'(-28960);
			1656: out = 24'(-51892);
			1657: out = 24'(-37492);
			1658: out = 24'(-21388);
			1659: out = 24'(-29716);
			1660: out = 24'(-37768);
			1661: out = 24'(-47204);
			1662: out = 24'(-50948);
			1663: out = 24'(-23132);
			1664: out = 24'(-13360);
			1665: out = 24'(-24504);
			1666: out = 24'(-25608);
			1667: out = 24'(-34240);
			1668: out = 24'(-46048);
			1669: out = 24'(-78176);
			1670: out = 24'(-94936);
			1671: out = 24'(-50548);
			1672: out = 24'(-10804);
			1673: out = 24'(-22644);
			1674: out = 24'(-13140);
			1675: out = 24'(-408);
			1676: out = 24'(2556);
			1677: out = 24'(-56024);
			1678: out = 24'(-92692);
			1679: out = 24'(-57140);
			1680: out = 24'(-53996);
			1681: out = 24'(-43392);
			1682: out = 24'(8240);
			1683: out = 24'(32788);
			1684: out = 24'(-48968);
			1685: out = 24'(-113712);
			1686: out = 24'(-86328);
			1687: out = 24'(-25408);
			1688: out = 24'(17364);
			1689: out = 24'(-23936);
			1690: out = 24'(-81456);
			1691: out = 24'(-72020);
			1692: out = 24'(-61020);
			1693: out = 24'(-16980);
			1694: out = 24'(-15272);
			1695: out = 24'(-61144);
			1696: out = 24'(-68032);
			1697: out = 24'(-63524);
			1698: out = 24'(-32956);
			1699: out = 24'(-56972);
			1700: out = 24'(-34028);
			1701: out = 24'(-9260);
			1702: out = 24'(-7956);
			1703: out = 24'(-1548);
			1704: out = 24'(-45844);
			1705: out = 24'(-44692);
			1706: out = 24'(-6384);
			1707: out = 24'(22696);
			1708: out = 24'(-1240);
			1709: out = 24'(-44472);
			1710: out = 24'(-70160);
			1711: out = 24'(-59740);
			1712: out = 24'(-54084);
			1713: out = 24'(-46468);
			1714: out = 24'(-59044);
			1715: out = 24'(-55184);
			1716: out = 24'(-41400);
			1717: out = 24'(-25124);
			1718: out = 24'(-77364);
			1719: out = 24'(-67148);
			1720: out = 24'(-19768);
			1721: out = 24'(-360);
			1722: out = 24'(-26408);
			1723: out = 24'(-52096);
			1724: out = 24'(-63616);
			1725: out = 24'(-76176);
			1726: out = 24'(-47300);
			1727: out = 24'(22860);
			1728: out = 24'(46816);
			1729: out = 24'(-8092);
			1730: out = 24'(-68396);
			1731: out = 24'(-60324);
			1732: out = 24'(9032);
			1733: out = 24'(30528);
			1734: out = 24'(-46036);
			1735: out = 24'(-79084);
			1736: out = 24'(-28144);
			1737: out = 24'(29320);
			1738: out = 24'(-24912);
			1739: out = 24'(-84508);
			1740: out = 24'(-37652);
			1741: out = 24'(27748);
			1742: out = 24'(31728);
			1743: out = 24'(-4944);
			1744: out = 24'(-10500);
			1745: out = 24'(-16000);
			1746: out = 24'(-33268);
			1747: out = 24'(-82252);
			1748: out = 24'(-54008);
			1749: out = 24'(7616);
			1750: out = 24'(-33448);
			1751: out = 24'(-115888);
			1752: out = 24'(-72616);
			1753: out = 24'(-20104);
			1754: out = 24'(5000);
			1755: out = 24'(26436);
			1756: out = 24'(36044);
			1757: out = 24'(-38944);
			1758: out = 24'(-88792);
			1759: out = 24'(-70964);
			1760: out = 24'(-31288);
			1761: out = 24'(40540);
			1762: out = 24'(49840);
			1763: out = 24'(-41388);
			1764: out = 24'(-84740);
			1765: out = 24'(-52976);
			1766: out = 24'(-1404);
			1767: out = 24'(17384);
			1768: out = 24'(-15384);
			1769: out = 24'(-30624);
			1770: out = 24'(5548);
			1771: out = 24'(41520);
			1772: out = 24'(14768);
			1773: out = 24'(-38520);
			1774: out = 24'(-66804);
			1775: out = 24'(-40552);
			1776: out = 24'(-12484);
			1777: out = 24'(-35336);
			1778: out = 24'(-2788);
			1779: out = 24'(3136);
			1780: out = 24'(12648);
			1781: out = 24'(35780);
			1782: out = 24'(40892);
			1783: out = 24'(-21836);
			1784: out = 24'(-65088);
			1785: out = 24'(-65064);
			1786: out = 24'(-9140);
			1787: out = 24'(84364);
			1788: out = 24'(43924);
			1789: out = 24'(-61280);
			1790: out = 24'(-35464);
			1791: out = 24'(3504);
			1792: out = 24'(7868);
			1793: out = 24'(656);
			1794: out = 24'(14828);
			1795: out = 24'(17088);
			1796: out = 24'(24120);
			1797: out = 24'(57208);
			1798: out = 24'(34588);
			1799: out = 24'(5636);
			1800: out = 24'(-23984);
			1801: out = 24'(-34124);
			1802: out = 24'(-9296);
			1803: out = 24'(56212);
			1804: out = 24'(70984);
			1805: out = 24'(-20404);
			1806: out = 24'(-38864);
			1807: out = 24'(19408);
			1808: out = 24'(42860);
			1809: out = 24'(22404);
			1810: out = 24'(-13652);
			1811: out = 24'(-26808);
			1812: out = 24'(-7788);
			1813: out = 24'(31704);
			1814: out = 24'(48096);
			1815: out = 24'(37964);
			1816: out = 24'(38868);
			1817: out = 24'(8144);
			1818: out = 24'(-696);
			1819: out = 24'(14760);
			1820: out = 24'(17012);
			1821: out = 24'(13932);
			1822: out = 24'(46660);
			1823: out = 24'(38944);
			1824: out = 24'(9408);
			1825: out = 24'(8300);
			1826: out = 24'(37696);
			1827: out = 24'(63448);
			1828: out = 24'(32564);
			1829: out = 24'(40944);
			1830: out = 24'(33212);
			1831: out = 24'(8036);
			1832: out = 24'(-13580);
			1833: out = 24'(4584);
			1834: out = 24'(20284);
			1835: out = 24'(39360);
			1836: out = 24'(51876);
			1837: out = 24'(35136);
			1838: out = 24'(-29584);
			1839: out = 24'(-43340);
			1840: out = 24'(-12876);
			1841: out = 24'(-1652);
			1842: out = 24'(41016);
			1843: out = 24'(88072);
			1844: out = 24'(74932);
			1845: out = 24'(3700);
			1846: out = 24'(-26464);
			1847: out = 24'(36064);
			1848: out = 24'(90980);
			1849: out = 24'(68296);
			1850: out = 24'(49448);
			1851: out = 24'(53396);
			1852: out = 24'(46756);
			1853: out = 24'(-4140);
			1854: out = 24'(-38492);
			1855: out = 24'(-18420);
			1856: out = 24'(1940);
			1857: out = 24'(19880);
			1858: out = 24'(51236);
			1859: out = 24'(52500);
			1860: out = 24'(15468);
			1861: out = 24'(30308);
			1862: out = 24'(41928);
			1863: out = 24'(62084);
			1864: out = 24'(69728);
			1865: out = 24'(69720);
			1866: out = 24'(30872);
			1867: out = 24'(-20948);
			1868: out = 24'(-42408);
			1869: out = 24'(-11172);
			1870: out = 24'(71708);
			1871: out = 24'(109484);
			1872: out = 24'(40128);
			1873: out = 24'(-21408);
			1874: out = 24'(9064);
			1875: out = 24'(47376);
			1876: out = 24'(62516);
			1877: out = 24'(46940);
			1878: out = 24'(2536);
			1879: out = 24'(-27864);
			1880: out = 24'(-23524);
			1881: out = 24'(-6348);
			1882: out = 24'(29816);
			1883: out = 24'(22096);
			1884: out = 24'(11984);
			1885: out = 24'(46652);
			1886: out = 24'(70680);
			1887: out = 24'(7176);
			1888: out = 24'(-44912);
			1889: out = 24'(-35236);
			1890: out = 24'(-1696);
			1891: out = 24'(52512);
			1892: out = 24'(107936);
			1893: out = 24'(53296);
			1894: out = 24'(-17032);
			1895: out = 24'(-12220);
			1896: out = 24'(5584);
			1897: out = 24'(7020);
			1898: out = 24'(8328);
			1899: out = 24'(-4564);
			1900: out = 24'(-17684);
			1901: out = 24'(20872);
			1902: out = 24'(3296);
			1903: out = 24'(-51296);
			1904: out = 24'(3092);
			1905: out = 24'(49716);
			1906: out = 24'(50464);
			1907: out = 24'(30604);
			1908: out = 24'(3152);
			1909: out = 24'(19916);
			1910: out = 24'(44388);
			1911: out = 24'(39228);
			1912: out = 24'(11892);
			1913: out = 24'(-23296);
			1914: out = 24'(-10316);
			1915: out = 24'(35492);
			1916: out = 24'(52100);
			1917: out = 24'(6852);
			1918: out = 24'(-11772);
			1919: out = 24'(2040);
			1920: out = 24'(17744);
			1921: out = 24'(-4768);
			1922: out = 24'(-25384);
			1923: out = 24'(30644);
			1924: out = 24'(72476);
			1925: out = 24'(22180);
			1926: out = 24'(-37184);
			1927: out = 24'(-46652);
			1928: out = 24'(9704);
			1929: out = 24'(23832);
			1930: out = 24'(-2776);
			1931: out = 24'(5248);
			1932: out = 24'(7944);
			1933: out = 24'(15432);
			1934: out = 24'(27508);
			1935: out = 24'(50172);
			1936: out = 24'(62080);
			1937: out = 24'(14788);
			1938: out = 24'(-36572);
			1939: out = 24'(-32876);
			1940: out = 24'(-23776);
			1941: out = 24'(7972);
			1942: out = 24'(27720);
			1943: out = 24'(-35036);
			1944: out = 24'(-61896);
			1945: out = 24'(6924);
			1946: out = 24'(63296);
			1947: out = 24'(39876);
			1948: out = 24'(44192);
			1949: out = 24'(60552);
			1950: out = 24'(24360);
			1951: out = 24'(-27868);
			1952: out = 24'(-61496);
			1953: out = 24'(-30360);
			1954: out = 24'(28804);
			1955: out = 24'(62068);
			1956: out = 24'(64);
			1957: out = 24'(-33396);
			1958: out = 24'(9164);
			1959: out = 24'(51172);
			1960: out = 24'(57404);
			1961: out = 24'(25856);
			1962: out = 24'(-19192);
			1963: out = 24'(-27536);
			1964: out = 24'(9328);
			1965: out = 24'(46188);
			1966: out = 24'(51356);
			1967: out = 24'(43096);
			1968: out = 24'(20732);
			1969: out = 24'(36392);
			1970: out = 24'(25608);
			1971: out = 24'(13868);
			1972: out = 24'(8056);
			1973: out = 24'(20152);
			1974: out = 24'(37484);
			1975: out = 24'(3852);
			1976: out = 24'(17524);
			1977: out = 24'(61656);
			1978: out = 24'(41092);
			1979: out = 24'(-42608);
			1980: out = 24'(-61128);
			1981: out = 24'(-27608);
			1982: out = 24'(-11124);
			1983: out = 24'(-3660);
			1984: out = 24'(11292);
			1985: out = 24'(-11784);
			1986: out = 24'(3376);
			1987: out = 24'(20424);
			1988: out = 24'(23052);
			1989: out = 24'(-23456);
			1990: out = 24'(-39156);
			1991: out = 24'(-11868);
			1992: out = 24'(-1048);
			1993: out = 24'(51916);
			1994: out = 24'(50872);
			1995: out = 24'(46796);
			1996: out = 24'(20864);
			1997: out = 24'(8080);
			1998: out = 24'(18940);
			1999: out = 24'(1608);
			2000: out = 24'(868);
			2001: out = 24'(22836);
			2002: out = 24'(10732);
			2003: out = 24'(-1500);
			2004: out = 24'(-18672);
			2005: out = 24'(-41392);
			2006: out = 24'(-15124);
			2007: out = 24'(-21280);
			2008: out = 24'(-33304);
			2009: out = 24'(8600);
			2010: out = 24'(12168);
			2011: out = 24'(-10144);
			2012: out = 24'(-29028);
			2013: out = 24'(-5824);
			2014: out = 24'(-3500);
			2015: out = 24'(-31592);
			2016: out = 24'(13284);
			2017: out = 24'(51908);
			2018: out = 24'(22124);
			2019: out = 24'(-21152);
			2020: out = 24'(-1856);
			2021: out = 24'(11360);
			2022: out = 24'(7544);
			2023: out = 24'(-50528);
			2024: out = 24'(-54396);
			2025: out = 24'(-33676);
			2026: out = 24'(-564);
			2027: out = 24'(-2696);
			2028: out = 24'(-42732);
			2029: out = 24'(-41636);
			2030: out = 24'(-19448);
			2031: out = 24'(-12756);
			2032: out = 24'(-51144);
			2033: out = 24'(-18392);
			2034: out = 24'(-9032);
			2035: out = 24'(-12124);
			2036: out = 24'(31932);
			2037: out = 24'(34208);
			2038: out = 24'(-2260);
			2039: out = 24'(-36744);
			2040: out = 24'(-41064);
			2041: out = 24'(-31868);
			2042: out = 24'(-51404);
			2043: out = 24'(-39076);
			2044: out = 24'(-18228);
			2045: out = 24'(-37372);
			2046: out = 24'(-40596);
			2047: out = 24'(-20804);
			2048: out = 24'(9008);
			2049: out = 24'(16704);
			2050: out = 24'(6340);
			2051: out = 24'(-18940);
			2052: out = 24'(-31880);
			2053: out = 24'(-13052);
			2054: out = 24'(-15932);
			2055: out = 24'(-16680);
			2056: out = 24'(-48912);
			2057: out = 24'(-79956);
			2058: out = 24'(-73292);
			2059: out = 24'(-56800);
			2060: out = 24'(-4280);
			2061: out = 24'(6384);
			2062: out = 24'(-15604);
			2063: out = 24'(212);
			2064: out = 24'(7036);
			2065: out = 24'(-41996);
			2066: out = 24'(-79848);
			2067: out = 24'(-55944);
			2068: out = 24'(-37872);
			2069: out = 24'(-20472);
			2070: out = 24'(-15092);
			2071: out = 24'(-2564);
			2072: out = 24'(3940);
			2073: out = 24'(-12312);
			2074: out = 24'(-48004);
			2075: out = 24'(-52188);
			2076: out = 24'(-51440);
			2077: out = 24'(-44900);
			2078: out = 24'(2276);
			2079: out = 24'(36004);
			2080: out = 24'(-31624);
			2081: out = 24'(-58088);
			2082: out = 24'(-45892);
			2083: out = 24'(-38856);
			2084: out = 24'(-66152);
			2085: out = 24'(-54216);
			2086: out = 24'(8156);
			2087: out = 24'(-3892);
			2088: out = 24'(-27388);
			2089: out = 24'(-50072);
			2090: out = 24'(-43960);
			2091: out = 24'(-21508);
			2092: out = 24'(-15528);
			2093: out = 24'(2044);
			2094: out = 24'(-18572);
			2095: out = 24'(-28460);
			2096: out = 24'(-46244);
			2097: out = 24'(-31968);
			2098: out = 24'(20404);
			2099: out = 24'(-11800);
			2100: out = 24'(-43272);
			2101: out = 24'(-35716);
			2102: out = 24'(-16872);
			2103: out = 24'(-31416);
			2104: out = 24'(-67180);
			2105: out = 24'(-61888);
			2106: out = 24'(-31080);
			2107: out = 24'(-10744);
			2108: out = 24'(-27124);
			2109: out = 24'(-15592);
			2110: out = 24'(-26764);
			2111: out = 24'(-26992);
			2112: out = 24'(-42164);
			2113: out = 24'(-33648);
			2114: out = 24'(-39372);
			2115: out = 24'(-56608);
			2116: out = 24'(-62568);
			2117: out = 24'(-62560);
			2118: out = 24'(-20328);
			2119: out = 24'(-20428);
			2120: out = 24'(-33468);
			2121: out = 24'(-53216);
			2122: out = 24'(-54472);
			2123: out = 24'(-45536);
			2124: out = 24'(-15840);
			2125: out = 24'(13324);
			2126: out = 24'(-31260);
			2127: out = 24'(-64636);
			2128: out = 24'(-38892);
			2129: out = 24'(20348);
			2130: out = 24'(-9920);
			2131: out = 24'(-34572);
			2132: out = 24'(-4172);
			2133: out = 24'(-5504);
			2134: out = 24'(-54640);
			2135: out = 24'(-88276);
			2136: out = 24'(-55468);
			2137: out = 24'(-6164);
			2138: out = 24'(-4868);
			2139: out = 24'(-50048);
			2140: out = 24'(-36968);
			2141: out = 24'(-44080);
			2142: out = 24'(-48436);
			2143: out = 24'(-26004);
			2144: out = 24'(-32304);
			2145: out = 24'(-11548);
			2146: out = 24'(-17160);
			2147: out = 24'(-12088);
			2148: out = 24'(-19040);
			2149: out = 24'(-32048);
			2150: out = 24'(-70520);
			2151: out = 24'(-46180);
			2152: out = 24'(-16532);
			2153: out = 24'(-52316);
			2154: out = 24'(-43700);
			2155: out = 24'(2492);
			2156: out = 24'(36584);
			2157: out = 24'(9144);
			2158: out = 24'(-8716);
			2159: out = 24'(-27836);
			2160: out = 24'(-14684);
			2161: out = 24'(-15312);
			2162: out = 24'(-43528);
			2163: out = 24'(-31568);
			2164: out = 24'(-35188);
			2165: out = 24'(18684);
			2166: out = 24'(38884);
			2167: out = 24'(4672);
			2168: out = 24'(-28344);
			2169: out = 24'(-29672);
			2170: out = 24'(-36856);
			2171: out = 24'(-26380);
			2172: out = 24'(14832);
			2173: out = 24'(-592);
			2174: out = 24'(-15304);
			2175: out = 24'(-8468);
			2176: out = 24'(38284);
			2177: out = 24'(35936);
			2178: out = 24'(19896);
			2179: out = 24'(5032);
			2180: out = 24'(-17516);
			2181: out = 24'(-43048);
			2182: out = 24'(-59008);
			2183: out = 24'(-6872);
			2184: out = 24'(53788);
			2185: out = 24'(51568);
			2186: out = 24'(3760);
			2187: out = 24'(-9784);
			2188: out = 24'(-13444);
			2189: out = 24'(7440);
			2190: out = 24'(51012);
			2191: out = 24'(31944);
			2192: out = 24'(-10568);
			2193: out = 24'(-31144);
			2194: out = 24'(10184);
			2195: out = 24'(61708);
			2196: out = 24'(63748);
			2197: out = 24'(-7852);
			2198: out = 24'(-27248);
			2199: out = 24'(-27544);
			2200: out = 24'(-6820);
			2201: out = 24'(51712);
			2202: out = 24'(58824);
			2203: out = 24'(35564);
			2204: out = 24'(16592);
			2205: out = 24'(17416);
			2206: out = 24'(15320);
			2207: out = 24'(-3648);
			2208: out = 24'(8956);
			2209: out = 24'(63908);
			2210: out = 24'(37612);
			2211: out = 24'(-18056);
			2212: out = 24'(-10648);
			2213: out = 24'(46100);
			2214: out = 24'(72808);
			2215: out = 24'(12368);
			2216: out = 24'(23176);
			2217: out = 24'(71148);
			2218: out = 24'(39648);
			2219: out = 24'(3456);
			2220: out = 24'(13060);
			2221: out = 24'(22924);
			2222: out = 24'(19144);
			2223: out = 24'(24548);
			2224: out = 24'(30288);
			2225: out = 24'(13172);
			2226: out = 24'(23720);
			2227: out = 24'(41836);
			2228: out = 24'(22532);
			2229: out = 24'(15876);
			2230: out = 24'(57712);
			2231: out = 24'(70276);
			2232: out = 24'(44660);
			2233: out = 24'(31136);
			2234: out = 24'(40204);
			2235: out = 24'(65004);
			2236: out = 24'(57568);
			2237: out = 24'(29868);
			2238: out = 24'(15884);
			2239: out = 24'(4088);
			2240: out = 24'(11156);
			2241: out = 24'(31584);
			2242: out = 24'(32740);
			2243: out = 24'(36304);
			2244: out = 24'(32620);
			2245: out = 24'(46904);
			2246: out = 24'(32240);
			2247: out = 24'(20384);
			2248: out = 24'(3176);
			2249: out = 24'(31112);
			2250: out = 24'(56480);
			2251: out = 24'(69436);
			2252: out = 24'(58476);
			2253: out = 24'(-720);
			2254: out = 24'(-16200);
			2255: out = 24'(30780);
			2256: out = 24'(84308);
			2257: out = 24'(61736);
			2258: out = 24'(14232);
			2259: out = 24'(-11672);
			2260: out = 24'(25476);
			2261: out = 24'(61496);
			2262: out = 24'(11200);
			2263: out = 24'(20352);
			2264: out = 24'(44920);
			2265: out = 24'(65948);
			2266: out = 24'(84172);
			2267: out = 24'(64524);
			2268: out = 24'(50904);
			2269: out = 24'(23344);
			2270: out = 24'(-6680);
			2271: out = 24'(-14572);
			2272: out = 24'(22716);
			2273: out = 24'(19380);
			2274: out = 24'(-15212);
			2275: out = 24'(19872);
			2276: out = 24'(64212);
			2277: out = 24'(50012);
			2278: out = 24'(29848);
			2279: out = 24'(-3544);
			2280: out = 24'(14552);
			2281: out = 24'(27368);
			2282: out = 24'(55280);
			2283: out = 24'(72852);
			2284: out = 24'(36596);
			2285: out = 24'(30736);
			2286: out = 24'(33940);
			2287: out = 24'(25156);
			2288: out = 24'(-9568);
			2289: out = 24'(-31304);
			2290: out = 24'(10516);
			2291: out = 24'(82484);
			2292: out = 24'(56336);
			2293: out = 24'(-19604);
			2294: out = 24'(-25544);
			2295: out = 24'(32664);
			2296: out = 24'(55940);
			2297: out = 24'(4244);
			2298: out = 24'(-8976);
			2299: out = 24'(40728);
			2300: out = 24'(53980);
			2301: out = 24'(41004);
			2302: out = 24'(45752);
			2303: out = 24'(23676);
			2304: out = 24'(5660);
			2305: out = 24'(4884);
			2306: out = 24'(51552);
			2307: out = 24'(79900);
			2308: out = 24'(17336);
			2309: out = 24'(-37272);
			2310: out = 24'(-26688);
			2311: out = 24'(-1128);
			2312: out = 24'(35976);
			2313: out = 24'(-1600);
			2314: out = 24'(-29524);
			2315: out = 24'(29768);
			2316: out = 24'(38832);
			2317: out = 24'(-29452);
			2318: out = 24'(-46832);
			2319: out = 24'(-21152);
			2320: out = 24'(22724);
			2321: out = 24'(74496);
			2322: out = 24'(78704);
			2323: out = 24'(23156);
			2324: out = 24'(-2740);
			2325: out = 24'(-28516);
			2326: out = 24'(-16304);
			2327: out = 24'(20372);
			2328: out = 24'(34388);
			2329: out = 24'(33352);
			2330: out = 24'(29616);
			2331: out = 24'(-3672);
			2332: out = 24'(-45236);
			2333: out = 24'(-27016);
			2334: out = 24'(18648);
			2335: out = 24'(37836);
			2336: out = 24'(45244);
			2337: out = 24'(5196);
			2338: out = 24'(-41284);
			2339: out = 24'(-41428);
			2340: out = 24'(-5536);
			2341: out = 24'(56936);
			2342: out = 24'(36676);
			2343: out = 24'(-12496);
			2344: out = 24'(-5084);
			2345: out = 24'(30240);
			2346: out = 24'(40192);
			2347: out = 24'(21648);
			2348: out = 24'(-2344);
			2349: out = 24'(9408);
			2350: out = 24'(-15392);
			2351: out = 24'(-30052);
			2352: out = 24'(-1796);
			2353: out = 24'(-12392);
			2354: out = 24'(-40560);
			2355: out = 24'(-33896);
			2356: out = 24'(13008);
			2357: out = 24'(9644);
			2358: out = 24'(13608);
			2359: out = 24'(47344);
			2360: out = 24'(36160);
			2361: out = 24'(-32664);
			2362: out = 24'(-75252);
			2363: out = 24'(-34160);
			2364: out = 24'(32240);
			2365: out = 24'(16692);
			2366: out = 24'(-3616);
			2367: out = 24'(-8984);
			2368: out = 24'(-28492);
			2369: out = 24'(-46840);
			2370: out = 24'(-46564);
			2371: out = 24'(-19920);
			2372: out = 24'(16520);
			2373: out = 24'(-1344);
			2374: out = 24'(-6032);
			2375: out = 24'(-14864);
			2376: out = 24'(-37488);
			2377: out = 24'(19092);
			2378: out = 24'(60876);
			2379: out = 24'(30336);
			2380: out = 24'(-26520);
			2381: out = 24'(-51448);
			2382: out = 24'(-42712);
			2383: out = 24'(-11004);
			2384: out = 24'(-21324);
			2385: out = 24'(-61500);
			2386: out = 24'(-42268);
			2387: out = 24'(9932);
			2388: out = 24'(-4356);
			2389: out = 24'(-15956);
			2390: out = 24'(-19736);
			2391: out = 24'(4720);
			2392: out = 24'(19016);
			2393: out = 24'(-16152);
			2394: out = 24'(-4632);
			2395: out = 24'(25788);
			2396: out = 24'(26696);
			2397: out = 24'(-23160);
			2398: out = 24'(-49192);
			2399: out = 24'(-19676);
			2400: out = 24'(-11288);
			2401: out = 24'(-73736);
			2402: out = 24'(-59616);
			2403: out = 24'(-580);
			2404: out = 24'(-15004);
			2405: out = 24'(-43732);
			2406: out = 24'(-27612);
			2407: out = 24'(-59936);
			2408: out = 24'(-38200);
			2409: out = 24'(22176);
			2410: out = 24'(37916);
			2411: out = 24'(-18468);
			2412: out = 24'(-82568);
			2413: out = 24'(-73168);
			2414: out = 24'(-15036);
			2415: out = 24'(33960);
			2416: out = 24'(-18244);
			2417: out = 24'(-51172);
			2418: out = 24'(-44228);
			2419: out = 24'(-24004);
			2420: out = 24'(34704);
			2421: out = 24'(14112);
			2422: out = 24'(-30736);
			2423: out = 24'(-20236);
			2424: out = 24'(-26736);
			2425: out = 24'(-24952);
			2426: out = 24'(-28668);
			2427: out = 24'(-36588);
			2428: out = 24'(-25800);
			2429: out = 24'(-40864);
			2430: out = 24'(-45364);
			2431: out = 24'(-17276);
			2432: out = 24'(-22028);
			2433: out = 24'(-61828);
			2434: out = 24'(-25200);
			2435: out = 24'(21028);
			2436: out = 24'(-19304);
			2437: out = 24'(-39936);
			2438: out = 24'(-61104);
			2439: out = 24'(-58624);
			2440: out = 24'(-19984);
			2441: out = 24'(28112);
			2442: out = 24'(43368);
			2443: out = 24'(-34568);
			2444: out = 24'(-103956);
			2445: out = 24'(-73724);
			2446: out = 24'(1024);
			2447: out = 24'(37536);
			2448: out = 24'(-13620);
			2449: out = 24'(-21432);
			2450: out = 24'(-23688);
			2451: out = 24'(-6964);
			2452: out = 24'(-3604);
			2453: out = 24'(-6928);
			2454: out = 24'(25612);
			2455: out = 24'(26160);
			2456: out = 24'(-16124);
			2457: out = 24'(-37280);
			2458: out = 24'(-36252);
			2459: out = 24'(-15684);
			2460: out = 24'(-22896);
			2461: out = 24'(-32468);
			2462: out = 24'(-39424);
			2463: out = 24'(-17424);
			2464: out = 24'(-16276);
			2465: out = 24'(-20776);
			2466: out = 24'(-26916);
			2467: out = 24'(-11360);
			2468: out = 24'(3316);
			2469: out = 24'(-9756);
			2470: out = 24'(-5944);
			2471: out = 24'(-18284);
			2472: out = 24'(-18260);
			2473: out = 24'(-15160);
			2474: out = 24'(-32672);
			2475: out = 24'(-41652);
			2476: out = 24'(-42280);
			2477: out = 24'(-59836);
			2478: out = 24'(-53468);
			2479: out = 24'(-28288);
			2480: out = 24'(-972);
			2481: out = 24'(-7272);
			2482: out = 24'(28956);
			2483: out = 24'(8432);
			2484: out = 24'(-13004);
			2485: out = 24'(-30488);
			2486: out = 24'(-16412);
			2487: out = 24'(9192);
			2488: out = 24'(-5288);
			2489: out = 24'(25216);
			2490: out = 24'(40480);
			2491: out = 24'(-19524);
			2492: out = 24'(-83412);
			2493: out = 24'(-82908);
			2494: out = 24'(-64368);
			2495: out = 24'(15604);
			2496: out = 24'(17720);
			2497: out = 24'(-47380);
			2498: out = 24'(-44432);
			2499: out = 24'(2144);
			2500: out = 24'(37764);
			2501: out = 24'(9348);
			2502: out = 24'(16292);
			2503: out = 24'(-3396);
			2504: out = 24'(-31444);
			2505: out = 24'(-35964);
			2506: out = 24'(-5208);
			2507: out = 24'(15868);
			2508: out = 24'(24896);
			2509: out = 24'(6368);
			2510: out = 24'(6092);
			2511: out = 24'(17640);
			2512: out = 24'(-20688);
			2513: out = 24'(-29144);
			2514: out = 24'(-10288);
			2515: out = 24'(5448);
			2516: out = 24'(13124);
			2517: out = 24'(-26232);
			2518: out = 24'(-35024);
			2519: out = 24'(1808);
			2520: out = 24'(16084);
			2521: out = 24'(13216);
			2522: out = 24'(-10448);
			2523: out = 24'(-44680);
			2524: out = 24'(-22732);
			2525: out = 24'(52);
			2526: out = 24'(26880);
			2527: out = 24'(29600);
			2528: out = 24'(16760);
			2529: out = 24'(-5288);
			2530: out = 24'(-1088);
			2531: out = 24'(39512);
			2532: out = 24'(24756);
			2533: out = 24'(-21020);
			2534: out = 24'(-27396);
			2535: out = 24'(-3720);
			2536: out = 24'(9132);
			2537: out = 24'(10900);
			2538: out = 24'(31180);
			2539: out = 24'(32184);
			2540: out = 24'(34644);
			2541: out = 24'(9616);
			2542: out = 24'(-33520);
			2543: out = 24'(-4580);
			2544: out = 24'(12080);
			2545: out = 24'(31036);
			2546: out = 24'(38776);
			2547: out = 24'(35308);
			2548: out = 24'(35424);
			2549: out = 24'(10720);
			2550: out = 24'(4820);
			2551: out = 24'(26960);
			2552: out = 24'(25700);
			2553: out = 24'(12168);
			2554: out = 24'(-7652);
			2555: out = 24'(-3660);
			2556: out = 24'(32880);
			2557: out = 24'(54120);
			2558: out = 24'(5536);
			2559: out = 24'(-38448);
			2560: out = 24'(-13084);
			2561: out = 24'(820);
			2562: out = 24'(14896);
			2563: out = 24'(12536);
			2564: out = 24'(13072);
			2565: out = 24'(7488);
			2566: out = 24'(44520);
			2567: out = 24'(71544);
			2568: out = 24'(24792);
			2569: out = 24'(-41984);
			2570: out = 24'(-47996);
			2571: out = 24'(-3164);
			2572: out = 24'(11144);
			2573: out = 24'(52668);
			2574: out = 24'(53456);
			2575: out = 24'(9148);
			2576: out = 24'(-16300);
			2577: out = 24'(10672);
			2578: out = 24'(20828);
			2579: out = 24'(-4524);
			2580: out = 24'(9260);
			2581: out = 24'(33740);
			2582: out = 24'(56780);
			2583: out = 24'(29808);
			2584: out = 24'(-7824);
			2585: out = 24'(-3860);
			2586: out = 24'(28388);
			2587: out = 24'(34628);
			2588: out = 24'(-9660);
			2589: out = 24'(-18024);
			2590: out = 24'(13344);
			2591: out = 24'(-12788);
			2592: out = 24'(17144);
			2593: out = 24'(76792);
			2594: out = 24'(44428);
			2595: out = 24'(-28236);
			2596: out = 24'(-26100);
			2597: out = 24'(23120);
			2598: out = 24'(34616);
			2599: out = 24'(47464);
			2600: out = 24'(22724);
			2601: out = 24'(-19184);
			2602: out = 24'(5688);
			2603: out = 24'(69068);
			2604: out = 24'(84240);
			2605: out = 24'(41156);
			2606: out = 24'(-16184);
			2607: out = 24'(-10968);
			2608: out = 24'(34892);
			2609: out = 24'(44440);
			2610: out = 24'(32376);
			2611: out = 24'(6796);
			2612: out = 24'(-8660);
			2613: out = 24'(3752);
			2614: out = 24'(19028);
			2615: out = 24'(-30940);
			2616: out = 24'(-32484);
			2617: out = 24'(8460);
			2618: out = 24'(7548);
			2619: out = 24'(38964);
			2620: out = 24'(63600);
			2621: out = 24'(-8240);
			2622: out = 24'(-57972);
			2623: out = 24'(-11388);
			2624: out = 24'(13468);
			2625: out = 24'(27188);
			2626: out = 24'(46592);
			2627: out = 24'(38360);
			2628: out = 24'(32864);
			2629: out = 24'(23760);
			2630: out = 24'(-7224);
			2631: out = 24'(-868);
			2632: out = 24'(32784);
			2633: out = 24'(36564);
			2634: out = 24'(-24580);
			2635: out = 24'(-51304);
			2636: out = 24'(-8212);
			2637: out = 24'(18296);
			2638: out = 24'(51392);
			2639: out = 24'(26540);
			2640: out = 24'(-6136);
			2641: out = 24'(31220);
			2642: out = 24'(34892);
			2643: out = 24'(1168);
			2644: out = 24'(-24328);
			2645: out = 24'(-23272);
			2646: out = 24'(-4072);
			2647: out = 24'(9968);
			2648: out = 24'(47620);
			2649: out = 24'(44256);
			2650: out = 24'(-14716);
			2651: out = 24'(-52468);
			2652: out = 24'(-9956);
			2653: out = 24'(14376);
			2654: out = 24'(20344);
			2655: out = 24'(1240);
			2656: out = 24'(-23736);
			2657: out = 24'(-14964);
			2658: out = 24'(-9636);
			2659: out = 24'(32068);
			2660: out = 24'(50568);
			2661: out = 24'(30848);
			2662: out = 24'(17840);
			2663: out = 24'(-20988);
			2664: out = 24'(-44284);
			2665: out = 24'(-4060);
			2666: out = 24'(11464);
			2667: out = 24'(42056);
			2668: out = 24'(45544);
			2669: out = 24'(7000);
			2670: out = 24'(-17380);
			2671: out = 24'(-23572);
			2672: out = 24'(-15212);
			2673: out = 24'(-15524);
			2674: out = 24'(-16028);
			2675: out = 24'(-2148);
			2676: out = 24'(15008);
			2677: out = 24'(41244);
			2678: out = 24'(27040);
			2679: out = 24'(40448);
			2680: out = 24'(47196);
			2681: out = 24'(-6072);
			2682: out = 24'(-24304);
			2683: out = 24'(-9268);
			2684: out = 24'(-10552);
			2685: out = 24'(-4012);
			2686: out = 24'(-2344);
			2687: out = 24'(3100);
			2688: out = 24'(5464);
			2689: out = 24'(-29704);
			2690: out = 24'(-50620);
			2691: out = 24'(-4572);
			2692: out = 24'(31384);
			2693: out = 24'(31260);
			2694: out = 24'(-48488);
			2695: out = 24'(-68972);
			2696: out = 24'(-4280);
			2697: out = 24'(78388);
			2698: out = 24'(88964);
			2699: out = 24'(-1664);
			2700: out = 24'(-19932);
			2701: out = 24'(3784);
			2702: out = 24'(11056);
			2703: out = 24'(23344);
			2704: out = 24'(21704);
			2705: out = 24'(-17624);
			2706: out = 24'(-39640);
			2707: out = 24'(-27968);
			2708: out = 24'(18264);
			2709: out = 24'(15804);
			2710: out = 24'(-44448);
			2711: out = 24'(-45640);
			2712: out = 24'(-7668);
			2713: out = 24'(25888);
			2714: out = 24'(16328);
			2715: out = 24'(-51804);
			2716: out = 24'(-13048);
			2717: out = 24'(18276);
			2718: out = 24'(35856);
			2719: out = 24'(64008);
			2720: out = 24'(51420);
			2721: out = 24'(-8536);
			2722: out = 24'(-58008);
			2723: out = 24'(-67184);
			2724: out = 24'(-14948);
			2725: out = 24'(23948);
			2726: out = 24'(-1032);
			2727: out = 24'(-19264);
			2728: out = 24'(-13776);
			2729: out = 24'(35636);
			2730: out = 24'(30028);
			2731: out = 24'(-12700);
			2732: out = 24'(-3028);
			2733: out = 24'(42880);
			2734: out = 24'(22296);
			2735: out = 24'(-27972);
			2736: out = 24'(-19232);
			2737: out = 24'(9252);
			2738: out = 24'(1588);
			2739: out = 24'(-29212);
			2740: out = 24'(-18584);
			2741: out = 24'(-6696);
			2742: out = 24'(-10968);
			2743: out = 24'(-4696);
			2744: out = 24'(11312);
			2745: out = 24'(-23848);
			2746: out = 24'(-23048);
			2747: out = 24'(-480);
			2748: out = 24'(-14572);
			2749: out = 24'(-15124);
			2750: out = 24'(16500);
			2751: out = 24'(14120);
			2752: out = 24'(-18452);
			2753: out = 24'(-3620);
			2754: out = 24'(-10324);
			2755: out = 24'(13068);
			2756: out = 24'(35860);
			2757: out = 24'(14172);
			2758: out = 24'(24620);
			2759: out = 24'(1640);
			2760: out = 24'(-16212);
			2761: out = 24'(-24112);
			2762: out = 24'(-16884);
			2763: out = 24'(19728);
			2764: out = 24'(11528);
			2765: out = 24'(-15620);
			2766: out = 24'(820);
			2767: out = 24'(-1940);
			2768: out = 24'(-12556);
			2769: out = 24'(10676);
			2770: out = 24'(3412);
			2771: out = 24'(-29508);
			2772: out = 24'(-75088);
			2773: out = 24'(-55016);
			2774: out = 24'(8676);
			2775: out = 24'(48800);
			2776: out = 24'(-5880);
			2777: out = 24'(-65120);
			2778: out = 24'(-28444);
			2779: out = 24'(-3140);
			2780: out = 24'(30028);
			2781: out = 24'(18964);
			2782: out = 24'(16036);
			2783: out = 24'(18012);
			2784: out = 24'(11596);
			2785: out = 24'(320);
			2786: out = 24'(-33548);
			2787: out = 24'(-47172);
			2788: out = 24'(-38044);
			2789: out = 24'(-22088);
			2790: out = 24'(-30000);
			2791: out = 24'(-17580);
			2792: out = 24'(-18896);
			2793: out = 24'(2520);
			2794: out = 24'(-27880);
			2795: out = 24'(-43532);
			2796: out = 24'(-13632);
			2797: out = 24'(-8308);
			2798: out = 24'(28368);
			2799: out = 24'(47428);
			2800: out = 24'(4404);
			2801: out = 24'(-56744);
			2802: out = 24'(-33280);
			2803: out = 24'(4440);
			2804: out = 24'(27240);
			2805: out = 24'(-19904);
			2806: out = 24'(-47816);
			2807: out = 24'(-34604);
			2808: out = 24'(-27884);
			2809: out = 24'(32);
			2810: out = 24'(-4924);
			2811: out = 24'(-43160);
			2812: out = 24'(-12400);
			2813: out = 24'(35444);
			2814: out = 24'(-3672);
			2815: out = 24'(-30696);
			2816: out = 24'(-23028);
			2817: out = 24'(24332);
			2818: out = 24'(1408);
			2819: out = 24'(-26936);
			2820: out = 24'(18024);
			2821: out = 24'(51368);
			2822: out = 24'(2420);
			2823: out = 24'(-60176);
			2824: out = 24'(-58072);
			2825: out = 24'(-11320);
			2826: out = 24'(-16152);
			2827: out = 24'(-43008);
			2828: out = 24'(-29936);
			2829: out = 24'(-31700);
			2830: out = 24'(-34280);
			2831: out = 24'(-15788);
			2832: out = 24'(-30372);
			2833: out = 24'(-16108);
			2834: out = 24'(30168);
			2835: out = 24'(31692);
			2836: out = 24'(-43860);
			2837: out = 24'(-82808);
			2838: out = 24'(-45968);
			2839: out = 24'(21552);
			2840: out = 24'(65960);
			2841: out = 24'(38248);
			2842: out = 24'(-3384);
			2843: out = 24'(-47440);
			2844: out = 24'(-50952);
			2845: out = 24'(-22072);
			2846: out = 24'(9844);
			2847: out = 24'(47836);
			2848: out = 24'(18464);
			2849: out = 24'(-65596);
			2850: out = 24'(-87156);
			2851: out = 24'(-37488);
			2852: out = 24'(5248);
			2853: out = 24'(18696);
			2854: out = 24'(10852);
			2855: out = 24'(-17264);
			2856: out = 24'(-72732);
			2857: out = 24'(-45796);
			2858: out = 24'(-1056);
			2859: out = 24'(27352);
			2860: out = 24'(40028);
			2861: out = 24'(-22540);
			2862: out = 24'(-79956);
			2863: out = 24'(-70876);
			2864: out = 24'(-1728);
			2865: out = 24'(46396);
			2866: out = 24'(27520);
			2867: out = 24'(27180);
			2868: out = 24'(15316);
			2869: out = 24'(-5032);
			2870: out = 24'(-31312);
			2871: out = 24'(-54984);
			2872: out = 24'(-33140);
			2873: out = 24'(5912);
			2874: out = 24'(34412);
			2875: out = 24'(-1220);
			2876: out = 24'(5296);
			2877: out = 24'(-6200);
			2878: out = 24'(22824);
			2879: out = 24'(6020);
			2880: out = 24'(-2424);
			2881: out = 24'(5964);
			2882: out = 24'(18212);
			2883: out = 24'(19192);
			2884: out = 24'(-13728);
			2885: out = 24'(-40504);
			2886: out = 24'(-27388);
			2887: out = 24'(-12420);
			2888: out = 24'(-27884);
			2889: out = 24'(-38596);
			2890: out = 24'(-24304);
			2891: out = 24'(6144);
			2892: out = 24'(-9196);
			2893: out = 24'(-63348);
			2894: out = 24'(-83092);
			2895: out = 24'(-22976);
			2896: out = 24'(24000);
			2897: out = 24'(42504);
			2898: out = 24'(25624);
			2899: out = 24'(-27636);
			2900: out = 24'(-38792);
			2901: out = 24'(-24948);
			2902: out = 24'(-9004);
			2903: out = 24'(23536);
			2904: out = 24'(-580);
			2905: out = 24'(-12824);
			2906: out = 24'(20416);
			2907: out = 24'(42792);
			2908: out = 24'(22256);
			2909: out = 24'(-16984);
			2910: out = 24'(-37440);
			2911: out = 24'(-1272);
			2912: out = 24'(14588);
			2913: out = 24'(-22648);
			2914: out = 24'(-26616);
			2915: out = 24'(-19524);
			2916: out = 24'(-26700);
			2917: out = 24'(-17976);
			2918: out = 24'(33356);
			2919: out = 24'(12556);
			2920: out = 24'(-27228);
			2921: out = 24'(31208);
			2922: out = 24'(59636);
			2923: out = 24'(33312);
			2924: out = 24'(-26968);
			2925: out = 24'(-39612);
			2926: out = 24'(2216);
			2927: out = 24'(26384);
			2928: out = 24'(-2736);
			2929: out = 24'(-32544);
			2930: out = 24'(-51336);
			2931: out = 24'(-60020);
			2932: out = 24'(-7596);
			2933: out = 24'(57208);
			2934: out = 24'(47436);
			2935: out = 24'(22240);
			2936: out = 24'(5148);
			2937: out = 24'(-36908);
			2938: out = 24'(-48472);
			2939: out = 24'(14300);
			2940: out = 24'(61624);
			2941: out = 24'(31884);
			2942: out = 24'(-11592);
			2943: out = 24'(-42108);
			2944: out = 24'(-23380);
			2945: out = 24'(31252);
			2946: out = 24'(45356);
			2947: out = 24'(16352);
			2948: out = 24'(25284);
			2949: out = 24'(9604);
			2950: out = 24'(-18108);
			2951: out = 24'(-20368);
			2952: out = 24'(32868);
			2953: out = 24'(66616);
			2954: out = 24'(42596);
			2955: out = 24'(-38336);
			2956: out = 24'(-44572);
			2957: out = 24'(8796);
			2958: out = 24'(72960);
			2959: out = 24'(65120);
			2960: out = 24'(3488);
			2961: out = 24'(-25848);
			2962: out = 24'(-24948);
			2963: out = 24'(18696);
			2964: out = 24'(47140);
			2965: out = 24'(28256);
			2966: out = 24'(-30548);
			2967: out = 24'(-51244);
			2968: out = 24'(-7604);
			2969: out = 24'(67008);
			2970: out = 24'(59228);
			2971: out = 24'(14948);
			2972: out = 24'(-9244);
			2973: out = 24'(42804);
			2974: out = 24'(56208);
			2975: out = 24'(17560);
			2976: out = 24'(-1884);
			2977: out = 24'(20352);
			2978: out = 24'(7004);
			2979: out = 24'(-14644);
			2980: out = 24'(3200);
			2981: out = 24'(4744);
			2982: out = 24'(1884);
			2983: out = 24'(-7748);
			2984: out = 24'(10000);
			2985: out = 24'(45388);
			2986: out = 24'(97908);
			2987: out = 24'(39916);
			2988: out = 24'(-26388);
			2989: out = 24'(-25348);
			2990: out = 24'(8432);
			2991: out = 24'(52720);
			2992: out = 24'(47716);
			2993: out = 24'(41772);
			2994: out = 24'(43988);
			2995: out = 24'(20628);
			2996: out = 24'(-41460);
			2997: out = 24'(-63852);
			2998: out = 24'(268);
			2999: out = 24'(34904);
			3000: out = 24'(11452);
			3001: out = 24'(33100);
			3002: out = 24'(30120);
			3003: out = 24'(-9092);
			3004: out = 24'(-10980);
			3005: out = 24'(-4112);
			3006: out = 24'(26800);
			3007: out = 24'(52992);
			3008: out = 24'(43556);
			3009: out = 24'(12596);
			3010: out = 24'(-4708);
			3011: out = 24'(36588);
			3012: out = 24'(78692);
			3013: out = 24'(52984);
			3014: out = 24'(-3852);
			3015: out = 24'(-20260);
			3016: out = 24'(-29568);
			3017: out = 24'(-27368);
			3018: out = 24'(-17576);
			3019: out = 24'(5384);
			3020: out = 24'(37072);
			3021: out = 24'(60088);
			3022: out = 24'(54712);
			3023: out = 24'(8000);
			3024: out = 24'(-860);
			3025: out = 24'(33984);
			3026: out = 24'(74836);
			3027: out = 24'(49720);
			3028: out = 24'(-20316);
			3029: out = 24'(-47292);
			3030: out = 24'(-22504);
			3031: out = 24'(20096);
			3032: out = 24'(49804);
			3033: out = 24'(-12416);
			3034: out = 24'(-30776);
			3035: out = 24'(29320);
			3036: out = 24'(92944);
			3037: out = 24'(53580);
			3038: out = 24'(-1800);
			3039: out = 24'(-19088);
			3040: out = 24'(496);
			3041: out = 24'(29748);
			3042: out = 24'(39444);
			3043: out = 24'(33456);
			3044: out = 24'(4892);
			3045: out = 24'(-17052);
			3046: out = 24'(528);
			3047: out = 24'(34856);
			3048: out = 24'(6588);
			3049: out = 24'(-70684);
			3050: out = 24'(-68472);
			3051: out = 24'(-6024);
			3052: out = 24'(42412);
			3053: out = 24'(62752);
			3054: out = 24'(50288);
			3055: out = 24'(21604);
			3056: out = 24'(-2484);
			3057: out = 24'(-32168);
			3058: out = 24'(-40364);
			3059: out = 24'(-16092);
			3060: out = 24'(43596);
			3061: out = 24'(58600);
			3062: out = 24'(33180);
			3063: out = 24'(46924);
			3064: out = 24'(48404);
			3065: out = 24'(30916);
			3066: out = 24'(-18232);
			3067: out = 24'(-39916);
			3068: out = 24'(-32012);
			3069: out = 24'(17372);
			3070: out = 24'(39728);
			3071: out = 24'(6700);
			3072: out = 24'(-732);
			3073: out = 24'(6696);
			3074: out = 24'(-13332);
			3075: out = 24'(-18600);
			3076: out = 24'(-9300);
			3077: out = 24'(10116);
			3078: out = 24'(25092);
			3079: out = 24'(22072);
			3080: out = 24'(-6656);
			3081: out = 24'(-7360);
			3082: out = 24'(7552);
			3083: out = 24'(-13456);
			3084: out = 24'(-5288);
			3085: out = 24'(17584);
			3086: out = 24'(-4952);
			3087: out = 24'(-18208);
			3088: out = 24'(-2324);
			3089: out = 24'(12336);
			3090: out = 24'(31344);
			3091: out = 24'(19748);
			3092: out = 24'(-24412);
			3093: out = 24'(-22476);
			3094: out = 24'(-16788);
			3095: out = 24'(12224);
			3096: out = 24'(30628);
			3097: out = 24'(6224);
			3098: out = 24'(28552);
			3099: out = 24'(49896);
			3100: out = 24'(29444);
			3101: out = 24'(-37068);
			3102: out = 24'(-78388);
			3103: out = 24'(-75320);
			3104: out = 24'(-17140);
			3105: out = 24'(47036);
			3106: out = 24'(27236);
			3107: out = 24'(13376);
			3108: out = 24'(32700);
			3109: out = 24'(22808);
			3110: out = 24'(668);
			3111: out = 24'(-22924);
			3112: out = 24'(7296);
			3113: out = 24'(52508);
			3114: out = 24'(43080);
			3115: out = 24'(-20512);
			3116: out = 24'(-59628);
			3117: out = 24'(-41144);
			3118: out = 24'(-35344);
			3119: out = 24'(-18864);
			3120: out = 24'(-1820);
			3121: out = 24'(-11276);
			3122: out = 24'(8228);
			3123: out = 24'(37820);
			3124: out = 24'(47972);
			3125: out = 24'(26016);
			3126: out = 24'(-34884);
			3127: out = 24'(-66324);
			3128: out = 24'(-46696);
			3129: out = 24'(-7340);
			3130: out = 24'(-1036);
			3131: out = 24'(-10000);
			3132: out = 24'(6508);
			3133: out = 24'(18796);
			3134: out = 24'(25964);
			3135: out = 24'(19340);
			3136: out = 24'(-18920);
			3137: out = 24'(-45556);
			3138: out = 24'(-13940);
			3139: out = 24'(-3972);
			3140: out = 24'(-34820);
			3141: out = 24'(-48832);
			3142: out = 24'(-53776);
			3143: out = 24'(6164);
			3144: out = 24'(42168);
			3145: out = 24'(6040);
			3146: out = 24'(22092);
			3147: out = 24'(35336);
			3148: out = 24'(9604);
			3149: out = 24'(-44300);
			3150: out = 24'(-72276);
			3151: out = 24'(-51300);
			3152: out = 24'(-40476);
			3153: out = 24'(-2624);
			3154: out = 24'(45384);
			3155: out = 24'(15960);
			3156: out = 24'(-9832);
			3157: out = 24'(-7392);
			3158: out = 24'(8024);
			3159: out = 24'(648);
			3160: out = 24'(-46448);
			3161: out = 24'(-74200);
			3162: out = 24'(-44208);
			3163: out = 24'(8884);
			3164: out = 24'(27016);
			3165: out = 24'(-23340);
			3166: out = 24'(-58132);
			3167: out = 24'(-25976);
			3168: out = 24'(42644);
			3169: out = 24'(40508);
			3170: out = 24'(-21436);
			3171: out = 24'(-79264);
			3172: out = 24'(-59468);
			3173: out = 24'(-12844);
			3174: out = 24'(15212);
			3175: out = 24'(33752);
			3176: out = 24'(-9908);
			3177: out = 24'(-47408);
			3178: out = 24'(-46180);
			3179: out = 24'(-39000);
			3180: out = 24'(14624);
			3181: out = 24'(51132);
			3182: out = 24'(4476);
			3183: out = 24'(-29496);
			3184: out = 24'(-29428);
			3185: out = 24'(-14336);
			3186: out = 24'(-12428);
			3187: out = 24'(-35716);
			3188: out = 24'(-70604);
			3189: out = 24'(-26956);
			3190: out = 24'(4748);
			3191: out = 24'(-2844);
			3192: out = 24'(39016);
			3193: out = 24'(38124);
			3194: out = 24'(-21616);
			3195: out = 24'(-38996);
			3196: out = 24'(-40084);
			3197: out = 24'(-36552);
			3198: out = 24'(-34460);
			3199: out = 24'(18780);
			3200: out = 24'(40680);
			3201: out = 24'(-21024);
			3202: out = 24'(-47240);
			3203: out = 24'(-18436);
			3204: out = 24'(37860);
			3205: out = 24'(53484);
			3206: out = 24'(-15856);
			3207: out = 24'(-47028);
			3208: out = 24'(-32276);
			3209: out = 24'(-14948);
			3210: out = 24'(21424);
			3211: out = 24'(8452);
			3212: out = 24'(-51136);
			3213: out = 24'(-45700);
			3214: out = 24'(-17736);
			3215: out = 24'(10220);
			3216: out = 24'(3080);
			3217: out = 24'(-30208);
			3218: out = 24'(-52016);
			3219: out = 24'(-34476);
			3220: out = 24'(-13032);
			3221: out = 24'(-2092);
			3222: out = 24'(-33576);
			3223: out = 24'(-49232);
			3224: out = 24'(12816);
			3225: out = 24'(18512);
			3226: out = 24'(3448);
			3227: out = 24'(-3284);
			3228: out = 24'(-20572);
			3229: out = 24'(-35416);
			3230: out = 24'(-16604);
			3231: out = 24'(-9108);
			3232: out = 24'(-7736);
			3233: out = 24'(38020);
			3234: out = 24'(1588);
			3235: out = 24'(-25608);
			3236: out = 24'(-8468);
			3237: out = 24'(8788);
			3238: out = 24'(9916);
			3239: out = 24'(-24528);
			3240: out = 24'(-3004);
			3241: out = 24'(27524);
			3242: out = 24'(6192);
			3243: out = 24'(-44968);
			3244: out = 24'(-30120);
			3245: out = 24'(-1012);
			3246: out = 24'(11872);
			3247: out = 24'(-5976);
			3248: out = 24'(-12668);
			3249: out = 24'(12620);
			3250: out = 24'(24180);
			3251: out = 24'(-6700);
			3252: out = 24'(-39712);
			3253: out = 24'(-38672);
			3254: out = 24'(-3236);
			3255: out = 24'(-2708);
			3256: out = 24'(-13440);
			3257: out = 24'(18568);
			3258: out = 24'(48672);
			3259: out = 24'(30080);
			3260: out = 24'(7640);
			3261: out = 24'(-23324);
			3262: out = 24'(-4324);
			3263: out = 24'(-2420);
			3264: out = 24'(17472);
			3265: out = 24'(36540);
			3266: out = 24'(13068);
			3267: out = 24'(7300);
			3268: out = 24'(10988);
			3269: out = 24'(-22108);
			3270: out = 24'(-28888);
			3271: out = 24'(-680);
			3272: out = 24'(7572);
			3273: out = 24'(-13908);
			3274: out = 24'(-37004);
			3275: out = 24'(11628);
			3276: out = 24'(12560);
			3277: out = 24'(-45712);
			3278: out = 24'(-23292);
			3279: out = 24'(33980);
			3280: out = 24'(16108);
			3281: out = 24'(-1992);
			3282: out = 24'(40092);
			3283: out = 24'(39580);
			3284: out = 24'(-27352);
			3285: out = 24'(-57668);
			3286: out = 24'(-50204);
			3287: out = 24'(-11388);
			3288: out = 24'(57304);
			3289: out = 24'(41596);
			3290: out = 24'(-15380);
			3291: out = 24'(3084);
			3292: out = 24'(48824);
			3293: out = 24'(69040);
			3294: out = 24'(13180);
			3295: out = 24'(-60808);
			3296: out = 24'(-40304);
			3297: out = 24'(32680);
			3298: out = 24'(57400);
			3299: out = 24'(12224);
			3300: out = 24'(-29040);
			3301: out = 24'(-13416);
			3302: out = 24'(42280);
			3303: out = 24'(51204);
			3304: out = 24'(42504);
			3305: out = 24'(22992);
			3306: out = 24'(-5332);
			3307: out = 24'(-18284);
			3308: out = 24'(-21564);
			3309: out = 24'(29816);
			3310: out = 24'(25016);
			3311: out = 24'(-22676);
			3312: out = 24'(-2408);
			3313: out = 24'(33984);
			3314: out = 24'(49320);
			3315: out = 24'(31964);
			3316: out = 24'(-8752);
			3317: out = 24'(2012);
			3318: out = 24'(20088);
			3319: out = 24'(37576);
			3320: out = 24'(-9384);
			3321: out = 24'(-40784);
			3322: out = 24'(-7912);
			3323: out = 24'(19528);
			3324: out = 24'(50124);
			3325: out = 24'(54044);
			3326: out = 24'(7252);
			3327: out = 24'(-23544);
			3328: out = 24'(-34436);
			3329: out = 24'(8788);
			3330: out = 24'(53636);
			3331: out = 24'(40232);
			3332: out = 24'(19380);
			3333: out = 24'(-2684);
			3334: out = 24'(-18776);
			3335: out = 24'(-61176);
			3336: out = 24'(-64172);
			3337: out = 24'(23860);
			3338: out = 24'(83024);
			3339: out = 24'(54772);
			3340: out = 24'(-3180);
			3341: out = 24'(-24684);
			3342: out = 24'(17468);
			3343: out = 24'(56684);
			3344: out = 24'(60020);
			3345: out = 24'(26968);
			3346: out = 24'(3900);
			3347: out = 24'(-17940);
			3348: out = 24'(8404);
			3349: out = 24'(17996);
			3350: out = 24'(2060);
			3351: out = 24'(-10536);
			3352: out = 24'(1740);
			3353: out = 24'(-4720);
			3354: out = 24'(12012);
			3355: out = 24'(49068);
			3356: out = 24'(20924);
			3357: out = 24'(-4244);
			3358: out = 24'(-20572);
			3359: out = 24'(-15232);
			3360: out = 24'(17052);
			3361: out = 24'(85512);
			3362: out = 24'(66040);
			3363: out = 24'(-11284);
			3364: out = 24'(-46848);
			3365: out = 24'(-8548);
			3366: out = 24'(33912);
			3367: out = 24'(46084);
			3368: out = 24'(-8656);
			3369: out = 24'(-21584);
			3370: out = 24'(14048);
			3371: out = 24'(35364);
			3372: out = 24'(36212);
			3373: out = 24'(16824);
			3374: out = 24'(-10964);
			3375: out = 24'(-20148);
			3376: out = 24'(-30352);
			3377: out = 24'(-25020);
			3378: out = 24'(3588);
			3379: out = 24'(21588);
			3380: out = 24'(38736);
			3381: out = 24'(-13196);
			3382: out = 24'(-27536);
			3383: out = 24'(-15728);
			3384: out = 24'(32944);
			3385: out = 24'(75172);
			3386: out = 24'(58224);
			3387: out = 24'(1812);
			3388: out = 24'(-36152);
			3389: out = 24'(-14996);
			3390: out = 24'(-12004);
			3391: out = 24'(16768);
			3392: out = 24'(26696);
			3393: out = 24'(5948);
			3394: out = 24'(-7588);
			3395: out = 24'(17116);
			3396: out = 24'(-13584);
			3397: out = 24'(-34800);
			3398: out = 24'(-4088);
			3399: out = 24'(18644);
			3400: out = 24'(-1416);
			3401: out = 24'(-24588);
			3402: out = 24'(-26896);
			3403: out = 24'(-32864);
			3404: out = 24'(15696);
			3405: out = 24'(34944);
			3406: out = 24'(20760);
			3407: out = 24'(23588);
			3408: out = 24'(14000);
			3409: out = 24'(-644);
			3410: out = 24'(10800);
			3411: out = 24'(3712);
			3412: out = 24'(-744);
			3413: out = 24'(33748);
			3414: out = 24'(46048);
			3415: out = 24'(-12916);
			3416: out = 24'(-58468);
			3417: out = 24'(-31764);
			3418: out = 24'(35292);
			3419: out = 24'(46000);
			3420: out = 24'(-6596);
			3421: out = 24'(-31252);
			3422: out = 24'(-2896);
			3423: out = 24'(21504);
			3424: out = 24'(6128);
			3425: out = 24'(-15760);
			3426: out = 24'(7932);
			3427: out = 24'(27560);
			3428: out = 24'(15940);
			3429: out = 24'(-17360);
			3430: out = 24'(-38328);
			3431: out = 24'(-42312);
			3432: out = 24'(-61852);
			3433: out = 24'(-13464);
			3434: out = 24'(33808);
			3435: out = 24'(28244);
			3436: out = 24'(6196);
			3437: out = 24'(11136);
			3438: out = 24'(22420);
			3439: out = 24'(11936);
			3440: out = 24'(-10540);
			3441: out = 24'(-33812);
			3442: out = 24'(-20916);
			3443: out = 24'(-3120);
			3444: out = 24'(13840);
			3445: out = 24'(10284);
			3446: out = 24'(-5276);
			3447: out = 24'(16516);
			3448: out = 24'(33808);
			3449: out = 24'(22436);
			3450: out = 24'(-29108);
			3451: out = 24'(-28180);
			3452: out = 24'(-27148);
			3453: out = 24'(21888);
			3454: out = 24'(19508);
			3455: out = 24'(-21132);
			3456: out = 24'(-11260);
			3457: out = 24'(26624);
			3458: out = 24'(49432);
			3459: out = 24'(11936);
			3460: out = 24'(-41256);
			3461: out = 24'(-40644);
			3462: out = 24'(-15332);
			3463: out = 24'(48884);
			3464: out = 24'(51096);
			3465: out = 24'(-18532);
			3466: out = 24'(-40400);
			3467: out = 24'(-18052);
			3468: out = 24'(-5672);
			3469: out = 24'(-6340);
			3470: out = 24'(-11076);
			3471: out = 24'(-28648);
			3472: out = 24'(-27272);
			3473: out = 24'(-45388);
			3474: out = 24'(8960);
			3475: out = 24'(17336);
			3476: out = 24'(-28044);
			3477: out = 24'(-2900);
			3478: out = 24'(55704);
			3479: out = 24'(26820);
			3480: out = 24'(-42224);
			3481: out = 24'(-37944);
			3482: out = 24'(-13096);
			3483: out = 24'(-13004);
			3484: out = 24'(4224);
			3485: out = 24'(14832);
			3486: out = 24'(-8196);
			3487: out = 24'(-38924);
			3488: out = 24'(-23968);
			3489: out = 24'(19624);
			3490: out = 24'(28912);
			3491: out = 24'(24152);
			3492: out = 24'(-26052);
			3493: out = 24'(-45948);
			3494: out = 24'(-27756);
			3495: out = 24'(11264);
			3496: out = 24'(4616);
			3497: out = 24'(-29492);
			3498: out = 24'(9692);
			3499: out = 24'(26660);
			3500: out = 24'(6924);
			3501: out = 24'(27692);
			3502: out = 24'(15980);
			3503: out = 24'(-492);
			3504: out = 24'(-28676);
			3505: out = 24'(-44216);
			3506: out = 24'(-14004);
			3507: out = 24'(32000);
			3508: out = 24'(12256);
			3509: out = 24'(-60148);
			3510: out = 24'(-68292);
			3511: out = 24'(-7396);
			3512: out = 24'(35696);
			3513: out = 24'(30076);
			3514: out = 24'(13640);
			3515: out = 24'(4160);
			3516: out = 24'(-3744);
			3517: out = 24'(-36416);
			3518: out = 24'(-7412);
			3519: out = 24'(47296);
			3520: out = 24'(7540);
			3521: out = 24'(-53528);
			3522: out = 24'(-41880);
			3523: out = 24'(2880);
			3524: out = 24'(-8000);
			3525: out = 24'(-35324);
			3526: out = 24'(-6176);
			3527: out = 24'(15376);
			3528: out = 24'(41176);
			3529: out = 24'(32888);
			3530: out = 24'(-12956);
			3531: out = 24'(-67676);
			3532: out = 24'(-80276);
			3533: out = 24'(-26052);
			3534: out = 24'(39336);
			3535: out = 24'(69800);
			3536: out = 24'(2736);
			3537: out = 24'(-47180);
			3538: out = 24'(-20988);
			3539: out = 24'(22928);
			3540: out = 24'(57708);
			3541: out = 24'(10736);
			3542: out = 24'(-24632);
			3543: out = 24'(-4628);
			3544: out = 24'(11568);
			3545: out = 24'(-940);
			3546: out = 24'(-32252);
			3547: out = 24'(-21972);
			3548: out = 24'(15384);
			3549: out = 24'(12184);
			3550: out = 24'(-5164);
			3551: out = 24'(-14208);
			3552: out = 24'(-1988);
			3553: out = 24'(-7704);
			3554: out = 24'(-6740);
			3555: out = 24'(-4680);
			3556: out = 24'(-30968);
			3557: out = 24'(-36704);
			3558: out = 24'(1060);
			3559: out = 24'(18876);
			3560: out = 24'(524);
			3561: out = 24'(-13756);
			3562: out = 24'(-44564);
			3563: out = 24'(-61064);
			3564: out = 24'(-12308);
			3565: out = 24'(-9168);
			3566: out = 24'(-5844);
			3567: out = 24'(24548);
			3568: out = 24'(8296);
			3569: out = 24'(12248);
			3570: out = 24'(22388);
			3571: out = 24'(32788);
			3572: out = 24'(12344);
			3573: out = 24'(-25500);
			3574: out = 24'(-12096);
			3575: out = 24'(-2448);
			3576: out = 24'(-1032);
			3577: out = 24'(-27504);
			3578: out = 24'(-29852);
			3579: out = 24'(-2052);
			3580: out = 24'(-3224);
			3581: out = 24'(-52236);
			3582: out = 24'(-45792);
			3583: out = 24'(9596);
			3584: out = 24'(26640);
			3585: out = 24'(-7208);
			3586: out = 24'(-25456);
			3587: out = 24'(-39440);
			3588: out = 24'(-18396);
			3589: out = 24'(43508);
			3590: out = 24'(65604);
			3591: out = 24'(8828);
			3592: out = 24'(-45276);
			3593: out = 24'(-47180);
			3594: out = 24'(-5972);
			3595: out = 24'(32092);
			3596: out = 24'(8804);
			3597: out = 24'(-7060);
			3598: out = 24'(17892);
			3599: out = 24'(-6032);
			3600: out = 24'(-40832);
			3601: out = 24'(-48148);
			3602: out = 24'(-36664);
			3603: out = 24'(30300);
			3604: out = 24'(78300);
			3605: out = 24'(20668);
			3606: out = 24'(-48576);
			3607: out = 24'(-43572);
			3608: out = 24'(-1332);
			3609: out = 24'(35604);
			3610: out = 24'(1808);
			3611: out = 24'(-17136);
			3612: out = 24'(420);
			3613: out = 24'(19176);
			3614: out = 24'(34412);
			3615: out = 24'(-3232);
			3616: out = 24'(-39764);
			3617: out = 24'(-14980);
			3618: out = 24'(2912);
			3619: out = 24'(18452);
			3620: out = 24'(13144);
			3621: out = 24'(-8200);
			3622: out = 24'(-736);
			3623: out = 24'(-27396);
			3624: out = 24'(-40752);
			3625: out = 24'(-26860);
			3626: out = 24'(2164);
			3627: out = 24'(25356);
			3628: out = 24'(-1040);
			3629: out = 24'(-6756);
			3630: out = 24'(-9676);
			3631: out = 24'(9240);
			3632: out = 24'(45336);
			3633: out = 24'(49112);
			3634: out = 24'(10544);
			3635: out = 24'(-31780);
			3636: out = 24'(-9304);
			3637: out = 24'(4976);
			3638: out = 24'(28988);
			3639: out = 24'(10736);
			3640: out = 24'(-6848);
			3641: out = 24'(-7988);
			3642: out = 24'(-13248);
			3643: out = 24'(30880);
			3644: out = 24'(45980);
			3645: out = 24'(-3560);
			3646: out = 24'(-41960);
			3647: out = 24'(-29028);
			3648: out = 24'(-26168);
			3649: out = 24'(-18116);
			3650: out = 24'(3244);
			3651: out = 24'(-12196);
			3652: out = 24'(-6072);
			3653: out = 24'(14988);
			3654: out = 24'(-4168);
			3655: out = 24'(-24016);
			3656: out = 24'(-36804);
			3657: out = 24'(-19600);
			3658: out = 24'(6960);
			3659: out = 24'(26728);
			3660: out = 24'(23036);
			3661: out = 24'(1568);
			3662: out = 24'(2888);
			3663: out = 24'(10464);
			3664: out = 24'(-5808);
			3665: out = 24'(-9512);
			3666: out = 24'(-172);
			3667: out = 24'(2280);
			3668: out = 24'(9520);
			3669: out = 24'(17268);
			3670: out = 24'(-27068);
			3671: out = 24'(-41876);
			3672: out = 24'(-2756);
			3673: out = 24'(26980);
			3674: out = 24'(31032);
			3675: out = 24'(24308);
			3676: out = 24'(15712);
			3677: out = 24'(-16996);
			3678: out = 24'(-37844);
			3679: out = 24'(-26008);
			3680: out = 24'(-2328);
			3681: out = 24'(9940);
			3682: out = 24'(43608);
			3683: out = 24'(27232);
			3684: out = 24'(-13612);
			3685: out = 24'(-38876);
			3686: out = 24'(-48440);
			3687: out = 24'(15580);
			3688: out = 24'(60644);
			3689: out = 24'(28056);
			3690: out = 24'(10300);
			3691: out = 24'(25520);
			3692: out = 24'(-5592);
			3693: out = 24'(-54136);
			3694: out = 24'(-76160);
			3695: out = 24'(-43656);
			3696: out = 24'(41872);
			3697: out = 24'(75724);
			3698: out = 24'(17364);
			3699: out = 24'(-18032);
			3700: out = 24'(-5552);
			3701: out = 24'(33416);
			3702: out = 24'(70660);
			3703: out = 24'(27056);
			3704: out = 24'(-17740);
			3705: out = 24'(-19620);
			3706: out = 24'(-11396);
			3707: out = 24'(-22456);
			3708: out = 24'(-17184);
			3709: out = 24'(-216);
			3710: out = 24'(17960);
			3711: out = 24'(30224);
			3712: out = 24'(33448);
			3713: out = 24'(-1144);
			3714: out = 24'(-17028);
			3715: out = 24'(22920);
			3716: out = 24'(12588);
			3717: out = 24'(16792);
			3718: out = 24'(11544);
			3719: out = 24'(21468);
			3720: out = 24'(17728);
			3721: out = 24'(6688);
			3722: out = 24'(20264);
			3723: out = 24'(10180);
			3724: out = 24'(-9728);
			3725: out = 24'(-32304);
			3726: out = 24'(-47584);
			3727: out = 24'(2368);
			3728: out = 24'(55688);
			3729: out = 24'(15044);
			3730: out = 24'(-36992);
			3731: out = 24'(-28604);
			3732: out = 24'(46232);
			3733: out = 24'(59124);
			3734: out = 24'(-14160);
			3735: out = 24'(-11468);
			3736: out = 24'(12660);
			3737: out = 24'(10868);
			3738: out = 24'(17916);
			3739: out = 24'(28796);
			3740: out = 24'(14396);
			3741: out = 24'(-2456);
			3742: out = 24'(-28772);
			3743: out = 24'(-58828);
			3744: out = 24'(-2960);
			3745: out = 24'(34820);
			3746: out = 24'(12568);
			3747: out = 24'(7268);
			3748: out = 24'(35744);
			3749: out = 24'(26552);
			3750: out = 24'(14060);
			3751: out = 24'(12496);
			3752: out = 24'(2772);
			3753: out = 24'(5008);
			3754: out = 24'(-32472);
			3755: out = 24'(-26600);
			3756: out = 24'(24716);
			3757: out = 24'(41508);
			3758: out = 24'(34012);
			3759: out = 24'(-7800);
			3760: out = 24'(-33700);
			3761: out = 24'(-10700);
			3762: out = 24'(16956);
			3763: out = 24'(51380);
			3764: out = 24'(56468);
			3765: out = 24'(17096);
			3766: out = 24'(4160);
			3767: out = 24'(16060);
			3768: out = 24'(-5504);
			3769: out = 24'(-2148);
			3770: out = 24'(-23308);
			3771: out = 24'(-24492);
			3772: out = 24'(26388);
			3773: out = 24'(53580);
			3774: out = 24'(22884);
			3775: out = 24'(-14092);
			3776: out = 24'(-21832);
			3777: out = 24'(38316);
			3778: out = 24'(52932);
			3779: out = 24'(14076);
			3780: out = 24'(-7072);
			3781: out = 24'(-1024);
			3782: out = 24'(-8144);
			3783: out = 24'(-34108);
			3784: out = 24'(-35068);
			3785: out = 24'(11780);
			3786: out = 24'(46804);
			3787: out = 24'(18060);
			3788: out = 24'(10352);
			3789: out = 24'(13976);
			3790: out = 24'(17368);
			3791: out = 24'(-10360);
			3792: out = 24'(-51084);
			3793: out = 24'(-35192);
			3794: out = 24'(-3236);
			3795: out = 24'(21000);
			3796: out = 24'(44856);
			3797: out = 24'(12736);
			3798: out = 24'(22808);
			3799: out = 24'(46332);
			3800: out = 24'(41160);
			3801: out = 24'(-8424);
			3802: out = 24'(-50452);
			3803: out = 24'(-41376);
			3804: out = 24'(-1436);
			3805: out = 24'(51656);
			3806: out = 24'(40896);
			3807: out = 24'(-11824);
			3808: out = 24'(1784);
			3809: out = 24'(43440);
			3810: out = 24'(55632);
			3811: out = 24'(-5296);
			3812: out = 24'(-22240);
			3813: out = 24'(-2768);
			3814: out = 24'(31232);
			3815: out = 24'(52620);
			3816: out = 24'(33960);
			3817: out = 24'(13676);
			3818: out = 24'(9692);
			3819: out = 24'(-4652);
			3820: out = 24'(-22588);
			3821: out = 24'(-18504);
			3822: out = 24'(-17096);
			3823: out = 24'(-31068);
			3824: out = 24'(-14680);
			3825: out = 24'(23968);
			3826: out = 24'(-7872);
			3827: out = 24'(-69704);
			3828: out = 24'(-58088);
			3829: out = 24'(-31628);
			3830: out = 24'(-12028);
			3831: out = 24'(57104);
			3832: out = 24'(57620);
			3833: out = 24'(-27704);
			3834: out = 24'(-73672);
			3835: out = 24'(-34416);
			3836: out = 24'(12492);
			3837: out = 24'(71664);
			3838: out = 24'(62644);
			3839: out = 24'(232);
			3840: out = 24'(-29856);
			3841: out = 24'(-10180);
			3842: out = 24'(29564);
			3843: out = 24'(5104);
			3844: out = 24'(-25704);
			3845: out = 24'(9212);
			3846: out = 24'(-3084);
			3847: out = 24'(-37692);
			3848: out = 24'(-13552);
			3849: out = 24'(-4888);
			3850: out = 24'(15464);
			3851: out = 24'(40884);
			3852: out = 24'(35392);
			3853: out = 24'(-10588);
			3854: out = 24'(-33072);
			3855: out = 24'(-12832);
			3856: out = 24'(49944);
			3857: out = 24'(46220);
			3858: out = 24'(-6148);
			3859: out = 24'(-26784);
			3860: out = 24'(1196);
			3861: out = 24'(25708);
			3862: out = 24'(3868);
			3863: out = 24'(-65664);
			3864: out = 24'(-56708);
			3865: out = 24'(-6060);
			3866: out = 24'(23980);
			3867: out = 24'(31556);
			3868: out = 24'(10760);
			3869: out = 24'(27864);
			3870: out = 24'(24776);
			3871: out = 24'(-4440);
			3872: out = 24'(-36760);
			3873: out = 24'(-53800);
			3874: out = 24'(-25824);
			3875: out = 24'(15052);
			3876: out = 24'(25704);
			3877: out = 24'(13728);
			3878: out = 24'(-25360);
			3879: out = 24'(-4432);
			3880: out = 24'(2528);
			3881: out = 24'(11416);
			3882: out = 24'(22440);
			3883: out = 24'(52972);
			3884: out = 24'(49144);
			3885: out = 24'(-13068);
			3886: out = 24'(-55660);
			3887: out = 24'(-48320);
			3888: out = 24'(-9616);
			3889: out = 24'(2140);
			3890: out = 24'(-24588);
			3891: out = 24'(-28632);
			3892: out = 24'(-1036);
			3893: out = 24'(-8732);
			3894: out = 24'(-20740);
			3895: out = 24'(-8784);
			3896: out = 24'(15964);
			3897: out = 24'(12768);
			3898: out = 24'(-33824);
			3899: out = 24'(-45624);
			3900: out = 24'(-23880);
			3901: out = 24'(28712);
			3902: out = 24'(45936);
			3903: out = 24'(-14224);
			3904: out = 24'(-26708);
			3905: out = 24'(-796);
			3906: out = 24'(1388);
			3907: out = 24'(9232);
			3908: out = 24'(-21368);
			3909: out = 24'(-39764);
			3910: out = 24'(1772);
			3911: out = 24'(4524);
			3912: out = 24'(-8512);
			3913: out = 24'(14156);
			3914: out = 24'(23328);
			3915: out = 24'(18124);
			3916: out = 24'(-17420);
			3917: out = 24'(-60692);
			3918: out = 24'(-27172);
			3919: out = 24'(17112);
			3920: out = 24'(15900);
			3921: out = 24'(-15892);
			3922: out = 24'(-12996);
			3923: out = 24'(-672);
			3924: out = 24'(-2008);
			3925: out = 24'(-13892);
			3926: out = 24'(-36844);
			3927: out = 24'(-7176);
			3928: out = 24'(6388);
			3929: out = 24'(8920);
			3930: out = 24'(5484);
			3931: out = 24'(-9212);
			3932: out = 24'(-3636);
			3933: out = 24'(7376);
			3934: out = 24'(-31824);
			3935: out = 24'(-27400);
			3936: out = 24'(-3780);
			3937: out = 24'(9292);
			3938: out = 24'(31048);
			3939: out = 24'(28836);
			3940: out = 24'(9332);
			3941: out = 24'(-28292);
			3942: out = 24'(-60396);
			3943: out = 24'(-44932);
			3944: out = 24'(-23336);
			3945: out = 24'(14480);
			3946: out = 24'(34440);
			3947: out = 24'(-29348);
			3948: out = 24'(-64020);
			3949: out = 24'(-58940);
			3950: out = 24'(-10064);
			3951: out = 24'(60216);
			3952: out = 24'(77408);
			3953: out = 24'(-8668);
			3954: out = 24'(-91164);
			3955: out = 24'(-78144);
			3956: out = 24'(-25984);
			3957: out = 24'(56400);
			3958: out = 24'(50612);
			3959: out = 24'(-21804);
			3960: out = 24'(-15892);
			3961: out = 24'(29876);
			3962: out = 24'(27032);
			3963: out = 24'(-1020);
			3964: out = 24'(-27856);
			3965: out = 24'(-15188);
			3966: out = 24'(-7908);
			3967: out = 24'(52);
			3968: out = 24'(-1936);
			3969: out = 24'(-27556);
			3970: out = 24'(-47924);
			3971: out = 24'(-28440);
			3972: out = 24'(5200);
			3973: out = 24'(17284);
			3974: out = 24'(-7676);
			3975: out = 24'(-18632);
			3976: out = 24'(8640);
			3977: out = 24'(-3548);
			3978: out = 24'(-29488);
			3979: out = 24'(-19360);
			3980: out = 24'(-9000);
			3981: out = 24'(13928);
			3982: out = 24'(32176);
			3983: out = 24'(20148);
			3984: out = 24'(-19168);
			3985: out = 24'(-39464);
			3986: out = 24'(-39468);
			3987: out = 24'(-30088);
			3988: out = 24'(6864);
			3989: out = 24'(47348);
			3990: out = 24'(31172);
			3991: out = 24'(12188);
			3992: out = 24'(8380);
			3993: out = 24'(-13516);
			3994: out = 24'(-28752);
			3995: out = 24'(-51328);
			3996: out = 24'(-23068);
			3997: out = 24'(19936);
			3998: out = 24'(13552);
			3999: out = 24'(6644);
			4000: out = 24'(4760);
			4001: out = 24'(43200);
			4002: out = 24'(54180);
			4003: out = 24'(26044);
			4004: out = 24'(-23688);
			4005: out = 24'(-32476);
			4006: out = 24'(-29644);
			4007: out = 24'(-27864);
			4008: out = 24'(-2500);
			4009: out = 24'(-8628);
			4010: out = 24'(-1228);
			4011: out = 24'(20928);
			4012: out = 24'(24204);
			4013: out = 24'(-13864);
			4014: out = 24'(15020);
			4015: out = 24'(33712);
			4016: out = 24'(8976);
			4017: out = 24'(-26236);
			4018: out = 24'(-39192);
			4019: out = 24'(-10772);
			4020: out = 24'(45272);
			4021: out = 24'(64720);
			4022: out = 24'(3244);
			4023: out = 24'(-44732);
			4024: out = 24'(-27896);
			4025: out = 24'(5564);
			4026: out = 24'(36084);
			4027: out = 24'(13328);
			4028: out = 24'(-25984);
			4029: out = 24'(560);
			4030: out = 24'(46684);
			4031: out = 24'(28824);
			4032: out = 24'(-16320);
			4033: out = 24'(-37816);
			4034: out = 24'(17220);
			4035: out = 24'(10304);
			4036: out = 24'(-16000);
			4037: out = 24'(15608);
			4038: out = 24'(43516);
			4039: out = 24'(-3112);
			4040: out = 24'(-58852);
			4041: out = 24'(-22420);
			4042: out = 24'(16868);
			4043: out = 24'(16612);
			4044: out = 24'(9252);
			4045: out = 24'(-4692);
			4046: out = 24'(-41552);
			4047: out = 24'(-40904);
			4048: out = 24'(6128);
			4049: out = 24'(39048);
			4050: out = 24'(58380);
			4051: out = 24'(34916);
			4052: out = 24'(-24812);
			4053: out = 24'(-34036);
			4054: out = 24'(-9684);
			4055: out = 24'(17308);
			4056: out = 24'(44212);
			4057: out = 24'(29384);
			4058: out = 24'(-10476);
			4059: out = 24'(2796);
			4060: out = 24'(18240);
			4061: out = 24'(6736);
			4062: out = 24'(18616);
			4063: out = 24'(23736);
			4064: out = 24'(-5592);
			4065: out = 24'(11216);
			4066: out = 24'(344);
			4067: out = 24'(-15684);
			4068: out = 24'(17188);
			4069: out = 24'(51956);
			4070: out = 24'(21360);
			4071: out = 24'(-15116);
			4072: out = 24'(8792);
			4073: out = 24'(22208);
			4074: out = 24'(36172);
			4075: out = 24'(32084);
			4076: out = 24'(28200);
			4077: out = 24'(7972);
			4078: out = 24'(-24128);
			4079: out = 24'(-37344);
			4080: out = 24'(-736);
			4081: out = 24'(39216);
			4082: out = 24'(-4);
			4083: out = 24'(-37540);
			4084: out = 24'(-18728);
			4085: out = 24'(-8040);
			4086: out = 24'(21888);
			4087: out = 24'(9420);
			4088: out = 24'(-10740);
			4089: out = 24'(-4368);
			4090: out = 24'(-1432);
			4091: out = 24'(27424);
			4092: out = 24'(2516);
			4093: out = 24'(14200);
			4094: out = 24'(22336);
			4095: out = 24'(32000);
			4096: out = 24'(18204);
			4097: out = 24'(-21244);
			4098: out = 24'(-1024);
			4099: out = 24'(25196);
			4100: out = 24'(18368);
			4101: out = 24'(-12872);
			4102: out = 24'(-7368);
			4103: out = 24'(29816);
			4104: out = 24'(29444);
			4105: out = 24'(-18456);
			4106: out = 24'(-15720);
			4107: out = 24'(1552);
			4108: out = 24'(-22144);
			4109: out = 24'(-10840);
			4110: out = 24'(25700);
			4111: out = 24'(12420);
			4112: out = 24'(-14888);
			4113: out = 24'(-8192);
			4114: out = 24'(-9252);
			4115: out = 24'(-17700);
			4116: out = 24'(-16264);
			4117: out = 24'(22944);
			4118: out = 24'(17992);
			4119: out = 24'(10140);
			4120: out = 24'(35516);
			4121: out = 24'(25820);
			4122: out = 24'(-6724);
			4123: out = 24'(-42424);
			4124: out = 24'(-28340);
			4125: out = 24'(9076);
			4126: out = 24'(45716);
			4127: out = 24'(50224);
			4128: out = 24'(21868);
			4129: out = 24'(11736);
			4130: out = 24'(-2340);
			4131: out = 24'(-3476);
			4132: out = 24'(1676);
			4133: out = 24'(27052);
			4134: out = 24'(46032);
			4135: out = 24'(20236);
			4136: out = 24'(-712);
			4137: out = 24'(7408);
			4138: out = 24'(-3412);
			4139: out = 24'(-23216);
			4140: out = 24'(-32404);
			4141: out = 24'(-19932);
			4142: out = 24'(4332);
			4143: out = 24'(39568);
			4144: out = 24'(11600);
			4145: out = 24'(-38084);
			4146: out = 24'(-59448);
			4147: out = 24'(-51968);
			4148: out = 24'(-30752);
			4149: out = 24'(38300);
			4150: out = 24'(83252);
			4151: out = 24'(-11788);
			4152: out = 24'(-50036);
			4153: out = 24'(-5836);
			4154: out = 24'(40424);
			4155: out = 24'(48336);
			4156: out = 24'(6572);
			4157: out = 24'(-14384);
			4158: out = 24'(3096);
			4159: out = 24'(12852);
			4160: out = 24'(12252);
			4161: out = 24'(-31472);
			4162: out = 24'(-34556);
			4163: out = 24'(11824);
			4164: out = 24'(7656);
			4165: out = 24'(12508);
			4166: out = 24'(12172);
			4167: out = 24'(2200);
			4168: out = 24'(-712);
			4169: out = 24'(5744);
			4170: out = 24'(4624);
			4171: out = 24'(-26188);
			4172: out = 24'(-1792);
			4173: out = 24'(43856);
			4174: out = 24'(17352);
			4175: out = 24'(-37408);
			4176: out = 24'(-44588);
			4177: out = 24'(5576);
			4178: out = 24'(53876);
			4179: out = 24'(9584);
			4180: out = 24'(-39064);
			4181: out = 24'(-28244);
			4182: out = 24'(9180);
			4183: out = 24'(14032);
			4184: out = 24'(-972);
			4185: out = 24'(-18072);
			4186: out = 24'(976);
			4187: out = 24'(35952);
			4188: out = 24'(37884);
			4189: out = 24'(33320);
			4190: out = 24'(-15168);
			4191: out = 24'(-28324);
			4192: out = 24'(-30508);
			4193: out = 24'(-11096);
			4194: out = 24'(31976);
			4195: out = 24'(37816);
			4196: out = 24'(-19828);
			4197: out = 24'(-37944);
			4198: out = 24'(-29696);
			4199: out = 24'(-28820);
			4200: out = 24'(11544);
			4201: out = 24'(14812);
			4202: out = 24'(-13888);
			4203: out = 24'(-12056);
			4204: out = 24'(21692);
			4205: out = 24'(-8204);
			4206: out = 24'(-32908);
			4207: out = 24'(-1376);
			4208: out = 24'(17500);
			4209: out = 24'(24232);
			4210: out = 24'(-18708);
			4211: out = 24'(-6576);
			4212: out = 24'(28524);
			4213: out = 24'(29540);
			4214: out = 24'(9804);
			4215: out = 24'(-24528);
			4216: out = 24'(-60892);
			4217: out = 24'(-60192);
			4218: out = 24'(-18936);
			4219: out = 24'(2912);
			4220: out = 24'(23924);
			4221: out = 24'(50252);
			4222: out = 24'(4820);
			4223: out = 24'(-40492);
			4224: out = 24'(-21376);
			4225: out = 24'(-7632);
			4226: out = 24'(21120);
			4227: out = 24'(35696);
			4228: out = 24'(4632);
			4229: out = 24'(-43644);
			4230: out = 24'(-45228);
			4231: out = 24'(18132);
			4232: out = 24'(34268);
			4233: out = 24'(30240);
			4234: out = 24'(6948);
			4235: out = 24'(-8392);
			4236: out = 24'(-3728);
			4237: out = 24'(-9380);
			4238: out = 24'(22168);
			4239: out = 24'(35284);
			4240: out = 24'(21904);
			4241: out = 24'(-17160);
			4242: out = 24'(-37364);
			4243: out = 24'(-32040);
			4244: out = 24'(5268);
			4245: out = 24'(3368);
			4246: out = 24'(-35748);
			4247: out = 24'(2008);
			4248: out = 24'(13816);
			4249: out = 24'(-15692);
			4250: out = 24'(-28000);
			4251: out = 24'(-13448);
			4252: out = 24'(23696);
			4253: out = 24'(31004);
			4254: out = 24'(16700);
			4255: out = 24'(-26236);
			4256: out = 24'(-53132);
			4257: out = 24'(-40252);
			4258: out = 24'(-17416);
			4259: out = 24'(12688);
			4260: out = 24'(-3776);
			4261: out = 24'(6732);
			4262: out = 24'(39260);
			4263: out = 24'(15800);
			4264: out = 24'(-2832);
			4265: out = 24'(-1688);
			4266: out = 24'(-12480);
			4267: out = 24'(-22552);
			4268: out = 24'(-20072);
			4269: out = 24'(-16224);
			4270: out = 24'(-11760);
			4271: out = 24'(-3252);
			4272: out = 24'(-14308);
			4273: out = 24'(6344);
			4274: out = 24'(3224);
			4275: out = 24'(-33288);
			4276: out = 24'(-15284);
			4277: out = 24'(36228);
			4278: out = 24'(25408);
			4279: out = 24'(-42568);
			4280: out = 24'(-58860);
			4281: out = 24'(-19756);
			4282: out = 24'(17140);
			4283: out = 24'(68344);
			4284: out = 24'(39000);
			4285: out = 24'(4904);
			4286: out = 24'(-1024);
			4287: out = 24'(-2964);
			4288: out = 24'(10844);
			4289: out = 24'(-12360);
			4290: out = 24'(-28896);
			4291: out = 24'(616);
			4292: out = 24'(37596);
			4293: out = 24'(2140);
			4294: out = 24'(-29268);
			4295: out = 24'(-16604);
			4296: out = 24'(-952);
			4297: out = 24'(21416);
			4298: out = 24'(14304);
			4299: out = 24'(-15664);
			4300: out = 24'(-10084);
			4301: out = 24'(3372);
			4302: out = 24'(3656);
			4303: out = 24'(-3420);
			4304: out = 24'(1780);
			4305: out = 24'(17372);
			4306: out = 24'(-5276);
			4307: out = 24'(-27440);
			4308: out = 24'(-23420);
			4309: out = 24'(-5140);
			4310: out = 24'(-22356);
			4311: out = 24'(-45508);
			4312: out = 24'(-45092);
			4313: out = 24'(-17292);
			4314: out = 24'(5864);
			4315: out = 24'(20504);
			4316: out = 24'(20860);
			4317: out = 24'(7384);
			4318: out = 24'(3216);
			4319: out = 24'(-8192);
			4320: out = 24'(-24392);
			4321: out = 24'(-4508);
			4322: out = 24'(17864);
			4323: out = 24'(17800);
			4324: out = 24'(3712);
			4325: out = 24'(19488);
			4326: out = 24'(44864);
			4327: out = 24'(8548);
			4328: out = 24'(-51988);
			4329: out = 24'(-60604);
			4330: out = 24'(-42872);
			4331: out = 24'(-19864);
			4332: out = 24'(25592);
			4333: out = 24'(4832);
			4334: out = 24'(-36960);
			4335: out = 24'(-24496);
			4336: out = 24'(-4936);
			4337: out = 24'(29332);
			4338: out = 24'(54660);
			4339: out = 24'(35840);
			4340: out = 24'(-14432);
			4341: out = 24'(-40020);
			4342: out = 24'(-21952);
			4343: out = 24'(4324);
			4344: out = 24'(16400);
			4345: out = 24'(2328);
			4346: out = 24'(-8756);
			4347: out = 24'(1212);
			4348: out = 24'(-14536);
			4349: out = 24'(-45192);
			4350: out = 24'(6356);
			4351: out = 24'(27912);
			4352: out = 24'(2740);
			4353: out = 24'(21688);
			4354: out = 24'(27768);
			4355: out = 24'(-25524);
			4356: out = 24'(-40320);
			4357: out = 24'(-19336);
			4358: out = 24'(12700);
			4359: out = 24'(22540);
			4360: out = 24'(36876);
			4361: out = 24'(22336);
			4362: out = 24'(12592);
			4363: out = 24'(20992);
			4364: out = 24'(32324);
			4365: out = 24'(30888);
			4366: out = 24'(-10332);
			4367: out = 24'(-45660);
			4368: out = 24'(-36292);
			4369: out = 24'(10308);
			4370: out = 24'(-11768);
			4371: out = 24'(-45080);
			4372: out = 24'(-26352);
			4373: out = 24'(-2052);
			4374: out = 24'(29388);
			4375: out = 24'(53712);
			4376: out = 24'(37620);
			4377: out = 24'(-3660);
			4378: out = 24'(-38420);
			4379: out = 24'(-23552);
			4380: out = 24'(11300);
			4381: out = 24'(48604);
			4382: out = 24'(23384);
			4383: out = 24'(4452);
			4384: out = 24'(29496);
			4385: out = 24'(40836);
			4386: out = 24'(-676);
			4387: out = 24'(-30892);
			4388: out = 24'(-26660);
			4389: out = 24'(4492);
			4390: out = 24'(20812);
			4391: out = 24'(8736);
			4392: out = 24'(6852);
			4393: out = 24'(10864);
			4394: out = 24'(21788);
			4395: out = 24'(-932);
			4396: out = 24'(-5676);
			4397: out = 24'(-460);
			4398: out = 24'(4864);
			4399: out = 24'(21964);
			4400: out = 24'(29284);
			4401: out = 24'(-12124);
			4402: out = 24'(-50048);
			4403: out = 24'(-47104);
			4404: out = 24'(-39344);
			4405: out = 24'(-4244);
			4406: out = 24'(19608);
			4407: out = 24'(4564);
			4408: out = 24'(-15168);
			4409: out = 24'(22868);
			4410: out = 24'(30236);
			4411: out = 24'(2624);
			4412: out = 24'(-12252);
			4413: out = 24'(-10372);
			4414: out = 24'(11192);
			4415: out = 24'(19992);
			4416: out = 24'(25108);
			4417: out = 24'(10592);
			4418: out = 24'(-17808);
			4419: out = 24'(-26628);
			4420: out = 24'(5448);
			4421: out = 24'(17760);
			4422: out = 24'(5036);
			4423: out = 24'(11484);
			4424: out = 24'(14688);
			4425: out = 24'(-7872);
			4426: out = 24'(-21312);
			4427: out = 24'(-14324);
			4428: out = 24'(11080);
			4429: out = 24'(12008);
			4430: out = 24'(2356);
			4431: out = 24'(5516);
			4432: out = 24'(128);
			4433: out = 24'(-3584);
			4434: out = 24'(-15320);
			4435: out = 24'(10100);
			4436: out = 24'(27900);
			4437: out = 24'(6840);
			4438: out = 24'(2396);
			4439: out = 24'(-2580);
			4440: out = 24'(16488);
			4441: out = 24'(17092);
			4442: out = 24'(2140);
			4443: out = 24'(-9552);
			4444: out = 24'(136);
			4445: out = 24'(5104);
			4446: out = 24'(-8076);
			4447: out = 24'(-1048);
			4448: out = 24'(-3500);
			4449: out = 24'(-4388);
			4450: out = 24'(-17984);
			4451: out = 24'(-3116);
			4452: out = 24'(35956);
			4453: out = 24'(17796);
			4454: out = 24'(-13904);
			4455: out = 24'(-9772);
			4456: out = 24'(-2876);
			4457: out = 24'(38336);
			4458: out = 24'(53360);
			4459: out = 24'(-8360);
			4460: out = 24'(-33348);
			4461: out = 24'(-35412);
			4462: out = 24'(9728);
			4463: out = 24'(19888);
			4464: out = 24'(-568);
			4465: out = 24'(22504);
			4466: out = 24'(53032);
			4467: out = 24'(39572);
			4468: out = 24'(-23728);
			4469: out = 24'(-62832);
			4470: out = 24'(-38704);
			4471: out = 24'(816);
			4472: out = 24'(34024);
			4473: out = 24'(47348);
			4474: out = 24'(19096);
			4475: out = 24'(-14660);
			4476: out = 24'(-680);
			4477: out = 24'(13444);
			4478: out = 24'(2588);
			4479: out = 24'(-6456);
			4480: out = 24'(-20480);
			4481: out = 24'(-3984);
			4482: out = 24'(14592);
			4483: out = 24'(20440);
			4484: out = 24'(5616);
			4485: out = 24'(-3356);
			4486: out = 24'(-33496);
			4487: out = 24'(-36680);
			4488: out = 24'(-36260);
			4489: out = 24'(7304);
			4490: out = 24'(46524);
			4491: out = 24'(6836);
			4492: out = 24'(-10212);
			4493: out = 24'(13428);
			4494: out = 24'(33820);
			4495: out = 24'(-3928);
			4496: out = 24'(-35244);
			4497: out = 24'(-17316);
			4498: out = 24'(19628);
			4499: out = 24'(19468);
			4500: out = 24'(7072);
			4501: out = 24'(-2848);
			4502: out = 24'(3952);
			4503: out = 24'(-10240);
			4504: out = 24'(-34544);
			4505: out = 24'(-15512);
			4506: out = 24'(23400);
			4507: out = 24'(18908);
			4508: out = 24'(1348);
			4509: out = 24'(-19300);
			4510: out = 24'(-19124);
			4511: out = 24'(23372);
			4512: out = 24'(25804);
			4513: out = 24'(-9420);
			4514: out = 24'(-44296);
			4515: out = 24'(-13668);
			4516: out = 24'(40760);
			4517: out = 24'(62024);
			4518: out = 24'(31996);
			4519: out = 24'(15404);
			4520: out = 24'(2092);
			4521: out = 24'(-15148);
			4522: out = 24'(-33420);
			4523: out = 24'(-49032);
			4524: out = 24'(1108);
			4525: out = 24'(58440);
			4526: out = 24'(15648);
			4527: out = 24'(-30792);
			4528: out = 24'(5392);
			4529: out = 24'(24524);
			4530: out = 24'(13956);
			4531: out = 24'(-17380);
			4532: out = 24'(-14708);
			4533: out = 24'(-11916);
			4534: out = 24'(412);
			4535: out = 24'(-3080);
			4536: out = 24'(13672);
			4537: out = 24'(42400);
			4538: out = 24'(44996);
			4539: out = 24'(-7296);
			4540: out = 24'(-24004);
			4541: out = 24'(-19044);
			4542: out = 24'(-6384);
			4543: out = 24'(3768);
			4544: out = 24'(12896);
			4545: out = 24'(10556);
			4546: out = 24'(10364);
			4547: out = 24'(-16680);
			4548: out = 24'(-37816);
			4549: out = 24'(-4692);
			4550: out = 24'(-1156);
			4551: out = 24'(17368);
			4552: out = 24'(23508);
			4553: out = 24'(20020);
			4554: out = 24'(-14344);
			4555: out = 24'(-28252);
			4556: out = 24'(-25272);
			4557: out = 24'(7260);
			4558: out = 24'(21184);
			4559: out = 24'(5980);
			4560: out = 24'(2100);
			4561: out = 24'(-3348);
			4562: out = 24'(-53288);
			4563: out = 24'(-61984);
			4564: out = 24'(-5280);
			4565: out = 24'(32948);
			4566: out = 24'(39472);
			4567: out = 24'(18328);
			4568: out = 24'(-1368);
			4569: out = 24'(-28504);
			4570: out = 24'(1956);
			4571: out = 24'(22568);
			4572: out = 24'(47100);
			4573: out = 24'(48304);
			4574: out = 24'(-5636);
			4575: out = 24'(-22156);
			4576: out = 24'(-12488);
			4577: out = 24'(7568);
			4578: out = 24'(6408);
			4579: out = 24'(-43672);
			4580: out = 24'(-20524);
			4581: out = 24'(21044);
			4582: out = 24'(22312);
			4583: out = 24'(27756);
			4584: out = 24'(28776);
			4585: out = 24'(18784);
			4586: out = 24'(-21856);
			4587: out = 24'(-54488);
			4588: out = 24'(-45732);
			4589: out = 24'(-4584);
			4590: out = 24'(-19340);
			4591: out = 24'(-18312);
			4592: out = 24'(36564);
			4593: out = 24'(26340);
			4594: out = 24'(-25740);
			4595: out = 24'(-19844);
			4596: out = 24'(-21308);
			4597: out = 24'(-4592);
			4598: out = 24'(18896);
			4599: out = 24'(29504);
			4600: out = 24'(-17360);
			4601: out = 24'(-39900);
			4602: out = 24'(-2352);
			4603: out = 24'(45408);
			4604: out = 24'(48224);
			4605: out = 24'(8968);
			4606: out = 24'(-10664);
			4607: out = 24'(5648);
			4608: out = 24'(9884);
			4609: out = 24'(-27160);
			4610: out = 24'(-38416);
			4611: out = 24'(-30332);
			4612: out = 24'(-9704);
			4613: out = 24'(11132);
			4614: out = 24'(13888);
			4615: out = 24'(-6660);
			4616: out = 24'(10376);
			4617: out = 24'(23820);
			4618: out = 24'(48);
			4619: out = 24'(-45708);
			4620: out = 24'(-51388);
			4621: out = 24'(-12160);
			4622: out = 24'(28156);
			4623: out = 24'(29200);
			4624: out = 24'(-15508);
			4625: out = 24'(-39200);
			4626: out = 24'(-39904);
			4627: out = 24'(10396);
			4628: out = 24'(58364);
			4629: out = 24'(22064);
			4630: out = 24'(-17252);
			4631: out = 24'(-17932);
			4632: out = 24'(-5896);
			4633: out = 24'(12188);
			4634: out = 24'(3088);
			4635: out = 24'(-23832);
			4636: out = 24'(-13588);
			4637: out = 24'(11696);
			4638: out = 24'(15808);
			4639: out = 24'(-15504);
			4640: out = 24'(-52932);
			4641: out = 24'(-41380);
			4642: out = 24'(26032);
			4643: out = 24'(42488);
			4644: out = 24'(28524);
			4645: out = 24'(13660);
			4646: out = 24'(-1312);
			4647: out = 24'(-6384);
			4648: out = 24'(-35764);
			4649: out = 24'(-14140);
			4650: out = 24'(31600);
			4651: out = 24'(-10448);
			4652: out = 24'(-36796);
			4653: out = 24'(8488);
			4654: out = 24'(1936);
			4655: out = 24'(-17612);
			4656: out = 24'(-24712);
			4657: out = 24'(-352);
			4658: out = 24'(7788);
			4659: out = 24'(-16460);
			4660: out = 24'(7136);
			4661: out = 24'(34904);
			4662: out = 24'(32036);
			4663: out = 24'(6684);
			4664: out = 24'(-14584);
			4665: out = 24'(-22136);
			4666: out = 24'(-26028);
			4667: out = 24'(-6408);
			4668: out = 24'(5620);
			4669: out = 24'(-6100);
			4670: out = 24'(-28556);
			4671: out = 24'(-24136);
			4672: out = 24'(41596);
			4673: out = 24'(43076);
			4674: out = 24'(-33648);
			4675: out = 24'(-45112);
			4676: out = 24'(-20704);
			4677: out = 24'(-12448);
			4678: out = 24'(324);
			4679: out = 24'(18588);
			4680: out = 24'(-6996);
			4681: out = 24'(-30392);
			4682: out = 24'(-608);
			4683: out = 24'(39280);
			4684: out = 24'(42880);
			4685: out = 24'(6060);
			4686: out = 24'(-27108);
			4687: out = 24'(2308);
			4688: out = 24'(26832);
			4689: out = 24'(-16292);
			4690: out = 24'(-56016);
			4691: out = 24'(-43276);
			4692: out = 24'(-2620);
			4693: out = 24'(21456);
			4694: out = 24'(5416);
			4695: out = 24'(-16040);
			4696: out = 24'(13032);
			4697: out = 24'(34224);
			4698: out = 24'(26440);
			4699: out = 24'(-7900);
			4700: out = 24'(-46492);
			4701: out = 24'(-35860);
			4702: out = 24'(-22436);
			4703: out = 24'(27360);
			4704: out = 24'(50532);
			4705: out = 24'(-2212);
			4706: out = 24'(-23072);
			4707: out = 24'(9072);
			4708: out = 24'(33036);
			4709: out = 24'(25560);
			4710: out = 24'(-21312);
			4711: out = 24'(-37876);
			4712: out = 24'(-25136);
			4713: out = 24'(-10932);
			4714: out = 24'(31512);
			4715: out = 24'(13932);
			4716: out = 24'(-33672);
			4717: out = 24'(-27036);
			4718: out = 24'(2980);
			4719: out = 24'(21232);
			4720: out = 24'(9772);
			4721: out = 24'(-18408);
			4722: out = 24'(-29308);
			4723: out = 24'(-37116);
			4724: out = 24'(1732);
			4725: out = 24'(53692);
			4726: out = 24'(25056);
			4727: out = 24'(-31620);
			4728: out = 24'(-37392);
			4729: out = 24'(-33908);
			4730: out = 24'(-10156);
			4731: out = 24'(17156);
			4732: out = 24'(-1432);
			4733: out = 24'(3736);
			4734: out = 24'(32116);
			4735: out = 24'(15720);
			4736: out = 24'(-2960);
			4737: out = 24'(-9556);
			4738: out = 24'(-15268);
			4739: out = 24'(16696);
			4740: out = 24'(25192);
			4741: out = 24'(21472);
			4742: out = 24'(-13308);
			4743: out = 24'(-10396);
			4744: out = 24'(27284);
			4745: out = 24'(35840);
			4746: out = 24'(-15672);
			4747: out = 24'(-34968);
			4748: out = 24'(-3564);
			4749: out = 24'(16380);
			4750: out = 24'(5556);
			4751: out = 24'(-10976);
			4752: out = 24'(19340);
			4753: out = 24'(49792);
			4754: out = 24'(28456);
			4755: out = 24'(-10900);
			4756: out = 24'(-26224);
			4757: out = 24'(-10224);
			4758: out = 24'(-1476);
			4759: out = 24'(-23280);
			4760: out = 24'(-16024);
			4761: out = 24'(14472);
			4762: out = 24'(18568);
			4763: out = 24'(6500);
			4764: out = 24'(4860);
			4765: out = 24'(2756);
			4766: out = 24'(4880);
			4767: out = 24'(-10856);
			4768: out = 24'(12100);
			4769: out = 24'(7336);
			4770: out = 24'(16876);
			4771: out = 24'(28712);
			4772: out = 24'(22732);
			4773: out = 24'(-21472);
			4774: out = 24'(-38848);
			4775: out = 24'(-23052);
			4776: out = 24'(-3680);
			4777: out = 24'(-8944);
			4778: out = 24'(-17700);
			4779: out = 24'(2012);
			4780: out = 24'(-1236);
			4781: out = 24'(-6168);
			4782: out = 24'(-264);
			4783: out = 24'(428);
			4784: out = 24'(7976);
			4785: out = 24'(52132);
			4786: out = 24'(69560);
			4787: out = 24'(3668);
			4788: out = 24'(-61220);
			4789: out = 24'(-53556);
			4790: out = 24'(-20044);
			4791: out = 24'(24692);
			4792: out = 24'(48000);
			4793: out = 24'(-14200);
			4794: out = 24'(-30380);
			4795: out = 24'(16548);
			4796: out = 24'(49572);
			4797: out = 24'(14748);
			4798: out = 24'(-36424);
			4799: out = 24'(-31380);
			4800: out = 24'(-9516);
			4801: out = 24'(31520);
			4802: out = 24'(45708);
			4803: out = 24'(-2308);
			4804: out = 24'(-33308);
			4805: out = 24'(3796);
			4806: out = 24'(10708);
			4807: out = 24'(18292);
			4808: out = 24'(19544);
			4809: out = 24'(11396);
			4810: out = 24'(-14804);
			4811: out = 24'(-37952);
			4812: out = 24'(-2032);
			4813: out = 24'(37028);
			4814: out = 24'(27224);
			4815: out = 24'(-20452);
			4816: out = 24'(-38248);
			4817: out = 24'(-26068);
			4818: out = 24'(26328);
			4819: out = 24'(63072);
			4820: out = 24'(19968);
			4821: out = 24'(-12604);
			4822: out = 24'(-8000);
			4823: out = 24'(24972);
			4824: out = 24'(7088);
			4825: out = 24'(-6864);
			4826: out = 24'(10136);
			4827: out = 24'(14372);
			4828: out = 24'(11748);
			4829: out = 24'(3452);
			4830: out = 24'(-2848);
			4831: out = 24'(-19184);
			4832: out = 24'(-30356);
			4833: out = 24'(-20088);
			4834: out = 24'(19420);
			4835: out = 24'(40388);
			4836: out = 24'(23716);
			4837: out = 24'(-17120);
			4838: out = 24'(-7348);
			4839: out = 24'(9100);
			4840: out = 24'(10536);
			4841: out = 24'(38400);
			4842: out = 24'(57016);
			4843: out = 24'(12848);
			4844: out = 24'(-45580);
			4845: out = 24'(-36176);
			4846: out = 24'(15124);
			4847: out = 24'(44248);
			4848: out = 24'(48);
			4849: out = 24'(-32580);
			4850: out = 24'(-10356);
			4851: out = 24'(10612);
			4852: out = 24'(18692);
			4853: out = 24'(-16512);
			4854: out = 24'(-43296);
			4855: out = 24'(-14184);
			4856: out = 24'(18368);
			4857: out = 24'(34412);
			4858: out = 24'(31612);
			4859: out = 24'(2280);
			4860: out = 24'(-3036);
			4861: out = 24'(-8472);
			4862: out = 24'(9676);
			4863: out = 24'(18656);
			4864: out = 24'(28816);
			4865: out = 24'(33656);
			4866: out = 24'(4252);
			4867: out = 24'(-52720);
			4868: out = 24'(-60384);
			4869: out = 24'(-14600);
			4870: out = 24'(5064);
			4871: out = 24'(2072);
			4872: out = 24'(12104);
			4873: out = 24'(31332);
			4874: out = 24'(7012);
			4875: out = 24'(-25728);
			4876: out = 24'(-3316);
			4877: out = 24'(40616);
			4878: out = 24'(41896);
			4879: out = 24'(4044);
			4880: out = 24'(-23140);
			4881: out = 24'(-23008);
			4882: out = 24'(-18368);
			4883: out = 24'(-13172);
			4884: out = 24'(-8720);
			4885: out = 24'(-156);
			4886: out = 24'(33968);
			4887: out = 24'(8132);
			4888: out = 24'(7936);
			4889: out = 24'(1668);
			4890: out = 24'(-8884);
			4891: out = 24'(23220);
			4892: out = 24'(30168);
			4893: out = 24'(13444);
			4894: out = 24'(-29288);
			4895: out = 24'(-33984);
			4896: out = 24'(3496);
			4897: out = 24'(22364);
			4898: out = 24'(10300);
			4899: out = 24'(-13664);
			4900: out = 24'(-32480);
			4901: out = 24'(824);
			4902: out = 24'(31872);
			4903: out = 24'(21152);
			4904: out = 24'(-16448);
			4905: out = 24'(-30928);
			4906: out = 24'(-9020);
			4907: out = 24'(19768);
			4908: out = 24'(46140);
			4909: out = 24'(14384);
			4910: out = 24'(-33332);
			4911: out = 24'(-45736);
			4912: out = 24'(-16928);
			4913: out = 24'(31892);
			4914: out = 24'(54320);
			4915: out = 24'(19960);
			4916: out = 24'(-25236);
			4917: out = 24'(-24864);
			4918: out = 24'(-16052);
			4919: out = 24'(10312);
			4920: out = 24'(21624);
			4921: out = 24'(-14844);
			4922: out = 24'(-47088);
			4923: out = 24'(-6988);
			4924: out = 24'(42300);
			4925: out = 24'(14304);
			4926: out = 24'(-20904);
			4927: out = 24'(-24624);
			4928: out = 24'(-2316);
			4929: out = 24'(40972);
			4930: out = 24'(40500);
			4931: out = 24'(25632);
			4932: out = 24'(-224);
			4933: out = 24'(-27460);
			4934: out = 24'(-23656);
			4935: out = 24'(-14084);
			4936: out = 24'(14980);
			4937: out = 24'(27948);
			4938: out = 24'(-14572);
			4939: out = 24'(-44292);
			4940: out = 24'(-28164);
			4941: out = 24'(-2112);
			4942: out = 24'(41448);
			4943: out = 24'(44072);
			4944: out = 24'(6228);
			4945: out = 24'(-38044);
			4946: out = 24'(-48012);
			4947: out = 24'(-32968);
			4948: out = 24'(-9912);
			4949: out = 24'(18280);
			4950: out = 24'(30724);
			4951: out = 24'(11108);
			4952: out = 24'(-20096);
			4953: out = 24'(-4360);
			4954: out = 24'(7452);
			4955: out = 24'(15832);
			4956: out = 24'(13184);
			4957: out = 24'(-4268);
			4958: out = 24'(-6864);
			4959: out = 24'(5440);
			4960: out = 24'(31332);
			4961: out = 24'(24896);
			4962: out = 24'(-11204);
			4963: out = 24'(-39384);
			4964: out = 24'(-11104);
			4965: out = 24'(-9968);
			4966: out = 24'(18584);
			4967: out = 24'(28068);
			4968: out = 24'(6352);
			4969: out = 24'(-8760);
			4970: out = 24'(4832);
			4971: out = 24'(2868);
			4972: out = 24'(-21516);
			4973: out = 24'(-26924);
			4974: out = 24'(5884);
			4975: out = 24'(7480);
			4976: out = 24'(-12068);
			4977: out = 24'(-15876);
			4978: out = 24'(-17280);
			4979: out = 24'(-16780);
			4980: out = 24'(-19680);
			4981: out = 24'(-4916);
			4982: out = 24'(-7412);
			4983: out = 24'(-8508);
			4984: out = 24'(15576);
			4985: out = 24'(27204);
			4986: out = 24'(-11696);
			4987: out = 24'(-69440);
			4988: out = 24'(-35676);
			4989: out = 24'(14684);
			4990: out = 24'(36304);
			4991: out = 24'(46744);
			4992: out = 24'(16232);
			4993: out = 24'(-19132);
			4994: out = 24'(-10116);
			4995: out = 24'(-10996);
			4996: out = 24'(-5396);
			4997: out = 24'(-28508);
			4998: out = 24'(-30068);
			4999: out = 24'(31768);
			5000: out = 24'(46284);
			5001: out = 24'(8104);
			5002: out = 24'(-1428);
			5003: out = 24'(4964);
			5004: out = 24'(-6076);
			5005: out = 24'(-38752);
			5006: out = 24'(-23592);
			5007: out = 24'(6068);
			5008: out = 24'(31428);
			5009: out = 24'(19084);
			5010: out = 24'(-38400);
			5011: out = 24'(-25512);
			5012: out = 24'(21360);
			5013: out = 24'(26976);
			5014: out = 24'(5016);
			5015: out = 24'(-15940);
			5016: out = 24'(-11232);
			5017: out = 24'(19268);
			5018: out = 24'(31132);
			5019: out = 24'(12208);
			5020: out = 24'(-17416);
			5021: out = 24'(-14524);
			5022: out = 24'(-1728);
			5023: out = 24'(-8316);
			5024: out = 24'(-33856);
			5025: out = 24'(-43648);
			5026: out = 24'(-16508);
			5027: out = 24'(33684);
			5028: out = 24'(20108);
			5029: out = 24'(-24100);
			5030: out = 24'(-34288);
			5031: out = 24'(-1636);
			5032: out = 24'(33416);
			5033: out = 24'(39484);
			5034: out = 24'(26836);
			5035: out = 24'(-4068);
			5036: out = 24'(-6200);
			5037: out = 24'(-10172);
			5038: out = 24'(-9700);
			5039: out = 24'(-15732);
			5040: out = 24'(-15832);
			5041: out = 24'(6124);
			5042: out = 24'(13864);
			5043: out = 24'(22436);
			5044: out = 24'(5700);
			5045: out = 24'(720);
			5046: out = 24'(-5864);
			5047: out = 24'(1188);
			5048: out = 24'(7232);
			5049: out = 24'(2388);
			5050: out = 24'(13496);
			5051: out = 24'(15004);
			5052: out = 24'(-19736);
			5053: out = 24'(-43404);
			5054: out = 24'(-37052);
			5055: out = 24'(-33256);
			5056: out = 24'(-9152);
			5057: out = 24'(18736);
			5058: out = 24'(16964);
			5059: out = 24'(-23816);
			5060: out = 24'(-43624);
			5061: out = 24'(-30428);
			5062: out = 24'(-4864);
			5063: out = 24'(12168);
			5064: out = 24'(15168);
			5065: out = 24'(22380);
			5066: out = 24'(-436);
			5067: out = 24'(-6624);
			5068: out = 24'(3888);
			5069: out = 24'(5940);
			5070: out = 24'(-6488);
			5071: out = 24'(1996);
			5072: out = 24'(-3728);
			5073: out = 24'(2596);
			5074: out = 24'(-20584);
			5075: out = 24'(-40872);
			5076: out = 24'(-6444);
			5077: out = 24'(15888);
			5078: out = 24'(22256);
			5079: out = 24'(940);
			5080: out = 24'(-15840);
			5081: out = 24'(-22728);
			5082: out = 24'(-10888);
			5083: out = 24'(34224);
			5084: out = 24'(35156);
			5085: out = 24'(19868);
			5086: out = 24'(-20440);
			5087: out = 24'(-19624);
			5088: out = 24'(13312);
			5089: out = 24'(33124);
			5090: out = 24'(36468);
			5091: out = 24'(256);
			5092: out = 24'(-15464);
			5093: out = 24'(-7564);
			5094: out = 24'(12280);
			5095: out = 24'(-2940);
			5096: out = 24'(-10832);
			5097: out = 24'(13868);
			5098: out = 24'(14912);
			5099: out = 24'(-21824);
			5100: out = 24'(-24916);
			5101: out = 24'(-2092);
			5102: out = 24'(6312);
			5103: out = 24'(19168);
			5104: out = 24'(15132);
			5105: out = 24'(-16564);
			5106: out = 24'(-32512);
			5107: out = 24'(-29000);
			5108: out = 24'(-23904);
			5109: out = 24'(-2700);
			5110: out = 24'(52204);
			5111: out = 24'(34860);
			5112: out = 24'(-8508);
			5113: out = 24'(-4980);
			5114: out = 24'(25908);
			5115: out = 24'(47604);
			5116: out = 24'(18440);
			5117: out = 24'(-30620);
			5118: out = 24'(-24892);
			5119: out = 24'(2580);
			5120: out = 24'(-17672);
			5121: out = 24'(-29988);
			5122: out = 24'(-22440);
			5123: out = 24'(7424);
			5124: out = 24'(23728);
			5125: out = 24'(26904);
			5126: out = 24'(21848);
			5127: out = 24'(-9204);
			5128: out = 24'(-18404);
			5129: out = 24'(-26852);
			5130: out = 24'(14984);
			5131: out = 24'(17200);
			5132: out = 24'(-4048);
			5133: out = 24'(16036);
			5134: out = 24'(30116);
			5135: out = 24'(8884);
			5136: out = 24'(-31872);
			5137: out = 24'(-26924);
			5138: out = 24'(10548);
			5139: out = 24'(35756);
			5140: out = 24'(8060);
			5141: out = 24'(-13612);
			5142: out = 24'(-26624);
			5143: out = 24'(11412);
			5144: out = 24'(29236);
			5145: out = 24'(-116);
			5146: out = 24'(-4284);
			5147: out = 24'(-1964);
			5148: out = 24'(-5920);
			5149: out = 24'(9180);
			5150: out = 24'(20860);
			5151: out = 24'(-14032);
			5152: out = 24'(-8476);
			5153: out = 24'(16096);
			5154: out = 24'(31008);
			5155: out = 24'(21168);
			5156: out = 24'(-5792);
			5157: out = 24'(-3592);
			5158: out = 24'(2152);
			5159: out = 24'(-10560);
			5160: out = 24'(-25172);
			5161: out = 24'(-1096);
			5162: out = 24'(6788);
			5163: out = 24'(-19728);
			5164: out = 24'(-17564);
			5165: out = 24'(-13164);
			5166: out = 24'(26376);
			5167: out = 24'(53724);
			5168: out = 24'(13992);
			5169: out = 24'(-7536);
			5170: out = 24'(-4236);
			5171: out = 24'(-5388);
			5172: out = 24'(18236);
			5173: out = 24'(21808);
			5174: out = 24'(16800);
			5175: out = 24'(-9096);
			5176: out = 24'(-33140);
			5177: out = 24'(-32800);
			5178: out = 24'(-33644);
			5179: out = 24'(2120);
			5180: out = 24'(45348);
			5181: out = 24'(32636);
			5182: out = 24'(-13476);
			5183: out = 24'(-53568);
			5184: out = 24'(-34888);
			5185: out = 24'(8592);
			5186: out = 24'(45132);
			5187: out = 24'(59348);
			5188: out = 24'(-8184);
			5189: out = 24'(-46508);
			5190: out = 24'(-21912);
			5191: out = 24'(37552);
			5192: out = 24'(49104);
			5193: out = 24'(-15748);
			5194: out = 24'(-23928);
			5195: out = 24'(2872);
			5196: out = 24'(24332);
			5197: out = 24'(33460);
			5198: out = 24'(-14664);
			5199: out = 24'(-26768);
			5200: out = 24'(14500);
			5201: out = 24'(32692);
			5202: out = 24'(20872);
			5203: out = 24'(-4544);
			5204: out = 24'(-3704);
			5205: out = 24'(16384);
			5206: out = 24'(-8556);
			5207: out = 24'(-22136);
			5208: out = 24'(-308);
			5209: out = 24'(13156);
			5210: out = 24'(9164);
			5211: out = 24'(-23212);
			5212: out = 24'(-14820);
			5213: out = 24'(5972);
			5214: out = 24'(-4724);
			5215: out = 24'(-9068);
			5216: out = 24'(13216);
			5217: out = 24'(1336);
			5218: out = 24'(-2960);
			5219: out = 24'(5008);
			5220: out = 24'(-8024);
			5221: out = 24'(-19208);
			5222: out = 24'(-23428);
			5223: out = 24'(10364);
			5224: out = 24'(21768);
			5225: out = 24'(6768);
			5226: out = 24'(9632);
			5227: out = 24'(11272);
			5228: out = 24'(-26112);
			5229: out = 24'(-40936);
			5230: out = 24'(-13708);
			5231: out = 24'(26580);
			5232: out = 24'(52812);
			5233: out = 24'(10692);
			5234: out = 24'(-50292);
			5235: out = 24'(-29544);
			5236: out = 24'(22200);
			5237: out = 24'(49512);
			5238: out = 24'(43440);
			5239: out = 24'(5968);
			5240: out = 24'(-16984);
			5241: out = 24'(-812);
			5242: out = 24'(-3640);
			5243: out = 24'(-11252);
			5244: out = 24'(-18432);
			5245: out = 24'(-34940);
			5246: out = 24'(1548);
			5247: out = 24'(32608);
			5248: out = 24'(23840);
			5249: out = 24'(380);
			5250: out = 24'(340);
			5251: out = 24'(-16376);
			5252: out = 24'(-11292);
			5253: out = 24'(-8384);
			5254: out = 24'(-1480);
			5255: out = 24'(14536);
			5256: out = 24'(5768);
			5257: out = 24'(13860);
			5258: out = 24'(15740);
			5259: out = 24'(1120);
			5260: out = 24'(-4916);
			5261: out = 24'(-13796);
			5262: out = 24'(-7544);
			5263: out = 24'(14820);
			5264: out = 24'(-3180);
			5265: out = 24'(-1996);
			5266: out = 24'(28136);
			5267: out = 24'(33880);
			5268: out = 24'(-1348);
			5269: out = 24'(-35704);
			5270: out = 24'(-41456);
			5271: out = 24'(-2128);
			5272: out = 24'(11704);
			5273: out = 24'(11816);
			5274: out = 24'(14572);
			5275: out = 24'(12272);
			5276: out = 24'(-2672);
			5277: out = 24'(-9144);
			5278: out = 24'(-160);
			5279: out = 24'(1408);
			5280: out = 24'(-3368);
			5281: out = 24'(1296);
			5282: out = 24'(-2452);
			5283: out = 24'(-13492);
			5284: out = 24'(-28848);
			5285: out = 24'(-12048);
			5286: out = 24'(18560);
			5287: out = 24'(28420);
			5288: out = 24'(10556);
			5289: out = 24'(8044);
			5290: out = 24'(11712);
			5291: out = 24'(-3088);
			5292: out = 24'(-30032);
			5293: out = 24'(-62260);
			5294: out = 24'(-48228);
			5295: out = 24'(10280);
			5296: out = 24'(54808);
			5297: out = 24'(26204);
			5298: out = 24'(-10300);
			5299: out = 24'(-6452);
			5300: out = 24'(19524);
			5301: out = 24'(27628);
			5302: out = 24'(-14968);
			5303: out = 24'(-52336);
			5304: out = 24'(-36804);
			5305: out = 24'(29008);
			5306: out = 24'(45620);
			5307: out = 24'(-3336);
			5308: out = 24'(7604);
			5309: out = 24'(29460);
			5310: out = 24'(29952);
			5311: out = 24'(-16368);
			5312: out = 24'(-27280);
			5313: out = 24'(-6640);
			5314: out = 24'(30920);
			5315: out = 24'(36076);
			5316: out = 24'(2336);
			5317: out = 24'(-13900);
			5318: out = 24'(7136);
			5319: out = 24'(7348);
			5320: out = 24'(-9852);
			5321: out = 24'(3032);
			5322: out = 24'(6168);
			5323: out = 24'(-17308);
			5324: out = 24'(-49952);
			5325: out = 24'(-24408);
			5326: out = 24'(-15076);
			5327: out = 24'(-18132);
			5328: out = 24'(-7572);
			5329: out = 24'(19704);
			5330: out = 24'(-3468);
			5331: out = 24'(-20796);
			5332: out = 24'(8328);
			5333: out = 24'(35896);
			5334: out = 24'(29216);
			5335: out = 24'(2692);
			5336: out = 24'(-12208);
			5337: out = 24'(-14116);
			5338: out = 24'(-12048);
			5339: out = 24'(-10068);
			5340: out = 24'(-33956);
			5341: out = 24'(-50356);
			5342: out = 24'(-672);
			5343: out = 24'(30100);
			5344: out = 24'(29156);
			5345: out = 24'(30544);
			5346: out = 24'(28500);
			5347: out = 24'(12120);
			5348: out = 24'(-33236);
			5349: out = 24'(-43792);
			5350: out = 24'(-26760);
			5351: out = 24'(-7612);
			5352: out = 24'(26348);
			5353: out = 24'(18648);
			5354: out = 24'(-11340);
			5355: out = 24'(-25084);
			5356: out = 24'(-12520);
			5357: out = 24'(49564);
			5358: out = 24'(67856);
			5359: out = 24'(2864);
			5360: out = 24'(-62344);
			5361: out = 24'(-47492);
			5362: out = 24'(-21524);
			5363: out = 24'(17616);
			5364: out = 24'(14224);
			5365: out = 24'(-15916);
			5366: out = 24'(-6912);
			5367: out = 24'(33364);
			5368: out = 24'(42908);
			5369: out = 24'(14600);
			5370: out = 24'(-30288);
			5371: out = 24'(-43036);
			5372: out = 24'(-14332);
			5373: out = 24'(28448);
			5374: out = 24'(34372);
			5375: out = 24'(-9544);
			5376: out = 24'(-35612);
			5377: out = 24'(-7296);
			5378: out = 24'(16232);
			5379: out = 24'(2068);
			5380: out = 24'(4784);
			5381: out = 24'(4808);
			5382: out = 24'(-17372);
			5383: out = 24'(-25564);
			5384: out = 24'(9136);
			5385: out = 24'(24516);
			5386: out = 24'(26016);
			5387: out = 24'(-26740);
			5388: out = 24'(-22040);
			5389: out = 24'(44);
			5390: out = 24'(-1968);
			5391: out = 24'(30060);
			5392: out = 24'(35480);
			5393: out = 24'(-12820);
			5394: out = 24'(-52880);
			5395: out = 24'(-51280);
			5396: out = 24'(-34616);
			5397: out = 24'(8196);
			5398: out = 24'(30204);
			5399: out = 24'(8380);
			5400: out = 24'(-15872);
			5401: out = 24'(10348);
			5402: out = 24'(6128);
			5403: out = 24'(-1580);
			5404: out = 24'(15804);
			5405: out = 24'(6184);
			5406: out = 24'(10224);
			5407: out = 24'(21028);
			5408: out = 24'(22656);
			5409: out = 24'(4800);
			5410: out = 24'(-35992);
			5411: out = 24'(-36536);
			5412: out = 24'(-23740);
			5413: out = 24'(-7364);
			5414: out = 24'(23432);
			5415: out = 24'(5592);
			5416: out = 24'(-20908);
			5417: out = 24'(2428);
			5418: out = 24'(1764);
			5419: out = 24'(5248);
			5420: out = 24'(14612);
			5421: out = 24'(-5316);
			5422: out = 24'(-36688);
			5423: out = 24'(-35572);
			5424: out = 24'(-864);
			5425: out = 24'(11584);
			5426: out = 24'(22292);
			5427: out = 24'(-5128);
			5428: out = 24'(-19420);
			5429: out = 24'(32148);
			5430: out = 24'(52256);
			5431: out = 24'(18540);
			5432: out = 24'(-18560);
			5433: out = 24'(-9128);
			5434: out = 24'(13260);
			5435: out = 24'(9868);
			5436: out = 24'(-4336);
			5437: out = 24'(5632);
			5438: out = 24'(-7216);
			5439: out = 24'(-16528);
			5440: out = 24'(820);
			5441: out = 24'(-11928);
			5442: out = 24'(-38628);
			5443: out = 24'(-32072);
			5444: out = 24'(-25256);
			5445: out = 24'(1924);
			5446: out = 24'(39220);
			5447: out = 24'(46384);
			5448: out = 24'(-6328);
			5449: out = 24'(-28004);
			5450: out = 24'(-12328);
			5451: out = 24'(7332);
			5452: out = 24'(14732);
			5453: out = 24'(6720);
			5454: out = 24'(22972);
			5455: out = 24'(9104);
			5456: out = 24'(5744);
			5457: out = 24'(22784);
			5458: out = 24'(15988);
			5459: out = 24'(-35432);
			5460: out = 24'(-64252);
			5461: out = 24'(-46852);
			5462: out = 24'(-13788);
			5463: out = 24'(45544);
			5464: out = 24'(36664);
			5465: out = 24'(-20912);
			5466: out = 24'(-28704);
			5467: out = 24'(-8932);
			5468: out = 24'(10132);
			5469: out = 24'(15984);
			5470: out = 24'(29904);
			5471: out = 24'(14004);
			5472: out = 24'(-10252);
			5473: out = 24'(6360);
			5474: out = 24'(15720);
			5475: out = 24'(7216);
			5476: out = 24'(-12224);
			5477: out = 24'(-18912);
			5478: out = 24'(-3492);
			5479: out = 24'(652);
			5480: out = 24'(18776);
			5481: out = 24'(16640);
			5482: out = 24'(-12404);
			5483: out = 24'(-52264);
			5484: out = 24'(-38348);
			5485: out = 24'(-5116);
			5486: out = 24'(25420);
			5487: out = 24'(38588);
			5488: out = 24'(21432);
			5489: out = 24'(2140);
			5490: out = 24'(-9812);
			5491: out = 24'(-28624);
			5492: out = 24'(-24532);
			5493: out = 24'(572);
			5494: out = 24'(-6300);
			5495: out = 24'(-19600);
			5496: out = 24'(-16064);
			5497: out = 24'(26708);
			5498: out = 24'(26916);
			5499: out = 24'(8668);
			5500: out = 24'(21712);
			5501: out = 24'(28256);
			5502: out = 24'(35120);
			5503: out = 24'(2616);
			5504: out = 24'(-9112);
			5505: out = 24'(-10608);
			5506: out = 24'(-8688);
			5507: out = 24'(-14420);
			5508: out = 24'(-7988);
			5509: out = 24'(-23332);
			5510: out = 24'(-28180);
			5511: out = 24'(-7384);
			5512: out = 24'(-1808);
			5513: out = 24'(6964);
			5514: out = 24'(26208);
			5515: out = 24'(2252);
			5516: out = 24'(-4044);
			5517: out = 24'(20712);
			5518: out = 24'(27148);
			5519: out = 24'(1644);
			5520: out = 24'(-30932);
			5521: out = 24'(-39648);
			5522: out = 24'(-20800);
			5523: out = 24'(33568);
			5524: out = 24'(37024);
			5525: out = 24'(-13188);
			5526: out = 24'(-20816);
			5527: out = 24'(-5468);
			5528: out = 24'(24576);
			5529: out = 24'(25080);
			5530: out = 24'(6152);
			5531: out = 24'(-6704);
			5532: out = 24'(-9864);
			5533: out = 24'(988);
			5534: out = 24'(-1180);
			5535: out = 24'(22240);
			5536: out = 24'(36996);
			5537: out = 24'(22716);
			5538: out = 24'(-8688);
			5539: out = 24'(-30372);
			5540: out = 24'(-13400);
			5541: out = 24'(5088);
			5542: out = 24'(10876);
			5543: out = 24'(6224);
			5544: out = 24'(12916);
			5545: out = 24'(26488);
			5546: out = 24'(40072);
			5547: out = 24'(23212);
			5548: out = 24'(-4024);
			5549: out = 24'(-18924);
			5550: out = 24'(-22480);
			5551: out = 24'(-33332);
			5552: out = 24'(-8856);
			5553: out = 24'(27244);
			5554: out = 24'(7472);
			5555: out = 24'(-24988);
			5556: out = 24'(-26752);
			5557: out = 24'(-7736);
			5558: out = 24'(25140);
			5559: out = 24'(20384);
			5560: out = 24'(-4364);
			5561: out = 24'(-14084);
			5562: out = 24'(-20368);
			5563: out = 24'(-10060);
			5564: out = 24'(32408);
			5565: out = 24'(22784);
			5566: out = 24'(-41192);
			5567: out = 24'(-26368);
			5568: out = 24'(-5516);
			5569: out = 24'(8092);
			5570: out = 24'(38000);
			5571: out = 24'(17480);
			5572: out = 24'(3888);
			5573: out = 24'(7784);
			5574: out = 24'(11588);
			5575: out = 24'(15812);
			5576: out = 24'(-16388);
			5577: out = 24'(-23780);
			5578: out = 24'(11592);
			5579: out = 24'(5004);
			5580: out = 24'(-3256);
			5581: out = 24'(29052);
			5582: out = 24'(24020);
			5583: out = 24'(-22288);
			5584: out = 24'(-59108);
			5585: out = 24'(-44472);
			5586: out = 24'(6496);
			5587: out = 24'(36976);
			5588: out = 24'(43228);
			5589: out = 24'(20704);
			5590: out = 24'(-14116);
			5591: out = 24'(-16652);
			5592: out = 24'(-2148);
			5593: out = 24'(4592);
			5594: out = 24'(-244);
			5595: out = 24'(4920);
			5596: out = 24'(33776);
			5597: out = 24'(2552);
			5598: out = 24'(10840);
			5599: out = 24'(35576);
			5600: out = 24'(39796);
			5601: out = 24'(8016);
			5602: out = 24'(-26776);
			5603: out = 24'(-34360);
			5604: out = 24'(-5240);
			5605: out = 24'(6992);
			5606: out = 24'(-15820);
			5607: out = 24'(-2320);
			5608: out = 24'(29148);
			5609: out = 24'(11972);
			5610: out = 24'(-31424);
			5611: out = 24'(-39372);
			5612: out = 24'(-29824);
			5613: out = 24'(1760);
			5614: out = 24'(60516);
			5615: out = 24'(25984);
			5616: out = 24'(-26948);
			5617: out = 24'(-35480);
			5618: out = 24'(6324);
			5619: out = 24'(52716);
			5620: out = 24'(39736);
			5621: out = 24'(9492);
			5622: out = 24'(-7600);
			5623: out = 24'(5408);
			5624: out = 24'(-3244);
			5625: out = 24'(-19584);
			5626: out = 24'(-15052);
			5627: out = 24'(-3288);
			5628: out = 24'(11080);
			5629: out = 24'(9380);
			5630: out = 24'(21740);
			5631: out = 24'(-612);
			5632: out = 24'(5628);
			5633: out = 24'(-6988);
			5634: out = 24'(3904);
			5635: out = 24'(20244);
			5636: out = 24'(10172);
			5637: out = 24'(5052);
			5638: out = 24'(8800);
			5639: out = 24'(6224);
			5640: out = 24'(-17788);
			5641: out = 24'(-33876);
			5642: out = 24'(-27400);
			5643: out = 24'(-18688);
			5644: out = 24'(-14816);
			5645: out = 24'(7252);
			5646: out = 24'(14212);
			5647: out = 24'(-37788);
			5648: out = 24'(-68516);
			5649: out = 24'(-14968);
			5650: out = 24'(13696);
			5651: out = 24'(43744);
			5652: out = 24'(45296);
			5653: out = 24'(14684);
			5654: out = 24'(-34900);
			5655: out = 24'(-60308);
			5656: out = 24'(-17928);
			5657: out = 24'(34016);
			5658: out = 24'(59572);
			5659: out = 24'(26276);
			5660: out = 24'(-36760);
			5661: out = 24'(-40216);
			5662: out = 24'(-11284);
			5663: out = 24'(23000);
			5664: out = 24'(26012);
			5665: out = 24'(15248);
			5666: out = 24'(-144);
			5667: out = 24'(-9004);
			5668: out = 24'(7180);
			5669: out = 24'(1396);
			5670: out = 24'(6256);
			5671: out = 24'(9840);
			5672: out = 24'(-2376);
			5673: out = 24'(2852);
			5674: out = 24'(23036);
			5675: out = 24'(32004);
			5676: out = 24'(26668);
			5677: out = 24'(5456);
			5678: out = 24'(-11264);
			5679: out = 24'(-16960);
			5680: out = 24'(-11472);
			5681: out = 24'(-27800);
			5682: out = 24'(-15544);
			5683: out = 24'(10304);
			5684: out = 24'(-868);
			5685: out = 24'(-23384);
			5686: out = 24'(-40680);
			5687: out = 24'(-34608);
			5688: out = 24'(3340);
			5689: out = 24'(37268);
			5690: out = 24'(40304);
			5691: out = 24'(-16008);
			5692: out = 24'(-54280);
			5693: out = 24'(-26316);
			5694: out = 24'(18844);
			5695: out = 24'(51692);
			5696: out = 24'(33416);
			5697: out = 24'(-1544);
			5698: out = 24'(-25000);
			5699: out = 24'(-40128);
			5700: out = 24'(-3352);
			5701: out = 24'(35756);
			5702: out = 24'(18904);
			5703: out = 24'(9736);
			5704: out = 24'(8560);
			5705: out = 24'(-5624);
			5706: out = 24'(-29576);
			5707: out = 24'(-40604);
			5708: out = 24'(4420);
			5709: out = 24'(45492);
			5710: out = 24'(6564);
			5711: out = 24'(-19612);
			5712: out = 24'(7048);
			5713: out = 24'(12560);
			5714: out = 24'(9456);
			5715: out = 24'(-11960);
			5716: out = 24'(-18524);
			5717: out = 24'(-6160);
			5718: out = 24'(-6228);
			5719: out = 24'(11920);
			5720: out = 24'(6900);
			5721: out = 24'(5420);
			5722: out = 24'(22976);
			5723: out = 24'(27864);
			5724: out = 24'(172);
			5725: out = 24'(-35300);
			5726: out = 24'(-25588);
			5727: out = 24'(2732);
			5728: out = 24'(29016);
			5729: out = 24'(33396);
			5730: out = 24'(16872);
			5731: out = 24'(6004);
			5732: out = 24'(4284);
			5733: out = 24'(-10092);
			5734: out = 24'(-12392);
			5735: out = 24'(-22224);
			5736: out = 24'(-18648);
			5737: out = 24'(-13884);
			5738: out = 24'(11656);
			5739: out = 24'(11672);
			5740: out = 24'(-17560);
			5741: out = 24'(-36620);
			5742: out = 24'(-21712);
			5743: out = 24'(-2172);
			5744: out = 24'(22616);
			5745: out = 24'(30140);
			5746: out = 24'(1676);
			5747: out = 24'(-23844);
			5748: out = 24'(-35012);
			5749: out = 24'(-9500);
			5750: out = 24'(-3200);
			5751: out = 24'(-5872);
			5752: out = 24'(2692);
			5753: out = 24'(7712);
			5754: out = 24'(1648);
			5755: out = 24'(-3172);
			5756: out = 24'(-14272);
			5757: out = 24'(-10880);
			5758: out = 24'(-3044);
			5759: out = 24'(-6592);
			5760: out = 24'(17644);
			5761: out = 24'(28260);
			5762: out = 24'(-6224);
			5763: out = 24'(-45896);
			5764: out = 24'(-51524);
			5765: out = 24'(-3156);
			5766: out = 24'(49192);
			5767: out = 24'(25776);
			5768: out = 24'(-22064);
			5769: out = 24'(-18228);
			5770: out = 24'(-18600);
			5771: out = 24'(-18884);
			5772: out = 24'(5544);
			5773: out = 24'(4056);
			5774: out = 24'(7160);
			5775: out = 24'(32008);
			5776: out = 24'(2784);
			5777: out = 24'(-33168);
			5778: out = 24'(-40500);
			5779: out = 24'(-18200);
			5780: out = 24'(29284);
			5781: out = 24'(54848);
			5782: out = 24'(37156);
			5783: out = 24'(-14820);
			5784: out = 24'(-44696);
			5785: out = 24'(-47768);
			5786: out = 24'(-20436);
			5787: out = 24'(19248);
			5788: out = 24'(45840);
			5789: out = 24'(6580);
			5790: out = 24'(-30868);
			5791: out = 24'(-22580);
			5792: out = 24'(9472);
			5793: out = 24'(38316);
			5794: out = 24'(17872);
			5795: out = 24'(-45600);
			5796: out = 24'(-40572);
			5797: out = 24'(6920);
			5798: out = 24'(28336);
			5799: out = 24'(21420);
			5800: out = 24'(2308);
			5801: out = 24'(-464);
			5802: out = 24'(24576);
			5803: out = 24'(29292);
			5804: out = 24'(8356);
			5805: out = 24'(-16868);
			5806: out = 24'(-13952);
			5807: out = 24'(4768);
			5808: out = 24'(23160);
			5809: out = 24'(31400);
			5810: out = 24'(5696);
			5811: out = 24'(-23956);
			5812: out = 24'(-19040);
			5813: out = 24'(2664);
			5814: out = 24'(-7840);
			5815: out = 24'(-32040);
			5816: out = 24'(-24544);
			5817: out = 24'(9204);
			5818: out = 24'(-9116);
			5819: out = 24'(-10920);
			5820: out = 24'(19820);
			5821: out = 24'(20060);
			5822: out = 24'(-15836);
			5823: out = 24'(-12616);
			5824: out = 24'(-11556);
			5825: out = 24'(-6028);
			5826: out = 24'(19100);
			5827: out = 24'(26016);
			5828: out = 24'(11292);
			5829: out = 24'(-29032);
			5830: out = 24'(-6832);
			5831: out = 24'(30460);
			5832: out = 24'(37464);
			5833: out = 24'(-20780);
			5834: out = 24'(-42200);
			5835: out = 24'(-21864);
			5836: out = 24'(4504);
			5837: out = 24'(48868);
			5838: out = 24'(38252);
			5839: out = 24'(1960);
			5840: out = 24'(-1880);
			5841: out = 24'(-1960);
			5842: out = 24'(-15872);
			5843: out = 24'(-25240);
			5844: out = 24'(-4120);
			5845: out = 24'(2336);
			5846: out = 24'(-2768);
			5847: out = 24'(23644);
			5848: out = 24'(10276);
			5849: out = 24'(-3412);
			5850: out = 24'(-9936);
			5851: out = 24'(-19464);
			5852: out = 24'(3228);
			5853: out = 24'(21300);
			5854: out = 24'(18564);
			5855: out = 24'(-9444);
			5856: out = 24'(-4180);
			5857: out = 24'(32268);
			5858: out = 24'(26512);
			5859: out = 24'(-12600);
			5860: out = 24'(-23928);
			5861: out = 24'(-3888);
			5862: out = 24'(-16880);
			5863: out = 24'(-12748);
			5864: out = 24'(-10124);
			5865: out = 24'(-20308);
			5866: out = 24'(-13944);
			5867: out = 24'(21988);
			5868: out = 24'(31616);
			5869: out = 24'(-7080);
			5870: out = 24'(-9884);
			5871: out = 24'(30140);
			5872: out = 24'(41672);
			5873: out = 24'(-1600);
			5874: out = 24'(-29292);
			5875: out = 24'(-12952);
			5876: out = 24'(14028);
			5877: out = 24'(14032);
			5878: out = 24'(-3556);
			5879: out = 24'(-24460);
			5880: out = 24'(-19388);
			5881: out = 24'(3600);
			5882: out = 24'(9312);
			5883: out = 24'(-13316);
			5884: out = 24'(-15256);
			5885: out = 24'(8456);
			5886: out = 24'(33024);
			5887: out = 24'(18360);
			5888: out = 24'(-4620);
			5889: out = 24'(14344);
			5890: out = 24'(16300);
			5891: out = 24'(2152);
			5892: out = 24'(2900);
			5893: out = 24'(-9964);
			5894: out = 24'(-33332);
			5895: out = 24'(-33912);
			5896: out = 24'(-2796);
			5897: out = 24'(24328);
			5898: out = 24'(6056);
			5899: out = 24'(-2508);
			5900: out = 24'(34692);
			5901: out = 24'(31952);
			5902: out = 24'(-14168);
			5903: out = 24'(-32576);
			5904: out = 24'(-24716);
			5905: out = 24'(6300);
			5906: out = 24'(29732);
			5907: out = 24'(13324);
			5908: out = 24'(-24316);
			5909: out = 24'(-21496);
			5910: out = 24'(10344);
			5911: out = 24'(44544);
			5912: out = 24'(7824);
			5913: out = 24'(-21992);
			5914: out = 24'(-1128);
			5915: out = 24'(15736);
			5916: out = 24'(21040);
			5917: out = 24'(9652);
			5918: out = 24'(-2616);
			5919: out = 24'(-13832);
			5920: out = 24'(-22116);
			5921: out = 24'(-49368);
			5922: out = 24'(-33172);
			5923: out = 24'(20104);
			5924: out = 24'(42312);
			5925: out = 24'(20936);
			5926: out = 24'(12540);
			5927: out = 24'(-13192);
			5928: out = 24'(-2516);
			5929: out = 24'(16620);
			5930: out = 24'(11184);
			5931: out = 24'(31664);
			5932: out = 24'(18724);
			5933: out = 24'(-1272);
			5934: out = 24'(-1496);
			5935: out = 24'(4344);
			5936: out = 24'(3096);
			5937: out = 24'(-24956);
			5938: out = 24'(-40136);
			5939: out = 24'(-2148);
			5940: out = 24'(7880);
			5941: out = 24'(1304);
			5942: out = 24'(10492);
			5943: out = 24'(14480);
			5944: out = 24'(-6484);
			5945: out = 24'(-41572);
			5946: out = 24'(-48268);
			5947: out = 24'(9528);
			5948: out = 24'(56060);
			5949: out = 24'(43036);
			5950: out = 24'(-22088);
			5951: out = 24'(-18452);
			5952: out = 24'(4632);
			5953: out = 24'(25700);
			5954: out = 24'(17820);
			5955: out = 24'(1972);
			5956: out = 24'(-5492);
			5957: out = 24'(-412);
			5958: out = 24'(11512);
			5959: out = 24'(6752);
			5960: out = 24'(3800);
			5961: out = 24'(6088);
			5962: out = 24'(-488);
			5963: out = 24'(-25632);
			5964: out = 24'(-30048);
			5965: out = 24'(-31140);
			5966: out = 24'(-34000);
			5967: out = 24'(2812);
			5968: out = 24'(37680);
			5969: out = 24'(15696);
			5970: out = 24'(4840);
			5971: out = 24'(-3520);
			5972: out = 24'(7360);
			5973: out = 24'(16812);
			5974: out = 24'(18684);
			5975: out = 24'(30540);
			5976: out = 24'(5460);
			5977: out = 24'(-7656);
			5978: out = 24'(-7356);
			5979: out = 24'(-10596);
			5980: out = 24'(-16392);
			5981: out = 24'(-20304);
			5982: out = 24'(-23176);
			5983: out = 24'(2156);
			5984: out = 24'(18928);
			5985: out = 24'(8180);
			5986: out = 24'(-6380);
			5987: out = 24'(-13080);
			5988: out = 24'(11072);
			5989: out = 24'(16472);
			5990: out = 24'(15396);
			5991: out = 24'(4928);
			5992: out = 24'(5820);
			5993: out = 24'(-3360);
			5994: out = 24'(-9164);
			5995: out = 24'(-104);
			5996: out = 24'(-15048);
			5997: out = 24'(-26668);
			5998: out = 24'(6364);
			5999: out = 24'(28228);
			6000: out = 24'(-10980);
			6001: out = 24'(-32608);
			6002: out = 24'(-12228);
			6003: out = 24'(8452);
			6004: out = 24'(21788);
			6005: out = 24'(26212);
			6006: out = 24'(-23668);
			6007: out = 24'(-28876);
			6008: out = 24'(-2724);
			6009: out = 24'(8000);
			6010: out = 24'(25956);
			6011: out = 24'(-6556);
			6012: out = 24'(-22496);
			6013: out = 24'(9164);
			6014: out = 24'(30728);
			6015: out = 24'(24400);
			6016: out = 24'(-24724);
			6017: out = 24'(-40500);
			6018: out = 24'(-13076);
			6019: out = 24'(16416);
			6020: out = 24'(32032);
			6021: out = 24'(31944);
			6022: out = 24'(12144);
			6023: out = 24'(-9084);
			6024: out = 24'(-12492);
			6025: out = 24'(-4204);
			6026: out = 24'(22196);
			6027: out = 24'(24848);
			6028: out = 24'(-10056);
			6029: out = 24'(-9912);
			6030: out = 24'(15700);
			6031: out = 24'(7924);
			6032: out = 24'(-9360);
			6033: out = 24'(-18612);
			6034: out = 24'(-15332);
			6035: out = 24'(-29284);
			6036: out = 24'(-5460);
			6037: out = 24'(20836);
			6038: out = 24'(12448);
			6039: out = 24'(-5836);
			6040: out = 24'(-4572);
			6041: out = 24'(-7040);
			6042: out = 24'(-6108);
			6043: out = 24'(-19784);
			6044: out = 24'(-20884);
			6045: out = 24'(-11816);
			6046: out = 24'(9580);
			6047: out = 24'(24180);
			6048: out = 24'(38020);
			6049: out = 24'(18496);
			6050: out = 24'(-9452);
			6051: out = 24'(-3468);
			6052: out = 24'(-3956);
			6053: out = 24'(12328);
			6054: out = 24'(24576);
			6055: out = 24'(7788);
			6056: out = 24'(-22808);
			6057: out = 24'(-26096);
			6058: out = 24'(-15812);
			6059: out = 24'(-6608);
			6060: out = 24'(-14280);
			6061: out = 24'(-24936);
			6062: out = 24'(3288);
			6063: out = 24'(10604);
			6064: out = 24'(16660);
			6065: out = 24'(4772);
			6066: out = 24'(13084);
			6067: out = 24'(11680);
			6068: out = 24'(6700);
			6069: out = 24'(7032);
			6070: out = 24'(8136);
			6071: out = 24'(7560);
			6072: out = 24'(-840);
			6073: out = 24'(8528);
			6074: out = 24'(5536);
			6075: out = 24'(-24528);
			6076: out = 24'(-45232);
			6077: out = 24'(-17656);
			6078: out = 24'(-4280);
			6079: out = 24'(-11540);
			6080: out = 24'(748);
			6081: out = 24'(12088);
			6082: out = 24'(-13416);
			6083: out = 24'(-28384);
			6084: out = 24'(-11572);
			6085: out = 24'(15000);
			6086: out = 24'(20996);
			6087: out = 24'(9580);
			6088: out = 24'(-716);
			6089: out = 24'(2260);
			6090: out = 24'(1892);
			6091: out = 24'(18700);
			6092: out = 24'(4800);
			6093: out = 24'(-15684);
			6094: out = 24'(-2508);
			6095: out = 24'(16928);
			6096: out = 24'(9484);
			6097: out = 24'(1648);
			6098: out = 24'(-3888);
			6099: out = 24'(-5084);
			6100: out = 24'(-41940);
			6101: out = 24'(-39628);
			6102: out = 24'(15448);
			6103: out = 24'(27932);
			6104: out = 24'(-5324);
			6105: out = 24'(-3796);
			6106: out = 24'(5600);
			6107: out = 24'(3116);
			6108: out = 24'(-6392);
			6109: out = 24'(-6520);
			6110: out = 24'(15788);
			6111: out = 24'(80);
			6112: out = 24'(-6540);
			6113: out = 24'(-2016);
			6114: out = 24'(11400);
			6115: out = 24'(18440);
			6116: out = 24'(3912);
			6117: out = 24'(-9360);
			6118: out = 24'(-3148);
			6119: out = 24'(-17888);
			6120: out = 24'(-20560);
			6121: out = 24'(-9112);
			6122: out = 24'(-25840);
			6123: out = 24'(-15072);
			6124: out = 24'(26644);
			6125: out = 24'(42112);
			6126: out = 24'(-4968);
			6127: out = 24'(-40108);
			6128: out = 24'(-6512);
			6129: out = 24'(21200);
			6130: out = 24'(43800);
			6131: out = 24'(15568);
			6132: out = 24'(-11688);
			6133: out = 24'(-17252);
			6134: out = 24'(-14420);
			6135: out = 24'(-1152);
			6136: out = 24'(21988);
			6137: out = 24'(22712);
			6138: out = 24'(-5032);
			6139: out = 24'(-37540);
			6140: out = 24'(-34456);
			6141: out = 24'(10604);
			6142: out = 24'(32128);
			6143: out = 24'(-6560);
			6144: out = 24'(-18360);
			6145: out = 24'(-128);
			6146: out = 24'(944);
			6147: out = 24'(4188);
			6148: out = 24'(4196);
			6149: out = 24'(20280);
			6150: out = 24'(8236);
			6151: out = 24'(-14672);
			6152: out = 24'(-17092);
			6153: out = 24'(636);
			6154: out = 24'(16684);
			6155: out = 24'(-23112);
			6156: out = 24'(-32696);
			6157: out = 24'(-4436);
			6158: out = 24'(7880);
			6159: out = 24'(27816);
			6160: out = 24'(15276);
			6161: out = 24'(-7388);
			6162: out = 24'(-8912);
			6163: out = 24'(10188);
			6164: out = 24'(13144);
			6165: out = 24'(-9052);
			6166: out = 24'(-29896);
			6167: out = 24'(-3240);
			6168: out = 24'(5708);
			6169: out = 24'(-17656);
			6170: out = 24'(-8264);
			6171: out = 24'(24044);
			6172: out = 24'(14596);
			6173: out = 24'(-14476);
			6174: out = 24'(-1360);
			6175: out = 24'(3716);
			6176: out = 24'(-20532);
			6177: out = 24'(-11576);
			6178: out = 24'(8336);
			6179: out = 24'(-10336);
			6180: out = 24'(-15900);
			6181: out = 24'(5736);
			6182: out = 24'(17388);
			6183: out = 24'(24128);
			6184: out = 24'(18176);
			6185: out = 24'(864);
			6186: out = 24'(1968);
			6187: out = 24'(4972);
			6188: out = 24'(-20168);
			6189: out = 24'(-24128);
			6190: out = 24'(-4508);
			6191: out = 24'(952);
			6192: out = 24'(16824);
			6193: out = 24'(-932);
			6194: out = 24'(-14568);
			6195: out = 24'(18816);
			6196: out = 24'(36772);
			6197: out = 24'(29568);
			6198: out = 24'(-15192);
			6199: out = 24'(-28140);
			6200: out = 24'(-18380);
			6201: out = 24'(-3656);
			6202: out = 24'(21680);
			6203: out = 24'(12364);
			6204: out = 24'(3016);
			6205: out = 24'(3272);
			6206: out = 24'(-20892);
			6207: out = 24'(-21148);
			6208: out = 24'(9264);
			6209: out = 24'(18900);
			6210: out = 24'(2520);
			6211: out = 24'(-25524);
			6212: out = 24'(-14520);
			6213: out = 24'(7200);
			6214: out = 24'(26748);
			6215: out = 24'(16916);
			6216: out = 24'(14428);
			6217: out = 24'(9268);
			6218: out = 24'(2372);
			6219: out = 24'(13872);
			6220: out = 24'(5772);
			6221: out = 24'(-3200);
			6222: out = 24'(-15008);
			6223: out = 24'(-24744);
			6224: out = 24'(-26712);
			6225: out = 24'(3380);
			6226: out = 24'(24844);
			6227: out = 24'(2900);
			6228: out = 24'(-2728);
			6229: out = 24'(52);
			6230: out = 24'(3848);
			6231: out = 24'(2564);
			6232: out = 24'(948);
			6233: out = 24'(4444);
			6234: out = 24'(13772);
			6235: out = 24'(3284);
			6236: out = 24'(-8380);
			6237: out = 24'(-21060);
			6238: out = 24'(-22924);
			6239: out = 24'(-26936);
			6240: out = 24'(-13284);
			6241: out = 24'(-4112);
			6242: out = 24'(12452);
			6243: out = 24'(2088);
			6244: out = 24'(-6976);
			6245: out = 24'(11452);
			6246: out = 24'(26100);
			6247: out = 24'(38276);
			6248: out = 24'(13808);
			6249: out = 24'(-21176);
			6250: out = 24'(-38672);
			6251: out = 24'(-27180);
			6252: out = 24'(-10012);
			6253: out = 24'(-9044);
			6254: out = 24'(-10952);
			6255: out = 24'(2056);
			6256: out = 24'(2776);
			6257: out = 24'(15552);
			6258: out = 24'(26588);
			6259: out = 24'(33264);
			6260: out = 24'(28956);
			6261: out = 24'(-504);
			6262: out = 24'(-24692);
			6263: out = 24'(-33508);
			6264: out = 24'(-34792);
			6265: out = 24'(-20728);
			6266: out = 24'(2244);
			6267: out = 24'(15504);
			6268: out = 24'(11776);
			6269: out = 24'(15272);
			6270: out = 24'(41288);
			6271: out = 24'(20740);
			6272: out = 24'(-4340);
			6273: out = 24'(-23236);
			6274: out = 24'(664);
			6275: out = 24'(10384);
			6276: out = 24'(-6480);
			6277: out = 24'(3788);
			6278: out = 24'(1588);
			6279: out = 24'(-12976);
			6280: out = 24'(-10272);
			6281: out = 24'(-32128);
			6282: out = 24'(-20968);
			6283: out = 24'(18688);
			6284: out = 24'(31128);
			6285: out = 24'(16732);
			6286: out = 24'(3328);
			6287: out = 24'(22536);
			6288: out = 24'(19912);
			6289: out = 24'(-6088);
			6290: out = 24'(-34144);
			6291: out = 24'(-19528);
			6292: out = 24'(3388);
			6293: out = 24'(9816);
			6294: out = 24'(6020);
			6295: out = 24'(4388);
			6296: out = 24'(17816);
			6297: out = 24'(11896);
			6298: out = 24'(-3560);
			6299: out = 24'(-6660);
			6300: out = 24'(-6332);
			6301: out = 24'(4620);
			6302: out = 24'(2348);
			6303: out = 24'(-7364);
			6304: out = 24'(-25372);
			6305: out = 24'(-12316);
			6306: out = 24'(17928);
			6307: out = 24'(6288);
			6308: out = 24'(6892);
			6309: out = 24'(14260);
			6310: out = 24'(17940);
			6311: out = 24'(17592);
			6312: out = 24'(-11324);
			6313: out = 24'(-31876);
			6314: out = 24'(-12664);
			6315: out = 24'(14396);
			6316: out = 24'(20936);
			6317: out = 24'(8668);
			6318: out = 24'(1676);
			6319: out = 24'(5288);
			6320: out = 24'(13652);
			6321: out = 24'(5136);
			6322: out = 24'(-13000);
			6323: out = 24'(-13788);
			6324: out = 24'(5824);
			6325: out = 24'(34360);
			6326: out = 24'(20412);
			6327: out = 24'(-7224);
			6328: out = 24'(-20696);
			6329: out = 24'(-5388);
			6330: out = 24'(26624);
			6331: out = 24'(28668);
			6332: out = 24'(-7676);
			6333: out = 24'(-26632);
			6334: out = 24'(-10992);
			6335: out = 24'(-12324);
			6336: out = 24'(12208);
			6337: out = 24'(27152);
			6338: out = 24'(4720);
			6339: out = 24'(-36180);
			6340: out = 24'(-32932);
			6341: out = 24'(-23860);
			6342: out = 24'(-17396);
			6343: out = 24'(12548);
			6344: out = 24'(9952);
			6345: out = 24'(-13884);
			6346: out = 24'(6092);
			6347: out = 24'(-2416);
			6348: out = 24'(10652);
			6349: out = 24'(13968);
			6350: out = 24'(10776);
			6351: out = 24'(6884);
			6352: out = 24'(5396);
			6353: out = 24'(22404);
			6354: out = 24'(10740);
			6355: out = 24'(-22188);
			6356: out = 24'(-22180);
			6357: out = 24'(-6412);
			6358: out = 24'(640);
			6359: out = 24'(23212);
			6360: out = 24'(24128);
			6361: out = 24'(-2528);
			6362: out = 24'(-26348);
			6363: out = 24'(-20400);
			6364: out = 24'(-2808);
			6365: out = 24'(-12184);
			6366: out = 24'(-4864);
			6367: out = 24'(8640);
			6368: out = 24'(7272);
			6369: out = 24'(7680);
			6370: out = 24'(21548);
			6371: out = 24'(46976);
			6372: out = 24'(23684);
			6373: out = 24'(-27636);
			6374: out = 24'(-46296);
			6375: out = 24'(-22968);
			6376: out = 24'(2744);
			6377: out = 24'(11276);
			6378: out = 24'(-8652);
			6379: out = 24'(-16008);
			6380: out = 24'(772);
			6381: out = 24'(15928);
			6382: out = 24'(24196);
			6383: out = 24'(11988);
			6384: out = 24'(-11880);
			6385: out = 24'(-1732);
			6386: out = 24'(-676);
			6387: out = 24'(-3912);
			6388: out = 24'(7560);
			6389: out = 24'(-11356);
			6390: out = 24'(-27288);
			6391: out = 24'(-10752);
			6392: out = 24'(13328);
			6393: out = 24'(17368);
			6394: out = 24'(10276);
			6395: out = 24'(13892);
			6396: out = 24'(18884);
			6397: out = 24'(19908);
			6398: out = 24'(8216);
			6399: out = 24'(-9672);
			6400: out = 24'(-17208);
			6401: out = 24'(-10664);
			6402: out = 24'(-7552);
			6403: out = 24'(-30872);
			6404: out = 24'(-17364);
			6405: out = 24'(16184);
			6406: out = 24'(18216);
			6407: out = 24'(13580);
			6408: out = 24'(5504);
			6409: out = 24'(3104);
			6410: out = 24'(11620);
			6411: out = 24'(12956);
			6412: out = 24'(-19768);
			6413: out = 24'(-52540);
			6414: out = 24'(-40764);
			6415: out = 24'(5668);
			6416: out = 24'(39140);
			6417: out = 24'(24688);
			6418: out = 24'(1492);
			6419: out = 24'(12660);
			6420: out = 24'(21932);
			6421: out = 24'(-492);
			6422: out = 24'(-31324);
			6423: out = 24'(-32264);
			6424: out = 24'(-3956);
			6425: out = 24'(33144);
			6426: out = 24'(29244);
			6427: out = 24'(-18300);
			6428: out = 24'(-27452);
			6429: out = 24'(9500);
			6430: out = 24'(35920);
			6431: out = 24'(20508);
			6432: out = 24'(5148);
			6433: out = 24'(-4004);
			6434: out = 24'(-11276);
			6435: out = 24'(-12288);
			6436: out = 24'(3360);
			6437: out = 24'(17112);
			6438: out = 24'(-15168);
			6439: out = 24'(-47024);
			6440: out = 24'(-16192);
			6441: out = 24'(10448);
			6442: out = 24'(21116);
			6443: out = 24'(9216);
			6444: out = 24'(-5728);
			6445: out = 24'(-11252);
			6446: out = 24'(160);
			6447: out = 24'(10524);
			6448: out = 24'(23128);
			6449: out = 24'(7556);
			6450: out = 24'(-15044);
			6451: out = 24'(-23252);
			6452: out = 24'(-9488);
			6453: out = 24'(13256);
			6454: out = 24'(28484);
			6455: out = 24'(-15892);
			6456: out = 24'(-26556);
			6457: out = 24'(-2712);
			6458: out = 24'(16860);
			6459: out = 24'(23760);
			6460: out = 24'(7648);
			6461: out = 24'(-9736);
			6462: out = 24'(-26284);
			6463: out = 24'(-32140);
			6464: out = 24'(-36416);
			6465: out = 24'(3336);
			6466: out = 24'(17636);
			6467: out = 24'(5508);
			6468: out = 24'(19532);
			6469: out = 24'(7488);
			6470: out = 24'(-4324);
			6471: out = 24'(-1176);
			6472: out = 24'(1864);
			6473: out = 24'(5420);
			6474: out = 24'(2808);
			6475: out = 24'(17032);
			6476: out = 24'(17900);
			6477: out = 24'(488);
			6478: out = 24'(-21216);
			6479: out = 24'(-7332);
			6480: out = 24'(13480);
			6481: out = 24'(8884);
			6482: out = 24'(124);
			6483: out = 24'(6532);
			6484: out = 24'(16484);
			6485: out = 24'(5336);
			6486: out = 24'(-31036);
			6487: out = 24'(-40988);
			6488: out = 24'(-4880);
			6489: out = 24'(14344);
			6490: out = 24'(-17300);
			6491: out = 24'(-15060);
			6492: out = 24'(14716);
			6493: out = 24'(12792);
			6494: out = 24'(-12268);
			6495: out = 24'(-11780);
			6496: out = 24'(2468);
			6497: out = 24'(13000);
			6498: out = 24'(27600);
			6499: out = 24'(-2652);
			6500: out = 24'(-17724);
			6501: out = 24'(-17388);
			6502: out = 24'(-4144);
			6503: out = 24'(9316);
			6504: out = 24'(-1424);
			6505: out = 24'(6220);
			6506: out = 24'(14828);
			6507: out = 24'(6124);
			6508: out = 24'(-27556);
			6509: out = 24'(-39616);
			6510: out = 24'(-13096);
			6511: out = 24'(20336);
			6512: out = 24'(25220);
			6513: out = 24'(2180);
			6514: out = 24'(6220);
			6515: out = 24'(11356);
			6516: out = 24'(1788);
			6517: out = 24'(-7660);
			6518: out = 24'(-12256);
			6519: out = 24'(2140);
			6520: out = 24'(16752);
			6521: out = 24'(16372);
			6522: out = 24'(2200);
			6523: out = 24'(1848);
			6524: out = 24'(1296);
			6525: out = 24'(7800);
			6526: out = 24'(-4172);
			6527: out = 24'(-22248);
			6528: out = 24'(-22796);
			6529: out = 24'(-4520);
			6530: out = 24'(9308);
			6531: out = 24'(780);
			6532: out = 24'(-22588);
			6533: out = 24'(-16752);
			6534: out = 24'(-14208);
			6535: out = 24'(-4476);
			6536: out = 24'(3924);
			6537: out = 24'(820);
			6538: out = 24'(-12676);
			6539: out = 24'(-8324);
			6540: out = 24'(1068);
			6541: out = 24'(3932);
			6542: out = 24'(6520);
			6543: out = 24'(-3072);
			6544: out = 24'(6992);
			6545: out = 24'(20272);
			6546: out = 24'(21252);
			6547: out = 24'(6128);
			6548: out = 24'(-12164);
			6549: out = 24'(-18152);
			6550: out = 24'(-8588);
			6551: out = 24'(-16208);
			6552: out = 24'(-20536);
			6553: out = 24'(-7032);
			6554: out = 24'(6740);
			6555: out = 24'(32468);
			6556: out = 24'(19404);
			6557: out = 24'(9652);
			6558: out = 24'(-13632);
			6559: out = 24'(-11152);
			6560: out = 24'(3244);
			6561: out = 24'(-616);
			6562: out = 24'(16892);
			6563: out = 24'(12240);
			6564: out = 24'(7660);
			6565: out = 24'(4776);
			6566: out = 24'(5584);
			6567: out = 24'(-21184);
			6568: out = 24'(-25496);
			6569: out = 24'(-8668);
			6570: out = 24'(-512);
			6571: out = 24'(-10540);
			6572: out = 24'(516);
			6573: out = 24'(-12260);
			6574: out = 24'(-26164);
			6575: out = 24'(-8388);
			6576: out = 24'(5004);
			6577: out = 24'(14784);
			6578: out = 24'(10468);
			6579: out = 24'(-5832);
			6580: out = 24'(-22880);
			6581: out = 24'(-21720);
			6582: out = 24'(10296);
			6583: out = 24'(31052);
			6584: out = 24'(31480);
			6585: out = 24'(-13520);
			6586: out = 24'(-46168);
			6587: out = 24'(-18492);
			6588: out = 24'(23744);
			6589: out = 24'(50512);
			6590: out = 24'(24508);
			6591: out = 24'(-11956);
			6592: out = 24'(-15796);
			6593: out = 24'(5384);
			6594: out = 24'(4244);
			6595: out = 24'(-27280);
			6596: out = 24'(-22720);
			6597: out = 24'(-12);
			6598: out = 24'(5760);
			6599: out = 24'(28540);
			6600: out = 24'(8956);
			6601: out = 24'(9892);
			6602: out = 24'(28092);
			6603: out = 24'(19140);
			6604: out = 24'(-9744);
			6605: out = 24'(-34240);
			6606: out = 24'(-27348);
			6607: out = 24'(-10032);
			6608: out = 24'(20152);
			6609: out = 24'(35552);
			6610: out = 24'(7380);
			6611: out = 24'(2228);
			6612: out = 24'(3356);
			6613: out = 24'(-620);
			6614: out = 24'(10520);
			6615: out = 24'(-5764);
			6616: out = 24'(-2200);
			6617: out = 24'(20412);
			6618: out = 24'(24860);
			6619: out = 24'(-17156);
			6620: out = 24'(-46096);
			6621: out = 24'(-43572);
			6622: out = 24'(-6652);
			6623: out = 24'(27184);
			6624: out = 24'(30772);
			6625: out = 24'(-7784);
			6626: out = 24'(-11168);
			6627: out = 24'(1620);
			6628: out = 24'(2736);
			6629: out = 24'(30008);
			6630: out = 24'(26088);
			6631: out = 24'(-2400);
			6632: out = 24'(-7184);
			6633: out = 24'(7956);
			6634: out = 24'(-4876);
			6635: out = 24'(-46404);
			6636: out = 24'(-43124);
			6637: out = 24'(428);
			6638: out = 24'(5132);
			6639: out = 24'(22616);
			6640: out = 24'(27252);
			6641: out = 24'(15876);
			6642: out = 24'(-1060);
			6643: out = 24'(-10364);
			6644: out = 24'(964);
			6645: out = 24'(9596);
			6646: out = 24'(1392);
			6647: out = 24'(-13844);
			6648: out = 24'(-8940);
			6649: out = 24'(-10524);
			6650: out = 24'(-11752);
			6651: out = 24'(12884);
			6652: out = 24'(19248);
			6653: out = 24'(2016);
			6654: out = 24'(8288);
			6655: out = 24'(9080);
			6656: out = 24'(4244);
			6657: out = 24'(3064);
			6658: out = 24'(-4648);
			6659: out = 24'(-20412);
			6660: out = 24'(-9136);
			6661: out = 24'(7504);
			6662: out = 24'(26488);
			6663: out = 24'(21208);
			6664: out = 24'(21236);
			6665: out = 24'(19580);
			6666: out = 24'(10652);
			6667: out = 24'(3236);
			6668: out = 24'(-9164);
			6669: out = 24'(-16984);
			6670: out = 24'(-22056);
			6671: out = 24'(-6336);
			6672: out = 24'(3460);
			6673: out = 24'(-2524);
			6674: out = 24'(-25396);
			6675: out = 24'(-19424);
			6676: out = 24'(-688);
			6677: out = 24'(28232);
			6678: out = 24'(32512);
			6679: out = 24'(5472);
			6680: out = 24'(-8392);
			6681: out = 24'(-17840);
			6682: out = 24'(-476);
			6683: out = 24'(-6396);
			6684: out = 24'(-4880);
			6685: out = 24'(23368);
			6686: out = 24'(20016);
			6687: out = 24'(-12712);
			6688: out = 24'(-36428);
			6689: out = 24'(-40616);
			6690: out = 24'(10240);
			6691: out = 24'(40956);
			6692: out = 24'(13552);
			6693: out = 24'(-9004);
			6694: out = 24'(-908);
			6695: out = 24'(13016);
			6696: out = 24'(1164);
			6697: out = 24'(-23604);
			6698: out = 24'(-13916);
			6699: out = 24'(22740);
			6700: out = 24'(32424);
			6701: out = 24'(17164);
			6702: out = 24'(6404);
			6703: out = 24'(-2528);
			6704: out = 24'(3500);
			6705: out = 24'(-5892);
			6706: out = 24'(-14356);
			6707: out = 24'(10800);
			6708: out = 24'(17432);
			6709: out = 24'(-19296);
			6710: out = 24'(-40316);
			6711: out = 24'(-18844);
			6712: out = 24'(10292);
			6713: out = 24'(7840);
			6714: out = 24'(6636);
			6715: out = 24'(12812);
			6716: out = 24'(-5152);
			6717: out = 24'(-16572);
			6718: out = 24'(-5900);
			6719: out = 24'(17712);
			6720: out = 24'(11804);
			6721: out = 24'(-16788);
			6722: out = 24'(-31992);
			6723: out = 24'(-8108);
			6724: out = 24'(33504);
			6725: out = 24'(19824);
			6726: out = 24'(-1340);
			6727: out = 24'(4536);
			6728: out = 24'(6664);
			6729: out = 24'(3616);
			6730: out = 24'(2520);
			6731: out = 24'(11848);
			6732: out = 24'(22016);
			6733: out = 24'(-3820);
			6734: out = 24'(-29932);
			6735: out = 24'(-26616);
			6736: out = 24'(-14604);
			6737: out = 24'(11568);
			6738: out = 24'(7692);
			6739: out = 24'(-11124);
			6740: out = 24'(5736);
			6741: out = 24'(22520);
			6742: out = 24'(4896);
			6743: out = 24'(-34972);
			6744: out = 24'(-43864);
			6745: out = 24'(-7036);
			6746: out = 24'(23640);
			6747: out = 24'(22680);
			6748: out = 24'(16032);
			6749: out = 24'(16048);
			6750: out = 24'(6508);
			6751: out = 24'(5608);
			6752: out = 24'(-4824);
			6753: out = 24'(-22812);
			6754: out = 24'(-32128);
			6755: out = 24'(2364);
			6756: out = 24'(25532);
			6757: out = 24'(2236);
			6758: out = 24'(-988);
			6759: out = 24'(11380);
			6760: out = 24'(21780);
			6761: out = 24'(4504);
			6762: out = 24'(-2456);
			6763: out = 24'(6384);
			6764: out = 24'(15416);
			6765: out = 24'(8016);
			6766: out = 24'(-8944);
			6767: out = 24'(-3456);
			6768: out = 24'(2364);
			6769: out = 24'(332);
			6770: out = 24'(-6012);
			6771: out = 24'(-10084);
			6772: out = 24'(-17012);
			6773: out = 24'(-9472);
			6774: out = 24'(-1436);
			6775: out = 24'(-3984);
			6776: out = 24'(-5164);
			6777: out = 24'(-10496);
			6778: out = 24'(-29184);
			6779: out = 24'(-17136);
			6780: out = 24'(25820);
			6781: out = 24'(43132);
			6782: out = 24'(-8064);
			6783: out = 24'(-54120);
			6784: out = 24'(-35704);
			6785: out = 24'(4440);
			6786: out = 24'(38264);
			6787: out = 24'(27216);
			6788: out = 24'(-12236);
			6789: out = 24'(-16420);
			6790: out = 24'(9668);
			6791: out = 24'(10244);
			6792: out = 24'(-4192);
			6793: out = 24'(-26540);
			6794: out = 24'(-15116);
			6795: out = 24'(18260);
			6796: out = 24'(10524);
			6797: out = 24'(10812);
			6798: out = 24'(12128);
			6799: out = 24'(15364);
			6800: out = 24'(10804);
			6801: out = 24'(-4288);
			6802: out = 24'(-35076);
			6803: out = 24'(-27320);
			6804: out = 24'(-16480);
			6805: out = 24'(-15576);
			6806: out = 24'(24012);
			6807: out = 24'(35984);
			6808: out = 24'(-3424);
			6809: out = 24'(-10552);
			6810: out = 24'(-10072);
			6811: out = 24'(4308);
			6812: out = 24'(11564);
			6813: out = 24'(16128);
			6814: out = 24'(17892);
			6815: out = 24'(440);
			6816: out = 24'(11968);
			6817: out = 24'(15212);
			6818: out = 24'(-2076);
			6819: out = 24'(-15296);
			6820: out = 24'(-9492);
			6821: out = 24'(-11112);
			6822: out = 24'(3548);
			6823: out = 24'(10508);
			6824: out = 24'(1436);
			6825: out = 24'(-5280);
			6826: out = 24'(2784);
			6827: out = 24'(21416);
			6828: out = 24'(15508);
			6829: out = 24'(-13596);
			6830: out = 24'(-13660);
			6831: out = 24'(-6588);
			6832: out = 24'(-15368);
			6833: out = 24'(-9328);
			6834: out = 24'(12952);
			6835: out = 24'(-3876);
			6836: out = 24'(-31664);
			6837: out = 24'(-18188);
			6838: out = 24'(3384);
			6839: out = 24'(15780);
			6840: out = 24'(9884);
			6841: out = 24'(-21212);
			6842: out = 24'(-21516);
			6843: out = 24'(-6772);
			6844: out = 24'(34616);
			6845: out = 24'(36904);
			6846: out = 24'(-944);
			6847: out = 24'(-16492);
			6848: out = 24'(-9436);
			6849: out = 24'(-3176);
			6850: out = 24'(-3564);
			6851: out = 24'(-9984);
			6852: out = 24'(-12576);
			6853: out = 24'(17708);
			6854: out = 24'(30672);
			6855: out = 24'(-7120);
			6856: out = 24'(-38860);
			6857: out = 24'(-28268);
			6858: out = 24'(8124);
			6859: out = 24'(18568);
			6860: out = 24'(30704);
			6861: out = 24'(18768);
			6862: out = 24'(-9160);
			6863: out = 24'(-29844);
			6864: out = 24'(-31080);
			6865: out = 24'(1560);
			6866: out = 24'(18708);
			6867: out = 24'(10296);
			6868: out = 24'(8560);
			6869: out = 24'(15016);
			6870: out = 24'(11112);
			6871: out = 24'(14052);
			6872: out = 24'(4792);
			6873: out = 24'(-4124);
			6874: out = 24'(-30592);
			6875: out = 24'(-26828);
			6876: out = 24'(-9800);
			6877: out = 24'(4432);
			6878: out = 24'(6800);
			6879: out = 24'(-11308);
			6880: out = 24'(-7444);
			6881: out = 24'(19468);
			6882: out = 24'(16772);
			6883: out = 24'(-14048);
			6884: out = 24'(-35420);
			6885: out = 24'(-28584);
			6886: out = 24'(3860);
			6887: out = 24'(44036);
			6888: out = 24'(33744);
			6889: out = 24'(-3724);
			6890: out = 24'(-19984);
			6891: out = 24'(-19288);
			6892: out = 24'(-7140);
			6893: out = 24'(13724);
			6894: out = 24'(23720);
			6895: out = 24'(1028);
			6896: out = 24'(1012);
			6897: out = 24'(-788);
			6898: out = 24'(-6368);
			6899: out = 24'(4060);
			6900: out = 24'(-11536);
			6901: out = 24'(4968);
			6902: out = 24'(22664);
			6903: out = 24'(252);
			6904: out = 24'(-2636);
			6905: out = 24'(3256);
			6906: out = 24'(-4400);
			6907: out = 24'(-18368);
			6908: out = 24'(-25860);
			6909: out = 24'(3816);
			6910: out = 24'(16256);
			6911: out = 24'(5868);
			6912: out = 24'(-1376);
			6913: out = 24'(-668);
			6914: out = 24'(-556);
			6915: out = 24'(-22276);
			6916: out = 24'(-15596);
			6917: out = 24'(10080);
			6918: out = 24'(16656);
			6919: out = 24'(17984);
			6920: out = 24'(16524);
			6921: out = 24'(7300);
			6922: out = 24'(-18280);
			6923: out = 24'(-30420);
			6924: out = 24'(-3896);
			6925: out = 24'(8584);
			6926: out = 24'(16692);
			6927: out = 24'(13428);
			6928: out = 24'(-8388);
			6929: out = 24'(-23148);
			6930: out = 24'(-16088);
			6931: out = 24'(13744);
			6932: out = 24'(6472);
			6933: out = 24'(-12920);
			6934: out = 24'(-12);
			6935: out = 24'(4220);
			6936: out = 24'(12656);
			6937: out = 24'(19464);
			6938: out = 24'(12044);
			6939: out = 24'(15648);
			6940: out = 24'(-1848);
			6941: out = 24'(-14004);
			6942: out = 24'(-10240);
			6943: out = 24'(-6632);
			6944: out = 24'(9272);
			6945: out = 24'(7952);
			6946: out = 24'(-8488);
			6947: out = 24'(-11556);
			6948: out = 24'(-5432);
			6949: out = 24'(-1864);
			6950: out = 24'(10240);
			6951: out = 24'(9728);
			6952: out = 24'(4316);
			6953: out = 24'(5980);
			6954: out = 24'(-15676);
			6955: out = 24'(-29356);
			6956: out = 24'(-4264);
			6957: out = 24'(13832);
			6958: out = 24'(-944);
			6959: out = 24'(7456);
			6960: out = 24'(12752);
			6961: out = 24'(4404);
			6962: out = 24'(180);
			6963: out = 24'(-5592);
			6964: out = 24'(-2292);
			6965: out = 24'(-696);
			6966: out = 24'(18244);
			6967: out = 24'(26644);
			6968: out = 24'(-6324);
			6969: out = 24'(-37336);
			6970: out = 24'(-24600);
			6971: out = 24'(2364);
			6972: out = 24'(19220);
			6973: out = 24'(7296);
			6974: out = 24'(15408);
			6975: out = 24'(5484);
			6976: out = 24'(-19200);
			6977: out = 24'(-1628);
			6978: out = 24'(27272);
			6979: out = 24'(17872);
			6980: out = 24'(-26016);
			6981: out = 24'(-40808);
			6982: out = 24'(-19096);
			6983: out = 24'(9836);
			6984: out = 24'(39872);
			6985: out = 24'(8184);
			6986: out = 24'(-27124);
			6987: out = 24'(-2904);
			6988: out = 24'(25240);
			6989: out = 24'(30412);
			6990: out = 24'(8976);
			6991: out = 24'(-9596);
			6992: out = 24'(-1348);
			6993: out = 24'(2276);
			6994: out = 24'(-2032);
			6995: out = 24'(-3912);
			6996: out = 24'(3412);
			6997: out = 24'(20932);
			6998: out = 24'(15268);
			6999: out = 24'(-25280);
			7000: out = 24'(-30752);
			7001: out = 24'(-4476);
			7002: out = 24'(12456);
			7003: out = 24'(4840);
			7004: out = 24'(8024);
			7005: out = 24'(16268);
			7006: out = 24'(-3368);
			7007: out = 24'(-16584);
			7008: out = 24'(-1888);
			7009: out = 24'(21160);
			7010: out = 24'(24272);
			7011: out = 24'(-15364);
			7012: out = 24'(-24728);
			7013: out = 24'(-9868);
			7014: out = 24'(-7552);
			7015: out = 24'(5452);
			7016: out = 24'(7484);
			7017: out = 24'(-10176);
			7018: out = 24'(-22724);
			7019: out = 24'(856);
			7020: out = 24'(17596);
			7021: out = 24'(12248);
			7022: out = 24'(10680);
			7023: out = 24'(6744);
			7024: out = 24'(-5952);
			7025: out = 24'(-812);
			7026: out = 24'(-3240);
			7027: out = 24'(-3456);
			7028: out = 24'(11392);
			7029: out = 24'(11816);
			7030: out = 24'(1416);
			7031: out = 24'(-6948);
			7032: out = 24'(-7940);
			7033: out = 24'(2552);
			7034: out = 24'(1876);
			7035: out = 24'(-14892);
			7036: out = 24'(-8804);
			7037: out = 24'(3284);
			7038: out = 24'(22640);
			7039: out = 24'(3588);
			7040: out = 24'(-3136);
			7041: out = 24'(13628);
			7042: out = 24'(7100);
			7043: out = 24'(-13508);
			7044: out = 24'(-2332);
			7045: out = 24'(8876);
			7046: out = 24'(-1088);
			7047: out = 24'(-22032);
			7048: out = 24'(-16920);
			7049: out = 24'(-11140);
			7050: out = 24'(-9320);
			7051: out = 24'(5828);
			7052: out = 24'(4124);
			7053: out = 24'(-1216);
			7054: out = 24'(-148);
			7055: out = 24'(6176);
			7056: out = 24'(1776);
			7057: out = 24'(-7404);
			7058: out = 24'(-1472);
			7059: out = 24'(7516);
			7060: out = 24'(16424);
			7061: out = 24'(5680);
			7062: out = 24'(-9596);
			7063: out = 24'(368);
			7064: out = 24'(23408);
			7065: out = 24'(14804);
			7066: out = 24'(-10264);
			7067: out = 24'(2068);
			7068: out = 24'(3452);
			7069: out = 24'(-7224);
			7070: out = 24'(-15792);
			7071: out = 24'(-20040);
			7072: out = 24'(4596);
			7073: out = 24'(12968);
			7074: out = 24'(-8656);
			7075: out = 24'(1168);
			7076: out = 24'(5580);
			7077: out = 24'(11180);
			7078: out = 24'(19404);
			7079: out = 24'(7836);
			7080: out = 24'(-7204);
			7081: out = 24'(-29204);
			7082: out = 24'(-19072);
			7083: out = 24'(-1544);
			7084: out = 24'(16964);
			7085: out = 24'(14124);
			7086: out = 24'(7424);
			7087: out = 24'(15604);
			7088: out = 24'(-352);
			7089: out = 24'(-25180);
			7090: out = 24'(-29396);
			7091: out = 24'(-7228);
			7092: out = 24'(11292);
			7093: out = 24'(14348);
			7094: out = 24'(20080);
			7095: out = 24'(19592);
			7096: out = 24'(-4148);
			7097: out = 24'(-23444);
			7098: out = 24'(-16348);
			7099: out = 24'(-4980);
			7100: out = 24'(-6104);
			7101: out = 24'(-4248);
			7102: out = 24'(14480);
			7103: out = 24'(19680);
			7104: out = 24'(-8536);
			7105: out = 24'(-12424);
			7106: out = 24'(-168);
			7107: out = 24'(4016);
			7108: out = 24'(5516);
			7109: out = 24'(4476);
			7110: out = 24'(-464);
			7111: out = 24'(-9908);
			7112: out = 24'(-16136);
			7113: out = 24'(-3736);
			7114: out = 24'(5128);
			7115: out = 24'(-1992);
			7116: out = 24'(8848);
			7117: out = 24'(27488);
			7118: out = 24'(11664);
			7119: out = 24'(-16488);
			7120: out = 24'(-31616);
			7121: out = 24'(-4120);
			7122: out = 24'(27728);
			7123: out = 24'(23584);
			7124: out = 24'(3060);
			7125: out = 24'(-6004);
			7126: out = 24'(-6492);
			7127: out = 24'(-16448);
			7128: out = 24'(-13928);
			7129: out = 24'(11844);
			7130: out = 24'(27656);
			7131: out = 24'(-5720);
			7132: out = 24'(-40456);
			7133: out = 24'(-20192);
			7134: out = 24'(9844);
			7135: out = 24'(22348);
			7136: out = 24'(9648);
			7137: out = 24'(-19548);
			7138: out = 24'(-28648);
			7139: out = 24'(-580);
			7140: out = 24'(31048);
			7141: out = 24'(27272);
			7142: out = 24'(-2228);
			7143: out = 24'(-14144);
			7144: out = 24'(6720);
			7145: out = 24'(14196);
			7146: out = 24'(17208);
			7147: out = 24'(9672);
			7148: out = 24'(5032);
			7149: out = 24'(1560);
			7150: out = 24'(-3480);
			7151: out = 24'(-8252);
			7152: out = 24'(-8964);
			7153: out = 24'(-6004);
			7154: out = 24'(-14068);
			7155: out = 24'(-5740);
			7156: out = 24'(1656);
			7157: out = 24'(7376);
			7158: out = 24'(-6992);
			7159: out = 24'(-23788);
			7160: out = 24'(-22228);
			7161: out = 24'(568);
			7162: out = 24'(24648);
			7163: out = 24'(13664);
			7164: out = 24'(316);
			7165: out = 24'(-4588);
			7166: out = 24'(4960);
			7167: out = 24'(16368);
			7168: out = 24'(1316);
			7169: out = 24'(464);
			7170: out = 24'(13840);
			7171: out = 24'(17192);
			7172: out = 24'(-16660);
			7173: out = 24'(-42508);
			7174: out = 24'(-17152);
			7175: out = 24'(14072);
			7176: out = 24'(7444);
			7177: out = 24'(-22456);
			7178: out = 24'(-15428);
			7179: out = 24'(4336);
			7180: out = 24'(14016);
			7181: out = 24'(26956);
			7182: out = 24'(12860);
			7183: out = 24'(-9800);
			7184: out = 24'(-26052);
			7185: out = 24'(-9644);
			7186: out = 24'(21616);
			7187: out = 24'(26888);
			7188: out = 24'(2528);
			7189: out = 24'(-24200);
			7190: out = 24'(-13348);
			7191: out = 24'(21060);
			7192: out = 24'(19324);
			7193: out = 24'(424);
			7194: out = 24'(-17716);
			7195: out = 24'(-8976);
			7196: out = 24'(2152);
			7197: out = 24'(-10648);
			7198: out = 24'(168);
			7199: out = 24'(15912);
			7200: out = 24'(13428);
			7201: out = 24'(-12496);
			7202: out = 24'(-19320);
			7203: out = 24'(-8744);
			7204: out = 24'(4024);
			7205: out = 24'(1312);
			7206: out = 24'(-7784);
			7207: out = 24'(-356);
			7208: out = 24'(7776);
			7209: out = 24'(-9648);
			7210: out = 24'(-13220);
			7211: out = 24'(-6512);
			7212: out = 24'(13508);
			7213: out = 24'(27952);
			7214: out = 24'(9696);
			7215: out = 24'(-12276);
			7216: out = 24'(-22928);
			7217: out = 24'(2376);
			7218: out = 24'(8260);
			7219: out = 24'(-912);
			7220: out = 24'(-5888);
			7221: out = 24'(10688);
			7222: out = 24'(26676);
			7223: out = 24'(7448);
			7224: out = 24'(3700);
			7225: out = 24'(3644);
			7226: out = 24'(3532);
			7227: out = 24'(-948);
			7228: out = 24'(-11072);
			7229: out = 24'(-3736);
			7230: out = 24'(12304);
			7231: out = 24'(10012);
			7232: out = 24'(-2300);
			7233: out = 24'(5124);
			7234: out = 24'(13808);
			7235: out = 24'(-2072);
			7236: out = 24'(-27884);
			7237: out = 24'(-24228);
			7238: out = 24'(-9068);
			7239: out = 24'(-7632);
			7240: out = 24'(4132);
			7241: out = 24'(2864);
			7242: out = 24'(-17908);
			7243: out = 24'(-22156);
			7244: out = 24'(-6212);
			7245: out = 24'(10460);
			7246: out = 24'(7908);
			7247: out = 24'(5452);
			7248: out = 24'(-14768);
			7249: out = 24'(-24988);
			7250: out = 24'(-17336);
			7251: out = 24'(-472);
			7252: out = 24'(12344);
			7253: out = 24'(220);
			7254: out = 24'(3012);
			7255: out = 24'(5232);
			7256: out = 24'(-2244);
			7257: out = 24'(1672);
			7258: out = 24'(7900);
			7259: out = 24'(1336);
			7260: out = 24'(3280);
			7261: out = 24'(-9964);
			7262: out = 24'(-8856);
			7263: out = 24'(-676);
			7264: out = 24'(-5492);
			7265: out = 24'(10772);
			7266: out = 24'(12072);
			7267: out = 24'(-16500);
			7268: out = 24'(-21308);
			7269: out = 24'(-1132);
			7270: out = 24'(-5272);
			7271: out = 24'(1680);
			7272: out = 24'(15848);
			7273: out = 24'(7908);
			7274: out = 24'(-24112);
			7275: out = 24'(-23720);
			7276: out = 24'(14232);
			7277: out = 24'(29188);
			7278: out = 24'(13864);
			7279: out = 24'(-7736);
			7280: out = 24'(-4476);
			7281: out = 24'(3572);
			7282: out = 24'(-6000);
			7283: out = 24'(-16860);
			7284: out = 24'(-21716);
			7285: out = 24'(-1608);
			7286: out = 24'(23120);
			7287: out = 24'(27380);
			7288: out = 24'(-2000);
			7289: out = 24'(-10348);
			7290: out = 24'(7052);
			7291: out = 24'(17732);
			7292: out = 24'(19824);
			7293: out = 24'(1860);
			7294: out = 24'(-20792);
			7295: out = 24'(-30304);
			7296: out = 24'(-14256);
			7297: out = 24'(-17204);
			7298: out = 24'(-6920);
			7299: out = 24'(14444);
			7300: out = 24'(21740);
			7301: out = 24'(13024);
			7302: out = 24'(-5204);
			7303: out = 24'(-18208);
			7304: out = 24'(-2552);
			7305: out = 24'(18288);
			7306: out = 24'(13076);
			7307: out = 24'(-4952);
			7308: out = 24'(-768);
			7309: out = 24'(1476);
			7310: out = 24'(-8156);
			7311: out = 24'(1844);
			7312: out = 24'(-10472);
			7313: out = 24'(-10588);
			7314: out = 24'(4496);
			7315: out = 24'(8872);
			7316: out = 24'(13568);
			7317: out = 24'(19212);
			7318: out = 24'(13356);
			7319: out = 24'(10476);
			7320: out = 24'(1928);
			7321: out = 24'(-3264);
			7322: out = 24'(-11508);
			7323: out = 24'(-15616);
			7324: out = 24'(6528);
			7325: out = 24'(7240);
			7326: out = 24'(-184);
			7327: out = 24'(11680);
			7328: out = 24'(12264);
			7329: out = 24'(-5468);
			7330: out = 24'(-27372);
			7331: out = 24'(-34580);
			7332: out = 24'(-12180);
			7333: out = 24'(676);
			7334: out = 24'(24316);
			7335: out = 24'(19420);
			7336: out = 24'(4092);
			7337: out = 24'(2532);
			7338: out = 24'(-968);
			7339: out = 24'(8932);
			7340: out = 24'(13824);
			7341: out = 24'(12244);
			7342: out = 24'(-2880);
			7343: out = 24'(-2464);
			7344: out = 24'(7776);
			7345: out = 24'(3996);
			7346: out = 24'(2372);
			7347: out = 24'(-3392);
			7348: out = 24'(-11500);
			7349: out = 24'(-17024);
			7350: out = 24'(9212);
			7351: out = 24'(4420);
			7352: out = 24'(-15748);
			7353: out = 24'(-2820);
			7354: out = 24'(12528);
			7355: out = 24'(12828);
			7356: out = 24'(-13040);
			7357: out = 24'(-2072);
			7358: out = 24'(11488);
			7359: out = 24'(23224);
			7360: out = 24'(17724);
			7361: out = 24'(2680);
			7362: out = 24'(-15820);
			7363: out = 24'(-23348);
			7364: out = 24'(-32432);
			7365: out = 24'(-9984);
			7366: out = 24'(23812);
			7367: out = 24'(-1784);
			7368: out = 24'(-34860);
			7369: out = 24'(-13728);
			7370: out = 24'(3044);
			7371: out = 24'(17460);
			7372: out = 24'(27020);
			7373: out = 24'(19336);
			7374: out = 24'(-6424);
			7375: out = 24'(-25796);
			7376: out = 24'(-23700);
			7377: out = 24'(-11316);
			7378: out = 24'(14488);
			7379: out = 24'(28088);
			7380: out = 24'(18780);
			7381: out = 24'(5376);
			7382: out = 24'(1856);
			7383: out = 24'(10732);
			7384: out = 24'(18308);
			7385: out = 24'(4500);
			7386: out = 24'(-14988);
			7387: out = 24'(-11688);
			7388: out = 24'(10460);
			7389: out = 24'(8084);
			7390: out = 24'(-19556);
			7391: out = 24'(-19724);
			7392: out = 24'(-1484);
			7393: out = 24'(2524);
			7394: out = 24'(-2280);
			7395: out = 24'(11040);
			7396: out = 24'(-7348);
			7397: out = 24'(-7624);
			7398: out = 24'(9716);
			7399: out = 24'(29268);
			7400: out = 24'(10972);
			7401: out = 24'(-24360);
			7402: out = 24'(-30916);
			7403: out = 24'(-4480);
			7404: out = 24'(16892);
			7405: out = 24'(-72);
			7406: out = 24'(-19204);
			7407: out = 24'(-10948);
			7408: out = 24'(160);
			7409: out = 24'(10632);
			7410: out = 24'(21548);
			7411: out = 24'(10080);
			7412: out = 24'(-1580);
			7413: out = 24'(-14680);
			7414: out = 24'(-16196);
			7415: out = 24'(2896);
			7416: out = 24'(10996);
			7417: out = 24'(19648);
			7418: out = 24'(30048);
			7419: out = 24'(7600);
			7420: out = 24'(-11820);
			7421: out = 24'(-23884);
			7422: out = 24'(-9572);
			7423: out = 24'(13408);
			7424: out = 24'(11756);
			7425: out = 24'(-620);
			7426: out = 24'(1044);
			7427: out = 24'(-15984);
			7428: out = 24'(-16404);
			7429: out = 24'(7688);
			7430: out = 24'(-1156);
			7431: out = 24'(5324);
			7432: out = 24'(21432);
			7433: out = 24'(17176);
			7434: out = 24'(-22168);
			7435: out = 24'(-37444);
			7436: out = 24'(-19808);
			7437: out = 24'(11104);
			7438: out = 24'(27408);
			7439: out = 24'(16584);
			7440: out = 24'(-11616);
			7441: out = 24'(-16876);
			7442: out = 24'(-16048);
			7443: out = 24'(-5016);
			7444: out = 24'(26784);
			7445: out = 24'(31044);
			7446: out = 24'(-8948);
			7447: out = 24'(-22664);
			7448: out = 24'(-16140);
			7449: out = 24'(-2184);
			7450: out = 24'(15408);
			7451: out = 24'(3268);
			7452: out = 24'(-3736);
			7453: out = 24'(7340);
			7454: out = 24'(31624);
			7455: out = 24'(22796);
			7456: out = 24'(-3820);
			7457: out = 24'(-13984);
			7458: out = 24'(-264);
			7459: out = 24'(12800);
			7460: out = 24'(17972);
			7461: out = 24'(9284);
			7462: out = 24'(3288);
			7463: out = 24'(-3620);
			7464: out = 24'(-15008);
			7465: out = 24'(-30300);
			7466: out = 24'(-18864);
			7467: out = 24'(5164);
			7468: out = 24'(-2968);
			7469: out = 24'(-18876);
			7470: out = 24'(3312);
			7471: out = 24'(14924);
			7472: out = 24'(7728);
			7473: out = 24'(-6344);
			7474: out = 24'(-4220);
			7475: out = 24'(-13432);
			7476: out = 24'(-17564);
			7477: out = 24'(9304);
			7478: out = 24'(24524);
			7479: out = 24'(6756);
			7480: out = 24'(-1996);
			7481: out = 24'(5748);
			7482: out = 24'(10360);
			7483: out = 24'(-4960);
			7484: out = 24'(-31416);
			7485: out = 24'(-26428);
			7486: out = 24'(-7492);
			7487: out = 24'(17308);
			7488: out = 24'(13996);
			7489: out = 24'(-3700);
			7490: out = 24'(-13960);
			7491: out = 24'(-3684);
			7492: out = 24'(24312);
			7493: out = 24'(25388);
			7494: out = 24'(424);
			7495: out = 24'(-17708);
			7496: out = 24'(-10860);
			7497: out = 24'(12100);
			7498: out = 24'(12324);
			7499: out = 24'(-9564);
			7500: out = 24'(-6664);
			7501: out = 24'(9976);
			7502: out = 24'(1916);
			7503: out = 24'(-3140);
			7504: out = 24'(-756);
			7505: out = 24'(4676);
			7506: out = 24'(19160);
			7507: out = 24'(5460);
			7508: out = 24'(-1028);
			7509: out = 24'(-1044);
			7510: out = 24'(-4792);
			7511: out = 24'(8856);
			7512: out = 24'(728);
			7513: out = 24'(-1316);
			7514: out = 24'(1692);
			7515: out = 24'(-7172);
			7516: out = 24'(-7736);
			7517: out = 24'(-6976);
			7518: out = 24'(-4056);
			7519: out = 24'(9144);
			7520: out = 24'(2224);
			7521: out = 24'(-3980);
			7522: out = 24'(5428);
			7523: out = 24'(10696);
			7524: out = 24'(5316);
			7525: out = 24'(-13192);
			7526: out = 24'(-20112);
			7527: out = 24'(-12500);
			7528: out = 24'(3236);
			7529: out = 24'(17264);
			7530: out = 24'(5808);
			7531: out = 24'(-8880);
			7532: out = 24'(-2228);
			7533: out = 24'(4532);
			7534: out = 24'(-14592);
			7535: out = 24'(-21280);
			7536: out = 24'(-5096);
			7537: out = 24'(-1944);
			7538: out = 24'(6784);
			7539: out = 24'(-1532);
			7540: out = 24'(-15676);
			7541: out = 24'(824);
			7542: out = 24'(21260);
			7543: out = 24'(14960);
			7544: out = 24'(-3924);
			7545: out = 24'(-13008);
			7546: out = 24'(-5640);
			7547: out = 24'(23420);
			7548: out = 24'(18512);
			7549: out = 24'(-10820);
			7550: out = 24'(-25812);
			7551: out = 24'(-8044);
			7552: out = 24'(22028);
			7553: out = 24'(18980);
			7554: out = 24'(-11300);
			7555: out = 24'(-6828);
			7556: out = 24'(6448);
			7557: out = 24'(9368);
			7558: out = 24'(6908);
			7559: out = 24'(68);
			7560: out = 24'(-13252);
			7561: out = 24'(-22272);
			7562: out = 24'(-25444);
			7563: out = 24'(796);
			7564: out = 24'(27080);
			7565: out = 24'(8576);
			7566: out = 24'(-24000);
			7567: out = 24'(-4924);
			7568: out = 24'(9316);
			7569: out = 24'(2900);
			7570: out = 24'(1620);
			7571: out = 24'(-1060);
			7572: out = 24'(-13404);
			7573: out = 24'(-7052);
			7574: out = 24'(-1116);
			7575: out = 24'(-12636);
			7576: out = 24'(7876);
			7577: out = 24'(11604);
			7578: out = 24'(14148);
			7579: out = 24'(1536);
			7580: out = 24'(-16680);
			7581: out = 24'(1392);
			7582: out = 24'(23104);
			7583: out = 24'(25656);
			7584: out = 24'(5104);
			7585: out = 24'(-20824);
			7586: out = 24'(-17944);
			7587: out = 24'(-11332);
			7588: out = 24'(-2248);
			7589: out = 24'(7172);
			7590: out = 24'(11304);
			7591: out = 24'(-8604);
			7592: out = 24'(-12852);
			7593: out = 24'(11656);
			7594: out = 24'(7352);
			7595: out = 24'(13864);
			7596: out = 24'(16816);
			7597: out = 24'(20948);
			7598: out = 24'(5436);
			7599: out = 24'(-14176);
			7600: out = 24'(-19024);
			7601: out = 24'(-3940);
			7602: out = 24'(9536);
			7603: out = 24'(-4524);
			7604: out = 24'(-15108);
			7605: out = 24'(-4156);
			7606: out = 24'(4688);
			7607: out = 24'(4984);
			7608: out = 24'(-2972);
			7609: out = 24'(6972);
			7610: out = 24'(9728);
			7611: out = 24'(11116);
			7612: out = 24'(3124);
			7613: out = 24'(-10192);
			7614: out = 24'(-18492);
			7615: out = 24'(-14880);
			7616: out = 24'(1524);
			7617: out = 24'(-4084);
			7618: out = 24'(-12056);
			7619: out = 24'(60);
			7620: out = 24'(11964);
			7621: out = 24'(13916);
			7622: out = 24'(-5808);
			7623: out = 24'(-14852);
			7624: out = 24'(-4132);
			7625: out = 24'(8208);
			7626: out = 24'(5272);
			7627: out = 24'(-412);
			7628: out = 24'(8872);
			7629: out = 24'(8124);
			7630: out = 24'(-1568);
			7631: out = 24'(5136);
			7632: out = 24'(1508);
			7633: out = 24'(-6800);
			7634: out = 24'(-8652);
			7635: out = 24'(4756);
			7636: out = 24'(14028);
			7637: out = 24'(-8444);
			7638: out = 24'(-14488);
			7639: out = 24'(-6760);
			7640: out = 24'(-2132);
			7641: out = 24'(6936);
			7642: out = 24'(3792);
			7643: out = 24'(-10784);
			7644: out = 24'(-11424);
			7645: out = 24'(3956);
			7646: out = 24'(-5840);
			7647: out = 24'(-18112);
			7648: out = 24'(-11608);
			7649: out = 24'(2944);
			7650: out = 24'(1084);
			7651: out = 24'(-1244);
			7652: out = 24'(8668);
			7653: out = 24'(23904);
			7654: out = 24'(11880);
			7655: out = 24'(-21128);
			7656: out = 24'(-39132);
			7657: out = 24'(-19548);
			7658: out = 24'(12348);
			7659: out = 24'(6136);
			7660: out = 24'(-5788);
			7661: out = 24'(3804);
			7662: out = 24'(16248);
			7663: out = 24'(24424);
			7664: out = 24'(-3880);
			7665: out = 24'(-19000);
			7666: out = 24'(-3748);
			7667: out = 24'(12016);
			7668: out = 24'(16996);
			7669: out = 24'(17892);
			7670: out = 24'(15048);
			7671: out = 24'(-1396);
			7672: out = 24'(-28484);
			7673: out = 24'(-35620);
			7674: out = 24'(-18764);
			7675: out = 24'(-1436);
			7676: out = 24'(11124);
			7677: out = 24'(9992);
			7678: out = 24'(-7560);
			7679: out = 24'(-8900);
			7680: out = 24'(12728);
			7681: out = 24'(27516);
			7682: out = 24'(24556);
			7683: out = 24'(-7712);
			7684: out = 24'(-19300);
			7685: out = 24'(-5772);
			7686: out = 24'(-4424);
			7687: out = 24'(11488);
			7688: out = 24'(16504);
			7689: out = 24'(3840);
			7690: out = 24'(-4876);
			7691: out = 24'(-1928);
			7692: out = 24'(1980);
			7693: out = 24'(-5480);
			7694: out = 24'(-1672);
			7695: out = 24'(5520);
			7696: out = 24'(17484);
			7697: out = 24'(26708);
			7698: out = 24'(4484);
			7699: out = 24'(-13968);
			7700: out = 24'(-16536);
			7701: out = 24'(-11620);
			7702: out = 24'(-3260);
			7703: out = 24'(7840);
			7704: out = 24'(13952);
			7705: out = 24'(-1208);
			7706: out = 24'(-21008);
			7707: out = 24'(-11184);
			7708: out = 24'(-112);
			7709: out = 24'(15296);
			7710: out = 24'(4060);
			7711: out = 24'(-9792);
			7712: out = 24'(-9640);
			7713: out = 24'(2068);
			7714: out = 24'(13604);
			7715: out = 24'(22176);
			7716: out = 24'(6708);
			7717: out = 24'(-12480);
			7718: out = 24'(-7864);
			7719: out = 24'(-4352);
			7720: out = 24'(1740);
			7721: out = 24'(9832);
			7722: out = 24'(7360);
			7723: out = 24'(-480);
			7724: out = 24'(-12040);
			7725: out = 24'(-8300);
			7726: out = 24'(-9080);
			7727: out = 24'(-10292);
			7728: out = 24'(2396);
			7729: out = 24'(19544);
			7730: out = 24'(9420);
			7731: out = 24'(-2536);
			7732: out = 24'(-3944);
			7733: out = 24'(10384);
			7734: out = 24'(14480);
			7735: out = 24'(2716);
			7736: out = 24'(8316);
			7737: out = 24'(5064);
			7738: out = 24'(-7368);
			7739: out = 24'(-15308);
			7740: out = 24'(-4380);
			7741: out = 24'(396);
			7742: out = 24'(-1408);
			7743: out = 24'(-2292);
			7744: out = 24'(-8160);
			7745: out = 24'(-27404);
			7746: out = 24'(-17712);
			7747: out = 24'(3960);
			7748: out = 24'(11752);
			7749: out = 24'(5904);
			7750: out = 24'(6028);
			7751: out = 24'(7068);
			7752: out = 24'(-5432);
			7753: out = 24'(3016);
			7754: out = 24'(-5648);
			7755: out = 24'(12256);
			7756: out = 24'(23704);
			7757: out = 24'(12988);
			7758: out = 24'(8660);
			7759: out = 24'(3632);
			7760: out = 24'(-656);
			7761: out = 24'(-5100);
			7762: out = 24'(-19124);
			7763: out = 24'(-13572);
			7764: out = 24'(9376);
			7765: out = 24'(8820);
			7766: out = 24'(-9412);
			7767: out = 24'(-4152);
			7768: out = 24'(712);
			7769: out = 24'(3172);
			7770: out = 24'(3600);
			7771: out = 24'(1224);
			7772: out = 24'(8844);
			7773: out = 24'(7532);
			7774: out = 24'(7084);
			7775: out = 24'(-5572);
			7776: out = 24'(-17744);
			7777: out = 24'(-14312);
			7778: out = 24'(-7400);
			7779: out = 24'(2656);
			7780: out = 24'(10592);
			7781: out = 24'(9884);
			7782: out = 24'(6724);
			7783: out = 24'(-5908);
			7784: out = 24'(3724);
			7785: out = 24'(11516);
			7786: out = 24'(-2360);
			7787: out = 24'(2768);
			7788: out = 24'(12200);
			7789: out = 24'(-5284);
			7790: out = 24'(-18692);
			7791: out = 24'(-6048);
			7792: out = 24'(4900);
			7793: out = 24'(-220);
			7794: out = 24'(-21188);
			7795: out = 24'(-18380);
			7796: out = 24'(760);
			7797: out = 24'(8776);
			7798: out = 24'(9908);
			7799: out = 24'(-10684);
			7800: out = 24'(-27500);
			7801: out = 24'(-1668);
			7802: out = 24'(14288);
			7803: out = 24'(16868);
			7804: out = 24'(6604);
			7805: out = 24'(-17524);
			7806: out = 24'(-5788);
			7807: out = 24'(664);
			7808: out = 24'(9136);
			7809: out = 24'(19512);
			7810: out = 24'(13148);
			7811: out = 24'(4304);
			7812: out = 24'(-13464);
			7813: out = 24'(-26924);
			7814: out = 24'(-22300);
			7815: out = 24'(-4648);
			7816: out = 24'(18440);
			7817: out = 24'(24488);
			7818: out = 24'(13404);
			7819: out = 24'(-4532);
			7820: out = 24'(-10776);
			7821: out = 24'(-356);
			7822: out = 24'(11552);
			7823: out = 24'(11564);
			7824: out = 24'(-7784);
			7825: out = 24'(-1876);
			7826: out = 24'(15784);
			7827: out = 24'(22680);
			7828: out = 24'(-3572);
			7829: out = 24'(-16252);
			7830: out = 24'(-16056);
			7831: out = 24'(-5084);
			7832: out = 24'(-4960);
			7833: out = 24'(1040);
			7834: out = 24'(-96);
			7835: out = 24'(-4984);
			7836: out = 24'(272);
			7837: out = 24'(15312);
			7838: out = 24'(31104);
			7839: out = 24'(9340);
			7840: out = 24'(-14564);
			7841: out = 24'(-18460);
			7842: out = 24'(-3260);
			7843: out = 24'(2460);
			7844: out = 24'(-18316);
			7845: out = 24'(-7612);
			7846: out = 24'(14720);
			7847: out = 24'(12540);
			7848: out = 24'(-6780);
			7849: out = 24'(-13496);
			7850: out = 24'(288);
			7851: out = 24'(4188);
			7852: out = 24'(11324);
			7853: out = 24'(21240);
			7854: out = 24'(3280);
			7855: out = 24'(-28612);
			7856: out = 24'(-36468);
			7857: out = 24'(-27208);
			7858: out = 24'(-2560);
			7859: out = 24'(24436);
			7860: out = 24'(916);
			7861: out = 24'(-13912);
			7862: out = 24'(5180);
			7863: out = 24'(25356);
			7864: out = 24'(18112);
			7865: out = 24'(-15016);
			7866: out = 24'(-21612);
			7867: out = 24'(-6984);
			7868: out = 24'(18388);
			7869: out = 24'(29188);
			7870: out = 24'(-4408);
			7871: out = 24'(-21332);
			7872: out = 24'(-6972);
			7873: out = 24'(-948);
			7874: out = 24'(13072);
			7875: out = 24'(8352);
			7876: out = 24'(-944);
			7877: out = 24'(-4240);
			7878: out = 24'(-3024);
			7879: out = 24'(-3660);
			7880: out = 24'(-2524);
			7881: out = 24'(-4408);
			7882: out = 24'(9588);
			7883: out = 24'(8096);
			7884: out = 24'(-568);
			7885: out = 24'(1976);
			7886: out = 24'(-1592);
			7887: out = 24'(-13740);
			7888: out = 24'(-23008);
			7889: out = 24'(-13924);
			7890: out = 24'(15264);
			7891: out = 24'(20428);
			7892: out = 24'(2904);
			7893: out = 24'(-5588);
			7894: out = 24'(-4692);
			7895: out = 24'(10068);
			7896: out = 24'(23080);
			7897: out = 24'(18208);
			7898: out = 24'(-2828);
			7899: out = 24'(-14816);
			7900: out = 24'(-6092);
			7901: out = 24'(-4332);
			7902: out = 24'(-3852);
			7903: out = 24'(-6252);
			7904: out = 24'(1616);
			7905: out = 24'(8584);
			7906: out = 24'(-732);
			7907: out = 24'(-8620);
			7908: out = 24'(-4292);
			7909: out = 24'(820);
			7910: out = 24'(-7612);
			7911: out = 24'(5640);
			7912: out = 24'(744);
			7913: out = 24'(-2192);
			7914: out = 24'(2188);
			7915: out = 24'(1648);
			7916: out = 24'(1768);
			7917: out = 24'(-1860);
			7918: out = 24'(3464);
			7919: out = 24'(16600);
			7920: out = 24'(20176);
			7921: out = 24'(2592);
			7922: out = 24'(-18672);
			7923: out = 24'(-21400);
			7924: out = 24'(840);
			7925: out = 24'(12584);
			7926: out = 24'(4216);
			7927: out = 24'(-13784);
			7928: out = 24'(-10356);
			7929: out = 24'(3136);
			7930: out = 24'(12748);
			7931: out = 24'(-10788);
			7932: out = 24'(-13468);
			7933: out = 24'(1784);
			7934: out = 24'(12120);
			7935: out = 24'(16376);
			7936: out = 24'(1968);
			7937: out = 24'(-980);
			7938: out = 24'(-2344);
			7939: out = 24'(-4192);
			7940: out = 24'(1984);
			7941: out = 24'(1460);
			7942: out = 24'(10456);
			7943: out = 24'(13796);
			7944: out = 24'(5132);
			7945: out = 24'(-3016);
			7946: out = 24'(-7652);
			7947: out = 24'(1324);
			7948: out = 24'(12308);
			7949: out = 24'(4888);
			7950: out = 24'(-13508);
			7951: out = 24'(-7352);
			7952: out = 24'(-4464);
			7953: out = 24'(-4176);
			7954: out = 24'(-14560);
			7955: out = 24'(-7532);
			7956: out = 24'(1664);
			7957: out = 24'(-2032);
			7958: out = 24'(9972);
			7959: out = 24'(9348);
			7960: out = 24'(3616);
			7961: out = 24'(-14132);
			7962: out = 24'(-9312);
			7963: out = 24'(-10880);
			7964: out = 24'(1656);
			7965: out = 24'(8752);
			7966: out = 24'(-1080);
			7967: out = 24'(-13320);
			7968: out = 24'(-968);
			7969: out = 24'(14504);
			7970: out = 24'(4000);
			7971: out = 24'(-14536);
			7972: out = 24'(-12412);
			7973: out = 24'(10308);
			7974: out = 24'(-3332);
			7975: out = 24'(-6264);
			7976: out = 24'(16640);
			7977: out = 24'(11356);
			7978: out = 24'(-10624);
			7979: out = 24'(-5600);
			7980: out = 24'(512);
			7981: out = 24'(-2632);
			7982: out = 24'(-7952);
			7983: out = 24'(-5152);
			7984: out = 24'(-4440);
			7985: out = 24'(2680);
			7986: out = 24'(5000);
			7987: out = 24'(-11428);
			7988: out = 24'(-5644);
			7989: out = 24'(-472);
			7990: out = 24'(4372);
			7991: out = 24'(19088);
			7992: out = 24'(10312);
			7993: out = 24'(-1644);
			7994: out = 24'(-7240);
			7995: out = 24'(-4488);
			7996: out = 24'(184);
			7997: out = 24'(-1044);
			7998: out = 24'(2896);
			7999: out = 24'(9176);
			8000: out = 24'(7724);
			8001: out = 24'(4948);
			8002: out = 24'(-5668);
			8003: out = 24'(-13548);
			8004: out = 24'(-25020);
			8005: out = 24'(-15712);
			8006: out = 24'(12672);
			8007: out = 24'(23028);
			8008: out = 24'(92);
			8009: out = 24'(-9760);
			8010: out = 24'(652);
			8011: out = 24'(7032);
			8012: out = 24'(3604);
			8013: out = 24'(-5172);
			8014: out = 24'(-17940);
			8015: out = 24'(-12248);
			8016: out = 24'(10380);
			8017: out = 24'(12964);
			8018: out = 24'(1592);
			8019: out = 24'(-10684);
			8020: out = 24'(-760);
			8021: out = 24'(22344);
			8022: out = 24'(23884);
			8023: out = 24'(2292);
			8024: out = 24'(-23196);
			8025: out = 24'(-20336);
			8026: out = 24'(-13340);
			8027: out = 24'(5508);
			8028: out = 24'(16724);
			8029: out = 24'(360);
			8030: out = 24'(-23460);
			8031: out = 24'(-14772);
			8032: out = 24'(-680);
			8033: out = 24'(6644);
			8034: out = 24'(16028);
			8035: out = 24'(5596);
			8036: out = 24'(-12236);
			8037: out = 24'(-7196);
			8038: out = 24'(-3892);
			8039: out = 24'(-4200);
			8040: out = 24'(860);
			8041: out = 24'(-3228);
			8042: out = 24'(4848);
			8043: out = 24'(9908);
			8044: out = 24'(7316);
			8045: out = 24'(2512);
			8046: out = 24'(6996);
			8047: out = 24'(-2248);
			8048: out = 24'(-11132);
			8049: out = 24'(-7816);
			8050: out = 24'(-9116);
			8051: out = 24'(15520);
			8052: out = 24'(28532);
			8053: out = 24'(4016);
			8054: out = 24'(-15544);
			8055: out = 24'(-17312);
			8056: out = 24'(-1136);
			8057: out = 24'(21968);
			8058: out = 24'(18308);
			8059: out = 24'(-6676);
			8060: out = 24'(-23932);
			8061: out = 24'(-16368);
			8062: out = 24'(14284);
			8063: out = 24'(23628);
			8064: out = 24'(6932);
			8065: out = 24'(-15012);
			8066: out = 24'(-10552);
			8067: out = 24'(-14868);
			8068: out = 24'(-9384);
			8069: out = 24'(5284);
			8070: out = 24'(10140);
			8071: out = 24'(14220);
			8072: out = 24'(5348);
			8073: out = 24'(-10444);
			8074: out = 24'(-6140);
			8075: out = 24'(10384);
			8076: out = 24'(12860);
			8077: out = 24'(6196);
			8078: out = 24'(-10824);
			8079: out = 24'(-18672);
			8080: out = 24'(-3240);
			8081: out = 24'(10800);
			8082: out = 24'(11672);
			8083: out = 24'(5384);
			8084: out = 24'(4660);
			8085: out = 24'(5156);
			8086: out = 24'(2120);
			8087: out = 24'(-4584);
			8088: out = 24'(-14524);
			8089: out = 24'(-10288);
			8090: out = 24'(14028);
			8091: out = 24'(10504);
			8092: out = 24'(-8840);
			8093: out = 24'(-4968);
			8094: out = 24'(13140);
			8095: out = 24'(24252);
			8096: out = 24'(5284);
			8097: out = 24'(-12684);
			8098: out = 24'(-7900);
			8099: out = 24'(3384);
			8100: out = 24'(11296);
			8101: out = 24'(2396);
			8102: out = 24'(-8652);
			8103: out = 24'(-3820);
			8104: out = 24'(9428);
			8105: out = 24'(6380);
			8106: out = 24'(9084);
			8107: out = 24'(9968);
			8108: out = 24'(7592);
			8109: out = 24'(-6336);
			8110: out = 24'(-13380);
			8111: out = 24'(-11312);
			8112: out = 24'(-14408);
			8113: out = 24'(-19836);
			8114: out = 24'(1524);
			8115: out = 24'(7408);
			8116: out = 24'(816);
			8117: out = 24'(-1328);
			8118: out = 24'(15244);
			8119: out = 24'(18920);
			8120: out = 24'(-8160);
			8121: out = 24'(-23736);
			8122: out = 24'(-14592);
			8123: out = 24'(-4076);
			8124: out = 24'(-2212);
			8125: out = 24'(2372);
			8126: out = 24'(-656);
			8127: out = 24'(-6748);
			8128: out = 24'(512);
			8129: out = 24'(-2076);
			8130: out = 24'(-8836);
			8131: out = 24'(7004);
			8132: out = 24'(18332);
			8133: out = 24'(13048);
			8134: out = 24'(-2280);
			8135: out = 24'(-7844);
			8136: out = 24'(1024);
			8137: out = 24'(4148);
			8138: out = 24'(-3904);
			8139: out = 24'(-8892);
			8140: out = 24'(-7076);
			8141: out = 24'(-2532);
			8142: out = 24'(11880);
			8143: out = 24'(14176);
			8144: out = 24'(-17832);
			8145: out = 24'(-28556);
			8146: out = 24'(-4204);
			8147: out = 24'(18000);
			8148: out = 24'(18392);
			8149: out = 24'(5180);
			8150: out = 24'(-1956);
			8151: out = 24'(-372);
			8152: out = 24'(12740);
			8153: out = 24'(13600);
			8154: out = 24'(2248);
			8155: out = 24'(-388);
			8156: out = 24'(-3124);
			8157: out = 24'(-2288);
			8158: out = 24'(668);
			8159: out = 24'(5056);
			8160: out = 24'(8908);
			8161: out = 24'(-672);
			8162: out = 24'(-11492);
			8163: out = 24'(-8272);
			8164: out = 24'(-9164);
			8165: out = 24'(-5304);
			8166: out = 24'(3460);
			8167: out = 24'(5368);
			8168: out = 24'(-3452);
			8169: out = 24'(4072);
			8170: out = 24'(12248);
			8171: out = 24'(-2476);
			8172: out = 24'(-13124);
			8173: out = 24'(-9092);
			8174: out = 24'(1420);
			8175: out = 24'(2296);
			8176: out = 24'(2888);
			8177: out = 24'(8112);
			8178: out = 24'(5392);
			8179: out = 24'(1912);
			8180: out = 24'(-8500);
			8181: out = 24'(-8464);
			8182: out = 24'(12260);
			8183: out = 24'(13404);
			8184: out = 24'(-3672);
			8185: out = 24'(-7540);
			8186: out = 24'(-1260);
			8187: out = 24'(1428);
			8188: out = 24'(8248);
			8189: out = 24'(16972);
			8190: out = 24'(4864);
			8191: out = 24'(-12496);
			8192: out = 24'(-13580);
			8193: out = 24'(-17528);
			8194: out = 24'(5940);
			8195: out = 24'(28564);
			8196: out = 24'(9960);
			8197: out = 24'(-9652);
			8198: out = 24'(-4000);
			8199: out = 24'(7024);
			8200: out = 24'(12172);
			8201: out = 24'(1296);
			8202: out = 24'(1884);
			8203: out = 24'(6972);
			8204: out = 24'(7476);
			8205: out = 24'(12904);
			8206: out = 24'(10700);
			8207: out = 24'(-5920);
			8208: out = 24'(-21776);
			8209: out = 24'(-22696);
			8210: out = 24'(-6588);
			8211: out = 24'(12596);
			8212: out = 24'(-4288);
			8213: out = 24'(-21812);
			8214: out = 24'(-10180);
			8215: out = 24'(6928);
			8216: out = 24'(6052);
			8217: out = 24'(1216);
			8218: out = 24'(-12);
			8219: out = 24'(-15580);
			8220: out = 24'(-14000);
			8221: out = 24'(-1408);
			8222: out = 24'(12400);
			8223: out = 24'(18096);
			8224: out = 24'(-320);
			8225: out = 24'(-21216);
			8226: out = 24'(-21280);
			8227: out = 24'(1196);
			8228: out = 24'(12880);
			8229: out = 24'(-11960);
			8230: out = 24'(-6984);
			8231: out = 24'(13072);
			8232: out = 24'(11212);
			8233: out = 24'(3960);
			8234: out = 24'(-536);
			8235: out = 24'(156);
			8236: out = 24'(4220);
			8237: out = 24'(1248);
			8238: out = 24'(-9976);
			8239: out = 24'(-7396);
			8240: out = 24'(12588);
			8241: out = 24'(20864);
			8242: out = 24'(2216);
			8243: out = 24'(-21396);
			8244: out = 24'(-12624);
			8245: out = 24'(6836);
			8246: out = 24'(15516);
			8247: out = 24'(-608);
			8248: out = 24'(-13292);
			8249: out = 24'(-4364);
			8250: out = 24'(-7072);
			8251: out = 24'(5244);
			8252: out = 24'(18264);
			8253: out = 24'(-1332);
			8254: out = 24'(-8468);
			8255: out = 24'(-2488);
			8256: out = 24'(-1792);
			8257: out = 24'(-12640);
			8258: out = 24'(-12584);
			8259: out = 24'(-4104);
			8260: out = 24'(11296);
			8261: out = 24'(27028);
			8262: out = 24'(18916);
			8263: out = 24'(-9036);
			8264: out = 24'(-18112);
			8265: out = 24'(-6124);
			8266: out = 24'(1216);
			8267: out = 24'(8920);
			8268: out = 24'(14804);
			8269: out = 24'(5432);
			8270: out = 24'(-15248);
			8271: out = 24'(-13256);
			8272: out = 24'(4408);
			8273: out = 24'(10180);
			8274: out = 24'(9888);
			8275: out = 24'(-9140);
			8276: out = 24'(-24400);
			8277: out = 24'(-8536);
			8278: out = 24'(8216);
			8279: out = 24'(13596);
			8280: out = 24'(-4136);
			8281: out = 24'(-6248);
			8282: out = 24'(7384);
			8283: out = 24'(4228);
			8284: out = 24'(532);
			8285: out = 24'(2856);
			8286: out = 24'(-2236);
			8287: out = 24'(-4848);
			8288: out = 24'(-1236);
			8289: out = 24'(136);
			8290: out = 24'(1828);
			8291: out = 24'(-10084);
			8292: out = 24'(-8192);
			8293: out = 24'(9780);
			8294: out = 24'(5796);
			8295: out = 24'(-2176);
			8296: out = 24'(5624);
			8297: out = 24'(4052);
			8298: out = 24'(-22512);
			8299: out = 24'(-32212);
			8300: out = 24'(-12324);
			8301: out = 24'(2764);
			8302: out = 24'(21540);
			8303: out = 24'(20752);
			8304: out = 24'(-2488);
			8305: out = 24'(-12140);
			8306: out = 24'(-4748);
			8307: out = 24'(15508);
			8308: out = 24'(22448);
			8309: out = 24'(8868);
			8310: out = 24'(-4516);
			8311: out = 24'(-2600);
			8312: out = 24'(-752);
			8313: out = 24'(-1944);
			8314: out = 24'(-13340);
			8315: out = 24'(-11724);
			8316: out = 24'(-1840);
			8317: out = 24'(3024);
			8318: out = 24'(8988);
			8319: out = 24'(6112);
			8320: out = 24'(-8612);
			8321: out = 24'(-7000);
			8322: out = 24'(1424);
			8323: out = 24'(-11448);
			8324: out = 24'(-11564);
			8325: out = 24'(-4988);
			8326: out = 24'(-292);
			8327: out = 24'(12944);
			8328: out = 24'(11620);
			8329: out = 24'(10416);
			8330: out = 24'(5532);
			8331: out = 24'(-4096);
			8332: out = 24'(-14104);
			8333: out = 24'(-8460);
			8334: out = 24'(1596);
			8335: out = 24'(6076);
			8336: out = 24'(11540);
			8337: out = 24'(2824);
			8338: out = 24'(7288);
			8339: out = 24'(7324);
			8340: out = 24'(-4884);
			8341: out = 24'(-2416);
			8342: out = 24'(2660);
			8343: out = 24'(7784);
			8344: out = 24'(9992);
			8345: out = 24'(1872);
			8346: out = 24'(-4204);
			8347: out = 24'(-4740);
			8348: out = 24'(-7960);
			8349: out = 24'(-8160);
			8350: out = 24'(-9532);
			8351: out = 24'(-7808);
			8352: out = 24'(-10352);
			8353: out = 24'(-10132);
			8354: out = 24'(6652);
			8355: out = 24'(15284);
			8356: out = 24'(5596);
			8357: out = 24'(-6532);
			8358: out = 24'(-5448);
			8359: out = 24'(-896);
			8360: out = 24'(1276);
			8361: out = 24'(3340);
			8362: out = 24'(9144);
			8363: out = 24'(2764);
			8364: out = 24'(1376);
			8365: out = 24'(-2164);
			8366: out = 24'(-3900);
			8367: out = 24'(-4988);
			8368: out = 24'(-6164);
			8369: out = 24'(-984);
			8370: out = 24'(4992);
			8371: out = 24'(13812);
			8372: out = 24'(1444);
			8373: out = 24'(-7844);
			8374: out = 24'(-14092);
			8375: out = 24'(-6044);
			8376: out = 24'(6032);
			8377: out = 24'(12676);
			8378: out = 24'(5932);
			8379: out = 24'(2936);
			8380: out = 24'(7144);
			8381: out = 24'(4572);
			8382: out = 24'(-3932);
			8383: out = 24'(-4972);
			8384: out = 24'(-9948);
			8385: out = 24'(-11976);
			8386: out = 24'(-1008);
			8387: out = 24'(14116);
			8388: out = 24'(3280);
			8389: out = 24'(-6788);
			8390: out = 24'(-2876);
			8391: out = 24'(-2340);
			8392: out = 24'(-12440);
			8393: out = 24'(-17976);
			8394: out = 24'(8564);
			8395: out = 24'(4480);
			8396: out = 24'(2612);
			8397: out = 24'(20220);
			8398: out = 24'(14124);
			8399: out = 24'(-2000);
			8400: out = 24'(-18580);
			8401: out = 24'(-8736);
			8402: out = 24'(15700);
			8403: out = 24'(19948);
			8404: out = 24'(724);
			8405: out = 24'(-13652);
			8406: out = 24'(-13900);
			8407: out = 24'(-5624);
			8408: out = 24'(820);
			8409: out = 24'(-1124);
			8410: out = 24'(-4228);
			8411: out = 24'(-160);
			8412: out = 24'(-4172);
			8413: out = 24'(-1356);
			8414: out = 24'(3484);
			8415: out = 24'(7412);
			8416: out = 24'(10172);
			8417: out = 24'(-4764);
			8418: out = 24'(-6096);
			8419: out = 24'(-3164);
			8420: out = 24'(6292);
			8421: out = 24'(2648);
			8422: out = 24'(-5444);
			8423: out = 24'(5948);
			8424: out = 24'(-268);
			8425: out = 24'(5364);
			8426: out = 24'(8504);
			8427: out = 24'(5560);
			8428: out = 24'(-508);
			8429: out = 24'(324);
			8430: out = 24'(-6040);
			8431: out = 24'(1852);
			8432: out = 24'(8876);
			8433: out = 24'(3500);
			8434: out = 24'(-2044);
			8435: out = 24'(-7008);
			8436: out = 24'(-2428);
			8437: out = 24'(-3396);
			8438: out = 24'(2856);
			8439: out = 24'(8964);
			8440: out = 24'(-7396);
			8441: out = 24'(-13868);
			8442: out = 24'(-1468);
			8443: out = 24'(16116);
			8444: out = 24'(-3428);
			8445: out = 24'(-19572);
			8446: out = 24'(-680);
			8447: out = 24'(15624);
			8448: out = 24'(13040);
			8449: out = 24'(3168);
			8450: out = 24'(-2424);
			8451: out = 24'(-648);
			8452: out = 24'(-4744);
			8453: out = 24'(-15136);
			8454: out = 24'(-616);
			8455: out = 24'(11420);
			8456: out = 24'(508);
			8457: out = 24'(-8704);
			8458: out = 24'(-6284);
			8459: out = 24'(-2540);
			8460: out = 24'(-880);
			8461: out = 24'(3860);
			8462: out = 24'(6556);
			8463: out = 24'(7236);
			8464: out = 24'(8852);
			8465: out = 24'(-2744);
			8466: out = 24'(-10380);
			8467: out = 24'(-9996);
			8468: out = 24'(-5828);
			8469: out = 24'(7152);
			8470: out = 24'(10412);
			8471: out = 24'(7600);
			8472: out = 24'(9536);
			8473: out = 24'(8768);
			8474: out = 24'(-11332);
			8475: out = 24'(-16408);
			8476: out = 24'(-19412);
			8477: out = 24'(2540);
			8478: out = 24'(23924);
			8479: out = 24'(14264);
			8480: out = 24'(-10340);
			8481: out = 24'(-7268);
			8482: out = 24'(-12);
			8483: out = 24'(6072);
			8484: out = 24'(7588);
			8485: out = 24'(-1792);
			8486: out = 24'(-6996);
			8487: out = 24'(-4460);
			8488: out = 24'(-5128);
			8489: out = 24'(-7580);
			8490: out = 24'(2356);
			8491: out = 24'(1776);
			8492: out = 24'(3228);
			8493: out = 24'(9492);
			8494: out = 24'(12384);
			8495: out = 24'(-1252);
			8496: out = 24'(-8904);
			8497: out = 24'(-5040);
			8498: out = 24'(2084);
			8499: out = 24'(7744);
			8500: out = 24'(924);
			8501: out = 24'(-12164);
			8502: out = 24'(2160);
			8503: out = 24'(8668);
			8504: out = 24'(2720);
			8505: out = 24'(-8516);
			8506: out = 24'(-4608);
			8507: out = 24'(-1336);
			8508: out = 24'(1088);
			8509: out = 24'(10512);
			8510: out = 24'(16016);
			8511: out = 24'(5308);
			8512: out = 24'(-11852);
			8513: out = 24'(-1240);
			8514: out = 24'(5900);
			8515: out = 24'(3512);
			8516: out = 24'(-8116);
			8517: out = 24'(-15144);
			8518: out = 24'(-5148);
			8519: out = 24'(4368);
			8520: out = 24'(4);
			8521: out = 24'(-3988);
			8522: out = 24'(2432);
			8523: out = 24'(2316);
			8524: out = 24'(1336);
			8525: out = 24'(1860);
			8526: out = 24'(10580);
			8527: out = 24'(4148);
			8528: out = 24'(-11204);
			8529: out = 24'(-1104);
			8530: out = 24'(7292);
			8531: out = 24'(6692);
			8532: out = 24'(-904);
			8533: out = 24'(-11608);
			8534: out = 24'(-14892);
			8535: out = 24'(-17260);
			8536: out = 24'(1512);
			8537: out = 24'(19156);
			8538: out = 24'(10784);
			8539: out = 24'(-9332);
			8540: out = 24'(-19336);
			8541: out = 24'(-13520);
			8542: out = 24'(-972);
			8543: out = 24'(18232);
			8544: out = 24'(8992);
			8545: out = 24'(-12844);
			8546: out = 24'(-5876);
			8547: out = 24'(2800);
			8548: out = 24'(9020);
			8549: out = 24'(7000);
			8550: out = 24'(-11800);
			8551: out = 24'(-4988);
			8552: out = 24'(14776);
			8553: out = 24'(14080);
			8554: out = 24'(-1524);
			8555: out = 24'(-16768);
			8556: out = 24'(-7072);
			8557: out = 24'(12388);
			8558: out = 24'(9108);
			8559: out = 24'(-6944);
			8560: out = 24'(-12276);
			8561: out = 24'(-2772);
			8562: out = 24'(9760);
			8563: out = 24'(12752);
			8564: out = 24'(2440);
			8565: out = 24'(28);
			8566: out = 24'(-344);
			8567: out = 24'(152);
			8568: out = 24'(2432);
			8569: out = 24'(-11400);
			8570: out = 24'(-10620);
			8571: out = 24'(3836);
			8572: out = 24'(9480);
			8573: out = 24'(948);
			8574: out = 24'(-8196);
			8575: out = 24'(-416);
			8576: out = 24'(18408);
			8577: out = 24'(7500);
			8578: out = 24'(-16852);
			8579: out = 24'(-17284);
			8580: out = 24'(-9392);
			8581: out = 24'(8456);
			8582: out = 24'(14112);
			8583: out = 24'(4368);
			8584: out = 24'(3632);
			8585: out = 24'(12904);
			8586: out = 24'(2872);
			8587: out = 24'(-15236);
			8588: out = 24'(-28456);
			8589: out = 24'(-11552);
			8590: out = 24'(4100);
			8591: out = 24'(2616);
			8592: out = 24'(11636);
			8593: out = 24'(11012);
			8594: out = 24'(2592);
			8595: out = 24'(-11612);
			8596: out = 24'(-8112);
			8597: out = 24'(-7452);
			8598: out = 24'(-1112);
			8599: out = 24'(15312);
			8600: out = 24'(15764);
			8601: out = 24'(2124);
			8602: out = 24'(-3596);
			8603: out = 24'(-1456);
			8604: out = 24'(8276);
			8605: out = 24'(1636);
			8606: out = 24'(-6704);
			8607: out = 24'(-1128);
			8608: out = 24'(-584);
			8609: out = 24'(-1640);
			8610: out = 24'(8348);
			8611: out = 24'(7548);
			8612: out = 24'(-10296);
			8613: out = 24'(-19844);
			8614: out = 24'(-5040);
			8615: out = 24'(9836);
			8616: out = 24'(1916);
			8617: out = 24'(-1512);
			8618: out = 24'(-4632);
			8619: out = 24'(-5196);
			8620: out = 24'(-2828);
			8621: out = 24'(-3392);
			8622: out = 24'(2516);
			8623: out = 24'(-288);
			8624: out = 24'(1140);
			8625: out = 24'(-1872);
			8626: out = 24'(-2536);
			8627: out = 24'(4788);
			8628: out = 24'(5992);
			8629: out = 24'(12728);
			8630: out = 24'(6512);
			8631: out = 24'(-15796);
			8632: out = 24'(-17012);
			8633: out = 24'(6248);
			8634: out = 24'(14216);
			8635: out = 24'(-360);
			8636: out = 24'(-25072);
			8637: out = 24'(-9752);
			8638: out = 24'(9964);
			8639: out = 24'(18264);
			8640: out = 24'(9148);
			8641: out = 24'(6268);
			8642: out = 24'(7152);
			8643: out = 24'(2324);
			8644: out = 24'(1660);
			8645: out = 24'(-3460);
			8646: out = 24'(-2748);
			8647: out = 24'(-3192);
			8648: out = 24'(-1792);
			8649: out = 24'(-7212);
			8650: out = 24'(-488);
			8651: out = 24'(-2448);
			8652: out = 24'(-4592);
			8653: out = 24'(-1676);
			8654: out = 24'(268);
			8655: out = 24'(-7336);
			8656: out = 24'(-8564);
			8657: out = 24'(6564);
			8658: out = 24'(7784);
			8659: out = 24'(14380);
			8660: out = 24'(9292);
			8661: out = 24'(4064);
			8662: out = 24'(-540);
			8663: out = 24'(-6176);
			8664: out = 24'(-13264);
			8665: out = 24'(-9872);
			8666: out = 24'(7236);
			8667: out = 24'(3448);
			8668: out = 24'(-1612);
			8669: out = 24'(8248);
			8670: out = 24'(5072);
			8671: out = 24'(-5888);
			8672: out = 24'(-11112);
			8673: out = 24'(-16616);
			8674: out = 24'(-2124);
			8675: out = 24'(13604);
			8676: out = 24'(17396);
			8677: out = 24'(-2388);
			8678: out = 24'(-14204);
			8679: out = 24'(-6772);
			8680: out = 24'(3744);
			8681: out = 24'(5688);
			8682: out = 24'(-3156);
			8683: out = 24'(-5148);
			8684: out = 24'(3884);
			8685: out = 24'(13360);
			8686: out = 24'(156);
			8687: out = 24'(-3852);
			8688: out = 24'(-7704);
			8689: out = 24'(3360);
			8690: out = 24'(2892);
			8691: out = 24'(176);
			8692: out = 24'(5784);
			8693: out = 24'(8416);
			8694: out = 24'(-2376);
			8695: out = 24'(-15896);
			8696: out = 24'(-13032);
			8697: out = 24'(1316);
			8698: out = 24'(5704);
			8699: out = 24'(5952);
			8700: out = 24'(11284);
			8701: out = 24'(8880);
			8702: out = 24'(-5184);
			8703: out = 24'(-17516);
			8704: out = 24'(-14076);
			8705: out = 24'(-17356);
			8706: out = 24'(-10024);
			8707: out = 24'(10348);
			8708: out = 24'(10408);
			8709: out = 24'(-2272);
			8710: out = 24'(-2132);
			8711: out = 24'(696);
			8712: out = 24'(6552);
			8713: out = 24'(20);
			8714: out = 24'(-5684);
			8715: out = 24'(-3792);
			8716: out = 24'(-2432);
			8717: out = 24'(3452);
			8718: out = 24'(8932);
			8719: out = 24'(1124);
			8720: out = 24'(-19264);
			8721: out = 24'(-15520);
			8722: out = 24'(-5308);
			8723: out = 24'(4044);
			8724: out = 24'(16604);
			8725: out = 24'(4608);
			8726: out = 24'(-2512);
			8727: out = 24'(6648);
			8728: out = 24'(9700);
			8729: out = 24'(9032);
			8730: out = 24'(672);
			8731: out = 24'(-13288);
			8732: out = 24'(-6064);
			8733: out = 24'(-7636);
			8734: out = 24'(-5496);
			8735: out = 24'(7440);
			8736: out = 24'(7440);
			8737: out = 24'(-264);
			8738: out = 24'(236);
			8739: out = 24'(12092);
			8740: out = 24'(580);
			8741: out = 24'(-18892);
			8742: out = 24'(-10404);
			8743: out = 24'(8780);
			8744: out = 24'(7488);
			8745: out = 24'(6128);
			8746: out = 24'(9756);
			8747: out = 24'(6276);
			8748: out = 24'(-8048);
			8749: out = 24'(-25192);
			8750: out = 24'(-19728);
			8751: out = 24'(5972);
			8752: out = 24'(15376);
			8753: out = 24'(-1808);
			8754: out = 24'(-6436);
			8755: out = 24'(-4220);
			8756: out = 24'(5004);
			8757: out = 24'(22324);
			8758: out = 24'(11756);
			8759: out = 24'(-6396);
			8760: out = 24'(-13772);
			8761: out = 24'(-8140);
			8762: out = 24'(-6040);
			8763: out = 24'(1824);
			8764: out = 24'(4900);
			8765: out = 24'(3152);
			8766: out = 24'(4376);
			8767: out = 24'(5828);
			8768: out = 24'(5460);
			8769: out = 24'(-568);
			8770: out = 24'(-556);
			8771: out = 24'(1208);
			8772: out = 24'(9216);
			8773: out = 24'(9692);
			8774: out = 24'(6128);
			8775: out = 24'(-1252);
			8776: out = 24'(-1876);
			8777: out = 24'(-7564);
			8778: out = 24'(-13584);
			8779: out = 24'(-7680);
			8780: out = 24'(-1728);
			8781: out = 24'(4);
			8782: out = 24'(7352);
			8783: out = 24'(852);
			8784: out = 24'(-10212);
			8785: out = 24'(-6892);
			8786: out = 24'(-5388);
			8787: out = 24'(4752);
			8788: out = 24'(5736);
			8789: out = 24'(4756);
			8790: out = 24'(3984);
			8791: out = 24'(8960);
			8792: out = 24'(6276);
			8793: out = 24'(-9904);
			8794: out = 24'(-15084);
			8795: out = 24'(-7504);
			8796: out = 24'(9256);
			8797: out = 24'(11800);
			8798: out = 24'(-1724);
			8799: out = 24'(-8004);
			8800: out = 24'(-5036);
			8801: out = 24'(-1396);
			8802: out = 24'(4600);
			8803: out = 24'(6076);
			8804: out = 24'(-672);
			8805: out = 24'(-20);
			8806: out = 24'(356);
			8807: out = 24'(-4396);
			8808: out = 24'(-10584);
			8809: out = 24'(-23040);
			8810: out = 24'(-4260);
			8811: out = 24'(14264);
			8812: out = 24'(13556);
			8813: out = 24'(8788);
			8814: out = 24'(5324);
			8815: out = 24'(-3760);
			8816: out = 24'(-8440);
			8817: out = 24'(-11316);
			8818: out = 24'(-12064);
			8819: out = 24'(-2512);
			8820: out = 24'(4500);
			8821: out = 24'(10464);
			8822: out = 24'(10288);
			8823: out = 24'(3352);
			8824: out = 24'(3832);
			8825: out = 24'(8632);
			8826: out = 24'(5960);
			8827: out = 24'(-2084);
			8828: out = 24'(-9188);
			8829: out = 24'(796);
			8830: out = 24'(15048);
			8831: out = 24'(11948);
			8832: out = 24'(-14044);
			8833: out = 24'(-13648);
			8834: out = 24'(692);
			8835: out = 24'(9252);
			8836: out = 24'(1024);
			8837: out = 24'(-6320);
			8838: out = 24'(6032);
			8839: out = 24'(12656);
			8840: out = 24'(7652);
			8841: out = 24'(1760);
			8842: out = 24'(280);
			8843: out = 24'(1596);
			8844: out = 24'(-3188);
			8845: out = 24'(-4228);
			8846: out = 24'(-184);
			8847: out = 24'(1860);
			8848: out = 24'(-8920);
			8849: out = 24'(-4220);
			8850: out = 24'(1104);
			8851: out = 24'(-7096);
			8852: out = 24'(-4684);
			8853: out = 24'(2332);
			8854: out = 24'(5016);
			8855: out = 24'(8040);
			8856: out = 24'(8576);
			8857: out = 24'(-2200);
			8858: out = 24'(-9692);
			8859: out = 24'(-10572);
			8860: out = 24'(-2388);
			8861: out = 24'(4460);
			8862: out = 24'(4188);
			8863: out = 24'(6700);
			8864: out = 24'(8488);
			8865: out = 24'(4040);
			8866: out = 24'(-6540);
			8867: out = 24'(-10732);
			8868: out = 24'(-3296);
			8869: out = 24'(-6196);
			8870: out = 24'(-2208);
			8871: out = 24'(11116);
			8872: out = 24'(10196);
			8873: out = 24'(-16316);
			8874: out = 24'(-28868);
			8875: out = 24'(-17140);
			8876: out = 24'(-1836);
			8877: out = 24'(20852);
			8878: out = 24'(19588);
			8879: out = 24'(-6236);
			8880: out = 24'(-24220);
			8881: out = 24'(-16608);
			8882: out = 24'(-1816);
			8883: out = 24'(9380);
			8884: out = 24'(16268);
			8885: out = 24'(6680);
			8886: out = 24'(-17820);
			8887: out = 24'(-22716);
			8888: out = 24'(-9884);
			8889: out = 24'(10664);
			8890: out = 24'(24852);
			8891: out = 24'(11092);
			8892: out = 24'(-4524);
			8893: out = 24'(-14504);
			8894: out = 24'(-1324);
			8895: out = 24'(15560);
			8896: out = 24'(14472);
			8897: out = 24'(5328);
			8898: out = 24'(-5100);
			8899: out = 24'(-10712);
			8900: out = 24'(-3776);
			8901: out = 24'(10584);
			8902: out = 24'(9064);
			8903: out = 24'(-2580);
			8904: out = 24'(2116);
			8905: out = 24'(1768);
			8906: out = 24'(-5588);
			8907: out = 24'(-8696);
			8908: out = 24'(-15424);
			8909: out = 24'(2584);
			8910: out = 24'(17960);
			8911: out = 24'(10368);
			8912: out = 24'(-4480);
			8913: out = 24'(-4416);
			8914: out = 24'(2652);
			8915: out = 24'(6896);
			8916: out = 24'(3476);
			8917: out = 24'(6144);
			8918: out = 24'(-2312);
			8919: out = 24'(-4276);
			8920: out = 24'(1584);
			8921: out = 24'(-1372);
			8922: out = 24'(-5376);
			8923: out = 24'(1188);
			8924: out = 24'(972);
			8925: out = 24'(1580);
			8926: out = 24'(6356);
			8927: out = 24'(8908);
			8928: out = 24'(5780);
			8929: out = 24'(-764);
			8930: out = 24'(-3996);
			8931: out = 24'(-880);
			8932: out = 24'(-6668);
			8933: out = 24'(-7068);
			8934: out = 24'(-8512);
			8935: out = 24'(-10952);
			8936: out = 24'(7772);
			8937: out = 24'(17924);
			8938: out = 24'(3392);
			8939: out = 24'(-9480);
			8940: out = 24'(-4424);
			8941: out = 24'(1868);
			8942: out = 24'(9404);
			8943: out = 24'(9852);
			8944: out = 24'(2276);
			8945: out = 24'(-412);
			8946: out = 24'(1228);
			8947: out = 24'(-264);
			8948: out = 24'(-2376);
			8949: out = 24'(-12120);
			8950: out = 24'(-10424);
			8951: out = 24'(3280);
			8952: out = 24'(10204);
			8953: out = 24'(-6352);
			8954: out = 24'(-15236);
			8955: out = 24'(-6496);
			8956: out = 24'(3184);
			8957: out = 24'(8748);
			8958: out = 24'(9548);
			8959: out = 24'(1440);
			8960: out = 24'(-10900);
			8961: out = 24'(-3256);
			8962: out = 24'(3544);
			8963: out = 24'(-260);
			8964: out = 24'(-7636);
			8965: out = 24'(-13528);
			8966: out = 24'(1036);
			8967: out = 24'(18092);
			8968: out = 24'(11964);
			8969: out = 24'(3180);
			8970: out = 24'(-892);
			8971: out = 24'(4668);
			8972: out = 24'(-1672);
			8973: out = 24'(-6792);
			8974: out = 24'(-3296);
			8975: out = 24'(9120);
			8976: out = 24'(11596);
			8977: out = 24'(-3332);
			8978: out = 24'(-5256);
			8979: out = 24'(-1984);
			8980: out = 24'(-3620);
			8981: out = 24'(2152);
			8982: out = 24'(5452);
			8983: out = 24'(-6648);
			8984: out = 24'(-2992);
			8985: out = 24'(-856);
			8986: out = 24'(3704);
			8987: out = 24'(13148);
			8988: out = 24'(6604);
			8989: out = 24'(-6308);
			8990: out = 24'(-6660);
			8991: out = 24'(-3584);
			8992: out = 24'(-8408);
			8993: out = 24'(-20436);
			8994: out = 24'(-2928);
			8995: out = 24'(8736);
			8996: out = 24'(10736);
			8997: out = 24'(8828);
			8998: out = 24'(7900);
			8999: out = 24'(6968);
			9000: out = 24'(1060);
			9001: out = 24'(-5156);
			9002: out = 24'(-8148);
			9003: out = 24'(-1296);
			9004: out = 24'(8760);
			9005: out = 24'(4100);
			9006: out = 24'(-11272);
			9007: out = 24'(-8664);
			9008: out = 24'(7528);
			9009: out = 24'(11764);
			9010: out = 24'(-8484);
			9011: out = 24'(-19748);
			9012: out = 24'(-11156);
			9013: out = 24'(-5016);
			9014: out = 24'(7768);
			9015: out = 24'(10860);
			9016: out = 24'(-184);
			9017: out = 24'(-7832);
			9018: out = 24'(428);
			9019: out = 24'(2088);
			9020: out = 24'(5668);
			9021: out = 24'(7076);
			9022: out = 24'(1584);
			9023: out = 24'(1516);
			9024: out = 24'(3616);
			9025: out = 24'(3016);
			9026: out = 24'(3240);
			9027: out = 24'(692);
			9028: out = 24'(5244);
			9029: out = 24'(-1232);
			9030: out = 24'(-7168);
			9031: out = 24'(-2512);
			9032: out = 24'(2428);
			9033: out = 24'(-8408);
			9034: out = 24'(-10740);
			9035: out = 24'(1512);
			9036: out = 24'(-2296);
			9037: out = 24'(784);
			9038: out = 24'(11868);
			9039: out = 24'(3260);
			9040: out = 24'(-18580);
			9041: out = 24'(-18688);
			9042: out = 24'(-5692);
			9043: out = 24'(9028);
			9044: out = 24'(14076);
			9045: out = 24'(-2300);
			9046: out = 24'(-22012);
			9047: out = 24'(-8088);
			9048: out = 24'(13248);
			9049: out = 24'(14532);
			9050: out = 24'(8204);
			9051: out = 24'(5404);
			9052: out = 24'(4328);
			9053: out = 24'(1988);
			9054: out = 24'(-7936);
			9055: out = 24'(-10568);
			9056: out = 24'(2388);
			9057: out = 24'(-972);
			9058: out = 24'(-3896);
			9059: out = 24'(-2148);
			9060: out = 24'(-3840);
			9061: out = 24'(3460);
			9062: out = 24'(4044);
			9063: out = 24'(-4548);
			9064: out = 24'(-3068);
			9065: out = 24'(1172);
			9066: out = 24'(8656);
			9067: out = 24'(7712);
			9068: out = 24'(2700);
			9069: out = 24'(2012);
			9070: out = 24'(-1660);
			9071: out = 24'(-12664);
			9072: out = 24'(-8144);
			9073: out = 24'(-1264);
			9074: out = 24'(4668);
			9075: out = 24'(7268);
			9076: out = 24'(-3168);
			9077: out = 24'(-13672);
			9078: out = 24'(-8348);
			9079: out = 24'(8860);
			9080: out = 24'(13792);
			9081: out = 24'(4052);
			9082: out = 24'(-4524);
			9083: out = 24'(-1416);
			9084: out = 24'(9428);
			9085: out = 24'(-3492);
			9086: out = 24'(-6856);
			9087: out = 24'(-1880);
			9088: out = 24'(-1064);
			9089: out = 24'(2756);
			9090: out = 24'(12184);
			9091: out = 24'(3964);
			9092: out = 24'(-7716);
			9093: out = 24'(-11836);
			9094: out = 24'(-932);
			9095: out = 24'(14168);
			9096: out = 24'(3448);
			9097: out = 24'(-9784);
			9098: out = 24'(-2252);
			9099: out = 24'(4216);
			9100: out = 24'(-5388);
			9101: out = 24'(-20800);
			9102: out = 24'(-12112);
			9103: out = 24'(-484);
			9104: out = 24'(316);
			9105: out = 24'(14608);
			9106: out = 24'(17452);
			9107: out = 24'(-1296);
			9108: out = 24'(-18388);
			9109: out = 24'(-13320);
			9110: out = 24'(1024);
			9111: out = 24'(3436);
			9112: out = 24'(-280);
			9113: out = 24'(5780);
			9114: out = 24'(-3300);
			9115: out = 24'(-5292);
			9116: out = 24'(2388);
			9117: out = 24'(6208);
			9118: out = 24'(11612);
			9119: out = 24'(7384);
			9120: out = 24'(-8948);
			9121: out = 24'(-15544);
			9122: out = 24'(-8312);
			9123: out = 24'(4004);
			9124: out = 24'(18228);
			9125: out = 24'(11848);
			9126: out = 24'(-5272);
			9127: out = 24'(-8948);
			9128: out = 24'(-2700);
			9129: out = 24'(4116);
			9130: out = 24'(-8996);
			9131: out = 24'(-2276);
			9132: out = 24'(9288);
			9133: out = 24'(8364);
			9134: out = 24'(-3128);
			9135: out = 24'(-4828);
			9136: out = 24'(6632);
			9137: out = 24'(8476);
			9138: out = 24'(4236);
			9139: out = 24'(-1896);
			9140: out = 24'(-3884);
			9141: out = 24'(-760);
			9142: out = 24'(-1964);
			9143: out = 24'(-3524);
			9144: out = 24'(3588);
			9145: out = 24'(10076);
			9146: out = 24'(-496);
			9147: out = 24'(-14608);
			9148: out = 24'(-10840);
			9149: out = 24'(-1416);
			9150: out = 24'(7508);
			9151: out = 24'(-1240);
			9152: out = 24'(-1004);
			9153: out = 24'(2536);
			9154: out = 24'(-1132);
			9155: out = 24'(-12808);
			9156: out = 24'(-1972);
			9157: out = 24'(6784);
			9158: out = 24'(-884);
			9159: out = 24'(2624);
			9160: out = 24'(4684);
			9161: out = 24'(-1028);
			9162: out = 24'(4568);
			9163: out = 24'(7400);
			9164: out = 24'(2032);
			9165: out = 24'(-8008);
			9166: out = 24'(-6596);
			9167: out = 24'(-292);
			9168: out = 24'(-924);
			9169: out = 24'(-1392);
			9170: out = 24'(756);
			9171: out = 24'(6900);
			9172: out = 24'(-1572);
			9173: out = 24'(4532);
			9174: out = 24'(12564);
			9175: out = 24'(7856);
			9176: out = 24'(-5836);
			9177: out = 24'(-9300);
			9178: out = 24'(-7512);
			9179: out = 24'(-5600);
			9180: out = 24'(304);
			9181: out = 24'(-4800);
			9182: out = 24'(-4756);
			9183: out = 24'(8380);
			9184: out = 24'(15128);
			9185: out = 24'(4400);
			9186: out = 24'(-12932);
			9187: out = 24'(-11712);
			9188: out = 24'(6104);
			9189: out = 24'(18840);
			9190: out = 24'(5796);
			9191: out = 24'(-7484);
			9192: out = 24'(-2736);
			9193: out = 24'(11616);
			9194: out = 24'(7800);
			9195: out = 24'(-3888);
			9196: out = 24'(-7348);
			9197: out = 24'(312);
			9198: out = 24'(2416);
			9199: out = 24'(5476);
			9200: out = 24'(3744);
			9201: out = 24'(744);
			9202: out = 24'(-14520);
			9203: out = 24'(-14424);
			9204: out = 24'(-2464);
			9205: out = 24'(-3788);
			9206: out = 24'(4156);
			9207: out = 24'(12096);
			9208: out = 24'(1892);
			9209: out = 24'(-10448);
			9210: out = 24'(-11196);
			9211: out = 24'(-7308);
			9212: out = 24'(8936);
			9213: out = 24'(12828);
			9214: out = 24'(7768);
			9215: out = 24'(-5640);
			9216: out = 24'(-5552);
			9217: out = 24'(-2052);
			9218: out = 24'(1708);
			9219: out = 24'(1976);
			9220: out = 24'(-3320);
			9221: out = 24'(2784);
			9222: out = 24'(2788);
			9223: out = 24'(10556);
			9224: out = 24'(8888);
			9225: out = 24'(6044);
			9226: out = 24'(1360);
			9227: out = 24'(-2220);
			9228: out = 24'(3376);
			9229: out = 24'(4468);
			9230: out = 24'(152);
			9231: out = 24'(-5372);
			9232: out = 24'(-8300);
			9233: out = 24'(-5184);
			9234: out = 24'(-3000);
			9235: out = 24'(-12544);
			9236: out = 24'(-14784);
			9237: out = 24'(-11136);
			9238: out = 24'(-6312);
			9239: out = 24'(8328);
			9240: out = 24'(19776);
			9241: out = 24'(10892);
			9242: out = 24'(-9876);
			9243: out = 24'(-17212);
			9244: out = 24'(-5912);
			9245: out = 24'(7628);
			9246: out = 24'(9836);
			9247: out = 24'(10964);
			9248: out = 24'(5272);
			9249: out = 24'(-11772);
			9250: out = 24'(-18424);
			9251: out = 24'(-10840);
			9252: out = 24'(3500);
			9253: out = 24'(10852);
			9254: out = 24'(9016);
			9255: out = 24'(-3100);
			9256: out = 24'(-10392);
			9257: out = 24'(-7856);
			9258: out = 24'(3904);
			9259: out = 24'(17364);
			9260: out = 24'(16916);
			9261: out = 24'(3160);
			9262: out = 24'(-6464);
			9263: out = 24'(-3180);
			9264: out = 24'(-5472);
			9265: out = 24'(-9060);
			9266: out = 24'(-6652);
			9267: out = 24'(884);
			9268: out = 24'(2652);
			9269: out = 24'(8968);
			9270: out = 24'(11992);
			9271: out = 24'(10588);
			9272: out = 24'(4468);
			9273: out = 24'(-688);
			9274: out = 24'(-4848);
			9275: out = 24'(-5232);
			9276: out = 24'(-5236);
			9277: out = 24'(-4420);
			9278: out = 24'(-2700);
			9279: out = 24'(524);
			9280: out = 24'(2672);
			9281: out = 24'(1852);
			9282: out = 24'(-5180);
			9283: out = 24'(-9256);
			9284: out = 24'(-5184);
			9285: out = 24'(976);
			9286: out = 24'(11204);
			9287: out = 24'(7028);
			9288: out = 24'(-2152);
			9289: out = 24'(-8916);
			9290: out = 24'(-3624);
			9291: out = 24'(6412);
			9292: out = 24'(-1328);
			9293: out = 24'(1148);
			9294: out = 24'(3160);
			9295: out = 24'(2880);
			9296: out = 24'(9916);
			9297: out = 24'(12376);
			9298: out = 24'(6020);
			9299: out = 24'(-3124);
			9300: out = 24'(-12444);
			9301: out = 24'(-8200);
			9302: out = 24'(-5420);
			9303: out = 24'(-6476);
			9304: out = 24'(-3028);
			9305: out = 24'(-16);
			9306: out = 24'(-40);
			9307: out = 24'(4704);
			9308: out = 24'(9708);
			9309: out = 24'(2552);
			9310: out = 24'(-8156);
			9311: out = 24'(-6668);
			9312: out = 24'(-6392);
			9313: out = 24'(-3004);
			9314: out = 24'(2968);
			9315: out = 24'(6952);
			9316: out = 24'(7192);
			9317: out = 24'(7668);
			9318: out = 24'(2172);
			9319: out = 24'(1496);
			9320: out = 24'(3656);
			9321: out = 24'(1808);
			9322: out = 24'(-1824);
			9323: out = 24'(-840);
			9324: out = 24'(9152);
			9325: out = 24'(4616);
			9326: out = 24'(-7136);
			9327: out = 24'(-10460);
			9328: out = 24'(-3880);
			9329: out = 24'(2788);
			9330: out = 24'(2964);
			9331: out = 24'(2196);
			9332: out = 24'(-4360);
			9333: out = 24'(-4464);
			9334: out = 24'(1912);
			9335: out = 24'(5188);
			9336: out = 24'(-10164);
			9337: out = 24'(-10044);
			9338: out = 24'(-1580);
			9339: out = 24'(6868);
			9340: out = 24'(5156);
			9341: out = 24'(1324);
			9342: out = 24'(5124);
			9343: out = 24'(4864);
			9344: out = 24'(2284);
			9345: out = 24'(-10316);
			9346: out = 24'(-11104);
			9347: out = 24'(-7124);
			9348: out = 24'(2132);
			9349: out = 24'(11468);
			9350: out = 24'(4844);
			9351: out = 24'(1812);
			9352: out = 24'(1752);
			9353: out = 24'(1556);
			9354: out = 24'(-5764);
			9355: out = 24'(-5792);
			9356: out = 24'(3616);
			9357: out = 24'(1068);
			9358: out = 24'(2036);
			9359: out = 24'(6456);
			9360: out = 24'(5148);
			9361: out = 24'(-484);
			9362: out = 24'(-6996);
			9363: out = 24'(-4204);
			9364: out = 24'(-6752);
			9365: out = 24'(-7632);
			9366: out = 24'(472);
			9367: out = 24'(5976);
			9368: out = 24'(88);
			9369: out = 24'(-5292);
			9370: out = 24'(-6792);
			9371: out = 24'(-1288);
			9372: out = 24'(-2712);
			9373: out = 24'(-3144);
			9374: out = 24'(9168);
			9375: out = 24'(4760);
			9376: out = 24'(1052);
			9377: out = 24'(7144);
			9378: out = 24'(5384);
			9379: out = 24'(-9740);
			9380: out = 24'(-13680);
			9381: out = 24'(-8728);
			9382: out = 24'(1992);
			9383: out = 24'(508);
			9384: out = 24'(-3112);
			9385: out = 24'(-468);
			9386: out = 24'(3076);
			9387: out = 24'(11492);
			9388: out = 24'(10452);
			9389: out = 24'(-740);
			9390: out = 24'(-15180);
			9391: out = 24'(-8044);
			9392: out = 24'(-7660);
			9393: out = 24'(-4720);
			9394: out = 24'(11320);
			9395: out = 24'(12652);
			9396: out = 24'(-2532);
			9397: out = 24'(-6936);
			9398: out = 24'(1720);
			9399: out = 24'(9476);
			9400: out = 24'(3332);
			9401: out = 24'(-6984);
			9402: out = 24'(-8832);
			9403: out = 24'(-5628);
			9404: out = 24'(5064);
			9405: out = 24'(10616);
			9406: out = 24'(-3816);
			9407: out = 24'(-21856);
			9408: out = 24'(-12152);
			9409: out = 24'(8204);
			9410: out = 24'(12500);
			9411: out = 24'(10152);
			9412: out = 24'(-28);
			9413: out = 24'(-8012);
			9414: out = 24'(-888);
			9415: out = 24'(736);
			9416: out = 24'(9096);
			9417: out = 24'(7292);
			9418: out = 24'(-1720);
			9419: out = 24'(-2280);
			9420: out = 24'(-2380);
			9421: out = 24'(380);
			9422: out = 24'(-1380);
			9423: out = 24'(-6556);
			9424: out = 24'(2852);
			9425: out = 24'(2884);
			9426: out = 24'(1780);
			9427: out = 24'(-1044);
			9428: out = 24'(-2012);
			9429: out = 24'(2728);
			9430: out = 24'(10220);
			9431: out = 24'(8640);
			9432: out = 24'(892);
			9433: out = 24'(-2108);
			9434: out = 24'(-1020);
			9435: out = 24'(1924);
			9436: out = 24'(-3960);
			9437: out = 24'(-5620);
			9438: out = 24'(-5288);
			9439: out = 24'(-592);
			9440: out = 24'(-4876);
			9441: out = 24'(-2816);
			9442: out = 24'(-8084);
			9443: out = 24'(-6604);
			9444: out = 24'(2816);
			9445: out = 24'(9176);
			9446: out = 24'(10044);
			9447: out = 24'(-1420);
			9448: out = 24'(-1444);
			9449: out = 24'(-2348);
			9450: out = 24'(-160);
			9451: out = 24'(1876);
			9452: out = 24'(-472);
			9453: out = 24'(6348);
			9454: out = 24'(9568);
			9455: out = 24'(-4260);
			9456: out = 24'(-12788);
			9457: out = 24'(-12296);
			9458: out = 24'(-6752);
			9459: out = 24'(5304);
			9460: out = 24'(9596);
			9461: out = 24'(876);
			9462: out = 24'(-2756);
			9463: out = 24'(-5036);
			9464: out = 24'(932);
			9465: out = 24'(6084);
			9466: out = 24'(-5088);
			9467: out = 24'(-5428);
			9468: out = 24'(5040);
			9469: out = 24'(4212);
			9470: out = 24'(-8176);
			9471: out = 24'(-9292);
			9472: out = 24'(-3796);
			9473: out = 24'(-636);
			9474: out = 24'(8200);
			9475: out = 24'(2548);
			9476: out = 24'(-7948);
			9477: out = 24'(-1492);
			9478: out = 24'(9352);
			9479: out = 24'(13544);
			9480: out = 24'(-584);
			9481: out = 24'(1392);
			9482: out = 24'(9084);
			9483: out = 24'(8512);
			9484: out = 24'(-9392);
			9485: out = 24'(-13408);
			9486: out = 24'(-4716);
			9487: out = 24'(-944);
			9488: out = 24'(936);
			9489: out = 24'(2248);
			9490: out = 24'(5160);
			9491: out = 24'(-420);
			9492: out = 24'(-3192);
			9493: out = 24'(-836);
			9494: out = 24'(1140);
			9495: out = 24'(4572);
			9496: out = 24'(2660);
			9497: out = 24'(-2984);
			9498: out = 24'(-5572);
			9499: out = 24'(-7684);
			9500: out = 24'(-6908);
			9501: out = 24'(7896);
			9502: out = 24'(13796);
			9503: out = 24'(-4016);
			9504: out = 24'(-14240);
			9505: out = 24'(-6836);
			9506: out = 24'(2060);
			9507: out = 24'(15180);
			9508: out = 24'(11080);
			9509: out = 24'(-1964);
			9510: out = 24'(-2828);
			9511: out = 24'(-2396);
			9512: out = 24'(3028);
			9513: out = 24'(-68);
			9514: out = 24'(-4556);
			9515: out = 24'(2460);
			9516: out = 24'(3892);
			9517: out = 24'(536);
			9518: out = 24'(-4872);
			9519: out = 24'(-9700);
			9520: out = 24'(-6928);
			9521: out = 24'(-1224);
			9522: out = 24'(-960);
			9523: out = 24'(5424);
			9524: out = 24'(4328);
			9525: out = 24'(-948);
			9526: out = 24'(-9852);
			9527: out = 24'(-13764);
			9528: out = 24'(3088);
			9529: out = 24'(12044);
			9530: out = 24'(9308);
			9531: out = 24'(4664);
			9532: out = 24'(2356);
			9533: out = 24'(-3260);
			9534: out = 24'(-8428);
			9535: out = 24'(-6320);
			9536: out = 24'(-2732);
			9537: out = 24'(-3220);
			9538: out = 24'(4864);
			9539: out = 24'(2444);
			9540: out = 24'(-2456);
			9541: out = 24'(7728);
			9542: out = 24'(9020);
			9543: out = 24'(4672);
			9544: out = 24'(-304);
			9545: out = 24'(52);
			9546: out = 24'(-3592);
			9547: out = 24'(-5120);
			9548: out = 24'(7376);
			9549: out = 24'(8584);
			9550: out = 24'(-180);
			9551: out = 24'(368);
			9552: out = 24'(-1676);
			9553: out = 24'(1404);
			9554: out = 24'(2792);
			9555: out = 24'(-2840);
			9556: out = 24'(972);
			9557: out = 24'(9500);
			9558: out = 24'(2292);
			9559: out = 24'(-12756);
			9560: out = 24'(-18232);
			9561: out = 24'(-2796);
			9562: out = 24'(4284);
			9563: out = 24'(-2080);
			9564: out = 24'(5548);
			9565: out = 24'(10676);
			9566: out = 24'(1628);
			9567: out = 24'(-17628);
			9568: out = 24'(-18928);
			9569: out = 24'(-5636);
			9570: out = 24'(6088);
			9571: out = 24'(12584);
			9572: out = 24'(9764);
			9573: out = 24'(-2416);
			9574: out = 24'(-15268);
			9575: out = 24'(-8572);
			9576: out = 24'(960);
			9577: out = 24'(13872);
			9578: out = 24'(8036);
			9579: out = 24'(-8452);
			9580: out = 24'(-9892);
			9581: out = 24'(1288);
			9582: out = 24'(15412);
			9583: out = 24'(7924);
			9584: out = 24'(-3504);
			9585: out = 24'(428);
			9586: out = 24'(4488);
			9587: out = 24'(4676);
			9588: out = 24'(6528);
			9589: out = 24'(-732);
			9590: out = 24'(-8144);
			9591: out = 24'(-15932);
			9592: out = 24'(-10816);
			9593: out = 24'(6224);
			9594: out = 24'(7284);
			9595: out = 24'(-5308);
			9596: out = 24'(-1588);
			9597: out = 24'(1260);
			9598: out = 24'(-5960);
			9599: out = 24'(-2624);
			9600: out = 24'(1992);
			9601: out = 24'(7120);
			9602: out = 24'(5044);
			9603: out = 24'(-3536);
			9604: out = 24'(-5396);
			9605: out = 24'(-660);
			9606: out = 24'(3788);
			9607: out = 24'(520);
			9608: out = 24'(-2288);
			9609: out = 24'(-280);
			9610: out = 24'(7992);
			9611: out = 24'(15716);
			9612: out = 24'(7128);
			9613: out = 24'(-8328);
			9614: out = 24'(-12080);
			9615: out = 24'(-4400);
			9616: out = 24'(2916);
			9617: out = 24'(9656);
			9618: out = 24'(4020);
			9619: out = 24'(-1272);
			9620: out = 24'(2244);
			9621: out = 24'(-576);
			9622: out = 24'(-9760);
			9623: out = 24'(-11424);
			9624: out = 24'(-9668);
			9625: out = 24'(1996);
			9626: out = 24'(10200);
			9627: out = 24'(9836);
			9628: out = 24'(-28);
			9629: out = 24'(-4032);
			9630: out = 24'(-6624);
			9631: out = 24'(3184);
			9632: out = 24'(11256);
			9633: out = 24'(4764);
			9634: out = 24'(-8016);
			9635: out = 24'(-7600);
			9636: out = 24'(664);
			9637: out = 24'(5424);
			9638: out = 24'(-4068);
			9639: out = 24'(-10644);
			9640: out = 24'(-2156);
			9641: out = 24'(4992);
			9642: out = 24'(9388);
			9643: out = 24'(4968);
			9644: out = 24'(-8056);
			9645: out = 24'(-7656);
			9646: out = 24'(1364);
			9647: out = 24'(7292);
			9648: out = 24'(3536);
			9649: out = 24'(-4040);
			9650: out = 24'(512);
			9651: out = 24'(3724);
			9652: out = 24'(-4056);
			9653: out = 24'(-4504);
			9654: out = 24'(712);
			9655: out = 24'(1524);
			9656: out = 24'(-3052);
			9657: out = 24'(-860);
			9658: out = 24'(4120);
			9659: out = 24'(2876);
			9660: out = 24'(-864);
			9661: out = 24'(-12740);
			9662: out = 24'(-17440);
			9663: out = 24'(1456);
			9664: out = 24'(16928);
			9665: out = 24'(11232);
			9666: out = 24'(-4704);
			9667: out = 24'(-9676);
			9668: out = 24'(2600);
			9669: out = 24'(13492);
			9670: out = 24'(7080);
			9671: out = 24'(144);
			9672: out = 24'(4140);
			9673: out = 24'(8688);
			9674: out = 24'(1784);
			9675: out = 24'(-11944);
			9676: out = 24'(-9008);
			9677: out = 24'(1188);
			9678: out = 24'(120);
			9679: out = 24'(-3624);
			9680: out = 24'(-636);
			9681: out = 24'(2464);
			9682: out = 24'(4252);
			9683: out = 24'(4748);
			9684: out = 24'(4092);
			9685: out = 24'(544);
			9686: out = 24'(2660);
			9687: out = 24'(2636);
			9688: out = 24'(4268);
			9689: out = 24'(2796);
			9690: out = 24'(-3480);
			9691: out = 24'(-2088);
			9692: out = 24'(1364);
			9693: out = 24'(-1984);
			9694: out = 24'(-8932);
			9695: out = 24'(-10656);
			9696: out = 24'(-3184);
			9697: out = 24'(3164);
			9698: out = 24'(4844);
			9699: out = 24'(-5856);
			9700: out = 24'(-8572);
			9701: out = 24'(1660);
			9702: out = 24'(3264);
			9703: out = 24'(272);
			9704: out = 24'(772);
			9705: out = 24'(6912);
			9706: out = 24'(5224);
			9707: out = 24'(136);
			9708: out = 24'(1152);
			9709: out = 24'(4424);
			9710: out = 24'(4400);
			9711: out = 24'(-5388);
			9712: out = 24'(-5864);
			9713: out = 24'(-2144);
			9714: out = 24'(5940);
			9715: out = 24'(2188);
			9716: out = 24'(-6608);
			9717: out = 24'(-8992);
			9718: out = 24'(904);
			9719: out = 24'(9180);
			9720: out = 24'(1608);
			9721: out = 24'(-2412);
			9722: out = 24'(2460);
			9723: out = 24'(8284);
			9724: out = 24'(-188);
			9725: out = 24'(-9704);
			9726: out = 24'(-5792);
			9727: out = 24'(-1640);
			9728: out = 24'(-6468);
			9729: out = 24'(-8496);
			9730: out = 24'(-892);
			9731: out = 24'(-1652);
			9732: out = 24'(1580);
			9733: out = 24'(2544);
			9734: out = 24'(-1592);
			9735: out = 24'(-11372);
			9736: out = 24'(-8196);
			9737: out = 24'(5552);
			9738: out = 24'(6456);
			9739: out = 24'(7600);
			9740: out = 24'(9612);
			9741: out = 24'(5236);
			9742: out = 24'(-9692);
			9743: out = 24'(-20504);
			9744: out = 24'(-18392);
			9745: out = 24'(-1736);
			9746: out = 24'(11968);
			9747: out = 24'(6300);
			9748: out = 24'(-1020);
			9749: out = 24'(1284);
			9750: out = 24'(5480);
			9751: out = 24'(7916);
			9752: out = 24'(1460);
			9753: out = 24'(4328);
			9754: out = 24'(11244);
			9755: out = 24'(5088);
			9756: out = 24'(-8036);
			9757: out = 24'(-11296);
			9758: out = 24'(-1440);
			9759: out = 24'(-824);
			9760: out = 24'(-14524);
			9761: out = 24'(-8504);
			9762: out = 24'(3540);
			9763: out = 24'(3344);
			9764: out = 24'(6400);
			9765: out = 24'(12824);
			9766: out = 24'(5224);
			9767: out = 24'(-9760);
			9768: out = 24'(-20644);
			9769: out = 24'(-10312);
			9770: out = 24'(5320);
			9771: out = 24'(8368);
			9772: out = 24'(3212);
			9773: out = 24'(-3936);
			9774: out = 24'(-7088);
			9775: out = 24'(-2368);
			9776: out = 24'(8036);
			9777: out = 24'(7276);
			9778: out = 24'(512);
			9779: out = 24'(-4992);
			9780: out = 24'(-9992);
			9781: out = 24'(-3680);
			9782: out = 24'(1228);
			9783: out = 24'(6748);
			9784: out = 24'(10692);
			9785: out = 24'(1244);
			9786: out = 24'(-9352);
			9787: out = 24'(-12024);
			9788: out = 24'(-4772);
			9789: out = 24'(11368);
			9790: out = 24'(11364);
			9791: out = 24'(280);
			9792: out = 24'(-7460);
			9793: out = 24'(-996);
			9794: out = 24'(9104);
			9795: out = 24'(9016);
			9796: out = 24'(-2752);
			9797: out = 24'(-3076);
			9798: out = 24'(-2008);
			9799: out = 24'(-2012);
			9800: out = 24'(2580);
			9801: out = 24'(1988);
			9802: out = 24'(-4724);
			9803: out = 24'(-6144);
			9804: out = 24'(-1500);
			9805: out = 24'(-1212);
			9806: out = 24'(-5396);
			9807: out = 24'(888);
			9808: out = 24'(4584);
			9809: out = 24'(7452);
			9810: out = 24'(1868);
			9811: out = 24'(1048);
			9812: out = 24'(5444);
			9813: out = 24'(4488);
			9814: out = 24'(-3828);
			9815: out = 24'(-8708);
			9816: out = 24'(-3548);
			9817: out = 24'(480);
			9818: out = 24'(1432);
			9819: out = 24'(2560);
			9820: out = 24'(6432);
			9821: out = 24'(1244);
			9822: out = 24'(-8192);
			9823: out = 24'(-8584);
			9824: out = 24'(-5392);
			9825: out = 24'(3056);
			9826: out = 24'(7948);
			9827: out = 24'(-484);
			9828: out = 24'(-8484);
			9829: out = 24'(-7316);
			9830: out = 24'(2612);
			9831: out = 24'(8452);
			9832: out = 24'(5488);
			9833: out = 24'(2168);
			9834: out = 24'(-7584);
			9835: out = 24'(-12896);
			9836: out = 24'(-8728);
			9837: out = 24'(4324);
			9838: out = 24'(14368);
			9839: out = 24'(704);
			9840: out = 24'(-5240);
			9841: out = 24'(5004);
			9842: out = 24'(6248);
			9843: out = 24'(4916);
			9844: out = 24'(-852);
			9845: out = 24'(-2320);
			9846: out = 24'(-5468);
			9847: out = 24'(-9688);
			9848: out = 24'(-488);
			9849: out = 24'(2776);
			9850: out = 24'(-156);
			9851: out = 24'(2320);
			9852: out = 24'(2072);
			9853: out = 24'(-2548);
			9854: out = 24'(-3892);
			9855: out = 24'(1456);
			9856: out = 24'(6364);
			9857: out = 24'(3448);
			9858: out = 24'(-3084);
			9859: out = 24'(-4700);
			9860: out = 24'(6524);
			9861: out = 24'(11340);
			9862: out = 24'(-3136);
			9863: out = 24'(-11864);
			9864: out = 24'(-6936);
			9865: out = 24'(2720);
			9866: out = 24'(4672);
			9867: out = 24'(6636);
			9868: out = 24'(4196);
			9869: out = 24'(1720);
			9870: out = 24'(-520);
			9871: out = 24'(520);
			9872: out = 24'(-328);
			9873: out = 24'(-6268);
			9874: out = 24'(-5480);
			9875: out = 24'(-2056);
			9876: out = 24'(1192);
			9877: out = 24'(1668);
			9878: out = 24'(2532);
			9879: out = 24'(-1292);
			9880: out = 24'(456);
			9881: out = 24'(4052);
			9882: out = 24'(2784);
			9883: out = 24'(-988);
			9884: out = 24'(-820);
			9885: out = 24'(-3000);
			9886: out = 24'(-4508);
			9887: out = 24'(-3388);
			9888: out = 24'(-5272);
			9889: out = 24'(4696);
			9890: out = 24'(9320);
			9891: out = 24'(-1900);
			9892: out = 24'(-7032);
			9893: out = 24'(-3860);
			9894: out = 24'(1784);
			9895: out = 24'(9796);
			9896: out = 24'(5228);
			9897: out = 24'(-6832);
			9898: out = 24'(-13364);
			9899: out = 24'(-3480);
			9900: out = 24'(12120);
			9901: out = 24'(8864);
			9902: out = 24'(-304);
			9903: out = 24'(-1396);
			9904: out = 24'(4320);
			9905: out = 24'(2416);
			9906: out = 24'(1544);
			9907: out = 24'(-1876);
			9908: out = 24'(-1004);
			9909: out = 24'(3124);
			9910: out = 24'(4056);
			9911: out = 24'(-1184);
			9912: out = 24'(-5468);
			9913: out = 24'(-1044);
			9914: out = 24'(2676);
			9915: out = 24'(312);
			9916: out = 24'(-3020);
			9917: out = 24'(-604);
			9918: out = 24'(2724);
			9919: out = 24'(3644);
			9920: out = 24'(-2860);
			9921: out = 24'(-8572);
			9922: out = 24'(-7792);
			9923: out = 24'(1192);
			9924: out = 24'(10204);
			9925: out = 24'(4424);
			9926: out = 24'(-2780);
			9927: out = 24'(-4240);
			9928: out = 24'(5188);
			9929: out = 24'(8324);
			9930: out = 24'(1292);
			9931: out = 24'(-7012);
			9932: out = 24'(-6100);
			9933: out = 24'(464);
			9934: out = 24'(1220);
			9935: out = 24'(-76);
			9936: out = 24'(-5864);
			9937: out = 24'(-8460);
			9938: out = 24'(-3744);
			9939: out = 24'(5436);
			9940: out = 24'(9036);
			9941: out = 24'(7032);
			9942: out = 24'(124);
			9943: out = 24'(-8884);
			9944: out = 24'(-4544);
			9945: out = 24'(-976);
			9946: out = 24'(3028);
			9947: out = 24'(8004);
			9948: out = 24'(1820);
			9949: out = 24'(196);
			9950: out = 24'(5004);
			9951: out = 24'(3240);
			9952: out = 24'(-1712);
			9953: out = 24'(-8028);
			9954: out = 24'(-7748);
			9955: out = 24'(-1668);
			9956: out = 24'(2836);
			9957: out = 24'(7584);
			9958: out = 24'(8844);
			9959: out = 24'(7288);
			9960: out = 24'(-1656);
			9961: out = 24'(-2872);
			9962: out = 24'(-1132);
			9963: out = 24'(3116);
			9964: out = 24'(-696);
			9965: out = 24'(588);
			9966: out = 24'(6796);
			9967: out = 24'(1932);
			9968: out = 24'(-8800);
			9969: out = 24'(-5144);
			9970: out = 24'(-4136);
			9971: out = 24'(-1088);
			9972: out = 24'(5068);
			9973: out = 24'(2532);
			9974: out = 24'(-6552);
			9975: out = 24'(-10260);
			9976: out = 24'(108);
			9977: out = 24'(4932);
			9978: out = 24'(5736);
			9979: out = 24'(4628);
			9980: out = 24'(4268);
			9981: out = 24'(-5700);
			9982: out = 24'(-9196);
			9983: out = 24'(-3644);
			9984: out = 24'(6856);
			9985: out = 24'(7688);
			9986: out = 24'(-6460);
			9987: out = 24'(-12012);
			9988: out = 24'(-4072);
			9989: out = 24'(2752);
			9990: out = 24'(2812);
			9991: out = 24'(724);
			9992: out = 24'(84);
			9993: out = 24'(3184);
			9994: out = 24'(5420);
			9995: out = 24'(-2512);
			9996: out = 24'(-7236);
			9997: out = 24'(-5372);
			9998: out = 24'(5340);
			9999: out = 24'(6152);
			10000: out = 24'(4060);
			10001: out = 24'(4732);
			10002: out = 24'(7992);
			10003: out = 24'(2948);
			10004: out = 24'(-7312);
			10005: out = 24'(-11384);
			10006: out = 24'(-5804);
			10007: out = 24'(1744);
			10008: out = 24'(5636);
			10009: out = 24'(4000);
			10010: out = 24'(-1564);
			10011: out = 24'(-2880);
			10012: out = 24'(1424);
			10013: out = 24'(5304);
			10014: out = 24'(-2328);
			10015: out = 24'(-13288);
			10016: out = 24'(-9072);
			10017: out = 24'(1500);
			10018: out = 24'(6064);
			10019: out = 24'(2680);
			10020: out = 24'(-7280);
			10021: out = 24'(-4592);
			10022: out = 24'(6808);
			10023: out = 24'(9816);
			10024: out = 24'(1208);
			10025: out = 24'(-12108);
			10026: out = 24'(-5544);
			10027: out = 24'(3888);
			10028: out = 24'(6568);
			10029: out = 24'(6772);
			10030: out = 24'(2096);
			10031: out = 24'(-2584);
			10032: out = 24'(-12);
			10033: out = 24'(-3740);
			10034: out = 24'(-6776);
			10035: out = 24'(-1264);
			10036: out = 24'(2816);
			10037: out = 24'(-3476);
			10038: out = 24'(-724);
			10039: out = 24'(-668);
			10040: out = 24'(1468);
			10041: out = 24'(7364);
			10042: out = 24'(152);
			10043: out = 24'(1680);
			10044: out = 24'(2280);
			10045: out = 24'(7652);
			10046: out = 24'(4140);
			10047: out = 24'(-772);
			10048: out = 24'(2044);
			10049: out = 24'(4420);
			10050: out = 24'(528);
			10051: out = 24'(-1572);
			10052: out = 24'(-380);
			10053: out = 24'(-672);
			10054: out = 24'(-5324);
			10055: out = 24'(-10240);
			10056: out = 24'(-6752);
			10057: out = 24'(-2160);
			10058: out = 24'(-352);
			10059: out = 24'(2800);
			10060: out = 24'(8828);
			10061: out = 24'(4144);
			10062: out = 24'(-4744);
			10063: out = 24'(-10564);
			10064: out = 24'(-8404);
			10065: out = 24'(2440);
			10066: out = 24'(-1392);
			10067: out = 24'(-36);
			10068: out = 24'(1796);
			10069: out = 24'(-552);
			10070: out = 24'(1060);
			10071: out = 24'(1868);
			10072: out = 24'(4276);
			10073: out = 24'(7516);
			10074: out = 24'(792);
			10075: out = 24'(-7124);
			10076: out = 24'(-10104);
			10077: out = 24'(-6956);
			10078: out = 24'(2892);
			10079: out = 24'(4524);
			10080: out = 24'(-7844);
			10081: out = 24'(-5516);
			10082: out = 24'(4832);
			10083: out = 24'(6356);
			10084: out = 24'(3588);
			10085: out = 24'(1268);
			10086: out = 24'(-1976);
			10087: out = 24'(-3832);
			10088: out = 24'(1484);
			10089: out = 24'(1792);
			10090: out = 24'(-2672);
			10091: out = 24'(-4080);
			10092: out = 24'(2796);
			10093: out = 24'(4092);
			10094: out = 24'(3856);
			10095: out = 24'(9104);
			10096: out = 24'(6136);
			10097: out = 24'(-3976);
			10098: out = 24'(-13884);
			10099: out = 24'(-10608);
			10100: out = 24'(-84);
			10101: out = 24'(10176);
			10102: out = 24'(4276);
			10103: out = 24'(-7660);
			10104: out = 24'(-5764);
			10105: out = 24'(124);
			10106: out = 24'(5796);
			10107: out = 24'(5384);
			10108: out = 24'(-5924);
			10109: out = 24'(-10256);
			10110: out = 24'(-4252);
			10111: out = 24'(4036);
			10112: out = 24'(6496);
			10113: out = 24'(4508);
			10114: out = 24'(1156);
			10115: out = 24'(-4672);
			10116: out = 24'(236);
			10117: out = 24'(5920);
			10118: out = 24'(5940);
			10119: out = 24'(2560);
			10120: out = 24'(-2276);
			10121: out = 24'(-4272);
			10122: out = 24'(-5448);
			10123: out = 24'(-356);
			10124: out = 24'(1872);
			10125: out = 24'(-5192);
			10126: out = 24'(-5528);
			10127: out = 24'(4704);
			10128: out = 24'(1436);
			10129: out = 24'(-7724);
			10130: out = 24'(-8200);
			10131: out = 24'(-28);
			10132: out = 24'(2816);
			10133: out = 24'(1356);
			10134: out = 24'(2348);
			10135: out = 24'(4012);
			10136: out = 24'(3616);
			10137: out = 24'(1964);
			10138: out = 24'(-2788);
			10139: out = 24'(-5760);
			10140: out = 24'(-3180);
			10141: out = 24'(-280);
			10142: out = 24'(6680);
			10143: out = 24'(11512);
			10144: out = 24'(6008);
			10145: out = 24'(-4784);
			10146: out = 24'(-8056);
			10147: out = 24'(-6080);
			10148: out = 24'(352);
			10149: out = 24'(356);
			10150: out = 24'(204);
			10151: out = 24'(2848);
			10152: out = 24'(3488);
			10153: out = 24'(-1312);
			10154: out = 24'(-2408);
			10155: out = 24'(2708);
			10156: out = 24'(3324);
			10157: out = 24'(-6388);
			10158: out = 24'(-6988);
			10159: out = 24'(2448);
			10160: out = 24'(-452);
			10161: out = 24'(-1540);
			10162: out = 24'(4884);
			10163: out = 24'(5036);
			10164: out = 24'(-5332);
			10165: out = 24'(-19764);
			10166: out = 24'(-17156);
			10167: out = 24'(1268);
			10168: out = 24'(14644);
			10169: out = 24'(10088);
			10170: out = 24'(-2456);
			10171: out = 24'(-4952);
			10172: out = 24'(-3548);
			10173: out = 24'(6736);
			10174: out = 24'(3788);
			10175: out = 24'(3476);
			10176: out = 24'(5868);
			10177: out = 24'(3200);
			10178: out = 24'(-164);
			10179: out = 24'(-2872);
			10180: out = 24'(-5200);
			10181: out = 24'(-2008);
			10182: out = 24'(-3128);
			10183: out = 24'(-2744);
			10184: out = 24'(-152);
			10185: out = 24'(1640);
			10186: out = 24'(3388);
			10187: out = 24'(-1432);
			10188: out = 24'(-7340);
			10189: out = 24'(-4840);
			10190: out = 24'(1508);
			10191: out = 24'(7196);
			10192: out = 24'(2440);
			10193: out = 24'(1216);
			10194: out = 24'(2836);
			10195: out = 24'(3740);
			10196: out = 24'(480);
			10197: out = 24'(-292);
			10198: out = 24'(-2840);
			10199: out = 24'(-1832);
			10200: out = 24'(-1240);
			10201: out = 24'(604);
			10202: out = 24'(5656);
			10203: out = 24'(2720);
			10204: out = 24'(-7928);
			10205: out = 24'(-12540);
			10206: out = 24'(-8640);
			10207: out = 24'(-2708);
			10208: out = 24'(6464);
			10209: out = 24'(4892);
			10210: out = 24'(-1008);
			10211: out = 24'(-4416);
			10212: out = 24'(-240);
			10213: out = 24'(3768);
			10214: out = 24'(4488);
			10215: out = 24'(1312);
			10216: out = 24'(-3240);
			10217: out = 24'(-3116);
			10218: out = 24'(-2592);
			10219: out = 24'(3332);
			10220: out = 24'(9148);
			10221: out = 24'(5208);
			10222: out = 24'(-2000);
			10223: out = 24'(-4380);
			10224: out = 24'(-3080);
			10225: out = 24'(2556);
			10226: out = 24'(4724);
			10227: out = 24'(-1008);
			10228: out = 24'(-4616);
			10229: out = 24'(-3028);
			10230: out = 24'(12);
			10231: out = 24'(2624);
			10232: out = 24'(2564);
			10233: out = 24'(-1872);
			10234: out = 24'(2228);
			10235: out = 24'(4216);
			10236: out = 24'(108);
			10237: out = 24'(-5500);
			10238: out = 24'(-7868);
			10239: out = 24'(-2944);
			10240: out = 24'(4460);
			10241: out = 24'(6280);
			10242: out = 24'(-1828);
			10243: out = 24'(-44);
			10244: out = 24'(6472);
			10245: out = 24'(5352);
			10246: out = 24'(-5216);
			10247: out = 24'(-13752);
			10248: out = 24'(-7232);
			10249: out = 24'(4728);
			10250: out = 24'(13052);
			10251: out = 24'(7352);
			10252: out = 24'(-3060);
			10253: out = 24'(-6196);
			10254: out = 24'(1328);
			10255: out = 24'(6672);
			10256: out = 24'(8820);
			10257: out = 24'(1752);
			10258: out = 24'(-2864);
			10259: out = 24'(-3752);
			10260: out = 24'(-3540);
			10261: out = 24'(-2164);
			10262: out = 24'(-5108);
			10263: out = 24'(-10244);
			10264: out = 24'(-5008);
			10265: out = 24'(3364);
			10266: out = 24'(1288);
			10267: out = 24'(2188);
			10268: out = 24'(8588);
			10269: out = 24'(6752);
			10270: out = 24'(-5052);
			10271: out = 24'(-12612);
			10272: out = 24'(-8036);
			10273: out = 24'(1276);
			10274: out = 24'(11192);
			10275: out = 24'(8552);
			10276: out = 24'(-4672);
			10277: out = 24'(-12680);
			10278: out = 24'(-7696);
			10279: out = 24'(5352);
			10280: out = 24'(6632);
			10281: out = 24'(2568);
			10282: out = 24'(1192);
			10283: out = 24'(-420);
			10284: out = 24'(-5688);
			10285: out = 24'(-5076);
			10286: out = 24'(1724);
			10287: out = 24'(5796);
			10288: out = 24'(8268);
			10289: out = 24'(1460);
			10290: out = 24'(-7120);
			10291: out = 24'(-6164);
			10292: out = 24'(2272);
			10293: out = 24'(8820);
			10294: out = 24'(4536);
			10295: out = 24'(-3636);
			10296: out = 24'(-4328);
			10297: out = 24'(952);
			10298: out = 24'(8908);
			10299: out = 24'(5616);
			10300: out = 24'(-4872);
			10301: out = 24'(-5628);
			10302: out = 24'(-2624);
			10303: out = 24'(-2456);
			10304: out = 24'(292);
			10305: out = 24'(1664);
			10306: out = 24'(944);
			10307: out = 24'(-260);
			10308: out = 24'(3032);
			10309: out = 24'(2848);
			10310: out = 24'(-628);
			10311: out = 24'(4228);
			10312: out = 24'(5964);
			10313: out = 24'(4668);
			10314: out = 24'(-1256);
			10315: out = 24'(-5104);
			10316: out = 24'(-3984);
			10317: out = 24'(2512);
			10318: out = 24'(1888);
			10319: out = 24'(-6140);
			10320: out = 24'(-8532);
			10321: out = 24'(-972);
			10322: out = 24'(5296);
			10323: out = 24'(-324);
			10324: out = 24'(-6744);
			10325: out = 24'(-784);
			10326: out = 24'(3700);
			10327: out = 24'(4544);
			10328: out = 24'(-4);
			10329: out = 24'(176);
			10330: out = 24'(4212);
			10331: out = 24'(2272);
			10332: out = 24'(-896);
			10333: out = 24'(-4144);
			10334: out = 24'(-488);
			10335: out = 24'(228);
			10336: out = 24'(-480);
			10337: out = 24'(2568);
			10338: out = 24'(-220);
			10339: out = 24'(-1928);
			10340: out = 24'(572);
			10341: out = 24'(1308);
			10342: out = 24'(28);
			10343: out = 24'(624);
			10344: out = 24'(524);
			10345: out = 24'(-2676);
			10346: out = 24'(-3516);
			10347: out = 24'(-4640);
			10348: out = 24'(-2540);
			10349: out = 24'(36);
			10350: out = 24'(1676);
			10351: out = 24'(-1560);
			10352: out = 24'(-4180);
			10353: out = 24'(-572);
			10354: out = 24'(1560);
			10355: out = 24'(2636);
			10356: out = 24'(-4560);
			10357: out = 24'(-120);
			10358: out = 24'(4076);
			10359: out = 24'(1436);
			10360: out = 24'(2436);
			10361: out = 24'(4760);
			10362: out = 24'(-1888);
			10363: out = 24'(-5168);
			10364: out = 24'(984);
			10365: out = 24'(480);
			10366: out = 24'(-2240);
			10367: out = 24'(-8664);
			10368: out = 24'(-5396);
			10369: out = 24'(3696);
			10370: out = 24'(9720);
			10371: out = 24'(8060);
			10372: out = 24'(-188);
			10373: out = 24'(-3360);
			10374: out = 24'(-4288);
			10375: out = 24'(464);
			10376: out = 24'(2176);
			10377: out = 24'(3204);
			10378: out = 24'(3128);
			10379: out = 24'(3868);
			10380: out = 24'(-3880);
			10381: out = 24'(-7060);
			10382: out = 24'(-492);
			10383: out = 24'(2588);
			10384: out = 24'(-936);
			10385: out = 24'(-84);
			10386: out = 24'(1948);
			10387: out = 24'(-5692);
			10388: out = 24'(-10072);
			10389: out = 24'(-5876);
			10390: out = 24'(1084);
			10391: out = 24'(6404);
			10392: out = 24'(6468);
			10393: out = 24'(620);
			10394: out = 24'(-7072);
			10395: out = 24'(-7336);
			10396: out = 24'(3780);
			10397: out = 24'(9888);
			10398: out = 24'(2444);
			10399: out = 24'(-7244);
			10400: out = 24'(-6184);
			10401: out = 24'(408);
			10402: out = 24'(4452);
			10403: out = 24'(2460);
			10404: out = 24'(4);
			10405: out = 24'(6080);
			10406: out = 24'(8860);
			10407: out = 24'(-576);
			10408: out = 24'(-4104);
			10409: out = 24'(-3540);
			10410: out = 24'(3472);
			10411: out = 24'(364);
			10412: out = 24'(-1564);
			10413: out = 24'(5416);
			10414: out = 24'(5092);
			10415: out = 24'(-1352);
			10416: out = 24'(-1172);
			10417: out = 24'(-612);
			10418: out = 24'(636);
			10419: out = 24'(-4216);
			10420: out = 24'(-5120);
			10421: out = 24'(1316);
			10422: out = 24'(136);
			10423: out = 24'(-4236);
			10424: out = 24'(-3056);
			10425: out = 24'(-2772);
			10426: out = 24'(-9652);
			10427: out = 24'(-3156);
			10428: out = 24'(3804);
			10429: out = 24'(1944);
			10430: out = 24'(4828);
			10431: out = 24'(3376);
			10432: out = 24'(-4368);
			10433: out = 24'(-7168);
			10434: out = 24'(-2268);
			10435: out = 24'(7464);
			10436: out = 24'(5192);
			10437: out = 24'(-856);
			10438: out = 24'(-272);
			10439: out = 24'(3768);
			10440: out = 24'(5620);
			10441: out = 24'(-1060);
			10442: out = 24'(-8760);
			10443: out = 24'(-3760);
			10444: out = 24'(3112);
			10445: out = 24'(2636);
			10446: out = 24'(-1104);
			10447: out = 24'(-2200);
			10448: out = 24'(80);
			10449: out = 24'(5672);
			10450: out = 24'(7092);
			10451: out = 24'(4732);
			10452: out = 24'(1900);
			10453: out = 24'(680);
			10454: out = 24'(-688);
			10455: out = 24'(868);
			10456: out = 24'(-1076);
			10457: out = 24'(-4588);
			10458: out = 24'(-6508);
			10459: out = 24'(-1796);
			10460: out = 24'(2524);
			10461: out = 24'(-2256);
			10462: out = 24'(-5664);
			10463: out = 24'(2536);
			10464: out = 24'(4640);
			10465: out = 24'(-304);
			10466: out = 24'(-5936);
			10467: out = 24'(-1900);
			10468: out = 24'(-472);
			10469: out = 24'(-144);
			10470: out = 24'(2884);
			10471: out = 24'(-608);
			10472: out = 24'(-5904);
			10473: out = 24'(-4880);
			10474: out = 24'(-436);
			10475: out = 24'(64);
			10476: out = 24'(2120);
			10477: out = 24'(3676);
			10478: out = 24'(4628);
			10479: out = 24'(1860);
			10480: out = 24'(-1088);
			10481: out = 24'(-2084);
			10482: out = 24'(212);
			10483: out = 24'(2792);
			10484: out = 24'(-1520);
			10485: out = 24'(-2452);
			10486: out = 24'(-2108);
			10487: out = 24'(-1708);
			10488: out = 24'(1616);
			10489: out = 24'(5176);
			10490: out = 24'(-1332);
			10491: out = 24'(-6352);
			10492: out = 24'(-328);
			10493: out = 24'(6340);
			10494: out = 24'(124);
			10495: out = 24'(-2788);
			10496: out = 24'(2168);
			10497: out = 24'(2080);
			10498: out = 24'(-2048);
			10499: out = 24'(1104);
			10500: out = 24'(1444);
			10501: out = 24'(960);
			10502: out = 24'(-684);
			10503: out = 24'(-4148);
			10504: out = 24'(1956);
			10505: out = 24'(3292);
			10506: out = 24'(-1932);
			10507: out = 24'(-3052);
			10508: out = 24'(-2476);
			10509: out = 24'(-3360);
			10510: out = 24'(-1272);
			10511: out = 24'(68);
			10512: out = 24'(2596);
			10513: out = 24'(2048);
			10514: out = 24'(2024);
			10515: out = 24'(-672);
			10516: out = 24'(-56);
			10517: out = 24'(-916);
			10518: out = 24'(-4708);
			10519: out = 24'(-596);
			10520: out = 24'(2952);
			10521: out = 24'(1220);
			10522: out = 24'(-6560);
			10523: out = 24'(-4480);
			10524: out = 24'(1196);
			10525: out = 24'(3744);
			10526: out = 24'(656);
			10527: out = 24'(-340);
			10528: out = 24'(-936);
			10529: out = 24'(-2256);
			10530: out = 24'(2520);
			10531: out = 24'(2956);
			10532: out = 24'(3080);
			10533: out = 24'(-2980);
			10534: out = 24'(-5708);
			10535: out = 24'(-1168);
			10536: out = 24'(1980);
			10537: out = 24'(4136);
			10538: out = 24'(2072);
			10539: out = 24'(-6120);
			10540: out = 24'(-8272);
			10541: out = 24'(-2096);
			10542: out = 24'(4248);
			10543: out = 24'(4248);
			10544: out = 24'(-556);
			10545: out = 24'(-1560);
			10546: out = 24'(-1544);
			10547: out = 24'(-1888);
			10548: out = 24'(692);
			10549: out = 24'(4572);
			10550: out = 24'(1436);
			10551: out = 24'(616);
			10552: out = 24'(-508);
			10553: out = 24'(1916);
			10554: out = 24'(2316);
			10555: out = 24'(-2864);
			10556: out = 24'(-6244);
			10557: out = 24'(-1528);
			10558: out = 24'(-172);
			10559: out = 24'(-3888);
			10560: out = 24'(-1684);
			10561: out = 24'(1428);
			10562: out = 24'(744);
			10563: out = 24'(2872);
			10564: out = 24'(3872);
			10565: out = 24'(-1920);
			10566: out = 24'(-8876);
			10567: out = 24'(-8012);
			10568: out = 24'(1176);
			10569: out = 24'(6428);
			10570: out = 24'(3684);
			10571: out = 24'(1144);
			10572: out = 24'(2940);
			10573: out = 24'(2664);
			10574: out = 24'(1412);
			10575: out = 24'(-2464);
			10576: out = 24'(-4520);
			10577: out = 24'(-2288);
			10578: out = 24'(4580);
			10579: out = 24'(2484);
			10580: out = 24'(-2436);
			10581: out = 24'(-3020);
			10582: out = 24'(-1916);
			10583: out = 24'(-1944);
			10584: out = 24'(1460);
			10585: out = 24'(7008);
			10586: out = 24'(3448);
			10587: out = 24'(-3128);
			10588: out = 24'(-6704);
			10589: out = 24'(-1468);
			10590: out = 24'(5708);
			10591: out = 24'(404);
			10592: out = 24'(-3148);
			10593: out = 24'(-636);
			10594: out = 24'(-460);
			10595: out = 24'(-3036);
			10596: out = 24'(-2224);
			10597: out = 24'(1348);
			10598: out = 24'(1648);
			10599: out = 24'(608);
			10600: out = 24'(2248);
			10601: out = 24'(-572);
			10602: out = 24'(-1744);
			10603: out = 24'(-5052);
			10604: out = 24'(-608);
			10605: out = 24'(2660);
			10606: out = 24'(1268);
			10607: out = 24'(4580);
			10608: out = 24'(1972);
			10609: out = 24'(-3728);
			10610: out = 24'(-4588);
			10611: out = 24'(-1324);
			10612: out = 24'(2328);
			10613: out = 24'(1616);
			10614: out = 24'(4528);
			10615: out = 24'(5536);
			10616: out = 24'(296);
			10617: out = 24'(-5896);
			10618: out = 24'(-6332);
			10619: out = 24'(-736);
			10620: out = 24'(3636);
			10621: out = 24'(272);
			10622: out = 24'(-3912);
			10623: out = 24'(-3204);
			10624: out = 24'(-4536);
			10625: out = 24'(-4472);
			10626: out = 24'(5636);
			10627: out = 24'(3556);
			10628: out = 24'(-2188);
			10629: out = 24'(1236);
			10630: out = 24'(4784);
			10631: out = 24'(-332);
			10632: out = 24'(-7628);
			10633: out = 24'(-7272);
			10634: out = 24'(-1968);
			10635: out = 24'(6108);
			10636: out = 24'(8248);
			10637: out = 24'(-1800);
			10638: out = 24'(-3428);
			10639: out = 24'(32);
			10640: out = 24'(7680);
			10641: out = 24'(7108);
			10642: out = 24'(1800);
			10643: out = 24'(-164);
			10644: out = 24'(2676);
			10645: out = 24'(1708);
			10646: out = 24'(-3296);
			10647: out = 24'(-6412);
			10648: out = 24'(-2176);
			10649: out = 24'(440);
			10650: out = 24'(-2448);
			10651: out = 24'(144);
			10652: out = 24'(3172);
			10653: out = 24'(384);
			10654: out = 24'(-4172);
			10655: out = 24'(-6632);
			10656: out = 24'(-4932);
			10657: out = 24'(-2524);
			10658: out = 24'(1808);
			10659: out = 24'(7128);
			10660: out = 24'(2664);
			10661: out = 24'(-1048);
			10662: out = 24'(1448);
			10663: out = 24'(3064);
			10664: out = 24'(1180);
			10665: out = 24'(-5700);
			10666: out = 24'(-5364);
			10667: out = 24'(2492);
			10668: out = 24'(1312);
			10669: out = 24'(-436);
			10670: out = 24'(3232);
			10671: out = 24'(3352);
			10672: out = 24'(3136);
			10673: out = 24'(-144);
			10674: out = 24'(-2076);
			10675: out = 24'(-680);
			10676: out = 24'(-2196);
			10677: out = 24'(2216);
			10678: out = 24'(2612);
			10679: out = 24'(-152);
			10680: out = 24'(-1772);
			10681: out = 24'(1424);
			10682: out = 24'(2108);
			10683: out = 24'(3024);
			10684: out = 24'(-1188);
			10685: out = 24'(-3088);
			10686: out = 24'(-664);
			10687: out = 24'(1236);
			10688: out = 24'(3044);
			10689: out = 24'(-276);
			10690: out = 24'(-3420);
			10691: out = 24'(-120);
			10692: out = 24'(3224);
			10693: out = 24'(2400);
			10694: out = 24'(-584);
			10695: out = 24'(-3500);
			10696: out = 24'(-1204);
			10697: out = 24'(-1564);
			10698: out = 24'(1932);
			10699: out = 24'(4188);
			10700: out = 24'(-1156);
			10701: out = 24'(-9596);
			10702: out = 24'(-7536);
			10703: out = 24'(-3368);
			10704: out = 24'(-448);
			10705: out = 24'(4472);
			10706: out = 24'(2748);
			10707: out = 24'(-1768);
			10708: out = 24'(-168);
			10709: out = 24'(3496);
			10710: out = 24'(2036);
			10711: out = 24'(-264);
			10712: out = 24'(-1816);
			10713: out = 24'(-168);
			10714: out = 24'(-3012);
			10715: out = 24'(-3740);
			10716: out = 24'(3480);
			10717: out = 24'(4928);
			10718: out = 24'(1164);
			10719: out = 24'(-2740);
			10720: out = 24'(-4052);
			10721: out = 24'(-1640);
			10722: out = 24'(5600);
			10723: out = 24'(7044);
			10724: out = 24'(-1776);
			10725: out = 24'(-8684);
			10726: out = 24'(-3772);
			10727: out = 24'(4656);
			10728: out = 24'(5452);
			10729: out = 24'(-1216);
			10730: out = 24'(-2656);
			10731: out = 24'(3720);
			10732: out = 24'(4380);
			10733: out = 24'(396);
			10734: out = 24'(-2928);
			10735: out = 24'(-512);
			10736: out = 24'(-448);
			10737: out = 24'(-2612);
			10738: out = 24'(-3432);
			10739: out = 24'(-460);
			10740: out = 24'(5228);
			10741: out = 24'(4516);
			10742: out = 24'(-3392);
			10743: out = 24'(-7900);
			10744: out = 24'(-6012);
			10745: out = 24'(4320);
			10746: out = 24'(10092);
			10747: out = 24'(3992);
			10748: out = 24'(-6124);
			10749: out = 24'(-8348);
			10750: out = 24'(-2548);
			10751: out = 24'(4988);
			10752: out = 24'(5876);
			10753: out = 24'(-1296);
			10754: out = 24'(-4272);
			10755: out = 24'(-1908);
			10756: out = 24'(-476);
			10757: out = 24'(3316);
			10758: out = 24'(564);
			10759: out = 24'(512);
			10760: out = 24'(3824);
			10761: out = 24'(1736);
			10762: out = 24'(-1324);
			10763: out = 24'(-5204);
			10764: out = 24'(-4436);
			10765: out = 24'(848);
			10766: out = 24'(5548);
			10767: out = 24'(-256);
			10768: out = 24'(-2664);
			10769: out = 24'(2116);
			10770: out = 24'(2840);
			10771: out = 24'(1048);
			10772: out = 24'(-2652);
			10773: out = 24'(-688);
			10774: out = 24'(1220);
			10775: out = 24'(5072);
			10776: out = 24'(4240);
			10777: out = 24'(-688);
			10778: out = 24'(-7080);
			10779: out = 24'(-6032);
			10780: out = 24'(-1540);
			10781: out = 24'(508);
			10782: out = 24'(980);
			10783: out = 24'(1916);
			10784: out = 24'(444);
			10785: out = 24'(588);
			10786: out = 24'(880);
			10787: out = 24'(64);
			10788: out = 24'(-1264);
			10789: out = 24'(-972);
			10790: out = 24'(1468);
			10791: out = 24'(-1728);
			10792: out = 24'(-4336);
			10793: out = 24'(-1464);
			10794: out = 24'(2372);
			10795: out = 24'(4156);
			10796: out = 24'(3156);
			10797: out = 24'(2488);
			10798: out = 24'(2848);
			10799: out = 24'(628);
			10800: out = 24'(-2888);
			10801: out = 24'(-5180);
			10802: out = 24'(-7544);
			10803: out = 24'(-5752);
			10804: out = 24'(416);
			10805: out = 24'(1860);
			10806: out = 24'(1664);
			10807: out = 24'(2916);
			10808: out = 24'(5592);
			10809: out = 24'(5136);
			10810: out = 24'(-1876);
			10811: out = 24'(-7296);
			10812: out = 24'(-7432);
			10813: out = 24'(-4168);
			10814: out = 24'(2760);
			10815: out = 24'(6852);
			10816: out = 24'(2664);
			10817: out = 24'(-652);
			10818: out = 24'(588);
			10819: out = 24'(1480);
			10820: out = 24'(8);
			10821: out = 24'(-4052);
			10822: out = 24'(-3048);
			10823: out = 24'(1004);
			10824: out = 24'(4644);
			10825: out = 24'(452);
			10826: out = 24'(-3524);
			10827: out = 24'(-804);
			10828: out = 24'(4696);
			10829: out = 24'(3812);
			10830: out = 24'(-1204);
			10831: out = 24'(-1312);
			10832: out = 24'(1068);
			10833: out = 24'(1180);
			10834: out = 24'(-820);
			10835: out = 24'(-1404);
			10836: out = 24'(-1088);
			10837: out = 24'(-2764);
			10838: out = 24'(-3676);
			10839: out = 24'(-1120);
			10840: out = 24'(-912);
			10841: out = 24'(-192);
			10842: out = 24'(2216);
			10843: out = 24'(2856);
			10844: out = 24'(-1192);
			10845: out = 24'(-7292);
			10846: out = 24'(-7112);
			10847: out = 24'(-32);
			10848: out = 24'(5304);
			10849: out = 24'(4356);
			10850: out = 24'(496);
			10851: out = 24'(-888);
			10852: out = 24'(-1080);
			10853: out = 24'(1652);
			10854: out = 24'(2328);
			10855: out = 24'(-1840);
			10856: out = 24'(-2464);
			10857: out = 24'(-628);
			10858: out = 24'(2880);
			10859: out = 24'(3944);
			10860: out = 24'(1820);
			10861: out = 24'(252);
			10862: out = 24'(32);
			10863: out = 24'(-996);
			10864: out = 24'(-5420);
			10865: out = 24'(-7736);
			10866: out = 24'(-1224);
			10867: out = 24'(3124);
			10868: out = 24'(-820);
			10869: out = 24'(-2872);
			10870: out = 24'(576);
			10871: out = 24'(3420);
			10872: out = 24'(1412);
			10873: out = 24'(-6660);
			10874: out = 24'(-5188);
			10875: out = 24'(-572);
			10876: out = 24'(2092);
			10877: out = 24'(4916);
			10878: out = 24'(4840);
			10879: out = 24'(548);
			10880: out = 24'(-3268);
			10881: out = 24'(-5768);
			10882: out = 24'(-5972);
			10883: out = 24'(-1328);
			10884: out = 24'(860);
			10885: out = 24'(2544);
			10886: out = 24'(3720);
			10887: out = 24'(2144);
			10888: out = 24'(-1916);
			10889: out = 24'(-1208);
			10890: out = 24'(1892);
			10891: out = 24'(856);
			10892: out = 24'(-296);
			10893: out = 24'(988);
			10894: out = 24'(2028);
			10895: out = 24'(-2328);
			10896: out = 24'(-3168);
			10897: out = 24'(-1356);
			10898: out = 24'(2240);
			10899: out = 24'(68);
			10900: out = 24'(-3184);
			10901: out = 24'(-360);
			10902: out = 24'(2096);
			10903: out = 24'(3572);
			10904: out = 24'(1712);
			10905: out = 24'(912);
			10906: out = 24'(-2376);
			10907: out = 24'(-4728);
			10908: out = 24'(-2848);
			10909: out = 24'(2876);
			10910: out = 24'(5924);
			10911: out = 24'(172);
			10912: out = 24'(-3864);
			10913: out = 24'(-1500);
			10914: out = 24'(1680);
			10915: out = 24'(1592);
			10916: out = 24'(-5032);
			10917: out = 24'(-5756);
			10918: out = 24'(-196);
			10919: out = 24'(2512);
			10920: out = 24'(2616);
			10921: out = 24'(628);
			10922: out = 24'(1004);
			10923: out = 24'(-284);
			10924: out = 24'(-4068);
			10925: out = 24'(-184);
			10926: out = 24'(2764);
			10927: out = 24'(-252);
			10928: out = 24'(-1156);
			10929: out = 24'(2296);
			10930: out = 24'(1244);
			10931: out = 24'(-6024);
			10932: out = 24'(-9748);
			10933: out = 24'(-4944);
			10934: out = 24'(828);
			10935: out = 24'(4316);
			10936: out = 24'(5556);
			10937: out = 24'(2028);
			10938: out = 24'(-3168);
			10939: out = 24'(-5080);
			10940: out = 24'(-1672);
			10941: out = 24'(4048);
			10942: out = 24'(6376);
			10943: out = 24'(-912);
			10944: out = 24'(-6092);
			10945: out = 24'(-5100);
			10946: out = 24'(2036);
			10947: out = 24'(5468);
			10948: out = 24'(340);
			10949: out = 24'(-1760);
			10950: out = 24'(3380);
			10951: out = 24'(4340);
			10952: out = 24'(-1204);
			10953: out = 24'(-7556);
			10954: out = 24'(-4328);
			10955: out = 24'(792);
			10956: out = 24'(1280);
			10957: out = 24'(3540);
			10958: out = 24'(2484);
			10959: out = 24'(-1036);
			10960: out = 24'(-1048);
			10961: out = 24'(-1584);
			10962: out = 24'(-3712);
			10963: out = 24'(-3068);
			10964: out = 24'(532);
			10965: out = 24'(2408);
			10966: out = 24'(732);
			10967: out = 24'(2332);
			10968: out = 24'(2968);
			10969: out = 24'(1964);
			10970: out = 24'(556);
			10971: out = 24'(-1384);
			10972: out = 24'(1680);
			10973: out = 24'(3420);
			10974: out = 24'(1624);
			10975: out = 24'(-2040);
			10976: out = 24'(-1876);
			10977: out = 24'(-252);
			10978: out = 24'(-704);
			10979: out = 24'(-5164);
			10980: out = 24'(-2524);
			10981: out = 24'(1128);
			10982: out = 24'(2084);
			10983: out = 24'(3536);
			10984: out = 24'(4100);
			10985: out = 24'(1396);
			10986: out = 24'(-4976);
			10987: out = 24'(-5292);
			10988: out = 24'(-756);
			10989: out = 24'(2096);
			10990: out = 24'(572);
			10991: out = 24'(-1868);
			10992: out = 24'(-248);
			10993: out = 24'(2376);
			10994: out = 24'(852);
			10995: out = 24'(720);
			10996: out = 24'(164);
			10997: out = 24'(-620);
			10998: out = 24'(-212);
			10999: out = 24'(-1524);
			11000: out = 24'(-3628);
			11001: out = 24'(-1956);
			11002: out = 24'(2020);
			11003: out = 24'(4504);
			11004: out = 24'(3264);
			11005: out = 24'(-424);
			11006: out = 24'(-1576);
			11007: out = 24'(-1532);
			11008: out = 24'(764);
			11009: out = 24'(5808);
			11010: out = 24'(2220);
			11011: out = 24'(-3204);
			11012: out = 24'(-2844);
			11013: out = 24'(740);
			11014: out = 24'(2924);
			11015: out = 24'(-708);
			11016: out = 24'(-6332);
			11017: out = 24'(-2776);
			11018: out = 24'(3140);
			11019: out = 24'(4348);
			11020: out = 24'(-2824);
			11021: out = 24'(-3088);
			11022: out = 24'(1132);
			11023: out = 24'(3164);
			11024: out = 24'(2632);
			11025: out = 24'(844);
			11026: out = 24'(-516);
			11027: out = 24'(1332);
			11028: out = 24'(3200);
			11029: out = 24'(240);
			11030: out = 24'(-4528);
			11031: out = 24'(-5952);
			11032: out = 24'(-1368);
			11033: out = 24'(-132);
			11034: out = 24'(1360);
			11035: out = 24'(716);
			11036: out = 24'(1820);
			11037: out = 24'(40);
			11038: out = 24'(-4884);
			11039: out = 24'(-2380);
			11040: out = 24'(1924);
			11041: out = 24'(5428);
			11042: out = 24'(2684);
			11043: out = 24'(-128);
			11044: out = 24'(-1104);
			11045: out = 24'(188);
			11046: out = 24'(568);
			11047: out = 24'(-504);
			11048: out = 24'(-28);
			11049: out = 24'(696);
			11050: out = 24'(292);
			11051: out = 24'(-1828);
			11052: out = 24'(-852);
			11053: out = 24'(-1864);
			11054: out = 24'(-1440);
			11055: out = 24'(-1436);
			11056: out = 24'(-3144);
			11057: out = 24'(-1232);
			11058: out = 24'(760);
			11059: out = 24'(1328);
			11060: out = 24'(1988);
			11061: out = 24'(1792);
			11062: out = 24'(3056);
			11063: out = 24'(-1284);
			11064: out = 24'(-3740);
			11065: out = 24'(1740);
			11066: out = 24'(4172);
			11067: out = 24'(932);
			11068: out = 24'(-2932);
			11069: out = 24'(-5404);
			11070: out = 24'(-396);
			11071: out = 24'(3572);
			11072: out = 24'(2268);
			11073: out = 24'(-448);
			11074: out = 24'(-144);
			11075: out = 24'(2412);
			11076: out = 24'(2128);
			11077: out = 24'(92);
			11078: out = 24'(-3632);
			11079: out = 24'(-3372);
			11080: out = 24'(1944);
			11081: out = 24'(1064);
			11082: out = 24'(-2384);
			11083: out = 24'(-3344);
			11084: out = 24'(-3648);
			11085: out = 24'(2088);
			11086: out = 24'(6924);
			11087: out = 24'(2752);
			11088: out = 24'(-6148);
			11089: out = 24'(-9164);
			11090: out = 24'(-6592);
			11091: out = 24'(2296);
			11092: out = 24'(8088);
			11093: out = 24'(1920);
			11094: out = 24'(-2408);
			11095: out = 24'(-204);
			11096: out = 24'(2000);
			11097: out = 24'(1084);
			11098: out = 24'(-1912);
			11099: out = 24'(-1828);
			11100: out = 24'(2948);
			11101: out = 24'(7076);
			11102: out = 24'(2292);
			11103: out = 24'(-4752);
			11104: out = 24'(-5392);
			11105: out = 24'(-1860);
			11106: out = 24'(764);
			11107: out = 24'(2644);
			11108: out = 24'(3292);
			11109: out = 24'(-1120);
			11110: out = 24'(-3612);
			11111: out = 24'(-708);
			11112: out = 24'(152);
			11113: out = 24'(-20);
			11114: out = 24'(-3036);
			11115: out = 24'(-2892);
			11116: out = 24'(668);
			11117: out = 24'(2192);
			11118: out = 24'(3540);
			11119: out = 24'(-116);
			11120: out = 24'(-3300);
			11121: out = 24'(-872);
			11122: out = 24'(1384);
			11123: out = 24'(2476);
			11124: out = 24'(2920);
			11125: out = 24'(2840);
			11126: out = 24'(-148);
			11127: out = 24'(-5192);
			11128: out = 24'(-7364);
			11129: out = 24'(-1764);
			11130: out = 24'(2912);
			11131: out = 24'(-120);
			11132: out = 24'(-2844);
			11133: out = 24'(-2788);
			11134: out = 24'(-924);
			11135: out = 24'(1552);
			11136: out = 24'(4336);
			11137: out = 24'(4472);
			11138: out = 24'(-1272);
			11139: out = 24'(-6160);
			11140: out = 24'(-6040);
			11141: out = 24'(1416);
			11142: out = 24'(5044);
			11143: out = 24'(1036);
			11144: out = 24'(-1548);
			11145: out = 24'(-1144);
			11146: out = 24'(-864);
			11147: out = 24'(3964);
			11148: out = 24'(2180);
			11149: out = 24'(-80);
			11150: out = 24'(-24);
			11151: out = 24'(24);
			11152: out = 24'(576);
			11153: out = 24'(-3136);
			11154: out = 24'(-2208);
			11155: out = 24'(2932);
			11156: out = 24'(3128);
			11157: out = 24'(1276);
			11158: out = 24'(388);
			11159: out = 24'(364);
			11160: out = 24'(-2024);
			11161: out = 24'(-3044);
			11162: out = 24'(-1876);
			11163: out = 24'(-288);
			11164: out = 24'(432);
			11165: out = 24'(-2212);
			11166: out = 24'(-2468);
			11167: out = 24'(508);
			11168: out = 24'(2520);
			11169: out = 24'(3056);
			11170: out = 24'(-4);
			11171: out = 24'(-5560);
			11172: out = 24'(-7428);
			11173: out = 24'(-1024);
			11174: out = 24'(4888);
			11175: out = 24'(3176);
			11176: out = 24'(1496);
			11177: out = 24'(256);
			11178: out = 24'(932);
			11179: out = 24'(-112);
			11180: out = 24'(588);
			11181: out = 24'(264);
			11182: out = 24'(-452);
			11183: out = 24'(-368);
			11184: out = 24'(-1868);
			11185: out = 24'(2760);
			11186: out = 24'(4188);
			11187: out = 24'(-472);
			11188: out = 24'(-2764);
			11189: out = 24'(-1292);
			11190: out = 24'(1532);
			11191: out = 24'(2740);
			11192: out = 24'(1888);
			11193: out = 24'(1084);
			11194: out = 24'(-636);
			11195: out = 24'(-1316);
			11196: out = 24'(-460);
			11197: out = 24'(1056);
			11198: out = 24'(1324);
			11199: out = 24'(-1696);
			11200: out = 24'(-3692);
			11201: out = 24'(-860);
			11202: out = 24'(2780);
			11203: out = 24'(796);
			11204: out = 24'(-5972);
			11205: out = 24'(-5552);
			11206: out = 24'(-596);
			11207: out = 24'(2536);
			11208: out = 24'(2560);
			11209: out = 24'(1268);
			11210: out = 24'(1492);
			11211: out = 24'(-4);
			11212: out = 24'(-1932);
			11213: out = 24'(-4764);
			11214: out = 24'(-4704);
			11215: out = 24'(-3544);
			11216: out = 24'(-192);
			11217: out = 24'(2976);
			11218: out = 24'(512);
			11219: out = 24'(-228);
			11220: out = 24'(2996);
			11221: out = 24'(2384);
			11222: out = 24'(348);
			11223: out = 24'(-1508);
			11224: out = 24'(-292);
			11225: out = 24'(-40);
			11226: out = 24'(340);
			11227: out = 24'(1644);
			11228: out = 24'(-404);
			11229: out = 24'(-4356);
			11230: out = 24'(-3400);
			11231: out = 24'(916);
			11232: out = 24'(2280);
			11233: out = 24'(2484);
			11234: out = 24'(-564);
			11235: out = 24'(112);
			11236: out = 24'(-448);
			11237: out = 24'(-1676);
			11238: out = 24'(88);
			11239: out = 24'(-832);
			11240: out = 24'(-1068);
			11241: out = 24'(1640);
			11242: out = 24'(-80);
			11243: out = 24'(-4372);
			11244: out = 24'(-5324);
			11245: out = 24'(-1624);
			11246: out = 24'(2092);
			11247: out = 24'(4104);
			11248: out = 24'(4472);
			11249: out = 24'(1452);
			11250: out = 24'(-2720);
			11251: out = 24'(-6040);
			11252: out = 24'(-4260);
			11253: out = 24'(-1784);
			11254: out = 24'(212);
			11255: out = 24'(3376);
			11256: out = 24'(1028);
			11257: out = 24'(-2640);
			11258: out = 24'(-928);
			11259: out = 24'(2888);
			11260: out = 24'(5268);
			11261: out = 24'(896);
			11262: out = 24'(-3428);
			11263: out = 24'(-3292);
			11264: out = 24'(-308);
			11265: out = 24'(2680);
			11266: out = 24'(1232);
			11267: out = 24'(-1008);
			11268: out = 24'(-2036);
			11269: out = 24'(372);
			11270: out = 24'(620);
			11271: out = 24'(-856);
			11272: out = 24'(1020);
			11273: out = 24'(692);
			11274: out = 24'(1924);
			11275: out = 24'(2180);
			11276: out = 24'(176);
			11277: out = 24'(1732);
			11278: out = 24'(1620);
			11279: out = 24'(-24);
			11280: out = 24'(-1540);
			11281: out = 24'(-2140);
			11282: out = 24'(-1052);
			11283: out = 24'(-908);
			11284: out = 24'(-236);
			11285: out = 24'(-64);
			11286: out = 24'(-352);
			11287: out = 24'(-164);
			11288: out = 24'(808);
			11289: out = 24'(460);
			11290: out = 24'(-344);
			11291: out = 24'(-2044);
			11292: out = 24'(880);
			11293: out = 24'(2532);
			11294: out = 24'(-1044);
			11295: out = 24'(-4828);
			11296: out = 24'(-2744);
			11297: out = 24'(52);
			11298: out = 24'(-644);
			11299: out = 24'(-1148);
			11300: out = 24'(1516);
			11301: out = 24'(1496);
			11302: out = 24'(-1688);
			11303: out = 24'(-2784);
			11304: out = 24'(-920);
			11305: out = 24'(-708);
			11306: out = 24'(1180);
			11307: out = 24'(3028);
			11308: out = 24'(896);
			11309: out = 24'(-2888);
			11310: out = 24'(-3120);
			11311: out = 24'(-56);
			11312: out = 24'(2168);
			11313: out = 24'(-44);
			11314: out = 24'(324);
			11315: out = 24'(448);
			11316: out = 24'(-860);
			11317: out = 24'(60);
			11318: out = 24'(244);
			11319: out = 24'(956);
			11320: out = 24'(1656);
			11321: out = 24'(-796);
			11322: out = 24'(-2340);
			11323: out = 24'(-2012);
			11324: out = 24'(-2668);
			11325: out = 24'(-612);
			11326: out = 24'(2536);
			11327: out = 24'(-644);
			11328: out = 24'(-3888);
			11329: out = 24'(-2252);
			11330: out = 24'(-1608);
			11331: out = 24'(2524);
			11332: out = 24'(5708);
			11333: out = 24'(2436);
			11334: out = 24'(-2808);
			11335: out = 24'(-5296);
			11336: out = 24'(-2452);
			11337: out = 24'(776);
			11338: out = 24'(2796);
			11339: out = 24'(1180);
			11340: out = 24'(244);
			11341: out = 24'(2084);
			11342: out = 24'(1736);
			11343: out = 24'(-468);
			11344: out = 24'(-508);
			11345: out = 24'(-860);
			11346: out = 24'(332);
			11347: out = 24'(480);
			11348: out = 24'(984);
			11349: out = 24'(-348);
			11350: out = 24'(-848);
			11351: out = 24'(-856);
			11352: out = 24'(1032);
			11353: out = 24'(2400);
			11354: out = 24'(-104);
			11355: out = 24'(-2940);
			11356: out = 24'(-972);
			11357: out = 24'(20);
			11358: out = 24'(-1684);
			11359: out = 24'(-2124);
			11360: out = 24'(-2072);
			11361: out = 24'(1480);
			11362: out = 24'(3392);
			11363: out = 24'(3244);
			11364: out = 24'(872);
			11365: out = 24'(-1396);
			11366: out = 24'(-1480);
			11367: out = 24'(-1612);
			11368: out = 24'(-72);
			11369: out = 24'(268);
			11370: out = 24'(-2296);
			11371: out = 24'(372);
			11372: out = 24'(3668);
			11373: out = 24'(-272);
			11374: out = 24'(-3212);
			11375: out = 24'(-2264);
			11376: out = 24'(1592);
			11377: out = 24'(2212);
			11378: out = 24'(-784);
			11379: out = 24'(532);
			11380: out = 24'(1536);
			11381: out = 24'(2116);
			11382: out = 24'(2244);
			11383: out = 24'(1440);
			11384: out = 24'(-716);
			11385: out = 24'(-1664);
			11386: out = 24'(-3144);
			11387: out = 24'(-1064);
			11388: out = 24'(1248);
			11389: out = 24'(-916);
			11390: out = 24'(-3932);
			11391: out = 24'(-2712);
			11392: out = 24'(-1092);
			11393: out = 24'(12);
			11394: out = 24'(2524);
			11395: out = 24'(2856);
			11396: out = 24'(-124);
			11397: out = 24'(-2252);
			11398: out = 24'(-4532);
			11399: out = 24'(-2724);
			11400: out = 24'(2168);
			11401: out = 24'(4248);
			11402: out = 24'(2144);
			11403: out = 24'(-1040);
			11404: out = 24'(-2664);
			11405: out = 24'(252);
			11406: out = 24'(3388);
			11407: out = 24'(3176);
			11408: out = 24'(652);
			11409: out = 24'(-1820);
			11410: out = 24'(-2392);
			11411: out = 24'(-2300);
			11412: out = 24'(-512);
			11413: out = 24'(268);
			11414: out = 24'(-1236);
			11415: out = 24'(-176);
			11416: out = 24'(276);
			11417: out = 24'(584);
			11418: out = 24'(776);
			11419: out = 24'(1624);
			11420: out = 24'(3156);
			11421: out = 24'(1720);
			11422: out = 24'(-248);
			11423: out = 24'(-1392);
			11424: out = 24'(-216);
			11425: out = 24'(1388);
			11426: out = 24'(-128);
			11427: out = 24'(-1736);
			11428: out = 24'(372);
			11429: out = 24'(556);
			11430: out = 24'(-1628);
			11431: out = 24'(-1800);
			11432: out = 24'(-1984);
			11433: out = 24'(-696);
			11434: out = 24'(-888);
			11435: out = 24'(424);
			11436: out = 24'(1824);
			11437: out = 24'(1224);
			11438: out = 24'(1132);
			11439: out = 24'(1628);
			11440: out = 24'(-232);
			11441: out = 24'(-2904);
			11442: out = 24'(-1344);
			11443: out = 24'(876);
			11444: out = 24'(1056);
			11445: out = 24'(-1588);
			11446: out = 24'(-1324);
			11447: out = 24'(652);
			11448: out = 24'(1112);
			11449: out = 24'(816);
			11450: out = 24'(-944);
			11451: out = 24'(-1112);
			11452: out = 24'(-216);
			11453: out = 24'(2484);
			11454: out = 24'(2188);
			11455: out = 24'(-1108);
			11456: out = 24'(-3192);
			11457: out = 24'(-288);
			11458: out = 24'(2216);
			11459: out = 24'(1580);
			11460: out = 24'(-2760);
			11461: out = 24'(-2092);
			11462: out = 24'(936);
			11463: out = 24'(724);
			11464: out = 24'(3400);
			11465: out = 24'(4328);
			11466: out = 24'(1312);
			11467: out = 24'(-3712);
			11468: out = 24'(-5200);
			11469: out = 24'(-3320);
			11470: out = 24'(1440);
			11471: out = 24'(2340);
			11472: out = 24'(-212);
			11473: out = 24'(-692);
			11474: out = 24'(544);
			11475: out = 24'(-752);
			11476: out = 24'(-1416);
			11477: out = 24'(-3128);
			11478: out = 24'(-2140);
			11479: out = 24'(848);
			11480: out = 24'(3112);
			11481: out = 24'(2684);
			11482: out = 24'(-48);
			11483: out = 24'(208);
			11484: out = 24'(1868);
			11485: out = 24'(1828);
			11486: out = 24'(-2012);
			11487: out = 24'(-4324);
			11488: out = 24'(-1344);
			11489: out = 24'(1752);
			11490: out = 24'(-92);
			11491: out = 24'(-2272);
			11492: out = 24'(-1440);
			11493: out = 24'(2360);
			11494: out = 24'(3424);
			11495: out = 24'(-40);
			11496: out = 24'(-1004);
			11497: out = 24'(196);
			11498: out = 24'(1848);
			11499: out = 24'(2240);
			11500: out = 24'(1448);
			11501: out = 24'(-192);
			11502: out = 24'(-2248);
			11503: out = 24'(-3976);
			11504: out = 24'(-3012);
			11505: out = 24'(884);
			11506: out = 24'(2420);
			11507: out = 24'(-1384);
			11508: out = 24'(-3124);
			11509: out = 24'(-432);
			11510: out = 24'(520);
			11511: out = 24'(1352);
			11512: out = 24'(2924);
			11513: out = 24'(2760);
			11514: out = 24'(-1340);
			11515: out = 24'(-3528);
			11516: out = 24'(-2568);
			11517: out = 24'(-96);
			11518: out = 24'(528);
			11519: out = 24'(-572);
			11520: out = 24'(-984);
			11521: out = 24'(608);
			11522: out = 24'(856);
			11523: out = 24'(-344);
			11524: out = 24'(-840);
			11525: out = 24'(-504);
			11526: out = 24'(1128);
			11527: out = 24'(1392);
			11528: out = 24'(-988);
			11529: out = 24'(-932);
			11530: out = 24'(-92);
			11531: out = 24'(1232);
			11532: out = 24'(1688);
			11533: out = 24'(-460);
			11534: out = 24'(-1160);
			11535: out = 24'(-736);
			11536: out = 24'(1648);
			11537: out = 24'(3176);
			11538: out = 24'(1308);
			11539: out = 24'(-2176);
			11540: out = 24'(-3344);
			11541: out = 24'(-1856);
			11542: out = 24'(1072);
			11543: out = 24'(2428);
			11544: out = 24'(1076);
			11545: out = 24'(-612);
			11546: out = 24'(-740);
			11547: out = 24'(-44);
			11548: out = 24'(-2428);
			11549: out = 24'(-3312);
			11550: out = 24'(-1568);
			11551: out = 24'(780);
			11552: out = 24'(1348);
			11553: out = 24'(2160);
			11554: out = 24'(3044);
			11555: out = 24'(1260);
			11556: out = 24'(-1468);
			11557: out = 24'(-3160);
			11558: out = 24'(-2572);
			11559: out = 24'(-876);
			11560: out = 24'(1172);
			11561: out = 24'(1928);
			11562: out = 24'(516);
			11563: out = 24'(744);
			11564: out = 24'(1496);
			11565: out = 24'(1940);
			11566: out = 24'(-680);
			11567: out = 24'(-2412);
			11568: out = 24'(-2620);
			11569: out = 24'(-532);
			11570: out = 24'(1256);
			11571: out = 24'(108);
			11572: out = 24'(-1972);
			11573: out = 24'(-1696);
			11574: out = 24'(352);
			11575: out = 24'(1112);
			11576: out = 24'(-960);
			11577: out = 24'(-2924);
			11578: out = 24'(-2248);
			11579: out = 24'(172);
			11580: out = 24'(1324);
			11581: out = 24'(884);
			11582: out = 24'(-832);
			11583: out = 24'(-2172);
			11584: out = 24'(-1528);
			11585: out = 24'(-1448);
			11586: out = 24'(512);
			11587: out = 24'(3576);
			11588: out = 24'(2092);
			11589: out = 24'(-760);
			11590: out = 24'(-2152);
			11591: out = 24'(-1016);
			11592: out = 24'(1064);
			11593: out = 24'(-440);
			11594: out = 24'(-876);
			11595: out = 24'(52);
			11596: out = 24'(1036);
			11597: out = 24'(504);
			11598: out = 24'(772);
			11599: out = 24'(660);
			11600: out = 24'(-1528);
			11601: out = 24'(-2872);
			11602: out = 24'(-1764);
			11603: out = 24'(-624);
			11604: out = 24'(1780);
			11605: out = 24'(1460);
			11606: out = 24'(392);
			11607: out = 24'(-164);
			11608: out = 24'(-388);
			11609: out = 24'(560);
			11610: out = 24'(-1188);
			11611: out = 24'(-2408);
			11612: out = 24'(-944);
			11613: out = 24'(1796);
			11614: out = 24'(1716);
			11615: out = 24'(176);
			11616: out = 24'(452);
			11617: out = 24'(312);
			11618: out = 24'(-1580);
			11619: out = 24'(-1472);
			11620: out = 24'(-1196);
			11621: out = 24'(-540);
			11622: out = 24'(-188);
			11623: out = 24'(-196);
			11624: out = 24'(-120);
			11625: out = 24'(-364);
			11626: out = 24'(1596);
			11627: out = 24'(2068);
			11628: out = 24'(-1172);
			11629: out = 24'(-4000);
			11630: out = 24'(-3240);
			11631: out = 24'(-1252);
			11632: out = 24'(1576);
			11633: out = 24'(2180);
			11634: out = 24'(556);
			11635: out = 24'(-1392);
			11636: out = 24'(-2256);
			11637: out = 24'(136);
			11638: out = 24'(652);
			11639: out = 24'(1932);
			11640: out = 24'(160);
			11641: out = 24'(-1260);
			11642: out = 24'(-1408);
			11643: out = 24'(-212);
			11644: out = 24'(1608);
			11645: out = 24'(864);
			11646: out = 24'(-516);
			11647: out = 24'(732);
			11648: out = 24'(720);
			11649: out = 24'(-436);
			11650: out = 24'(-1484);
			11651: out = 24'(-1940);
			11652: out = 24'(-1756);
			11653: out = 24'(-2348);
			11654: out = 24'(-428);
			11655: out = 24'(1664);
			11656: out = 24'(-188);
			11657: out = 24'(-808);
			11658: out = 24'(1188);
			11659: out = 24'(224);
			11660: out = 24'(-2836);
			11661: out = 24'(-4444);
			11662: out = 24'(-2084);
			11663: out = 24'(-120);
			11664: out = 24'(2040);
			11665: out = 24'(2132);
			11666: out = 24'(-488);
			11667: out = 24'(-372);
			11668: out = 24'(-748);
			11669: out = 24'(1016);
			11670: out = 24'(1136);
			11671: out = 24'(76);
			11672: out = 24'(-40);
			11673: out = 24'(-720);
			11674: out = 24'(-608);
			11675: out = 24'(148);
			11676: out = 24'(-48);
			11677: out = 24'(-2132);
			11678: out = 24'(-1900);
			11679: out = 24'(-764);
			11680: out = 24'(-844);
			11681: out = 24'(392);
			11682: out = 24'(1680);
			11683: out = 24'(-124);
			11684: out = 24'(-912);
			11685: out = 24'(136);
			11686: out = 24'(-492);
			11687: out = 24'(676);
			11688: out = 24'(-924);
			11689: out = 24'(-228);
			11690: out = 24'(720);
			11691: out = 24'(568);
			11692: out = 24'(1876);
			11693: out = 24'(1784);
			11694: out = 24'(144);
			11695: out = 24'(-2264);
			11696: out = 24'(-2248);
			11697: out = 24'(-2588);
			11698: out = 24'(-248);
			11699: out = 24'(692);
			11700: out = 24'(192);
			11701: out = 24'(960);
			11702: out = 24'(1120);
			11703: out = 24'(104);
			11704: out = 24'(-844);
			11705: out = 24'(240);
			11706: out = 24'(396);
			11707: out = 24'(808);
			11708: out = 24'(-404);
			11709: out = 24'(-1168);
			11710: out = 24'(636);
			11711: out = 24'(2524);
			11712: out = 24'(1176);
			11713: out = 24'(-772);
			11714: out = 24'(192);
			11715: out = 24'(956);
			11716: out = 24'(-560);
			11717: out = 24'(-1348);
			11718: out = 24'(-1272);
			11719: out = 24'(-868);
			11720: out = 24'(264);
			11721: out = 24'(-652);
			11722: out = 24'(-1068);
			11723: out = 24'(656);
			11724: out = 24'(2212);
			11725: out = 24'(1128);
			11726: out = 24'(-1724);
			11727: out = 24'(-1844);
			11728: out = 24'(-96);
			11729: out = 24'(812);
			11730: out = 24'(-160);
			11731: out = 24'(1156);
			11732: out = 24'(2660);
			11733: out = 24'(1184);
			11734: out = 24'(-1812);
			11735: out = 24'(-2292);
			11736: out = 24'(-264);
			11737: out = 24'(2444);
			11738: out = 24'(352);
			11739: out = 24'(-2116);
			11740: out = 24'(-812);
			11741: out = 24'(228);
			11742: out = 24'(-1668);
			11743: out = 24'(-2684);
			11744: out = 24'(-1196);
			default: out = 0;
		endcase
	end
endmodule
