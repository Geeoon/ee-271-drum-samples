module ride_lookup(index, out);
	input logic unsigned [13:0] index;
	output logic signed [15:0] out;
	always_comb begin
		case(index)
			0: out = 16'(0);
			1: out = 16'(16);
			2: out = 16'(71);
			3: out = 16'(21);
			4: out = 16'(8299);
			5: out = 16'(-26790);
			6: out = 16'(-624);
			7: out = 16'(3163);
			8: out = 16'(-5883);
			9: out = 16'(5972);
			10: out = 16'(-31196);
			11: out = 16'(21790);
			12: out = 16'(-25864);
			13: out = 16'(2007);
			14: out = 16'(-13956);
			15: out = 16'(4175);
			16: out = 16'(9642);
			17: out = 16'(-26317);
			18: out = 16'(19007);
			19: out = 16'(-29177);
			20: out = 16'(22250);
			21: out = 16'(-2054);
			22: out = 16'(-4989);
			23: out = 16'(-15057);
			24: out = 16'(-17665);
			25: out = 16'(-20738);
			26: out = 16'(8190);
			27: out = 16'(17093);
			28: out = 16'(-18636);
			29: out = 16'(13564);
			30: out = 16'(2697);
			31: out = 16'(8495);
			32: out = 16'(-5795);
			33: out = 16'(-2613);
			34: out = 16'(-23140);
			35: out = 16'(-5300);
			36: out = 16'(-680);
			37: out = 16'(26018);
			38: out = 16'(-23367);
			39: out = 16'(8175);
			40: out = 16'(-16412);
			41: out = 16'(6340);
			42: out = 16'(-7810);
			43: out = 16'(5297);
			44: out = 16'(7519);
			45: out = 16'(20595);
			46: out = 16'(16147);
			47: out = 16'(-14115);
			48: out = 16'(22248);
			49: out = 16'(6750);
			50: out = 16'(25234);
			51: out = 16'(-17694);
			52: out = 16'(24999);
			53: out = 16'(3398);
			54: out = 16'(22641);
			55: out = 16'(6667);
			56: out = 16'(-22748);
			57: out = 16'(14724);
			58: out = 16'(10078);
			59: out = 16'(2614);
			60: out = 16'(-1320);
			61: out = 16'(-4799);
			62: out = 16'(13238);
			63: out = 16'(16612);
			64: out = 16'(-28277);
			65: out = 16'(8771);
			66: out = 16'(-10863);
			67: out = 16'(1468);
			68: out = 16'(-1343);
			69: out = 16'(-2697);
			70: out = 16'(-2719);
			71: out = 16'(1543);
			72: out = 16'(7963);
			73: out = 16'(408);
			74: out = 16'(8816);
			75: out = 16'(10841);
			76: out = 16'(7575);
			77: out = 16'(-27354);
			78: out = 16'(20557);
			79: out = 16'(-29317);
			80: out = 16'(-3562);
			81: out = 16'(-26384);
			82: out = 16'(17278);
			83: out = 16'(-11522);
			84: out = 16'(-15799);
			85: out = 16'(-7166);
			86: out = 16'(20210);
			87: out = 16'(38);
			88: out = 16'(-14457);
			89: out = 16'(11991);
			90: out = 16'(10189);
			91: out = 16'(-5812);
			92: out = 16'(-6526);
			93: out = 16'(379);
			94: out = 16'(-5247);
			95: out = 16'(3098);
			96: out = 16'(-1144);
			97: out = 16'(-6261);
			98: out = 16'(-2194);
			99: out = 16'(-11106);
			100: out = 16'(10982);
			101: out = 16'(-16645);
			102: out = 16'(-16832);
			103: out = 16'(13351);
			104: out = 16'(2838);
			105: out = 16'(4317);
			106: out = 16'(1395);
			107: out = 16'(-1717);
			108: out = 16'(21583);
			109: out = 16'(3234);
			110: out = 16'(-425);
			111: out = 16'(19207);
			112: out = 16'(5406);
			113: out = 16'(-22000);
			114: out = 16'(-24067);
			115: out = 16'(6810);
			116: out = 16'(-24610);
			117: out = 16'(13427);
			118: out = 16'(-1911);
			119: out = 16'(9847);
			120: out = 16'(-18364);
			121: out = 16'(23047);
			122: out = 16'(2101);
			123: out = 16'(26178);
			124: out = 16'(3243);
			125: out = 16'(3066);
			126: out = 16'(-1511);
			127: out = 16'(5066);
			128: out = 16'(10461);
			129: out = 16'(14004);
			130: out = 16'(-15568);
			131: out = 16'(8341);
			132: out = 16'(-5789);
			133: out = 16'(-26587);
			134: out = 16'(8926);
			135: out = 16'(-2664);
			136: out = 16'(5126);
			137: out = 16'(-15759);
			138: out = 16'(3539);
			139: out = 16'(-5895);
			140: out = 16'(5436);
			141: out = 16'(15857);
			142: out = 16'(10115);
			143: out = 16'(-16394);
			144: out = 16'(-4470);
			145: out = 16'(15123);
			146: out = 16'(-16935);
			147: out = 16'(1738);
			148: out = 16'(592);
			149: out = 16'(8633);
			150: out = 16'(-934);
			151: out = 16'(-6663);
			152: out = 16'(2574);
			153: out = 16'(11477);
			154: out = 16'(6832);
			155: out = 16'(3368);
			156: out = 16'(-17527);
			157: out = 16'(1880);
			158: out = 16'(8037);
			159: out = 16'(-16673);
			160: out = 16'(1525);
			161: out = 16'(-9438);
			162: out = 16'(-8661);
			163: out = 16'(-9745);
			164: out = 16'(3644);
			165: out = 16'(15444);
			166: out = 16'(15004);
			167: out = 16'(15153);
			168: out = 16'(-1898);
			169: out = 16'(-3315);
			170: out = 16'(-4293);
			171: out = 16'(-14807);
			172: out = 16'(5719);
			173: out = 16'(-12136);
			174: out = 16'(6608);
			175: out = 16'(5395);
			176: out = 16'(-10127);
			177: out = 16'(13928);
			178: out = 16'(2518);
			179: out = 16'(15536);
			180: out = 16'(-3612);
			181: out = 16'(9514);
			182: out = 16'(-6249);
			183: out = 16'(-4763);
			184: out = 16'(-1265);
			185: out = 16'(9949);
			186: out = 16'(7851);
			187: out = 16'(18575);
			188: out = 16'(-7106);
			189: out = 16'(-2613);
			190: out = 16'(13732);
			191: out = 16'(9462);
			192: out = 16'(-12435);
			193: out = 16'(-10320);
			194: out = 16'(942);
			195: out = 16'(-4916);
			196: out = 16'(-11603);
			197: out = 16'(-5399);
			198: out = 16'(7638);
			199: out = 16'(-7220);
			200: out = 16'(13479);
			201: out = 16'(10165);
			202: out = 16'(-4084);
			203: out = 16'(-9470);
			204: out = 16'(17842);
			205: out = 16'(213);
			206: out = 16'(4766);
			207: out = 16'(100);
			208: out = 16'(4089);
			209: out = 16'(14373);
			210: out = 16'(15055);
			211: out = 16'(-8000);
			212: out = 16'(-1741);
			213: out = 16'(-2928);
			214: out = 16'(-23796);
			215: out = 16'(-3763);
			216: out = 16'(-11123);
			217: out = 16'(-8922);
			218: out = 16'(-17469);
			219: out = 16'(-6098);
			220: out = 16'(-4962);
			221: out = 16'(-438);
			222: out = 16'(-13367);
			223: out = 16'(6107);
			224: out = 16'(7171);
			225: out = 16'(-13454);
			226: out = 16'(-3973);
			227: out = 16'(864);
			228: out = 16'(-7920);
			229: out = 16'(-862);
			230: out = 16'(11608);
			231: out = 16'(7396);
			232: out = 16'(-20754);
			233: out = 16'(1958);
			234: out = 16'(11791);
			235: out = 16'(-10101);
			236: out = 16'(17616);
			237: out = 16'(-6445);
			238: out = 16'(-10599);
			239: out = 16'(6415);
			240: out = 16'(4301);
			241: out = 16'(19293);
			242: out = 16'(-11795);
			243: out = 16'(-5051);
			244: out = 16'(19978);
			245: out = 16'(-797);
			246: out = 16'(-7121);
			247: out = 16'(5121);
			248: out = 16'(-10038);
			249: out = 16'(12218);
			250: out = 16'(-4155);
			251: out = 16'(4287);
			252: out = 16'(-3429);
			253: out = 16'(14223);
			254: out = 16'(-1789);
			255: out = 16'(1775);
			256: out = 16'(-8838);
			257: out = 16'(9355);
			258: out = 16'(-7934);
			259: out = 16'(3395);
			260: out = 16'(14954);
			261: out = 16'(-11827);
			262: out = 16'(7552);
			263: out = 16'(-15894);
			264: out = 16'(1968);
			265: out = 16'(-8344);
			266: out = 16'(18115);
			267: out = 16'(1903);
			268: out = 16'(-25387);
			269: out = 16'(-26572);
			270: out = 16'(9608);
			271: out = 16'(-14714);
			272: out = 16'(-6426);
			273: out = 16'(-26374);
			274: out = 16'(3319);
			275: out = 16'(-16895);
			276: out = 16'(-2066);
			277: out = 16'(-9452);
			278: out = 16'(18652);
			279: out = 16'(10183);
			280: out = 16'(-10286);
			281: out = 16'(-9852);
			282: out = 16'(-483);
			283: out = 16'(4106);
			284: out = 16'(9405);
			285: out = 16'(-2773);
			286: out = 16'(22000);
			287: out = 16'(-15447);
			288: out = 16'(829);
			289: out = 16'(12452);
			290: out = 16'(3841);
			291: out = 16'(-12384);
			292: out = 16'(9983);
			293: out = 16'(429);
			294: out = 16'(1236);
			295: out = 16'(-8672);
			296: out = 16'(-3202);
			297: out = 16'(3180);
			298: out = 16'(487);
			299: out = 16'(13238);
			300: out = 16'(2931);
			301: out = 16'(726);
			302: out = 16'(7078);
			303: out = 16'(19172);
			304: out = 16'(-6171);
			305: out = 16'(311);
			306: out = 16'(10211);
			307: out = 16'(6824);
			308: out = 16'(22907);
			309: out = 16'(-8337);
			310: out = 16'(14548);
			311: out = 16'(-11988);
			312: out = 16'(19937);
			313: out = 16'(2006);
			314: out = 16'(-2294);
			315: out = 16'(-21186);
			316: out = 16'(8355);
			317: out = 16'(-15239);
			318: out = 16'(-7797);
			319: out = 16'(71);
			320: out = 16'(5813);
			321: out = 16'(9924);
			322: out = 16'(1432);
			323: out = 16'(7952);
			324: out = 16'(-1327);
			325: out = 16'(-8255);
			326: out = 16'(1994);
			327: out = 16'(1910);
			328: out = 16'(4175);
			329: out = 16'(19753);
			330: out = 16'(6695);
			331: out = 16'(16644);
			332: out = 16'(-20723);
			333: out = 16'(-18481);
			334: out = 16'(5426);
			335: out = 16'(6100);
			336: out = 16'(1203);
			337: out = 16'(1599);
			338: out = 16'(644);
			339: out = 16'(-10383);
			340: out = 16'(-14369);
			341: out = 16'(-2462);
			342: out = 16'(10091);
			343: out = 16'(-4111);
			344: out = 16'(-20100);
			345: out = 16'(-10525);
			346: out = 16'(9599);
			347: out = 16'(-22061);
			348: out = 16'(4942);
			349: out = 16'(13672);
			350: out = 16'(-7404);
			351: out = 16'(-15913);
			352: out = 16'(23318);
			353: out = 16'(6640);
			354: out = 16'(-18560);
			355: out = 16'(1756);
			356: out = 16'(10927);
			357: out = 16'(9011);
			358: out = 16'(-3473);
			359: out = 16'(19700);
			360: out = 16'(-3979);
			361: out = 16'(-3137);
			362: out = 16'(6288);
			363: out = 16'(8843);
			364: out = 16'(10369);
			365: out = 16'(-9938);
			366: out = 16'(11808);
			367: out = 16'(22725);
			368: out = 16'(-8998);
			369: out = 16'(-4456);
			370: out = 16'(4462);
			371: out = 16'(9595);
			372: out = 16'(-10354);
			373: out = 16'(-816);
			374: out = 16'(6469);
			375: out = 16'(5488);
			376: out = 16'(-15375);
			377: out = 16'(356);
			378: out = 16'(4082);
			379: out = 16'(9221);
			380: out = 16'(2850);
			381: out = 16'(23304);
			382: out = 16'(15399);
			383: out = 16'(-15062);
			384: out = 16'(6733);
			385: out = 16'(5822);
			386: out = 16'(17050);
			387: out = 16'(-15988);
			388: out = 16'(7047);
			389: out = 16'(875);
			390: out = 16'(5381);
			391: out = 16'(-21712);
			392: out = 16'(17929);
			393: out = 16'(-12730);
			394: out = 16'(-9079);
			395: out = 16'(641);
			396: out = 16'(-30798);
			397: out = 16'(-14805);
			398: out = 16'(1387);
			399: out = 16'(-1355);
			400: out = 16'(1610);
			401: out = 16'(-18833);
			402: out = 16'(-5325);
			403: out = 16'(-463);
			404: out = 16'(11268);
			405: out = 16'(4708);
			406: out = 16'(-19594);
			407: out = 16'(12449);
			408: out = 16'(-7167);
			409: out = 16'(-10177);
			410: out = 16'(-10382);
			411: out = 16'(20044);
			412: out = 16'(6817);
			413: out = 16'(-22538);
			414: out = 16'(-22101);
			415: out = 16'(2897);
			416: out = 16'(-245);
			417: out = 16'(-16608);
			418: out = 16'(11247);
			419: out = 16'(-13641);
			420: out = 16'(9033);
			421: out = 16'(1748);
			422: out = 16'(15412);
			423: out = 16'(-8702);
			424: out = 16'(-1481);
			425: out = 16'(-730);
			426: out = 16'(21765);
			427: out = 16'(218);
			428: out = 16'(-8273);
			429: out = 16'(8303);
			430: out = 16'(-1095);
			431: out = 16'(16990);
			432: out = 16'(-16108);
			433: out = 16'(20580);
			434: out = 16'(-6309);
			435: out = 16'(6341);
			436: out = 16'(-10621);
			437: out = 16'(15980);
			438: out = 16'(4616);
			439: out = 16'(3196);
			440: out = 16'(12762);
			441: out = 16'(4864);
			442: out = 16'(-7383);
			443: out = 16'(5483);
			444: out = 16'(17524);
			445: out = 16'(914);
			446: out = 16'(-21651);
			447: out = 16'(2565);
			448: out = 16'(11365);
			449: out = 16'(9486);
			450: out = 16'(-4675);
			451: out = 16'(3047);
			452: out = 16'(-2099);
			453: out = 16'(-18384);
			454: out = 16'(6909);
			455: out = 16'(5053);
			456: out = 16'(9189);
			457: out = 16'(-314);
			458: out = 16'(9463);
			459: out = 16'(4399);
			460: out = 16'(-17743);
			461: out = 16'(5998);
			462: out = 16'(7373);
			463: out = 16'(12385);
			464: out = 16'(-9601);
			465: out = 16'(-2934);
			466: out = 16'(-1816);
			467: out = 16'(-6713);
			468: out = 16'(-31592);
			469: out = 16'(1913);
			470: out = 16'(15132);
			471: out = 16'(-6562);
			472: out = 16'(-8799);
			473: out = 16'(-22498);
			474: out = 16'(-13891);
			475: out = 16'(-18650);
			476: out = 16'(1420);
			477: out = 16'(-12668);
			478: out = 16'(-4103);
			479: out = 16'(-5713);
			480: out = 16'(-15720);
			481: out = 16'(-5340);
			482: out = 16'(10055);
			483: out = 16'(-12640);
			484: out = 16'(91);
			485: out = 16'(19498);
			486: out = 16'(-2298);
			487: out = 16'(3609);
			488: out = 16'(-18464);
			489: out = 16'(16123);
			490: out = 16'(-6193);
			491: out = 16'(4307);
			492: out = 16'(11468);
			493: out = 16'(-267);
			494: out = 16'(12505);
			495: out = 16'(-22211);
			496: out = 16'(6954);
			497: out = 16'(-23619);
			498: out = 16'(-9827);
			499: out = 16'(-2817);
			500: out = 16'(932);
			501: out = 16'(4156);
			502: out = 16'(11225);
			503: out = 16'(12055);
			504: out = 16'(5360);
			505: out = 16'(8666);
			506: out = 16'(-6108);
			507: out = 16'(16460);
			508: out = 16'(19950);
			509: out = 16'(7450);
			510: out = 16'(24082);
			511: out = 16'(-13752);
			512: out = 16'(19656);
			513: out = 16'(9456);
			514: out = 16'(11341);
			515: out = 16'(12773);
			516: out = 16'(-1073);
			517: out = 16'(6840);
			518: out = 16'(-3053);
			519: out = 16'(21417);
			520: out = 16'(-3949);
			521: out = 16'(4004);
			522: out = 16'(-1219);
			523: out = 16'(-1996);
			524: out = 16'(9105);
			525: out = 16'(3187);
			526: out = 16'(-653);
			527: out = 16'(12759);
			528: out = 16'(7951);
			529: out = 16'(6346);
			530: out = 16'(16607);
			531: out = 16'(639);
			532: out = 16'(-4467);
			533: out = 16'(5699);
			534: out = 16'(5772);
			535: out = 16'(-5589);
			536: out = 16'(253);
			537: out = 16'(15591);
			538: out = 16'(-10365);
			539: out = 16'(-20685);
			540: out = 16'(-11674);
			541: out = 16'(3338);
			542: out = 16'(5253);
			543: out = 16'(-6163);
			544: out = 16'(813);
			545: out = 16'(-2781);
			546: out = 16'(-9373);
			547: out = 16'(727);
			548: out = 16'(2321);
			549: out = 16'(182);
			550: out = 16'(3881);
			551: out = 16'(-25128);
			552: out = 16'(9157);
			553: out = 16'(-5851);
			554: out = 16'(10475);
			555: out = 16'(3987);
			556: out = 16'(-17033);
			557: out = 16'(-24525);
			558: out = 16'(-2721);
			559: out = 16'(15281);
			560: out = 16'(-19814);
			561: out = 16'(635);
			562: out = 16'(-25361);
			563: out = 16'(1949);
			564: out = 16'(9158);
			565: out = 16'(-3412);
			566: out = 16'(-882);
			567: out = 16'(-14287);
			568: out = 16'(13223);
			569: out = 16'(10600);
			570: out = 16'(-4030);
			571: out = 16'(-16992);
			572: out = 16'(5781);
			573: out = 16'(10848);
			574: out = 16'(-9213);
			575: out = 16'(7443);
			576: out = 16'(-5009);
			577: out = 16'(-12760);
			578: out = 16'(-5841);
			579: out = 16'(2473);
			580: out = 16'(9815);
			581: out = 16'(-31086);
			582: out = 16'(4347);
			583: out = 16'(-27819);
			584: out = 16'(-2405);
			585: out = 16'(-8684);
			586: out = 16'(17069);
			587: out = 16'(1729);
			588: out = 16'(-26619);
			589: out = 16'(-10043);
			590: out = 16'(6829);
			591: out = 16'(-13657);
			592: out = 16'(1830);
			593: out = 16'(20733);
			594: out = 16'(935);
			595: out = 16'(6686);
			596: out = 16'(3815);
			597: out = 16'(13057);
			598: out = 16'(-15);
			599: out = 16'(8363);
			600: out = 16'(6563);
			601: out = 16'(15483);
			602: out = 16'(-7020);
			603: out = 16'(3840);
			604: out = 16'(14787);
			605: out = 16'(6430);
			606: out = 16'(1805);
			607: out = 16'(-11154);
			608: out = 16'(-14473);
			609: out = 16'(-7581);
			610: out = 16'(2069);
			611: out = 16'(17230);
			612: out = 16'(-6297);
			613: out = 16'(-304);
			614: out = 16'(17644);
			615: out = 16'(-8767);
			616: out = 16'(-11502);
			617: out = 16'(-476);
			618: out = 16'(2632);
			619: out = 16'(8411);
			620: out = 16'(21261);
			621: out = 16'(13600);
			622: out = 16'(-2350);
			623: out = 16'(-3907);
			624: out = 16'(-6399);
			625: out = 16'(21894);
			626: out = 16'(-896);
			627: out = 16'(-1865);
			628: out = 16'(-13861);
			629: out = 16'(11500);
			630: out = 16'(-24005);
			631: out = 16'(-8360);
			632: out = 16'(19535);
			633: out = 16'(5894);
			634: out = 16'(-882);
			635: out = 16'(17910);
			636: out = 16'(7267);
			637: out = 16'(-7870);
			638: out = 16'(8727);
			639: out = 16'(5724);
			640: out = 16'(21220);
			641: out = 16'(-16089);
			642: out = 16'(17518);
			643: out = 16'(10187);
			644: out = 16'(9575);
			645: out = 16'(4508);
			646: out = 16'(12807);
			647: out = 16'(382);
			648: out = 16'(-8005);
			649: out = 16'(9);
			650: out = 16'(9930);
			651: out = 16'(4844);
			652: out = 16'(-28756);
			653: out = 16'(15781);
			654: out = 16'(-5473);
			655: out = 16'(3994);
			656: out = 16'(2675);
			657: out = 16'(12760);
			658: out = 16'(6779);
			659: out = 16'(2798);
			660: out = 16'(-48);
			661: out = 16'(-1970);
			662: out = 16'(176);
			663: out = 16'(836);
			664: out = 16'(-7536);
			665: out = 16'(12546);
			666: out = 16'(7557);
			667: out = 16'(5992);
			668: out = 16'(-2236);
			669: out = 16'(-26132);
			670: out = 16'(24747);
			671: out = 16'(-8887);
			672: out = 16'(457);
			673: out = 16'(1523);
			674: out = 16'(-18409);
			675: out = 16'(4916);
			676: out = 16'(-13429);
			677: out = 16'(14324);
			678: out = 16'(-13322);
			679: out = 16'(88);
			680: out = 16'(-1945);
			681: out = 16'(13420);
			682: out = 16'(-1776);
			683: out = 16'(-19325);
			684: out = 16'(14136);
			685: out = 16'(-22242);
			686: out = 16'(8204);
			687: out = 16'(-7696);
			688: out = 16'(12698);
			689: out = 16'(-30438);
			690: out = 16'(-21775);
			691: out = 16'(17142);
			692: out = 16'(10560);
			693: out = 16'(8288);
			694: out = 16'(-1150);
			695: out = 16'(-9332);
			696: out = 16'(2659);
			697: out = 16'(11664);
			698: out = 16'(-8517);
			699: out = 16'(4886);
			700: out = 16'(-4142);
			701: out = 16'(-7677);
			702: out = 16'(-2436);
			703: out = 16'(-6758);
			704: out = 16'(-7659);
			705: out = 16'(17795);
			706: out = 16'(-15387);
			707: out = 16'(1760);
			708: out = 16'(-6013);
			709: out = 16'(-16355);
			710: out = 16'(9837);
			711: out = 16'(2222);
			712: out = 16'(-2496);
			713: out = 16'(-3902);
			714: out = 16'(8232);
			715: out = 16'(7048);
			716: out = 16'(-5463);
			717: out = 16'(1717);
			718: out = 16'(10839);
			719: out = 16'(-9128);
			720: out = 16'(1482);
			721: out = 16'(8684);
			722: out = 16'(5829);
			723: out = 16'(-3130);
			724: out = 16'(1104);
			725: out = 16'(-1264);
			726: out = 16'(-7981);
			727: out = 16'(-1860);
			728: out = 16'(-15574);
			729: out = 16'(12805);
			730: out = 16'(-19872);
			731: out = 16'(11417);
			732: out = 16'(3170);
			733: out = 16'(8008);
			734: out = 16'(-2589);
			735: out = 16'(-13677);
			736: out = 16'(-2446);
			737: out = 16'(1147);
			738: out = 16'(13682);
			739: out = 16'(-14708);
			740: out = 16'(13185);
			741: out = 16'(-19884);
			742: out = 16'(6577);
			743: out = 16'(4097);
			744: out = 16'(-4046);
			745: out = 16'(8538);
			746: out = 16'(-11811);
			747: out = 16'(3541);
			748: out = 16'(-2718);
			749: out = 16'(-1971);
			750: out = 16'(-12155);
			751: out = 16'(-22547);
			752: out = 16'(412);
			753: out = 16'(-2281);
			754: out = 16'(-9750);
			755: out = 16'(1857);
			756: out = 16'(2877);
			757: out = 16'(6734);
			758: out = 16'(1311);
			759: out = 16'(3804);
			760: out = 16'(3975);
			761: out = 16'(6078);
			762: out = 16'(-2869);
			763: out = 16'(542);
			764: out = 16'(8188);
			765: out = 16'(-3945);
			766: out = 16'(16399);
			767: out = 16'(-2570);
			768: out = 16'(-8);
			769: out = 16'(-5271);
			770: out = 16'(6581);
			771: out = 16'(18639);
			772: out = 16'(110);
			773: out = 16'(-10731);
			774: out = 16'(1512);
			775: out = 16'(-2217);
			776: out = 16'(12305);
			777: out = 16'(-3451);
			778: out = 16'(20794);
			779: out = 16'(-13428);
			780: out = 16'(3941);
			781: out = 16'(11381);
			782: out = 16'(3324);
			783: out = 16'(5173);
			784: out = 16'(-7381);
			785: out = 16'(-1780);
			786: out = 16'(-5443);
			787: out = 16'(3036);
			788: out = 16'(8215);
			789: out = 16'(-2249);
			790: out = 16'(6606);
			791: out = 16'(-15644);
			792: out = 16'(5349);
			793: out = 16'(18737);
			794: out = 16'(-1954);
			795: out = 16'(3137);
			796: out = 16'(-10146);
			797: out = 16'(6782);
			798: out = 16'(-4234);
			799: out = 16'(11698);
			800: out = 16'(-4046);
			801: out = 16'(5096);
			802: out = 16'(-18663);
			803: out = 16'(-22796);
			804: out = 16'(4791);
			805: out = 16'(3112);
			806: out = 16'(1426);
			807: out = 16'(-4161);
			808: out = 16'(12876);
			809: out = 16'(7274);
			810: out = 16'(-21087);
			811: out = 16'(-6188);
			812: out = 16'(7343);
			813: out = 16'(18198);
			814: out = 16'(-14689);
			815: out = 16'(-11827);
			816: out = 16'(11883);
			817: out = 16'(-9856);
			818: out = 16'(14);
			819: out = 16'(350);
			820: out = 16'(1514);
			821: out = 16'(-12387);
			822: out = 16'(6565);
			823: out = 16'(10592);
			824: out = 16'(-11363);
			825: out = 16'(-12398);
			826: out = 16'(-9010);
			827: out = 16'(14204);
			828: out = 16'(-6073);
			829: out = 16'(-930);
			830: out = 16'(4576);
			831: out = 16'(-11768);
			832: out = 16'(278);
			833: out = 16'(13324);
			834: out = 16'(-10946);
			835: out = 16'(4601);
			836: out = 16'(-9211);
			837: out = 16'(12825);
			838: out = 16'(-7540);
			839: out = 16'(3594);
			840: out = 16'(14877);
			841: out = 16'(-6946);
			842: out = 16'(-17800);
			843: out = 16'(2632);
			844: out = 16'(9316);
			845: out = 16'(-23480);
			846: out = 16'(16086);
			847: out = 16'(8345);
			848: out = 16'(-2453);
			849: out = 16'(-11408);
			850: out = 16'(-6372);
			851: out = 16'(6307);
			852: out = 16'(-14610);
			853: out = 16'(-12158);
			854: out = 16'(17428);
			855: out = 16'(5415);
			856: out = 16'(-266);
			857: out = 16'(-10534);
			858: out = 16'(9850);
			859: out = 16'(1968);
			860: out = 16'(2503);
			861: out = 16'(8851);
			862: out = 16'(-30402);
			863: out = 16'(3471);
			864: out = 16'(-30113);
			865: out = 16'(11943);
			866: out = 16'(-7762);
			867: out = 16'(20133);
			868: out = 16'(14270);
			869: out = 16'(-9025);
			870: out = 16'(13611);
			871: out = 16'(-12015);
			872: out = 16'(13600);
			873: out = 16'(-6615);
			874: out = 16'(15809);
			875: out = 16'(-5295);
			876: out = 16'(-3080);
			877: out = 16'(1168);
			878: out = 16'(6081);
			879: out = 16'(-1770);
			880: out = 16'(-8810);
			881: out = 16'(-5294);
			882: out = 16'(-6957);
			883: out = 16'(4062);
			884: out = 16'(1926);
			885: out = 16'(7139);
			886: out = 16'(-7839);
			887: out = 16'(-12493);
			888: out = 16'(-2091);
			889: out = 16'(11178);
			890: out = 16'(-13500);
			891: out = 16'(-1793);
			892: out = 16'(-546);
			893: out = 16'(7874);
			894: out = 16'(9381);
			895: out = 16'(-4419);
			896: out = 16'(6531);
			897: out = 16'(-8697);
			898: out = 16'(-3734);
			899: out = 16'(7568);
			900: out = 16'(11477);
			901: out = 16'(-3713);
			902: out = 16'(-12466);
			903: out = 16'(11389);
			904: out = 16'(10415);
			905: out = 16'(-2341);
			906: out = 16'(-548);
			907: out = 16'(9016);
			908: out = 16'(271);
			909: out = 16'(-25927);
			910: out = 16'(5547);
			911: out = 16'(22104);
			912: out = 16'(-1985);
			913: out = 16'(2205);
			914: out = 16'(17699);
			915: out = 16'(-7);
			916: out = 16'(-6544);
			917: out = 16'(5002);
			918: out = 16'(3720);
			919: out = 16'(12381);
			920: out = 16'(-7358);
			921: out = 16'(3073);
			922: out = 16'(953);
			923: out = 16'(114);
			924: out = 16'(1120);
			925: out = 16'(982);
			926: out = 16'(6330);
			927: out = 16'(-5451);
			928: out = 16'(4205);
			929: out = 16'(3494);
			930: out = 16'(-7885);
			931: out = 16'(7799);
			932: out = 16'(-12044);
			933: out = 16'(5066);
			934: out = 16'(-364);
			935: out = 16'(908);
			936: out = 16'(-10784);
			937: out = 16'(-3511);
			938: out = 16'(20504);
			939: out = 16'(7778);
			940: out = 16'(-2457);
			941: out = 16'(12645);
			942: out = 16'(-364);
			943: out = 16'(-30979);
			944: out = 16'(177);
			945: out = 16'(19182);
			946: out = 16'(14795);
			947: out = 16'(-5918);
			948: out = 16'(-6613);
			949: out = 16'(-2075);
			950: out = 16'(5511);
			951: out = 16'(-16378);
			952: out = 16'(1598);
			953: out = 16'(288);
			954: out = 16'(-17302);
			955: out = 16'(2276);
			956: out = 16'(13202);
			957: out = 16'(-4267);
			958: out = 16'(-567);
			959: out = 16'(4840);
			960: out = 16'(-8932);
			961: out = 16'(-860);
			962: out = 16'(-7838);
			963: out = 16'(-583);
			964: out = 16'(1132);
			965: out = 16'(6148);
			966: out = 16'(-5794);
			967: out = 16'(3920);
			968: out = 16'(8791);
			969: out = 16'(-8629);
			970: out = 16'(-24579);
			971: out = 16'(-12391);
			972: out = 16'(14098);
			973: out = 16'(-3064);
			974: out = 16'(3165);
			975: out = 16'(-4926);
			976: out = 16'(2215);
			977: out = 16'(-18710);
			978: out = 16'(-5812);
			979: out = 16'(3165);
			980: out = 16'(-1823);
			981: out = 16'(-11056);
			982: out = 16'(10496);
			983: out = 16'(-12746);
			984: out = 16'(7975);
			985: out = 16'(696);
			986: out = 16'(997);
			987: out = 16'(-2890);
			988: out = 16'(-15781);
			989: out = 16'(3581);
			990: out = 16'(9885);
			991: out = 16'(13181);
			992: out = 16'(-6105);
			993: out = 16'(7903);
			994: out = 16'(-3079);
			995: out = 16'(4789);
			996: out = 16'(-1965);
			997: out = 16'(6713);
			998: out = 16'(9108);
			999: out = 16'(-3336);
			1000: out = 16'(-10797);
			1001: out = 16'(8777);
			1002: out = 16'(5032);
			1003: out = 16'(-3095);
			1004: out = 16'(369);
			1005: out = 16'(21599);
			1006: out = 16'(9020);
			1007: out = 16'(-21228);
			1008: out = 16'(-3579);
			1009: out = 16'(-2543);
			1010: out = 16'(2297);
			1011: out = 16'(2061);
			1012: out = 16'(14054);
			1013: out = 16'(-328);
			1014: out = 16'(-9038);
			1015: out = 16'(-1096);
			1016: out = 16'(-7202);
			1017: out = 16'(13327);
			1018: out = 16'(-12445);
			1019: out = 16'(3776);
			1020: out = 16'(-3817);
			1021: out = 16'(2321);
			1022: out = 16'(-17872);
			1023: out = 16'(-9400);
			1024: out = 16'(2958);
			1025: out = 16'(186);
			1026: out = 16'(-751);
			1027: out = 16'(-47);
			1028: out = 16'(5146);
			1029: out = 16'(2101);
			1030: out = 16'(-4506);
			1031: out = 16'(566);
			1032: out = 16'(14339);
			1033: out = 16'(-8134);
			1034: out = 16'(4705);
			1035: out = 16'(11667);
			1036: out = 16'(99);
			1037: out = 16'(-3605);
			1038: out = 16'(-502);
			1039: out = 16'(10810);
			1040: out = 16'(3899);
			1041: out = 16'(-6142);
			1042: out = 16'(-1457);
			1043: out = 16'(5144);
			1044: out = 16'(-1675);
			1045: out = 16'(4344);
			1046: out = 16'(2974);
			1047: out = 16'(-86);
			1048: out = 16'(-10727);
			1049: out = 16'(2852);
			1050: out = 16'(-5643);
			1051: out = 16'(9854);
			1052: out = 16'(12652);
			1053: out = 16'(-9778);
			1054: out = 16'(6763);
			1055: out = 16'(-22420);
			1056: out = 16'(7730);
			1057: out = 16'(9199);
			1058: out = 16'(10777);
			1059: out = 16'(-12260);
			1060: out = 16'(-4309);
			1061: out = 16'(2775);
			1062: out = 16'(7396);
			1063: out = 16'(606);
			1064: out = 16'(-2104);
			1065: out = 16'(-5539);
			1066: out = 16'(13896);
			1067: out = 16'(13579);
			1068: out = 16'(-8919);
			1069: out = 16'(381);
			1070: out = 16'(-3593);
			1071: out = 16'(4151);
			1072: out = 16'(-8981);
			1073: out = 16'(3808);
			1074: out = 16'(-17645);
			1075: out = 16'(-1417);
			1076: out = 16'(2958);
			1077: out = 16'(334);
			1078: out = 16'(8529);
			1079: out = 16'(-2024);
			1080: out = 16'(1490);
			1081: out = 16'(900);
			1082: out = 16'(9079);
			1083: out = 16'(-5826);
			1084: out = 16'(8365);
			1085: out = 16'(1168);
			1086: out = 16'(-9447);
			1087: out = 16'(-1865);
			1088: out = 16'(-4625);
			1089: out = 16'(-283);
			1090: out = 16'(-7328);
			1091: out = 16'(17750);
			1092: out = 16'(-6966);
			1093: out = 16'(10650);
			1094: out = 16'(-2511);
			1095: out = 16'(3274);
			1096: out = 16'(-22625);
			1097: out = 16'(12562);
			1098: out = 16'(-20747);
			1099: out = 16'(1668);
			1100: out = 16'(26);
			1101: out = 16'(2471);
			1102: out = 16'(3761);
			1103: out = 16'(-17698);
			1104: out = 16'(8128);
			1105: out = 16'(-3940);
			1106: out = 16'(-12164);
			1107: out = 16'(-5831);
			1108: out = 16'(5070);
			1109: out = 16'(-17297);
			1110: out = 16'(10563);
			1111: out = 16'(-16678);
			1112: out = 16'(7493);
			1113: out = 16'(-800);
			1114: out = 16'(-496);
			1115: out = 16'(-836);
			1116: out = 16'(-3661);
			1117: out = 16'(-7839);
			1118: out = 16'(3153);
			1119: out = 16'(17759);
			1120: out = 16'(-16345);
			1121: out = 16'(-15135);
			1122: out = 16'(284);
			1123: out = 16'(17536);
			1124: out = 16'(-5090);
			1125: out = 16'(9852);
			1126: out = 16'(1681);
			1127: out = 16'(-1052);
			1128: out = 16'(223);
			1129: out = 16'(1467);
			1130: out = 16'(6929);
			1131: out = 16'(-2308);
			1132: out = 16'(11132);
			1133: out = 16'(-13239);
			1134: out = 16'(3379);
			1135: out = 16'(-4494);
			1136: out = 16'(9739);
			1137: out = 16'(-6081);
			1138: out = 16'(8086);
			1139: out = 16'(9523);
			1140: out = 16'(11703);
			1141: out = 16'(4907);
			1142: out = 16'(1365);
			1143: out = 16'(15327);
			1144: out = 16'(-11949);
			1145: out = 16'(-19866);
			1146: out = 16'(8961);
			1147: out = 16'(7314);
			1148: out = 16'(-449);
			1149: out = 16'(235);
			1150: out = 16'(1595);
			1151: out = 16'(-13309);
			1152: out = 16'(-1817);
			1153: out = 16'(14409);
			1154: out = 16'(-8223);
			1155: out = 16'(-4355);
			1156: out = 16'(1251);
			1157: out = 16'(2561);
			1158: out = 16'(4339);
			1159: out = 16'(-5564);
			1160: out = 16'(12067);
			1161: out = 16'(-2460);
			1162: out = 16'(969);
			1163: out = 16'(-560);
			1164: out = 16'(3374);
			1165: out = 16'(5541);
			1166: out = 16'(-3603);
			1167: out = 16'(558);
			1168: out = 16'(-7873);
			1169: out = 16'(7176);
			1170: out = 16'(1526);
			1171: out = 16'(9101);
			1172: out = 16'(12161);
			1173: out = 16'(1319);
			1174: out = 16'(-3214);
			1175: out = 16'(4746);
			1176: out = 16'(-2433);
			1177: out = 16'(-14152);
			1178: out = 16'(701);
			1179: out = 16'(5106);
			1180: out = 16'(3977);
			1181: out = 16'(-5751);
			1182: out = 16'(3550);
			1183: out = 16'(-16693);
			1184: out = 16'(-1894);
			1185: out = 16'(1764);
			1186: out = 16'(4424);
			1187: out = 16'(2949);
			1188: out = 16'(4269);
			1189: out = 16'(560);
			1190: out = 16'(-3732);
			1191: out = 16'(1078);
			1192: out = 16'(-50);
			1193: out = 16'(6690);
			1194: out = 16'(-16070);
			1195: out = 16'(7578);
			1196: out = 16'(7820);
			1197: out = 16'(-9166);
			1198: out = 16'(-16736);
			1199: out = 16'(18200);
			1200: out = 16'(12134);
			1201: out = 16'(-14842);
			1202: out = 16'(11683);
			1203: out = 16'(5815);
			1204: out = 16'(-9856);
			1205: out = 16'(-4522);
			1206: out = 16'(11584);
			1207: out = 16'(-3656);
			1208: out = 16'(-14142);
			1209: out = 16'(11616);
			1210: out = 16'(4000);
			1211: out = 16'(-5977);
			1212: out = 16'(-902);
			1213: out = 16'(4682);
			1214: out = 16'(7674);
			1215: out = 16'(-12119);
			1216: out = 16'(1938);
			1217: out = 16'(395);
			1218: out = 16'(3147);
			1219: out = 16'(2402);
			1220: out = 16'(3994);
			1221: out = 16'(3037);
			1222: out = 16'(-21580);
			1223: out = 16'(5868);
			1224: out = 16'(-12819);
			1225: out = 16'(-3213);
			1226: out = 16'(1128);
			1227: out = 16'(15682);
			1228: out = 16'(-7141);
			1229: out = 16'(-13623);
			1230: out = 16'(6255);
			1231: out = 16'(747);
			1232: out = 16'(402);
			1233: out = 16'(7204);
			1234: out = 16'(-6631);
			1235: out = 16'(-4755);
			1236: out = 16'(1910);
			1237: out = 16'(10100);
			1238: out = 16'(7094);
			1239: out = 16'(-22080);
			1240: out = 16'(12581);
			1241: out = 16'(-24792);
			1242: out = 16'(-8170);
			1243: out = 16'(-6480);
			1244: out = 16'(-9156);
			1245: out = 16'(-1857);
			1246: out = 16'(219);
			1247: out = 16'(7693);
			1248: out = 16'(-5519);
			1249: out = 16'(-462);
			1250: out = 16'(-9651);
			1251: out = 16'(-243);
			1252: out = 16'(-9639);
			1253: out = 16'(1886);
			1254: out = 16'(-1817);
			1255: out = 16'(-107);
			1256: out = 16'(-10759);
			1257: out = 16'(-8541);
			1258: out = 16'(9480);
			1259: out = 16'(7917);
			1260: out = 16'(-731);
			1261: out = 16'(4901);
			1262: out = 16'(852);
			1263: out = 16'(1412);
			1264: out = 16'(8966);
			1265: out = 16'(-828);
			1266: out = 16'(163);
			1267: out = 16'(-1076);
			1268: out = 16'(1093);
			1269: out = 16'(-20643);
			1270: out = 16'(12496);
			1271: out = 16'(-12986);
			1272: out = 16'(-5055);
			1273: out = 16'(18545);
			1274: out = 16'(6061);
			1275: out = 16'(-11553);
			1276: out = 16'(-3786);
			1277: out = 16'(10160);
			1278: out = 16'(-8933);
			1279: out = 16'(11732);
			1280: out = 16'(-6360);
			1281: out = 16'(-1532);
			1282: out = 16'(-5238);
			1283: out = 16'(5876);
			1284: out = 16'(4450);
			1285: out = 16'(5110);
			1286: out = 16'(5547);
			1287: out = 16'(1298);
			1288: out = 16'(434);
			1289: out = 16'(863);
			1290: out = 16'(5330);
			1291: out = 16'(9278);
			1292: out = 16'(1955);
			1293: out = 16'(14146);
			1294: out = 16'(5176);
			1295: out = 16'(-21859);
			1296: out = 16'(-636);
			1297: out = 16'(2032);
			1298: out = 16'(14050);
			1299: out = 16'(-4816);
			1300: out = 16'(5946);
			1301: out = 16'(-2897);
			1302: out = 16'(-11872);
			1303: out = 16'(17753);
			1304: out = 16'(-5648);
			1305: out = 16'(7293);
			1306: out = 16'(-2716);
			1307: out = 16'(7331);
			1308: out = 16'(-12236);
			1309: out = 16'(-10860);
			1310: out = 16'(18126);
			1311: out = 16'(-5452);
			1312: out = 16'(-604);
			1313: out = 16'(-6162);
			1314: out = 16'(12482);
			1315: out = 16'(-18245);
			1316: out = 16'(-157);
			1317: out = 16'(2994);
			1318: out = 16'(-7637);
			1319: out = 16'(-8168);
			1320: out = 16'(14713);
			1321: out = 16'(-3969);
			1322: out = 16'(-1740);
			1323: out = 16'(4398);
			1324: out = 16'(12946);
			1325: out = 16'(1839);
			1326: out = 16'(-1997);
			1327: out = 16'(-4450);
			1328: out = 16'(-14012);
			1329: out = 16'(1945);
			1330: out = 16'(3207);
			1331: out = 16'(13544);
			1332: out = 16'(-14185);
			1333: out = 16'(12279);
			1334: out = 16'(4014);
			1335: out = 16'(-4190);
			1336: out = 16'(-698);
			1337: out = 16'(3849);
			1338: out = 16'(10759);
			1339: out = 16'(-12498);
			1340: out = 16'(3031);
			1341: out = 16'(-5087);
			1342: out = 16'(-512);
			1343: out = 16'(-1193);
			1344: out = 16'(12984);
			1345: out = 16'(1568);
			1346: out = 16'(-7631);
			1347: out = 16'(-5358);
			1348: out = 16'(1995);
			1349: out = 16'(749);
			1350: out = 16'(18660);
			1351: out = 16'(2939);
			1352: out = 16'(-15737);
			1353: out = 16'(-9181);
			1354: out = 16'(-9931);
			1355: out = 16'(716);
			1356: out = 16'(-9032);
			1357: out = 16'(-617);
			1358: out = 16'(-220);
			1359: out = 16'(11788);
			1360: out = 16'(-9231);
			1361: out = 16'(6892);
			1362: out = 16'(-18799);
			1363: out = 16'(4937);
			1364: out = 16'(-3735);
			1365: out = 16'(-1567);
			1366: out = 16'(2395);
			1367: out = 16'(-4268);
			1368: out = 16'(-1109);
			1369: out = 16'(374);
			1370: out = 16'(4759);
			1371: out = 16'(-7602);
			1372: out = 16'(-16558);
			1373: out = 16'(-3453);
			1374: out = 16'(332);
			1375: out = 16'(6369);
			1376: out = 16'(9395);
			1377: out = 16'(-12116);
			1378: out = 16'(185);
			1379: out = 16'(7114);
			1380: out = 16'(2246);
			1381: out = 16'(1269);
			1382: out = 16'(-11200);
			1383: out = 16'(11951);
			1384: out = 16'(-4319);
			1385: out = 16'(6233);
			1386: out = 16'(-3504);
			1387: out = 16'(8381);
			1388: out = 16'(-12160);
			1389: out = 16'(6800);
			1390: out = 16'(13015);
			1391: out = 16'(-9486);
			1392: out = 16'(-167);
			1393: out = 16'(1200);
			1394: out = 16'(11503);
			1395: out = 16'(-202);
			1396: out = 16'(-752);
			1397: out = 16'(1180);
			1398: out = 16'(-2286);
			1399: out = 16'(-14462);
			1400: out = 16'(10340);
			1401: out = 16'(-10837);
			1402: out = 16'(-17474);
			1403: out = 16'(940);
			1404: out = 16'(13506);
			1405: out = 16'(-11601);
			1406: out = 16'(-5658);
			1407: out = 16'(-6821);
			1408: out = 16'(5877);
			1409: out = 16'(-4033);
			1410: out = 16'(-408);
			1411: out = 16'(8993);
			1412: out = 16'(-17039);
			1413: out = 16'(4090);
			1414: out = 16'(3853);
			1415: out = 16'(4141);
			1416: out = 16'(-6601);
			1417: out = 16'(2709);
			1418: out = 16'(5120);
			1419: out = 16'(87);
			1420: out = 16'(960);
			1421: out = 16'(7514);
			1422: out = 16'(3416);
			1423: out = 16'(-1742);
			1424: out = 16'(-1350);
			1425: out = 16'(2825);
			1426: out = 16'(-9441);
			1427: out = 16'(-21836);
			1428: out = 16'(7936);
			1429: out = 16'(-25647);
			1430: out = 16'(12463);
			1431: out = 16'(-10798);
			1432: out = 16'(10140);
			1433: out = 16'(-1803);
			1434: out = 16'(-482);
			1435: out = 16'(9019);
			1436: out = 16'(-2819);
			1437: out = 16'(-5386);
			1438: out = 16'(-3628);
			1439: out = 16'(6062);
			1440: out = 16'(1427);
			1441: out = 16'(3984);
			1442: out = 16'(-5830);
			1443: out = 16'(3900);
			1444: out = 16'(-17686);
			1445: out = 16'(2357);
			1446: out = 16'(5252);
			1447: out = 16'(2292);
			1448: out = 16'(-7415);
			1449: out = 16'(8287);
			1450: out = 16'(8974);
			1451: out = 16'(7018);
			1452: out = 16'(-11737);
			1453: out = 16'(11849);
			1454: out = 16'(1277);
			1455: out = 16'(-763);
			1456: out = 16'(14401);
			1457: out = 16'(2289);
			1458: out = 16'(-735);
			1459: out = 16'(-12617);
			1460: out = 16'(10582);
			1461: out = 16'(-1055);
			1462: out = 16'(-4578);
			1463: out = 16'(5634);
			1464: out = 16'(13904);
			1465: out = 16'(-3302);
			1466: out = 16'(-12181);
			1467: out = 16'(5742);
			1468: out = 16'(4589);
			1469: out = 16'(13267);
			1470: out = 16'(-5101);
			1471: out = 16'(-11529);
			1472: out = 16'(-5832);
			1473: out = 16'(11146);
			1474: out = 16'(3047);
			1475: out = 16'(8940);
			1476: out = 16'(183);
			1477: out = 16'(-1754);
			1478: out = 16'(-10634);
			1479: out = 16'(-13996);
			1480: out = 16'(3640);
			1481: out = 16'(-3580);
			1482: out = 16'(-1835);
			1483: out = 16'(2640);
			1484: out = 16'(5988);
			1485: out = 16'(-2983);
			1486: out = 16'(7167);
			1487: out = 16'(-6990);
			1488: out = 16'(480);
			1489: out = 16'(-8599);
			1490: out = 16'(8564);
			1491: out = 16'(3261);
			1492: out = 16'(-4036);
			1493: out = 16'(12757);
			1494: out = 16'(-15247);
			1495: out = 16'(15146);
			1496: out = 16'(-6803);
			1497: out = 16'(-683);
			1498: out = 16'(-5085);
			1499: out = 16'(2194);
			1500: out = 16'(-1726);
			1501: out = 16'(-9879);
			1502: out = 16'(12677);
			1503: out = 16'(2621);
			1504: out = 16'(-1599);
			1505: out = 16'(1873);
			1506: out = 16'(2592);
			1507: out = 16'(8095);
			1508: out = 16'(686);
			1509: out = 16'(4772);
			1510: out = 16'(12624);
			1511: out = 16'(-6333);
			1512: out = 16'(3890);
			1513: out = 16'(1400);
			1514: out = 16'(6489);
			1515: out = 16'(-24481);
			1516: out = 16'(-896);
			1517: out = 16'(-2431);
			1518: out = 16'(-14365);
			1519: out = 16'(5561);
			1520: out = 16'(16093);
			1521: out = 16'(5780);
			1522: out = 16'(-23520);
			1523: out = 16'(9332);
			1524: out = 16'(-13737);
			1525: out = 16'(15777);
			1526: out = 16'(-1840);
			1527: out = 16'(7153);
			1528: out = 16'(10149);
			1529: out = 16'(4633);
			1530: out = 16'(-924);
			1531: out = 16'(970);
			1532: out = 16'(-4168);
			1533: out = 16'(5473);
			1534: out = 16'(-3656);
			1535: out = 16'(3749);
			1536: out = 16'(6962);
			1537: out = 16'(-23111);
			1538: out = 16'(-7005);
			1539: out = 16'(8915);
			1540: out = 16'(10317);
			1541: out = 16'(-12865);
			1542: out = 16'(3666);
			1543: out = 16'(-493);
			1544: out = 16'(68);
			1545: out = 16'(-6835);
			1546: out = 16'(-1640);
			1547: out = 16'(6699);
			1548: out = 16'(-5694);
			1549: out = 16'(-3706);
			1550: out = 16'(1567);
			1551: out = 16'(4085);
			1552: out = 16'(-13134);
			1553: out = 16'(2318);
			1554: out = 16'(360);
			1555: out = 16'(-13293);
			1556: out = 16'(-6);
			1557: out = 16'(12482);
			1558: out = 16'(973);
			1559: out = 16'(-126);
			1560: out = 16'(12548);
			1561: out = 16'(-2725);
			1562: out = 16'(5186);
			1563: out = 16'(4237);
			1564: out = 16'(-8148);
			1565: out = 16'(8453);
			1566: out = 16'(6025);
			1567: out = 16'(-540);
			1568: out = 16'(5963);
			1569: out = 16'(1742);
			1570: out = 16'(9431);
			1571: out = 16'(-6834);
			1572: out = 16'(15021);
			1573: out = 16'(2072);
			1574: out = 16'(-9891);
			1575: out = 16'(1583);
			1576: out = 16'(-6902);
			1577: out = 16'(-3355);
			1578: out = 16'(-4570);
			1579: out = 16'(15894);
			1580: out = 16'(-504);
			1581: out = 16'(-1384);
			1582: out = 16'(-13456);
			1583: out = 16'(-1995);
			1584: out = 16'(2825);
			1585: out = 16'(-1400);
			1586: out = 16'(1565);
			1587: out = 16'(-21238);
			1588: out = 16'(1730);
			1589: out = 16'(6778);
			1590: out = 16'(1641);
			1591: out = 16'(-3702);
			1592: out = 16'(5953);
			1593: out = 16'(157);
			1594: out = 16'(-10012);
			1595: out = 16'(-8745);
			1596: out = 16'(10228);
			1597: out = 16'(-8157);
			1598: out = 16'(-1391);
			1599: out = 16'(-3779);
			1600: out = 16'(2082);
			1601: out = 16'(-21193);
			1602: out = 16'(-18390);
			1603: out = 16'(15064);
			1604: out = 16'(-10344);
			1605: out = 16'(971);
			1606: out = 16'(-828);
			1607: out = 16'(4901);
			1608: out = 16'(-7696);
			1609: out = 16'(1591);
			1610: out = 16'(1870);
			1611: out = 16'(-13959);
			1612: out = 16'(510);
			1613: out = 16'(4560);
			1614: out = 16'(-2804);
			1615: out = 16'(4124);
			1616: out = 16'(5555);
			1617: out = 16'(8647);
			1618: out = 16'(3486);
			1619: out = 16'(2973);
			1620: out = 16'(-3708);
			1621: out = 16'(-17647);
			1622: out = 16'(3099);
			1623: out = 16'(-9536);
			1624: out = 16'(8634);
			1625: out = 16'(-5274);
			1626: out = 16'(2046);
			1627: out = 16'(-5506);
			1628: out = 16'(2084);
			1629: out = 16'(-4437);
			1630: out = 16'(814);
			1631: out = 16'(-362);
			1632: out = 16'(-9637);
			1633: out = 16'(13202);
			1634: out = 16'(-131);
			1635: out = 16'(2756);
			1636: out = 16'(2180);
			1637: out = 16'(4740);
			1638: out = 16'(-539);
			1639: out = 16'(1082);
			1640: out = 16'(2726);
			1641: out = 16'(-6127);
			1642: out = 16'(1061);
			1643: out = 16'(5078);
			1644: out = 16'(11542);
			1645: out = 16'(-523);
			1646: out = 16'(-15564);
			1647: out = 16'(-2765);
			1648: out = 16'(1280);
			1649: out = 16'(-4992);
			1650: out = 16'(6473);
			1651: out = 16'(-18838);
			1652: out = 16'(11183);
			1653: out = 16'(-17382);
			1654: out = 16'(-3593);
			1655: out = 16'(3861);
			1656: out = 16'(8204);
			1657: out = 16'(-8197);
			1658: out = 16'(-644);
			1659: out = 16'(7601);
			1660: out = 16'(-7729);
			1661: out = 16'(-4440);
			1662: out = 16'(-1470);
			1663: out = 16'(12170);
			1664: out = 16'(-2854);
			1665: out = 16'(810);
			1666: out = 16'(578);
			1667: out = 16'(4815);
			1668: out = 16'(2078);
			1669: out = 16'(4167);
			1670: out = 16'(4067);
			1671: out = 16'(7842);
			1672: out = 16'(-7161);
			1673: out = 16'(14403);
			1674: out = 16'(-1491);
			1675: out = 16'(-1062);
			1676: out = 16'(8961);
			1677: out = 16'(-7452);
			1678: out = 16'(-397);
			1679: out = 16'(-8022);
			1680: out = 16'(9004);
			1681: out = 16'(-19860);
			1682: out = 16'(7642);
			1683: out = 16'(7594);
			1684: out = 16'(158);
			1685: out = 16'(-2020);
			1686: out = 16'(-2867);
			1687: out = 16'(6358);
			1688: out = 16'(-10944);
			1689: out = 16'(11528);
			1690: out = 16'(9789);
			1691: out = 16'(-3375);
			1692: out = 16'(-10921);
			1693: out = 16'(4998);
			1694: out = 16'(-15622);
			1695: out = 16'(-606);
			1696: out = 16'(-8041);
			1697: out = 16'(3022);
			1698: out = 16'(-20284);
			1699: out = 16'(-1193);
			1700: out = 16'(5331);
			1701: out = 16'(2273);
			1702: out = 16'(-5525);
			1703: out = 16'(-10081);
			1704: out = 16'(10308);
			1705: out = 16'(-12956);
			1706: out = 16'(4332);
			1707: out = 16'(-7999);
			1708: out = 16'(11768);
			1709: out = 16'(-3896);
			1710: out = 16'(2365);
			1711: out = 16'(-3076);
			1712: out = 16'(-8154);
			1713: out = 16'(-4033);
			1714: out = 16'(1155);
			1715: out = 16'(9675);
			1716: out = 16'(-941);
			1717: out = 16'(-3751);
			1718: out = 16'(-11884);
			1719: out = 16'(12651);
			1720: out = 16'(1971);
			1721: out = 16'(-877);
			1722: out = 16'(12922);
			1723: out = 16'(11003);
			1724: out = 16'(-4559);
			1725: out = 16'(3447);
			1726: out = 16'(4695);
			1727: out = 16'(6333);
			1728: out = 16'(4003);
			1729: out = 16'(2626);
			1730: out = 16'(5594);
			1731: out = 16'(-12575);
			1732: out = 16'(9733);
			1733: out = 16'(-4789);
			1734: out = 16'(7261);
			1735: out = 16'(3792);
			1736: out = 16'(-2429);
			1737: out = 16'(-9866);
			1738: out = 16'(-211);
			1739: out = 16'(-1294);
			1740: out = 16'(196);
			1741: out = 16'(1891);
			1742: out = 16'(2329);
			1743: out = 16'(8582);
			1744: out = 16'(-8242);
			1745: out = 16'(13588);
			1746: out = 16'(-8631);
			1747: out = 16'(7706);
			1748: out = 16'(-3081);
			1749: out = 16'(5975);
			1750: out = 16'(-5404);
			1751: out = 16'(-1324);
			1752: out = 16'(-4239);
			1753: out = 16'(2982);
			1754: out = 16'(1748);
			1755: out = 16'(1691);
			1756: out = 16'(2694);
			1757: out = 16'(-7635);
			1758: out = 16'(3928);
			1759: out = 16'(-8);
			1760: out = 16'(10953);
			1761: out = 16'(-9195);
			1762: out = 16'(-6550);
			1763: out = 16'(-9363);
			1764: out = 16'(4203);
			1765: out = 16'(6185);
			1766: out = 16'(-7703);
			1767: out = 16'(74);
			1768: out = 16'(-834);
			1769: out = 16'(-4536);
			1770: out = 16'(-9603);
			1771: out = 16'(3061);
			1772: out = 16'(4626);
			1773: out = 16'(-1448);
			1774: out = 16'(11040);
			1775: out = 16'(8129);
			1776: out = 16'(-2743);
			1777: out = 16'(-8779);
			1778: out = 16'(2358);
			1779: out = 16'(12740);
			1780: out = 16'(-5757);
			1781: out = 16'(1759);
			1782: out = 16'(-2522);
			1783: out = 16'(4054);
			1784: out = 16'(1064);
			1785: out = 16'(-185);
			1786: out = 16'(1952);
			1787: out = 16'(418);
			1788: out = 16'(1939);
			1789: out = 16'(-7750);
			1790: out = 16'(2386);
			1791: out = 16'(1954);
			1792: out = 16'(-348);
			1793: out = 16'(12490);
			1794: out = 16'(325);
			1795: out = 16'(-2718);
			1796: out = 16'(-5926);
			1797: out = 16'(2659);
			1798: out = 16'(1200);
			1799: out = 16'(-5928);
			1800: out = 16'(6360);
			1801: out = 16'(-6246);
			1802: out = 16'(-3480);
			1803: out = 16'(8928);
			1804: out = 16'(1032);
			1805: out = 16'(-1412);
			1806: out = 16'(236);
			1807: out = 16'(2771);
			1808: out = 16'(-9863);
			1809: out = 16'(4096);
			1810: out = 16'(-1578);
			1811: out = 16'(-6955);
			1812: out = 16'(1714);
			1813: out = 16'(-2398);
			1814: out = 16'(12038);
			1815: out = 16'(-5890);
			1816: out = 16'(3542);
			1817: out = 16'(4459);
			1818: out = 16'(-3499);
			1819: out = 16'(11245);
			1820: out = 16'(4378);
			1821: out = 16'(1043);
			1822: out = 16'(-8674);
			1823: out = 16'(927);
			1824: out = 16'(981);
			1825: out = 16'(8239);
			1826: out = 16'(1630);
			1827: out = 16'(-2007);
			1828: out = 16'(9529);
			1829: out = 16'(4393);
			1830: out = 16'(4266);
			1831: out = 16'(8614);
			1832: out = 16'(-5960);
			1833: out = 16'(3113);
			1834: out = 16'(-997);
			1835: out = 16'(8124);
			1836: out = 16'(-7324);
			1837: out = 16'(4273);
			1838: out = 16'(-1358);
			1839: out = 16'(-2115);
			1840: out = 16'(3205);
			1841: out = 16'(-16902);
			1842: out = 16'(3135);
			1843: out = 16'(1054);
			1844: out = 16'(6628);
			1845: out = 16'(-15896);
			1846: out = 16'(4126);
			1847: out = 16'(-15962);
			1848: out = 16'(6033);
			1849: out = 16'(4787);
			1850: out = 16'(130);
			1851: out = 16'(-338);
			1852: out = 16'(199);
			1853: out = 16'(-2289);
			1854: out = 16'(650);
			1855: out = 16'(1523);
			1856: out = 16'(-16489);
			1857: out = 16'(4935);
			1858: out = 16'(11402);
			1859: out = 16'(8981);
			1860: out = 16'(-14696);
			1861: out = 16'(9174);
			1862: out = 16'(-3540);
			1863: out = 16'(-12781);
			1864: out = 16'(1332);
			1865: out = 16'(9523);
			1866: out = 16'(-8816);
			1867: out = 16'(2212);
			1868: out = 16'(2435);
			1869: out = 16'(-6771);
			1870: out = 16'(2194);
			1871: out = 16'(-10295);
			1872: out = 16'(13924);
			1873: out = 16'(-17445);
			1874: out = 16'(2105);
			1875: out = 16'(11794);
			1876: out = 16'(5089);
			1877: out = 16'(-6783);
			1878: out = 16'(-217);
			1879: out = 16'(-1851);
			1880: out = 16'(296);
			1881: out = 16'(1490);
			1882: out = 16'(-2226);
			1883: out = 16'(709);
			1884: out = 16'(-1875);
			1885: out = 16'(6251);
			1886: out = 16'(-410);
			1887: out = 16'(4359);
			1888: out = 16'(-16084);
			1889: out = 16'(5352);
			1890: out = 16'(9412);
			1891: out = 16'(5198);
			1892: out = 16'(-1025);
			1893: out = 16'(1996);
			1894: out = 16'(-42);
			1895: out = 16'(-1045);
			1896: out = 16'(-151);
			1897: out = 16'(-904);
			1898: out = 16'(8226);
			1899: out = 16'(-8390);
			1900: out = 16'(-905);
			1901: out = 16'(-3648);
			1902: out = 16'(334);
			1903: out = 16'(-16373);
			1904: out = 16'(10305);
			1905: out = 16'(778);
			1906: out = 16'(-10299);
			1907: out = 16'(1527);
			1908: out = 16'(-1994);
			1909: out = 16'(1695);
			1910: out = 16'(4485);
			1911: out = 16'(3469);
			1912: out = 16'(-411);
			1913: out = 16'(8441);
			1914: out = 16'(-47);
			1915: out = 16'(-7);
			1916: out = 16'(-8702);
			1917: out = 16'(6966);
			1918: out = 16'(-1592);
			1919: out = 16'(-8222);
			1920: out = 16'(7640);
			1921: out = 16'(-2973);
			1922: out = 16'(9);
			1923: out = 16'(-1885);
			1924: out = 16'(7687);
			1925: out = 16'(342);
			1926: out = 16'(-1695);
			1927: out = 16'(-3157);
			1928: out = 16'(9683);
			1929: out = 16'(-13779);
			1930: out = 16'(13654);
			1931: out = 16'(-1849);
			1932: out = 16'(-2672);
			1933: out = 16'(-3234);
			1934: out = 16'(5982);
			1935: out = 16'(310);
			1936: out = 16'(332);
			1937: out = 16'(9054);
			1938: out = 16'(-5484);
			1939: out = 16'(685);
			1940: out = 16'(-12312);
			1941: out = 16'(9210);
			1942: out = 16'(2888);
			1943: out = 16'(-682);
			1944: out = 16'(7766);
			1945: out = 16'(540);
			1946: out = 16'(-6570);
			1947: out = 16'(3556);
			1948: out = 16'(-463);
			1949: out = 16'(1306);
			1950: out = 16'(-4003);
			1951: out = 16'(-895);
			1952: out = 16'(-5335);
			1953: out = 16'(-2372);
			1954: out = 16'(998);
			1955: out = 16'(-1164);
			1956: out = 16'(-235);
			1957: out = 16'(-69);
			1958: out = 16'(-3347);
			1959: out = 16'(-11316);
			1960: out = 16'(10431);
			1961: out = 16'(-15294);
			1962: out = 16'(4238);
			1963: out = 16'(2214);
			1964: out = 16'(-12385);
			1965: out = 16'(-33);
			1966: out = 16'(-8456);
			1967: out = 16'(460);
			1968: out = 16'(-5531);
			1969: out = 16'(13317);
			1970: out = 16'(-8171);
			1971: out = 16'(711);
			1972: out = 16'(-13034);
			1973: out = 16'(8323);
			1974: out = 16'(554);
			1975: out = 16'(2184);
			1976: out = 16'(2600);
			1977: out = 16'(1055);
			1978: out = 16'(419);
			1979: out = 16'(-2947);
			1980: out = 16'(487);
			1981: out = 16'(6764);
			1982: out = 16'(435);
			1983: out = 16'(-3742);
			1984: out = 16'(6671);
			1985: out = 16'(-9374);
			1986: out = 16'(1283);
			1987: out = 16'(-689);
			1988: out = 16'(4665);
			1989: out = 16'(-2678);
			1990: out = 16'(4451);
			1991: out = 16'(2471);
			1992: out = 16'(-2238);
			1993: out = 16'(-427);
			1994: out = 16'(-230);
			1995: out = 16'(6963);
			1996: out = 16'(-8648);
			1997: out = 16'(1629);
			1998: out = 16'(2480);
			1999: out = 16'(1589);
			2000: out = 16'(4407);
			2001: out = 16'(2234);
			2002: out = 16'(5127);
			2003: out = 16'(-4820);
			2004: out = 16'(-16903);
			2005: out = 16'(6434);
			2006: out = 16'(5322);
			2007: out = 16'(-1039);
			2008: out = 16'(8091);
			2009: out = 16'(7682);
			2010: out = 16'(-4524);
			2011: out = 16'(1641);
			2012: out = 16'(10784);
			2013: out = 16'(855);
			2014: out = 16'(7185);
			2015: out = 16'(-2439);
			2016: out = 16'(1956);
			2017: out = 16'(-3655);
			2018: out = 16'(2771);
			2019: out = 16'(6839);
			2020: out = 16'(-2700);
			2021: out = 16'(13556);
			2022: out = 16'(-4055);
			2023: out = 16'(-1741);
			2024: out = 16'(-355);
			2025: out = 16'(81);
			2026: out = 16'(-1953);
			2027: out = 16'(3009);
			2028: out = 16'(2744);
			2029: out = 16'(59);
			2030: out = 16'(1729);
			2031: out = 16'(2230);
			2032: out = 16'(-6747);
			2033: out = 16'(-2693);
			2034: out = 16'(4457);
			2035: out = 16'(-12419);
			2036: out = 16'(-538);
			2037: out = 16'(-925);
			2038: out = 16'(-642);
			2039: out = 16'(-5546);
			2040: out = 16'(8658);
			2041: out = 16'(3423);
			2042: out = 16'(-7289);
			2043: out = 16'(3436);
			2044: out = 16'(-7143);
			2045: out = 16'(3244);
			2046: out = 16'(-10322);
			2047: out = 16'(4439);
			2048: out = 16'(8964);
			2049: out = 16'(-2077);
			2050: out = 16'(-4595);
			2051: out = 16'(464);
			2052: out = 16'(1258);
			2053: out = 16'(1048);
			2054: out = 16'(5977);
			2055: out = 16'(1642);
			2056: out = 16'(-8444);
			2057: out = 16'(3717);
			2058: out = 16'(5156);
			2059: out = 16'(-1296);
			2060: out = 16'(-7062);
			2061: out = 16'(-2513);
			2062: out = 16'(4290);
			2063: out = 16'(-8795);
			2064: out = 16'(5680);
			2065: out = 16'(-2204);
			2066: out = 16'(2548);
			2067: out = 16'(-4095);
			2068: out = 16'(-510);
			2069: out = 16'(-8587);
			2070: out = 16'(340);
			2071: out = 16'(-236);
			2072: out = 16'(-2498);
			2073: out = 16'(5838);
			2074: out = 16'(5853);
			2075: out = 16'(-3112);
			2076: out = 16'(-462);
			2077: out = 16'(2005);
			2078: out = 16'(-5846);
			2079: out = 16'(1259);
			2080: out = 16'(3652);
			2081: out = 16'(-2881);
			2082: out = 16'(-5923);
			2083: out = 16'(-4890);
			2084: out = 16'(-6746);
			2085: out = 16'(11044);
			2086: out = 16'(-4741);
			2087: out = 16'(5067);
			2088: out = 16'(-1675);
			2089: out = 16'(-1728);
			2090: out = 16'(13181);
			2091: out = 16'(-11216);
			2092: out = 16'(11559);
			2093: out = 16'(-375);
			2094: out = 16'(2816);
			2095: out = 16'(-5558);
			2096: out = 16'(2165);
			2097: out = 16'(9911);
			2098: out = 16'(-2536);
			2099: out = 16'(7196);
			2100: out = 16'(8513);
			2101: out = 16'(5523);
			2102: out = 16'(-17784);
			2103: out = 16'(-2520);
			2104: out = 16'(4037);
			2105: out = 16'(-405);
			2106: out = 16'(-2585);
			2107: out = 16'(10836);
			2108: out = 16'(3775);
			2109: out = 16'(-66);
			2110: out = 16'(919);
			2111: out = 16'(6340);
			2112: out = 16'(-5123);
			2113: out = 16'(-671);
			2114: out = 16'(1012);
			2115: out = 16'(4767);
			2116: out = 16'(-3152);
			2117: out = 16'(545);
			2118: out = 16'(4784);
			2119: out = 16'(-6955);
			2120: out = 16'(11703);
			2121: out = 16'(-15646);
			2122: out = 16'(4670);
			2123: out = 16'(4293);
			2124: out = 16'(-1619);
			2125: out = 16'(-1383);
			2126: out = 16'(6645);
			2127: out = 16'(11243);
			2128: out = 16'(-12460);
			2129: out = 16'(5739);
			2130: out = 16'(4162);
			2131: out = 16'(5363);
			2132: out = 16'(-649);
			2133: out = 16'(5500);
			2134: out = 16'(1521);
			2135: out = 16'(10722);
			2136: out = 16'(-13617);
			2137: out = 16'(7908);
			2138: out = 16'(-7162);
			2139: out = 16'(-629);
			2140: out = 16'(167);
			2141: out = 16'(2113);
			2142: out = 16'(-3226);
			2143: out = 16'(-8525);
			2144: out = 16'(10446);
			2145: out = 16'(-3027);
			2146: out = 16'(609);
			2147: out = 16'(-12590);
			2148: out = 16'(11331);
			2149: out = 16'(-16230);
			2150: out = 16'(7061);
			2151: out = 16'(-1807);
			2152: out = 16'(-5469);
			2153: out = 16'(883);
			2154: out = 16'(3281);
			2155: out = 16'(3189);
			2156: out = 16'(-8610);
			2157: out = 16'(-1191);
			2158: out = 16'(-4643);
			2159: out = 16'(506);
			2160: out = 16'(-1656);
			2161: out = 16'(-3888);
			2162: out = 16'(-1053);
			2163: out = 16'(-2595);
			2164: out = 16'(2643);
			2165: out = 16'(2009);
			2166: out = 16'(-13470);
			2167: out = 16'(-7028);
			2168: out = 16'(3758);
			2169: out = 16'(112);
			2170: out = 16'(-4606);
			2171: out = 16'(3541);
			2172: out = 16'(5708);
			2173: out = 16'(4602);
			2174: out = 16'(5610);
			2175: out = 16'(4713);
			2176: out = 16'(-1943);
			2177: out = 16'(-6258);
			2178: out = 16'(-147);
			2179: out = 16'(-48);
			2180: out = 16'(-35);
			2181: out = 16'(-5200);
			2182: out = 16'(-8536);
			2183: out = 16'(7802);
			2184: out = 16'(1851);
			2185: out = 16'(1471);
			2186: out = 16'(-269);
			2187: out = 16'(1378);
			2188: out = 16'(-5194);
			2189: out = 16'(-18467);
			2190: out = 16'(8501);
			2191: out = 16'(14216);
			2192: out = 16'(-2719);
			2193: out = 16'(655);
			2194: out = 16'(9370);
			2195: out = 16'(-2572);
			2196: out = 16'(3094);
			2197: out = 16'(873);
			2198: out = 16'(11385);
			2199: out = 16'(-3125);
			2200: out = 16'(8610);
			2201: out = 16'(2735);
			2202: out = 16'(-3784);
			2203: out = 16'(-1514);
			2204: out = 16'(-3575);
			2205: out = 16'(6361);
			2206: out = 16'(1938);
			2207: out = 16'(8306);
			2208: out = 16'(-8204);
			2209: out = 16'(119);
			2210: out = 16'(4949);
			2211: out = 16'(6295);
			2212: out = 16'(-1205);
			2213: out = 16'(-10964);
			2214: out = 16'(-4022);
			2215: out = 16'(1405);
			2216: out = 16'(-10787);
			2217: out = 16'(8481);
			2218: out = 16'(3845);
			2219: out = 16'(-6150);
			2220: out = 16'(4374);
			2221: out = 16'(14468);
			2222: out = 16'(-8737);
			2223: out = 16'(-14469);
			2224: out = 16'(10328);
			2225: out = 16'(-2842);
			2226: out = 16'(-876);
			2227: out = 16'(23);
			2228: out = 16'(9540);
			2229: out = 16'(-4921);
			2230: out = 16'(-809);
			2231: out = 16'(7820);
			2232: out = 16'(-4267);
			2233: out = 16'(-5096);
			2234: out = 16'(-5740);
			2235: out = 16'(11042);
			2236: out = 16'(-590);
			2237: out = 16'(-3274);
			2238: out = 16'(8718);
			2239: out = 16'(-8777);
			2240: out = 16'(305);
			2241: out = 16'(-3368);
			2242: out = 16'(6012);
			2243: out = 16'(-4089);
			2244: out = 16'(1764);
			2245: out = 16'(10856);
			2246: out = 16'(-3190);
			2247: out = 16'(3396);
			2248: out = 16'(-1883);
			2249: out = 16'(2923);
			2250: out = 16'(6743);
			2251: out = 16'(-5033);
			2252: out = 16'(10426);
			2253: out = 16'(-1539);
			2254: out = 16'(-2485);
			2255: out = 16'(4082);
			2256: out = 16'(-7246);
			2257: out = 16'(1197);
			2258: out = 16'(-943);
			2259: out = 16'(4715);
			2260: out = 16'(-1626);
			2261: out = 16'(-2738);
			2262: out = 16'(3460);
			2263: out = 16'(5893);
			2264: out = 16'(201);
			2265: out = 16'(4658);
			2266: out = 16'(2125);
			2267: out = 16'(479);
			2268: out = 16'(1972);
			2269: out = 16'(779);
			2270: out = 16'(-9678);
			2271: out = 16'(3894);
			2272: out = 16'(-8629);
			2273: out = 16'(4533);
			2274: out = 16'(-3434);
			2275: out = 16'(-308);
			2276: out = 16'(-2057);
			2277: out = 16'(-526);
			2278: out = 16'(6493);
			2279: out = 16'(-17909);
			2280: out = 16'(8909);
			2281: out = 16'(-9450);
			2282: out = 16'(4244);
			2283: out = 16'(-10986);
			2284: out = 16'(5084);
			2285: out = 16'(9277);
			2286: out = 16'(-9822);
			2287: out = 16'(3110);
			2288: out = 16'(-1597);
			2289: out = 16'(-9385);
			2290: out = 16'(-5879);
			2291: out = 16'(5976);
			2292: out = 16'(6353);
			2293: out = 16'(-1538);
			2294: out = 16'(2809);
			2295: out = 16'(-625);
			2296: out = 16'(-6049);
			2297: out = 16'(6413);
			2298: out = 16'(773);
			2299: out = 16'(-2270);
			2300: out = 16'(-2886);
			2301: out = 16'(12151);
			2302: out = 16'(-5315);
			2303: out = 16'(-8259);
			2304: out = 16'(11474);
			2305: out = 16'(8609);
			2306: out = 16'(-5062);
			2307: out = 16'(-12608);
			2308: out = 16'(11587);
			2309: out = 16'(-14827);
			2310: out = 16'(-360);
			2311: out = 16'(4057);
			2312: out = 16'(1559);
			2313: out = 16'(-9978);
			2314: out = 16'(-4193);
			2315: out = 16'(6808);
			2316: out = 16'(-7488);
			2317: out = 16'(-26);
			2318: out = 16'(7185);
			2319: out = 16'(3693);
			2320: out = 16'(-9361);
			2321: out = 16'(4552);
			2322: out = 16'(6537);
			2323: out = 16'(2978);
			2324: out = 16'(-1676);
			2325: out = 16'(9031);
			2326: out = 16'(-4203);
			2327: out = 16'(4529);
			2328: out = 16'(-1076);
			2329: out = 16'(-1017);
			2330: out = 16'(636);
			2331: out = 16'(1063);
			2332: out = 16'(2320);
			2333: out = 16'(-1477);
			2334: out = 16'(4647);
			2335: out = 16'(-2022);
			2336: out = 16'(6026);
			2337: out = 16'(5419);
			2338: out = 16'(5278);
			2339: out = 16'(1942);
			2340: out = 16'(-4516);
			2341: out = 16'(6858);
			2342: out = 16'(-5007);
			2343: out = 16'(3297);
			2344: out = 16'(1307);
			2345: out = 16'(6464);
			2346: out = 16'(-7400);
			2347: out = 16'(-2315);
			2348: out = 16'(-2738);
			2349: out = 16'(2128);
			2350: out = 16'(1764);
			2351: out = 16'(-163);
			2352: out = 16'(1528);
			2353: out = 16'(965);
			2354: out = 16'(2474);
			2355: out = 16'(-5373);
			2356: out = 16'(7532);
			2357: out = 16'(-4219);
			2358: out = 16'(3209);
			2359: out = 16'(-9562);
			2360: out = 16'(147);
			2361: out = 16'(6992);
			2362: out = 16'(2209);
			2363: out = 16'(5582);
			2364: out = 16'(10950);
			2365: out = 16'(-1763);
			2366: out = 16'(-16358);
			2367: out = 16'(-1176);
			2368: out = 16'(-128);
			2369: out = 16'(3489);
			2370: out = 16'(2647);
			2371: out = 16'(13166);
			2372: out = 16'(-5135);
			2373: out = 16'(-556);
			2374: out = 16'(1473);
			2375: out = 16'(-537);
			2376: out = 16'(1450);
			2377: out = 16'(-2828);
			2378: out = 16'(8909);
			2379: out = 16'(-1999);
			2380: out = 16'(2035);
			2381: out = 16'(-206);
			2382: out = 16'(-2592);
			2383: out = 16'(-2572);
			2384: out = 16'(11078);
			2385: out = 16'(-5100);
			2386: out = 16'(-4196);
			2387: out = 16'(-6922);
			2388: out = 16'(4914);
			2389: out = 16'(-5135);
			2390: out = 16'(-263);
			2391: out = 16'(12232);
			2392: out = 16'(-1373);
			2393: out = 16'(-4444);
			2394: out = 16'(584);
			2395: out = 16'(4629);
			2396: out = 16'(-12049);
			2397: out = 16'(1111);
			2398: out = 16'(-2327);
			2399: out = 16'(3884);
			2400: out = 16'(-14009);
			2401: out = 16'(3280);
			2402: out = 16'(4265);
			2403: out = 16'(-12414);
			2404: out = 16'(-13800);
			2405: out = 16'(1939);
			2406: out = 16'(-7773);
			2407: out = 16'(-6393);
			2408: out = 16'(1663);
			2409: out = 16'(3190);
			2410: out = 16'(3330);
			2411: out = 16'(-6827);
			2412: out = 16'(7787);
			2413: out = 16'(-10969);
			2414: out = 16'(-1530);
			2415: out = 16'(883);
			2416: out = 16'(1468);
			2417: out = 16'(49);
			2418: out = 16'(-2651);
			2419: out = 16'(1475);
			2420: out = 16'(-2750);
			2421: out = 16'(-1055);
			2422: out = 16'(1830);
			2423: out = 16'(589);
			2424: out = 16'(-4412);
			2425: out = 16'(-253);
			2426: out = 16'(2243);
			2427: out = 16'(-3527);
			2428: out = 16'(922);
			2429: out = 16'(7153);
			2430: out = 16'(-4250);
			2431: out = 16'(-7936);
			2432: out = 16'(2776);
			2433: out = 16'(-7214);
			2434: out = 16'(-8308);
			2435: out = 16'(11839);
			2436: out = 16'(8130);
			2437: out = 16'(2026);
			2438: out = 16'(8939);
			2439: out = 16'(-5295);
			2440: out = 16'(3918);
			2441: out = 16'(-3146);
			2442: out = 16'(4365);
			2443: out = 16'(-3839);
			2444: out = 16'(1270);
			2445: out = 16'(-10358);
			2446: out = 16'(-2477);
			2447: out = 16'(10905);
			2448: out = 16'(6994);
			2449: out = 16'(-1467);
			2450: out = 16'(2813);
			2451: out = 16'(6807);
			2452: out = 16'(-814);
			2453: out = 16'(-4477);
			2454: out = 16'(3396);
			2455: out = 16'(13234);
			2456: out = 16'(-5326);
			2457: out = 16'(289);
			2458: out = 16'(9901);
			2459: out = 16'(-3707);
			2460: out = 16'(-10692);
			2461: out = 16'(10449);
			2462: out = 16'(-449);
			2463: out = 16'(1066);
			2464: out = 16'(921);
			2465: out = 16'(1620);
			2466: out = 16'(-969);
			2467: out = 16'(-4802);
			2468: out = 16'(9988);
			2469: out = 16'(-3710);
			2470: out = 16'(-13073);
			2471: out = 16'(827);
			2472: out = 16'(4427);
			2473: out = 16'(-6001);
			2474: out = 16'(-2713);
			2475: out = 16'(11496);
			2476: out = 16'(-6531);
			2477: out = 16'(-16353);
			2478: out = 16'(4024);
			2479: out = 16'(606);
			2480: out = 16'(-17331);
			2481: out = 16'(8203);
			2482: out = 16'(2228);
			2483: out = 16'(-3120);
			2484: out = 16'(-5047);
			2485: out = 16'(10723);
			2486: out = 16'(-8538);
			2487: out = 16'(3142);
			2488: out = 16'(7085);
			2489: out = 16'(1356);
			2490: out = 16'(-10577);
			2491: out = 16'(6971);
			2492: out = 16'(-4989);
			2493: out = 16'(-3212);
			2494: out = 16'(3108);
			2495: out = 16'(1956);
			2496: out = 16'(1946);
			2497: out = 16'(-3612);
			2498: out = 16'(2795);
			2499: out = 16'(2922);
			2500: out = 16'(-500);
			2501: out = 16'(-5506);
			2502: out = 16'(1126);
			2503: out = 16'(-3737);
			2504: out = 16'(-1014);
			2505: out = 16'(-128);
			2506: out = 16'(7206);
			2507: out = 16'(-5527);
			2508: out = 16'(3374);
			2509: out = 16'(-1736);
			2510: out = 16'(-9746);
			2511: out = 16'(4334);
			2512: out = 16'(347);
			2513: out = 16'(379);
			2514: out = 16'(601);
			2515: out = 16'(-1397);
			2516: out = 16'(-754);
			2517: out = 16'(-54);
			2518: out = 16'(-764);
			2519: out = 16'(-2874);
			2520: out = 16'(-88);
			2521: out = 16'(-2036);
			2522: out = 16'(-3043);
			2523: out = 16'(2879);
			2524: out = 16'(-520);
			2525: out = 16'(-3877);
			2526: out = 16'(3685);
			2527: out = 16'(-2860);
			2528: out = 16'(7656);
			2529: out = 16'(-11308);
			2530: out = 16'(-4320);
			2531: out = 16'(8358);
			2532: out = 16'(-7146);
			2533: out = 16'(3061);
			2534: out = 16'(5963);
			2535: out = 16'(2158);
			2536: out = 16'(-5943);
			2537: out = 16'(9763);
			2538: out = 16'(-1537);
			2539: out = 16'(-1969);
			2540: out = 16'(-590);
			2541: out = 16'(4906);
			2542: out = 16'(6951);
			2543: out = 16'(-5730);
			2544: out = 16'(-1465);
			2545: out = 16'(1840);
			2546: out = 16'(1557);
			2547: out = 16'(-5488);
			2548: out = 16'(10116);
			2549: out = 16'(-1185);
			2550: out = 16'(-4404);
			2551: out = 16'(10206);
			2552: out = 16'(8242);
			2553: out = 16'(622);
			2554: out = 16'(-5622);
			2555: out = 16'(5190);
			2556: out = 16'(6351);
			2557: out = 16'(-6727);
			2558: out = 16'(2071);
			2559: out = 16'(407);
			2560: out = 16'(-9951);
			2561: out = 16'(4570);
			2562: out = 16'(-20);
			2563: out = 16'(4067);
			2564: out = 16'(-9434);
			2565: out = 16'(7425);
			2566: out = 16'(-305);
			2567: out = 16'(2242);
			2568: out = 16'(469);
			2569: out = 16'(4426);
			2570: out = 16'(-3845);
			2571: out = 16'(-329);
			2572: out = 16'(5778);
			2573: out = 16'(-5057);
			2574: out = 16'(5160);
			2575: out = 16'(-7884);
			2576: out = 16'(-4405);
			2577: out = 16'(-10631);
			2578: out = 16'(9146);
			2579: out = 16'(662);
			2580: out = 16'(170);
			2581: out = 16'(-1563);
			2582: out = 16'(-1564);
			2583: out = 16'(-2249);
			2584: out = 16'(-3957);
			2585: out = 16'(561);
			2586: out = 16'(-4226);
			2587: out = 16'(102);
			2588: out = 16'(7569);
			2589: out = 16'(2656);
			2590: out = 16'(-4965);
			2591: out = 16'(-9937);
			2592: out = 16'(661);
			2593: out = 16'(-958);
			2594: out = 16'(-8369);
			2595: out = 16'(6058);
			2596: out = 16'(-4498);
			2597: out = 16'(-4925);
			2598: out = 16'(12878);
			2599: out = 16'(-392);
			2600: out = 16'(-4592);
			2601: out = 16'(-10075);
			2602: out = 16'(2344);
			2603: out = 16'(-12132);
			2604: out = 16'(-1791);
			2605: out = 16'(2704);
			2606: out = 16'(-1344);
			2607: out = 16'(4735);
			2608: out = 16'(8893);
			2609: out = 16'(3210);
			2610: out = 16'(-11258);
			2611: out = 16'(4097);
			2612: out = 16'(4719);
			2613: out = 16'(1473);
			2614: out = 16'(2739);
			2615: out = 16'(-4133);
			2616: out = 16'(-828);
			2617: out = 16'(-1693);
			2618: out = 16'(3513);
			2619: out = 16'(321);
			2620: out = 16'(-3269);
			2621: out = 16'(156);
			2622: out = 16'(-3948);
			2623: out = 16'(-272);
			2624: out = 16'(-1932);
			2625: out = 16'(8563);
			2626: out = 16'(-3704);
			2627: out = 16'(323);
			2628: out = 16'(5345);
			2629: out = 16'(-7854);
			2630: out = 16'(7597);
			2631: out = 16'(-4083);
			2632: out = 16'(1542);
			2633: out = 16'(-2122);
			2634: out = 16'(1297);
			2635: out = 16'(5155);
			2636: out = 16'(-7538);
			2637: out = 16'(3654);
			2638: out = 16'(5648);
			2639: out = 16'(3278);
			2640: out = 16'(-3803);
			2641: out = 16'(6640);
			2642: out = 16'(-4831);
			2643: out = 16'(-811);
			2644: out = 16'(756);
			2645: out = 16'(1012);
			2646: out = 16'(-5659);
			2647: out = 16'(-567);
			2648: out = 16'(717);
			2649: out = 16'(955);
			2650: out = 16'(-5697);
			2651: out = 16'(5565);
			2652: out = 16'(1189);
			2653: out = 16'(7017);
			2654: out = 16'(-7700);
			2655: out = 16'(-4675);
			2656: out = 16'(741);
			2657: out = 16'(951);
			2658: out = 16'(6200);
			2659: out = 16'(-9917);
			2660: out = 16'(222);
			2661: out = 16'(-5905);
			2662: out = 16'(3583);
			2663: out = 16'(-2016);
			2664: out = 16'(8561);
			2665: out = 16'(4167);
			2666: out = 16'(-279);
			2667: out = 16'(4597);
			2668: out = 16'(-2051);
			2669: out = 16'(-11375);
			2670: out = 16'(2515);
			2671: out = 16'(-2395);
			2672: out = 16'(5944);
			2673: out = 16'(4082);
			2674: out = 16'(2348);
			2675: out = 16'(2357);
			2676: out = 16'(-4052);
			2677: out = 16'(3349);
			2678: out = 16'(-3808);
			2679: out = 16'(-5177);
			2680: out = 16'(-9848);
			2681: out = 16'(8727);
			2682: out = 16'(-5899);
			2683: out = 16'(7599);
			2684: out = 16'(1625);
			2685: out = 16'(3063);
			2686: out = 16'(-1607);
			2687: out = 16'(-10458);
			2688: out = 16'(8009);
			2689: out = 16'(-7535);
			2690: out = 16'(3418);
			2691: out = 16'(-1997);
			2692: out = 16'(1571);
			2693: out = 16'(247);
			2694: out = 16'(2070);
			2695: out = 16'(-1210);
			2696: out = 16'(-2247);
			2697: out = 16'(4149);
			2698: out = 16'(3392);
			2699: out = 16'(-7629);
			2700: out = 16'(-8040);
			2701: out = 16'(573);
			2702: out = 16'(-4590);
			2703: out = 16'(-323);
			2704: out = 16'(77);
			2705: out = 16'(2712);
			2706: out = 16'(-10239);
			2707: out = 16'(-9644);
			2708: out = 16'(-1271);
			2709: out = 16'(7290);
			2710: out = 16'(-2639);
			2711: out = 16'(3576);
			2712: out = 16'(3507);
			2713: out = 16'(4387);
			2714: out = 16'(-9153);
			2715: out = 16'(1675);
			2716: out = 16'(3893);
			2717: out = 16'(-11675);
			2718: out = 16'(4608);
			2719: out = 16'(488);
			2720: out = 16'(833);
			2721: out = 16'(500);
			2722: out = 16'(-1925);
			2723: out = 16'(5464);
			2724: out = 16'(-33);
			2725: out = 16'(-1724);
			2726: out = 16'(1808);
			2727: out = 16'(1583);
			2728: out = 16'(1338);
			2729: out = 16'(888);
			2730: out = 16'(6041);
			2731: out = 16'(693);
			2732: out = 16'(-1982);
			2733: out = 16'(-984);
			2734: out = 16'(7120);
			2735: out = 16'(545);
			2736: out = 16'(-590);
			2737: out = 16'(4793);
			2738: out = 16'(113);
			2739: out = 16'(1857);
			2740: out = 16'(5507);
			2741: out = 16'(5882);
			2742: out = 16'(1388);
			2743: out = 16'(-2670);
			2744: out = 16'(5928);
			2745: out = 16'(-8602);
			2746: out = 16'(-620);
			2747: out = 16'(-9950);
			2748: out = 16'(7204);
			2749: out = 16'(1412);
			2750: out = 16'(169);
			2751: out = 16'(1141);
			2752: out = 16'(-2995);
			2753: out = 16'(4622);
			2754: out = 16'(344);
			2755: out = 16'(1407);
			2756: out = 16'(-1565);
			2757: out = 16'(1999);
			2758: out = 16'(444);
			2759: out = 16'(-13386);
			2760: out = 16'(-3732);
			2761: out = 16'(9755);
			2762: out = 16'(1474);
			2763: out = 16'(-10028);
			2764: out = 16'(3267);
			2765: out = 16'(-639);
			2766: out = 16'(-9169);
			2767: out = 16'(-597);
			2768: out = 16'(11305);
			2769: out = 16'(-2166);
			2770: out = 16'(3503);
			2771: out = 16'(7578);
			2772: out = 16'(5414);
			2773: out = 16'(-5439);
			2774: out = 16'(-3395);
			2775: out = 16'(1766);
			2776: out = 16'(3345);
			2777: out = 16'(-4586);
			2778: out = 16'(-702);
			2779: out = 16'(-8885);
			2780: out = 16'(2119);
			2781: out = 16'(796);
			2782: out = 16'(-318);
			2783: out = 16'(6891);
			2784: out = 16'(-1550);
			2785: out = 16'(604);
			2786: out = 16'(-311);
			2787: out = 16'(1367);
			2788: out = 16'(190);
			2789: out = 16'(1271);
			2790: out = 16'(-426);
			2791: out = 16'(3031);
			2792: out = 16'(-1834);
			2793: out = 16'(3422);
			2794: out = 16'(1387);
			2795: out = 16'(2163);
			2796: out = 16'(-11755);
			2797: out = 16'(3625);
			2798: out = 16'(-2339);
			2799: out = 16'(417);
			2800: out = 16'(859);
			2801: out = 16'(3593);
			2802: out = 16'(3195);
			2803: out = 16'(-8188);
			2804: out = 16'(-3303);
			2805: out = 16'(-16);
			2806: out = 16'(-931);
			2807: out = 16'(1082);
			2808: out = 16'(-390);
			2809: out = 16'(2194);
			2810: out = 16'(-4641);
			2811: out = 16'(-831);
			2812: out = 16'(-3106);
			2813: out = 16'(7506);
			2814: out = 16'(2554);
			2815: out = 16'(-5572);
			2816: out = 16'(-4095);
			2817: out = 16'(1498);
			2818: out = 16'(-7262);
			2819: out = 16'(-11488);
			2820: out = 16'(11246);
			2821: out = 16'(1441);
			2822: out = 16'(-5249);
			2823: out = 16'(881);
			2824: out = 16'(5200);
			2825: out = 16'(-5921);
			2826: out = 16'(717);
			2827: out = 16'(2363);
			2828: out = 16'(6258);
			2829: out = 16'(1621);
			2830: out = 16'(-8194);
			2831: out = 16'(694);
			2832: out = 16'(-26);
			2833: out = 16'(1061);
			2834: out = 16'(1788);
			2835: out = 16'(573);
			2836: out = 16'(205);
			2837: out = 16'(1853);
			2838: out = 16'(972);
			2839: out = 16'(4499);
			2840: out = 16'(1092);
			2841: out = 16'(993);
			2842: out = 16'(4094);
			2843: out = 16'(-678);
			2844: out = 16'(-535);
			2845: out = 16'(8087);
			2846: out = 16'(-2494);
			2847: out = 16'(6611);
			2848: out = 16'(4144);
			2849: out = 16'(-10659);
			2850: out = 16'(2291);
			2851: out = 16'(-4028);
			2852: out = 16'(-3382);
			2853: out = 16'(-4958);
			2854: out = 16'(888);
			2855: out = 16'(-6566);
			2856: out = 16'(-1460);
			2857: out = 16'(-232);
			2858: out = 16'(503);
			2859: out = 16'(-2207);
			2860: out = 16'(-4711);
			2861: out = 16'(-692);
			2862: out = 16'(-5762);
			2863: out = 16'(-3754);
			2864: out = 16'(707);
			2865: out = 16'(-570);
			2866: out = 16'(-2935);
			2867: out = 16'(6209);
			2868: out = 16'(-4315);
			2869: out = 16'(4518);
			2870: out = 16'(-5945);
			2871: out = 16'(5631);
			2872: out = 16'(-2057);
			2873: out = 16'(4432);
			2874: out = 16'(-5145);
			2875: out = 16'(-616);
			2876: out = 16'(-1591);
			2877: out = 16'(-627);
			2878: out = 16'(-898);
			2879: out = 16'(-578);
			2880: out = 16'(-4711);
			2881: out = 16'(5684);
			2882: out = 16'(-207);
			2883: out = 16'(-7024);
			2884: out = 16'(397);
			2885: out = 16'(2769);
			2886: out = 16'(-2540);
			2887: out = 16'(6731);
			2888: out = 16'(2754);
			2889: out = 16'(-5095);
			2890: out = 16'(613);
			2891: out = 16'(-426);
			2892: out = 16'(4443);
			2893: out = 16'(-1573);
			2894: out = 16'(-1892);
			2895: out = 16'(-6915);
			2896: out = 16'(3984);
			2897: out = 16'(307);
			2898: out = 16'(1159);
			2899: out = 16'(2903);
			2900: out = 16'(2477);
			2901: out = 16'(623);
			2902: out = 16'(-3932);
			2903: out = 16'(5977);
			2904: out = 16'(-3127);
			2905: out = 16'(-6563);
			2906: out = 16'(2376);
			2907: out = 16'(668);
			2908: out = 16'(1251);
			2909: out = 16'(-1467);
			2910: out = 16'(276);
			2911: out = 16'(1959);
			2912: out = 16'(-1338);
			2913: out = 16'(846);
			2914: out = 16'(4288);
			2915: out = 16'(-676);
			2916: out = 16'(-740);
			2917: out = 16'(-705);
			2918: out = 16'(8058);
			2919: out = 16'(-2770);
			2920: out = 16'(1159);
			2921: out = 16'(96);
			2922: out = 16'(402);
			2923: out = 16'(-1432);
			2924: out = 16'(-1443);
			2925: out = 16'(3616);
			2926: out = 16'(-2943);
			2927: out = 16'(3134);
			2928: out = 16'(-4742);
			2929: out = 16'(-280);
			2930: out = 16'(-796);
			2931: out = 16'(148);
			2932: out = 16'(-88);
			2933: out = 16'(-889);
			2934: out = 16'(4873);
			2935: out = 16'(-8614);
			2936: out = 16'(6504);
			2937: out = 16'(2970);
			2938: out = 16'(2670);
			2939: out = 16'(-3921);
			2940: out = 16'(1642);
			2941: out = 16'(-3881);
			2942: out = 16'(-2987);
			2943: out = 16'(2810);
			2944: out = 16'(-126);
			2945: out = 16'(874);
			2946: out = 16'(1663);
			2947: out = 16'(-2987);
			2948: out = 16'(5701);
			2949: out = 16'(287);
			2950: out = 16'(-6748);
			2951: out = 16'(113);
			2952: out = 16'(-4089);
			2953: out = 16'(7634);
			2954: out = 16'(-7314);
			2955: out = 16'(7051);
			2956: out = 16'(2024);
			2957: out = 16'(3064);
			2958: out = 16'(1328);
			2959: out = 16'(9263);
			2960: out = 16'(-3269);
			2961: out = 16'(-4257);
			2962: out = 16'(-4602);
			2963: out = 16'(426);
			2964: out = 16'(6804);
			2965: out = 16'(-6998);
			2966: out = 16'(-634);
			2967: out = 16'(-1498);
			2968: out = 16'(173);
			2969: out = 16'(-9301);
			2970: out = 16'(8141);
			2971: out = 16'(89);
			2972: out = 16'(16);
			2973: out = 16'(1196);
			2974: out = 16'(10442);
			2975: out = 16'(-5179);
			2976: out = 16'(-8330);
			2977: out = 16'(2389);
			2978: out = 16'(5710);
			2979: out = 16'(-2593);
			2980: out = 16'(-6891);
			2981: out = 16'(4896);
			2982: out = 16'(145);
			2983: out = 16'(-1027);
			2984: out = 16'(-5012);
			2985: out = 16'(4621);
			2986: out = 16'(3001);
			2987: out = 16'(-6386);
			2988: out = 16'(9224);
			2989: out = 16'(-220);
			2990: out = 16'(-1383);
			2991: out = 16'(-537);
			2992: out = 16'(3218);
			2993: out = 16'(96);
			2994: out = 16'(-3514);
			2995: out = 16'(5383);
			2996: out = 16'(-2376);
			2997: out = 16'(3342);
			2998: out = 16'(3662);
			2999: out = 16'(2172);
			3000: out = 16'(-1137);
			3001: out = 16'(-2318);
			3002: out = 16'(-1475);
			3003: out = 16'(890);
			3004: out = 16'(2439);
			3005: out = 16'(1470);
			3006: out = 16'(627);
			3007: out = 16'(268);
			3008: out = 16'(1558);
			3009: out = 16'(3022);
			3010: out = 16'(702);
			3011: out = 16'(-7087);
			3012: out = 16'(3856);
			3013: out = 16'(-2313);
			3014: out = 16'(2297);
			3015: out = 16'(-1400);
			3016: out = 16'(4596);
			3017: out = 16'(875);
			3018: out = 16'(783);
			3019: out = 16'(3276);
			3020: out = 16'(-626);
			3021: out = 16'(-5842);
			3022: out = 16'(-1727);
			3023: out = 16'(10202);
			3024: out = 16'(-2866);
			3025: out = 16'(-2857);
			3026: out = 16'(2811);
			3027: out = 16'(2679);
			3028: out = 16'(869);
			3029: out = 16'(-538);
			3030: out = 16'(8265);
			3031: out = 16'(4281);
			3032: out = 16'(-7764);
			3033: out = 16'(1419);
			3034: out = 16'(-762);
			3035: out = 16'(2826);
			3036: out = 16'(-9066);
			3037: out = 16'(9550);
			3038: out = 16'(2920);
			3039: out = 16'(-8354);
			3040: out = 16'(1802);
			3041: out = 16'(-5746);
			3042: out = 16'(570);
			3043: out = 16'(3476);
			3044: out = 16'(2500);
			3045: out = 16'(-244);
			3046: out = 16'(-3551);
			3047: out = 16'(276);
			3048: out = 16'(-3776);
			3049: out = 16'(3152);
			3050: out = 16'(-1162);
			3051: out = 16'(-430);
			3052: out = 16'(-6675);
			3053: out = 16'(-4720);
			3054: out = 16'(4665);
			3055: out = 16'(-8733);
			3056: out = 16'(2871);
			3057: out = 16'(-2946);
			3058: out = 16'(524);
			3059: out = 16'(523);
			3060: out = 16'(-4676);
			3061: out = 16'(1014);
			3062: out = 16'(2891);
			3063: out = 16'(9245);
			3064: out = 16'(-1346);
			3065: out = 16'(3940);
			3066: out = 16'(-3544);
			3067: out = 16'(-911);
			3068: out = 16'(220);
			3069: out = 16'(2148);
			3070: out = 16'(189);
			3071: out = 16'(-2877);
			3072: out = 16'(3777);
			3073: out = 16'(5505);
			3074: out = 16'(-6323);
			3075: out = 16'(5996);
			3076: out = 16'(-2290);
			3077: out = 16'(-8311);
			3078: out = 16'(-1389);
			3079: out = 16'(2745);
			3080: out = 16'(695);
			3081: out = 16'(-1461);
			3082: out = 16'(10297);
			3083: out = 16'(320);
			3084: out = 16'(-4795);
			3085: out = 16'(-9481);
			3086: out = 16'(3335);
			3087: out = 16'(-2588);
			3088: out = 16'(-1389);
			3089: out = 16'(3960);
			3090: out = 16'(1389);
			3091: out = 16'(-915);
			3092: out = 16'(-11641);
			3093: out = 16'(7200);
			3094: out = 16'(-8868);
			3095: out = 16'(-2443);
			3096: out = 16'(8048);
			3097: out = 16'(-5967);
			3098: out = 16'(-2781);
			3099: out = 16'(-7);
			3100: out = 16'(4161);
			3101: out = 16'(-6273);
			3102: out = 16'(5177);
			3103: out = 16'(2427);
			3104: out = 16'(-3963);
			3105: out = 16'(3640);
			3106: out = 16'(-690);
			3107: out = 16'(2402);
			3108: out = 16'(-2014);
			3109: out = 16'(250);
			3110: out = 16'(5777);
			3111: out = 16'(-7009);
			3112: out = 16'(-6453);
			3113: out = 16'(5315);
			3114: out = 16'(3434);
			3115: out = 16'(3644);
			3116: out = 16'(-894);
			3117: out = 16'(6575);
			3118: out = 16'(-71);
			3119: out = 16'(5696);
			3120: out = 16'(938);
			3121: out = 16'(4459);
			3122: out = 16'(-7178);
			3123: out = 16'(3439);
			3124: out = 16'(298);
			3125: out = 16'(-2555);
			3126: out = 16'(3639);
			3127: out = 16'(-84);
			3128: out = 16'(1729);
			3129: out = 16'(-5048);
			3130: out = 16'(-2130);
			3131: out = 16'(-1327);
			3132: out = 16'(-4249);
			3133: out = 16'(1105);
			3134: out = 16'(3651);
			3135: out = 16'(1708);
			3136: out = 16'(2154);
			3137: out = 16'(-788);
			3138: out = 16'(6093);
			3139: out = 16'(-223);
			3140: out = 16'(2939);
			3141: out = 16'(1244);
			3142: out = 16'(3976);
			3143: out = 16'(4466);
			3144: out = 16'(-6497);
			3145: out = 16'(2096);
			3146: out = 16'(-2401);
			3147: out = 16'(-1340);
			3148: out = 16'(5003);
			3149: out = 16'(79);
			3150: out = 16'(-2682);
			3151: out = 16'(-1275);
			3152: out = 16'(-2649);
			3153: out = 16'(1713);
			3154: out = 16'(6974);
			3155: out = 16'(-6809);
			3156: out = 16'(2344);
			3157: out = 16'(-2460);
			3158: out = 16'(4085);
			3159: out = 16'(-680);
			3160: out = 16'(5800);
			3161: out = 16'(-7474);
			3162: out = 16'(584);
			3163: out = 16'(1202);
			3164: out = 16'(789);
			3165: out = 16'(-2453);
			3166: out = 16'(1405);
			3167: out = 16'(-3885);
			3168: out = 16'(-464);
			3169: out = 16'(-5643);
			3170: out = 16'(930);
			3171: out = 16'(-10090);
			3172: out = 16'(1310);
			3173: out = 16'(4106);
			3174: out = 16'(-480);
			3175: out = 16'(4212);
			3176: out = 16'(3138);
			3177: out = 16'(696);
			3178: out = 16'(-1760);
			3179: out = 16'(407);
			3180: out = 16'(830);
			3181: out = 16'(3021);
			3182: out = 16'(-3473);
			3183: out = 16'(7073);
			3184: out = 16'(-245);
			3185: out = 16'(-7695);
			3186: out = 16'(762);
			3187: out = 16'(4684);
			3188: out = 16'(-7012);
			3189: out = 16'(-1195);
			3190: out = 16'(5408);
			3191: out = 16'(-2152);
			3192: out = 16'(93);
			3193: out = 16'(9454);
			3194: out = 16'(1428);
			3195: out = 16'(-606);
			3196: out = 16'(-1606);
			3197: out = 16'(2219);
			3198: out = 16'(-6669);
			3199: out = 16'(-699);
			3200: out = 16'(3744);
			3201: out = 16'(-125);
			3202: out = 16'(-1212);
			3203: out = 16'(1109);
			3204: out = 16'(2653);
			3205: out = 16'(-3061);
			3206: out = 16'(-1272);
			3207: out = 16'(4280);
			3208: out = 16'(-4899);
			3209: out = 16'(548);
			3210: out = 16'(4103);
			3211: out = 16'(3862);
			3212: out = 16'(162);
			3213: out = 16'(5495);
			3214: out = 16'(-624);
			3215: out = 16'(-7237);
			3216: out = 16'(288);
			3217: out = 16'(75);
			3218: out = 16'(-190);
			3219: out = 16'(-1596);
			3220: out = 16'(3595);
			3221: out = 16'(6209);
			3222: out = 16'(-2731);
			3223: out = 16'(1905);
			3224: out = 16'(-1020);
			3225: out = 16'(-896);
			3226: out = 16'(-3049);
			3227: out = 16'(-3919);
			3228: out = 16'(392);
			3229: out = 16'(-4974);
			3230: out = 16'(2233);
			3231: out = 16'(-7282);
			3232: out = 16'(6375);
			3233: out = 16'(6154);
			3234: out = 16'(-1074);
			3235: out = 16'(-1794);
			3236: out = 16'(343);
			3237: out = 16'(130);
			3238: out = 16'(183);
			3239: out = 16'(3759);
			3240: out = 16'(3888);
			3241: out = 16'(-6635);
			3242: out = 16'(6225);
			3243: out = 16'(-2777);
			3244: out = 16'(1300);
			3245: out = 16'(-1120);
			3246: out = 16'(1884);
			3247: out = 16'(-488);
			3248: out = 16'(-795);
			3249: out = 16'(3586);
			3250: out = 16'(-918);
			3251: out = 16'(-3855);
			3252: out = 16'(1315);
			3253: out = 16'(6688);
			3254: out = 16'(-2225);
			3255: out = 16'(-6480);
			3256: out = 16'(4277);
			3257: out = 16'(-1002);
			3258: out = 16'(-4444);
			3259: out = 16'(4226);
			3260: out = 16'(94);
			3261: out = 16'(330);
			3262: out = 16'(-4081);
			3263: out = 16'(8359);
			3264: out = 16'(-5448);
			3265: out = 16'(-274);
			3266: out = 16'(649);
			3267: out = 16'(7547);
			3268: out = 16'(-440);
			3269: out = 16'(-3176);
			3270: out = 16'(-217);
			3271: out = 16'(1121);
			3272: out = 16'(-4169);
			3273: out = 16'(746);
			3274: out = 16'(1872);
			3275: out = 16'(-4964);
			3276: out = 16'(-4772);
			3277: out = 16'(7124);
			3278: out = 16'(-1657);
			3279: out = 16'(1665);
			3280: out = 16'(-1212);
			3281: out = 16'(2779);
			3282: out = 16'(-10973);
			3283: out = 16'(-3804);
			3284: out = 16'(1068);
			3285: out = 16'(511);
			3286: out = 16'(-2428);
			3287: out = 16'(-10094);
			3288: out = 16'(6320);
			3289: out = 16'(1558);
			3290: out = 16'(-2081);
			3291: out = 16'(1418);
			3292: out = 16'(772);
			3293: out = 16'(-1538);
			3294: out = 16'(-3440);
			3295: out = 16'(1854);
			3296: out = 16'(-1);
			3297: out = 16'(-4676);
			3298: out = 16'(5459);
			3299: out = 16'(6350);
			3300: out = 16'(4577);
			3301: out = 16'(-5411);
			3302: out = 16'(-1926);
			3303: out = 16'(902);
			3304: out = 16'(2933);
			3305: out = 16'(249);
			3306: out = 16'(-1563);
			3307: out = 16'(1336);
			3308: out = 16'(3393);
			3309: out = 16'(1680);
			3310: out = 16'(1695);
			3311: out = 16'(175);
			3312: out = 16'(-2268);
			3313: out = 16'(1911);
			3314: out = 16'(-1625);
			3315: out = 16'(-4393);
			3316: out = 16'(330);
			3317: out = 16'(-2152);
			3318: out = 16'(4559);
			3319: out = 16'(883);
			3320: out = 16'(316);
			3321: out = 16'(-1043);
			3322: out = 16'(2849);
			3323: out = 16'(-436);
			3324: out = 16'(5156);
			3325: out = 16'(-4668);
			3326: out = 16'(2407);
			3327: out = 16'(-5698);
			3328: out = 16'(-422);
			3329: out = 16'(-511);
			3330: out = 16'(687);
			3331: out = 16'(-1724);
			3332: out = 16'(-4741);
			3333: out = 16'(6641);
			3334: out = 16'(-1131);
			3335: out = 16'(407);
			3336: out = 16'(-3687);
			3337: out = 16'(1628);
			3338: out = 16'(-3522);
			3339: out = 16'(-775);
			3340: out = 16'(2382);
			3341: out = 16'(7342);
			3342: out = 16'(-9809);
			3343: out = 16'(7552);
			3344: out = 16'(5362);
			3345: out = 16'(818);
			3346: out = 16'(-5117);
			3347: out = 16'(-1347);
			3348: out = 16'(753);
			3349: out = 16'(774);
			3350: out = 16'(-3435);
			3351: out = 16'(2450);
			3352: out = 16'(-1798);
			3353: out = 16'(12);
			3354: out = 16'(1440);
			3355: out = 16'(-230);
			3356: out = 16'(-552);
			3357: out = 16'(-823);
			3358: out = 16'(-550);
			3359: out = 16'(69);
			3360: out = 16'(2712);
			3361: out = 16'(-7977);
			3362: out = 16'(651);
			3363: out = 16'(2201);
			3364: out = 16'(-235);
			3365: out = 16'(4475);
			3366: out = 16'(4760);
			3367: out = 16'(-2369);
			3368: out = 16'(979);
			3369: out = 16'(2353);
			3370: out = 16'(1606);
			3371: out = 16'(653);
			3372: out = 16'(-5180);
			3373: out = 16'(4339);
			3374: out = 16'(-1339);
			3375: out = 16'(-967);
			3376: out = 16'(4481);
			3377: out = 16'(-1924);
			3378: out = 16'(4700);
			3379: out = 16'(6319);
			3380: out = 16'(-840);
			3381: out = 16'(-7728);
			3382: out = 16'(2456);
			3383: out = 16'(159);
			3384: out = 16'(594);
			3385: out = 16'(1424);
			3386: out = 16'(6149);
			3387: out = 16'(-3017);
			3388: out = 16'(-3599);
			3389: out = 16'(2645);
			3390: out = 16'(422);
			3391: out = 16'(-7370);
			3392: out = 16'(-157);
			3393: out = 16'(2247);
			3394: out = 16'(-642);
			3395: out = 16'(-1363);
			3396: out = 16'(-117);
			3397: out = 16'(2216);
			3398: out = 16'(-2973);
			3399: out = 16'(223);
			3400: out = 16'(2656);
			3401: out = 16'(-6655);
			3402: out = 16'(-655);
			3403: out = 16'(892);
			3404: out = 16'(1677);
			3405: out = 16'(-5316);
			3406: out = 16'(2761);
			3407: out = 16'(-2994);
			3408: out = 16'(-6864);
			3409: out = 16'(-1015);
			3410: out = 16'(1619);
			3411: out = 16'(2257);
			3412: out = 16'(-1904);
			3413: out = 16'(2681);
			3414: out = 16'(-5241);
			3415: out = 16'(1344);
			3416: out = 16'(1878);
			3417: out = 16'(1635);
			3418: out = 16'(-998);
			3419: out = 16'(138);
			3420: out = 16'(659);
			3421: out = 16'(1822);
			3422: out = 16'(-1244);
			3423: out = 16'(2946);
			3424: out = 16'(-536);
			3425: out = 16'(-483);
			3426: out = 16'(1556);
			3427: out = 16'(212);
			3428: out = 16'(-7550);
			3429: out = 16'(3857);
			3430: out = 16'(5813);
			3431: out = 16'(-1993);
			3432: out = 16'(996);
			3433: out = 16'(1077);
			3434: out = 16'(-169);
			3435: out = 16'(3504);
			3436: out = 16'(3553);
			3437: out = 16'(-211);
			3438: out = 16'(-2544);
			3439: out = 16'(4176);
			3440: out = 16'(3113);
			3441: out = 16'(-2665);
			3442: out = 16'(-1232);
			3443: out = 16'(5249);
			3444: out = 16'(-2761);
			3445: out = 16'(446);
			3446: out = 16'(-351);
			3447: out = 16'(-4989);
			3448: out = 16'(-5428);
			3449: out = 16'(917);
			3450: out = 16'(2547);
			3451: out = 16'(-1608);
			3452: out = 16'(-1176);
			3453: out = 16'(-4530);
			3454: out = 16'(2308);
			3455: out = 16'(1261);
			3456: out = 16'(3666);
			3457: out = 16'(-7687);
			3458: out = 16'(95);
			3459: out = 16'(-241);
			3460: out = 16'(-3727);
			3461: out = 16'(4557);
			3462: out = 16'(1054);
			3463: out = 16'(2298);
			3464: out = 16'(-11717);
			3465: out = 16'(-7396);
			3466: out = 16'(4152);
			3467: out = 16'(-3470);
			3468: out = 16'(-2639);
			3469: out = 16'(4097);
			3470: out = 16'(3080);
			3471: out = 16'(-6179);
			3472: out = 16'(-690);
			3473: out = 16'(2988);
			3474: out = 16'(-4290);
			3475: out = 16'(-148);
			3476: out = 16'(4471);
			3477: out = 16'(-8347);
			3478: out = 16'(190);
			3479: out = 16'(-3244);
			3480: out = 16'(8271);
			3481: out = 16'(-8823);
			3482: out = 16'(966);
			3483: out = 16'(5227);
			3484: out = 16'(-949);
			3485: out = 16'(-541);
			3486: out = 16'(2574);
			3487: out = 16'(-6041);
			3488: out = 16'(-436);
			3489: out = 16'(5666);
			3490: out = 16'(6160);
			3491: out = 16'(-2909);
			3492: out = 16'(471);
			3493: out = 16'(2434);
			3494: out = 16'(5562);
			3495: out = 16'(-224);
			3496: out = 16'(3785);
			3497: out = 16'(-227);
			3498: out = 16'(-3710);
			3499: out = 16'(-214);
			3500: out = 16'(650);
			3501: out = 16'(2003);
			3502: out = 16'(-5548);
			3503: out = 16'(5196);
			3504: out = 16'(-7510);
			3505: out = 16'(-5685);
			3506: out = 16'(4607);
			3507: out = 16'(7113);
			3508: out = 16'(727);
			3509: out = 16'(-11424);
			3510: out = 16'(3909);
			3511: out = 16'(3628);
			3512: out = 16'(-11031);
			3513: out = 16'(2676);
			3514: out = 16'(5381);
			3515: out = 16'(-3279);
			3516: out = 16'(-1101);
			3517: out = 16'(3008);
			3518: out = 16'(300);
			3519: out = 16'(-1547);
			3520: out = 16'(2025);
			3521: out = 16'(-1746);
			3522: out = 16'(647);
			3523: out = 16'(-4713);
			3524: out = 16'(-2862);
			3525: out = 16'(1417);
			3526: out = 16'(938);
			3527: out = 16'(4402);
			3528: out = 16'(-679);
			3529: out = 16'(8367);
			3530: out = 16'(-4521);
			3531: out = 16'(-2153);
			3532: out = 16'(-4771);
			3533: out = 16'(6642);
			3534: out = 16'(-5958);
			3535: out = 16'(6083);
			3536: out = 16'(5849);
			3537: out = 16'(-10491);
			3538: out = 16'(3060);
			3539: out = 16'(1043);
			3540: out = 16'(1402);
			3541: out = 16'(-2540);
			3542: out = 16'(-1231);
			3543: out = 16'(4240);
			3544: out = 16'(2137);
			3545: out = 16'(-1245);
			3546: out = 16'(9075);
			3547: out = 16'(-809);
			3548: out = 16'(-2118);
			3549: out = 16'(-6276);
			3550: out = 16'(6708);
			3551: out = 16'(-8448);
			3552: out = 16'(207);
			3553: out = 16'(3795);
			3554: out = 16'(-32);
			3555: out = 16'(-1883);
			3556: out = 16'(826);
			3557: out = 16'(5323);
			3558: out = 16'(-6133);
			3559: out = 16'(5382);
			3560: out = 16'(3289);
			3561: out = 16'(-8835);
			3562: out = 16'(-2251);
			3563: out = 16'(6327);
			3564: out = 16'(-265);
			3565: out = 16'(-3117);
			3566: out = 16'(4989);
			3567: out = 16'(3824);
			3568: out = 16'(-2439);
			3569: out = 16'(-3389);
			3570: out = 16'(3887);
			3571: out = 16'(-628);
			3572: out = 16'(-2563);
			3573: out = 16'(8439);
			3574: out = 16'(2304);
			3575: out = 16'(-4622);
			3576: out = 16'(-3561);
			3577: out = 16'(395);
			3578: out = 16'(-1548);
			3579: out = 16'(-729);
			3580: out = 16'(-1425);
			3581: out = 16'(1589);
			3582: out = 16'(5);
			3583: out = 16'(7952);
			3584: out = 16'(2112);
			3585: out = 16'(322);
			3586: out = 16'(-2696);
			3587: out = 16'(-846);
			3588: out = 16'(-1962);
			3589: out = 16'(-161);
			3590: out = 16'(2904);
			3591: out = 16'(3818);
			3592: out = 16'(1209);
			3593: out = 16'(606);
			3594: out = 16'(2231);
			3595: out = 16'(-5057);
			3596: out = 16'(688);
			3597: out = 16'(-1075);
			3598: out = 16'(-8806);
			3599: out = 16'(1632);
			3600: out = 16'(1813);
			3601: out = 16'(-386);
			3602: out = 16'(-1471);
			3603: out = 16'(6055);
			3604: out = 16'(-2037);
			3605: out = 16'(834);
			3606: out = 16'(2757);
			3607: out = 16'(51);
			3608: out = 16'(-3400);
			3609: out = 16'(2412);
			3610: out = 16'(-65);
			3611: out = 16'(1721);
			3612: out = 16'(-323);
			3613: out = 16'(2212);
			3614: out = 16'(-198);
			3615: out = 16'(2874);
			3616: out = 16'(4716);
			3617: out = 16'(-1158);
			3618: out = 16'(-1805);
			3619: out = 16'(849);
			3620: out = 16'(6745);
			3621: out = 16'(-3495);
			3622: out = 16'(1728);
			3623: out = 16'(525);
			3624: out = 16'(871);
			3625: out = 16'(-3104);
			3626: out = 16'(310);
			3627: out = 16'(-2345);
			3628: out = 16'(544);
			3629: out = 16'(-1748);
			3630: out = 16'(-859);
			3631: out = 16'(-382);
			3632: out = 16'(-2406);
			3633: out = 16'(596);
			3634: out = 16'(2462);
			3635: out = 16'(-4145);
			3636: out = 16'(-4230);
			3637: out = 16'(-806);
			3638: out = 16'(2865);
			3639: out = 16'(-2640);
			3640: out = 16'(927);
			3641: out = 16'(-2349);
			3642: out = 16'(1764);
			3643: out = 16'(-3077);
			3644: out = 16'(-719);
			3645: out = 16'(852);
			3646: out = 16'(1883);
			3647: out = 16'(822);
			3648: out = 16'(-9319);
			3649: out = 16'(5955);
			3650: out = 16'(-1126);
			3651: out = 16'(687);
			3652: out = 16'(1217);
			3653: out = 16'(-268);
			3654: out = 16'(-1026);
			3655: out = 16'(3349);
			3656: out = 16'(3050);
			3657: out = 16'(-1987);
			3658: out = 16'(19);
			3659: out = 16'(4110);
			3660: out = 16'(3855);
			3661: out = 16'(3532);
			3662: out = 16'(-10242);
			3663: out = 16'(323);
			3664: out = 16'(-476);
			3665: out = 16'(1348);
			3666: out = 16'(-504);
			3667: out = 16'(-1154);
			3668: out = 16'(3584);
			3669: out = 16'(-4791);
			3670: out = 16'(7781);
			3671: out = 16'(-3906);
			3672: out = 16'(-4969);
			3673: out = 16'(4879);
			3674: out = 16'(1181);
			3675: out = 16'(-934);
			3676: out = 16'(3882);
			3677: out = 16'(-1412);
			3678: out = 16'(2726);
			3679: out = 16'(2990);
			3680: out = 16'(4370);
			3681: out = 16'(-6576);
			3682: out = 16'(-5269);
			3683: out = 16'(1991);
			3684: out = 16'(2957);
			3685: out = 16'(-39);
			3686: out = 16'(-2876);
			3687: out = 16'(-517);
			3688: out = 16'(-4798);
			3689: out = 16'(4843);
			3690: out = 16'(-2062);
			3691: out = 16'(1706);
			3692: out = 16'(-369);
			3693: out = 16'(584);
			3694: out = 16'(1673);
			3695: out = 16'(-97);
			3696: out = 16'(-562);
			3697: out = 16'(-6395);
			3698: out = 16'(517);
			3699: out = 16'(-2749);
			3700: out = 16'(748);
			3701: out = 16'(1218);
			3702: out = 16'(-1734);
			3703: out = 16'(-473);
			3704: out = 16'(-3384);
			3705: out = 16'(-1668);
			3706: out = 16'(2816);
			3707: out = 16'(-10165);
			3708: out = 16'(6867);
			3709: out = 16'(-7698);
			3710: out = 16'(8964);
			3711: out = 16'(-4256);
			3712: out = 16'(-166);
			3713: out = 16'(-1148);
			3714: out = 16'(1079);
			3715: out = 16'(-2335);
			3716: out = 16'(1264);
			3717: out = 16'(2022);
			3718: out = 16'(-2248);
			3719: out = 16'(5909);
			3720: out = 16'(-166);
			3721: out = 16'(1907);
			3722: out = 16'(-1864);
			3723: out = 16'(707);
			3724: out = 16'(887);
			3725: out = 16'(2732);
			3726: out = 16'(-1606);
			3727: out = 16'(-4836);
			3728: out = 16'(-1294);
			3729: out = 16'(8938);
			3730: out = 16'(575);
			3731: out = 16'(1483);
			3732: out = 16'(73);
			3733: out = 16'(367);
			3734: out = 16'(-3169);
			3735: out = 16'(-1299);
			3736: out = 16'(9164);
			3737: out = 16'(-1705);
			3738: out = 16'(-522);
			3739: out = 16'(1059);
			3740: out = 16'(4305);
			3741: out = 16'(-1563);
			3742: out = 16'(-5615);
			3743: out = 16'(2473);
			3744: out = 16'(55);
			3745: out = 16'(1743);
			3746: out = 16'(-2123);
			3747: out = 16'(1350);
			3748: out = 16'(-2224);
			3749: out = 16'(-4949);
			3750: out = 16'(1488);
			3751: out = 16'(-151);
			3752: out = 16'(392);
			3753: out = 16'(-2482);
			3754: out = 16'(-367);
			3755: out = 16'(1823);
			3756: out = 16'(546);
			3757: out = 16'(1321);
			3758: out = 16'(-588);
			3759: out = 16'(-2820);
			3760: out = 16'(-693);
			3761: out = 16'(-1878);
			3762: out = 16'(1326);
			3763: out = 16'(-1124);
			3764: out = 16'(-329);
			3765: out = 16'(-1014);
			3766: out = 16'(10336);
			3767: out = 16'(-4497);
			3768: out = 16'(-3961);
			3769: out = 16'(10119);
			3770: out = 16'(-2044);
			3771: out = 16'(-6180);
			3772: out = 16'(-1437);
			3773: out = 16'(4143);
			3774: out = 16'(-4465);
			3775: out = 16'(3467);
			3776: out = 16'(5406);
			3777: out = 16'(-297);
			3778: out = 16'(-5831);
			3779: out = 16'(6634);
			3780: out = 16'(-648);
			3781: out = 16'(-53);
			3782: out = 16'(-993);
			3783: out = 16'(862);
			3784: out = 16'(84);
			3785: out = 16'(165);
			3786: out = 16'(1797);
			3787: out = 16'(545);
			3788: out = 16'(4491);
			3789: out = 16'(-1307);
			3790: out = 16'(7339);
			3791: out = 16'(-7108);
			3792: out = 16'(2402);
			3793: out = 16'(242);
			3794: out = 16'(1570);
			3795: out = 16'(843);
			3796: out = 16'(-351);
			3797: out = 16'(2560);
			3798: out = 16'(-7134);
			3799: out = 16'(848);
			3800: out = 16'(-166);
			3801: out = 16'(-74);
			3802: out = 16'(-1026);
			3803: out = 16'(3485);
			3804: out = 16'(496);
			3805: out = 16'(-2351);
			3806: out = 16'(4235);
			3807: out = 16'(1569);
			3808: out = 16'(-1900);
			3809: out = 16'(3121);
			3810: out = 16'(1816);
			3811: out = 16'(5718);
			3812: out = 16'(-1022);
			3813: out = 16'(-4104);
			3814: out = 16'(83);
			3815: out = 16'(55);
			3816: out = 16'(518);
			3817: out = 16'(-2284);
			3818: out = 16'(2224);
			3819: out = 16'(-892);
			3820: out = 16'(-359);
			3821: out = 16'(-750);
			3822: out = 16'(1809);
			3823: out = 16'(-9819);
			3824: out = 16'(-3861);
			3825: out = 16'(7738);
			3826: out = 16'(-2484);
			3827: out = 16'(-1320);
			3828: out = 16'(3267);
			3829: out = 16'(1625);
			3830: out = 16'(-2248);
			3831: out = 16'(-5272);
			3832: out = 16'(2482);
			3833: out = 16'(1197);
			3834: out = 16'(-5571);
			3835: out = 16'(132);
			3836: out = 16'(7337);
			3837: out = 16'(104);
			3838: out = 16'(-6294);
			3839: out = 16'(4534);
			3840: out = 16'(2240);
			3841: out = 16'(-2485);
			3842: out = 16'(2178);
			3843: out = 16'(3352);
			3844: out = 16'(-2629);
			3845: out = 16'(-8239);
			3846: out = 16'(7516);
			3847: out = 16'(-330);
			3848: out = 16'(-8418);
			3849: out = 16'(4194);
			3850: out = 16'(447);
			3851: out = 16'(2232);
			3852: out = 16'(-9396);
			3853: out = 16'(8995);
			3854: out = 16'(-4505);
			3855: out = 16'(796);
			3856: out = 16'(4719);
			3857: out = 16'(-4827);
			3858: out = 16'(-6893);
			3859: out = 16'(-241);
			3860: out = 16'(2279);
			3861: out = 16'(-1459);
			3862: out = 16'(1896);
			3863: out = 16'(4441);
			3864: out = 16'(1047);
			3865: out = 16'(-3729);
			3866: out = 16'(575);
			3867: out = 16'(-1568);
			3868: out = 16'(754);
			3869: out = 16'(-3263);
			3870: out = 16'(6844);
			3871: out = 16'(-4909);
			3872: out = 16'(187);
			3873: out = 16'(-985);
			3874: out = 16'(3767);
			3875: out = 16'(-3813);
			3876: out = 16'(-2864);
			3877: out = 16'(154);
			3878: out = 16'(-2560);
			3879: out = 16'(-163);
			3880: out = 16'(882);
			3881: out = 16'(4152);
			3882: out = 16'(-7374);
			3883: out = 16'(-2568);
			3884: out = 16'(472);
			3885: out = 16'(713);
			3886: out = 16'(1468);
			3887: out = 16'(4141);
			3888: out = 16'(-99);
			3889: out = 16'(4149);
			3890: out = 16'(-1209);
			3891: out = 16'(182);
			3892: out = 16'(-696);
			3893: out = 16'(2059);
			3894: out = 16'(1419);
			3895: out = 16'(5117);
			3896: out = 16'(4763);
			3897: out = 16'(-4640);
			3898: out = 16'(1618);
			3899: out = 16'(511);
			3900: out = 16'(-248);
			3901: out = 16'(-4737);
			3902: out = 16'(-411);
			3903: out = 16'(-2201);
			3904: out = 16'(1823);
			3905: out = 16'(2374);
			3906: out = 16'(3218);
			3907: out = 16'(139);
			3908: out = 16'(-1216);
			3909: out = 16'(2618);
			3910: out = 16'(-647);
			3911: out = 16'(-632);
			3912: out = 16'(-5667);
			3913: out = 16'(6147);
			3914: out = 16'(746);
			3915: out = 16'(2164);
			3916: out = 16'(-5105);
			3917: out = 16'(920);
			3918: out = 16'(-5665);
			3919: out = 16'(3200);
			3920: out = 16'(4720);
			3921: out = 16'(-3958);
			3922: out = 16'(-2617);
			3923: out = 16'(2547);
			3924: out = 16'(4578);
			3925: out = 16'(-1393);
			3926: out = 16'(969);
			3927: out = 16'(83);
			3928: out = 16'(-789);
			3929: out = 16'(-2887);
			3930: out = 16'(823);
			3931: out = 16'(-3081);
			3932: out = 16'(-5323);
			3933: out = 16'(1079);
			3934: out = 16'(-3960);
			3935: out = 16'(-4104);
			3936: out = 16'(7433);
			3937: out = 16'(548);
			3938: out = 16'(122);
			3939: out = 16'(4951);
			3940: out = 16'(507);
			3941: out = 16'(-2385);
			3942: out = 16'(-334);
			3943: out = 16'(484);
			3944: out = 16'(-1771);
			3945: out = 16'(-2247);
			3946: out = 16'(3411);
			3947: out = 16'(2594);
			3948: out = 16'(-4843);
			3949: out = 16'(-10801);
			3950: out = 16'(3020);
			3951: out = 16'(-4552);
			3952: out = 16'(2786);
			3953: out = 16'(-1857);
			3954: out = 16'(4695);
			3955: out = 16'(-5739);
			3956: out = 16'(1873);
			3957: out = 16'(3590);
			3958: out = 16'(-1293);
			3959: out = 16'(-4432);
			3960: out = 16'(3358);
			3961: out = 16'(791);
			3962: out = 16'(-796);
			3963: out = 16'(2148);
			3964: out = 16'(2911);
			3965: out = 16'(480);
			3966: out = 16'(-765);
			3967: out = 16'(1878);
			3968: out = 16'(-7278);
			3969: out = 16'(5999);
			3970: out = 16'(-6543);
			3971: out = 16'(8074);
			3972: out = 16'(-1748);
			3973: out = 16'(3345);
			3974: out = 16'(2148);
			3975: out = 16'(894);
			3976: out = 16'(571);
			3977: out = 16'(-6498);
			3978: out = 16'(-696);
			3979: out = 16'(803);
			3980: out = 16'(2214);
			3981: out = 16'(3038);
			3982: out = 16'(711);
			3983: out = 16'(690);
			3984: out = 16'(-3864);
			3985: out = 16'(2947);
			3986: out = 16'(-160);
			3987: out = 16'(-192);
			3988: out = 16'(-5123);
			3989: out = 16'(869);
			3990: out = 16'(2743);
			3991: out = 16'(1861);
			3992: out = 16'(-208);
			3993: out = 16'(-749);
			3994: out = 16'(-420);
			3995: out = 16'(3942);
			3996: out = 16'(-5750);
			3997: out = 16'(4301);
			3998: out = 16'(1745);
			3999: out = 16'(3771);
			4000: out = 16'(-3556);
			4001: out = 16'(2054);
			4002: out = 16'(-2260);
			4003: out = 16'(514);
			4004: out = 16'(2266);
			4005: out = 16'(-3452);
			4006: out = 16'(3068);
			4007: out = 16'(-7611);
			4008: out = 16'(2416);
			4009: out = 16'(2266);
			4010: out = 16'(-1148);
			4011: out = 16'(-6021);
			4012: out = 16'(3817);
			4013: out = 16'(3014);
			4014: out = 16'(-1457);
			4015: out = 16'(2992);
			4016: out = 16'(7695);
			4017: out = 16'(-10506);
			4018: out = 16'(-1120);
			4019: out = 16'(580);
			4020: out = 16'(2795);
			4021: out = 16'(-3123);
			4022: out = 16'(-17);
			4023: out = 16'(459);
			4024: out = 16'(749);
			4025: out = 16'(3049);
			4026: out = 16'(783);
			4027: out = 16'(-161);
			4028: out = 16'(-1701);
			4029: out = 16'(-2615);
			4030: out = 16'(7539);
			4031: out = 16'(4614);
			4032: out = 16'(-3842);
			4033: out = 16'(-9330);
			4034: out = 16'(6941);
			4035: out = 16'(-4778);
			4036: out = 16'(-2061);
			4037: out = 16'(1969);
			4038: out = 16'(2384);
			4039: out = 16'(-2653);
			4040: out = 16'(-3276);
			4041: out = 16'(7342);
			4042: out = 16'(-7688);
			4043: out = 16'(512);
			4044: out = 16'(739);
			4045: out = 16'(619);
			4046: out = 16'(-360);
			4047: out = 16'(-5851);
			4048: out = 16'(169);
			4049: out = 16'(500);
			4050: out = 16'(-712);
			4051: out = 16'(3776);
			4052: out = 16'(-2426);
			4053: out = 16'(3659);
			4054: out = 16'(-2083);
			4055: out = 16'(4523);
			4056: out = 16'(272);
			4057: out = 16'(-1888);
			4058: out = 16'(5737);
			4059: out = 16'(2104);
			4060: out = 16'(-2630);
			4061: out = 16'(-2280);
			4062: out = 16'(1495);
			4063: out = 16'(-7512);
			4064: out = 16'(-1431);
			4065: out = 16'(3814);
			4066: out = 16'(-385);
			4067: out = 16'(-2993);
			4068: out = 16'(1089);
			4069: out = 16'(431);
			4070: out = 16'(-1203);
			4071: out = 16'(4798);
			4072: out = 16'(-1320);
			4073: out = 16'(541);
			4074: out = 16'(-2336);
			4075: out = 16'(2755);
			4076: out = 16'(3160);
			4077: out = 16'(284);
			4078: out = 16'(-6754);
			4079: out = 16'(780);
			4080: out = 16'(5892);
			4081: out = 16'(-735);
			4082: out = 16'(-6659);
			4083: out = 16'(6725);
			4084: out = 16'(1210);
			4085: out = 16'(-4686);
			4086: out = 16'(6561);
			4087: out = 16'(261);
			4088: out = 16'(-2569);
			4089: out = 16'(-5302);
			4090: out = 16'(10173);
			4091: out = 16'(-3729);
			4092: out = 16'(-2795);
			4093: out = 16'(1110);
			4094: out = 16'(1020);
			4095: out = 16'(-357);
			4096: out = 16'(-421);
			4097: out = 16'(-7174);
			4098: out = 16'(4483);
			4099: out = 16'(-4362);
			4100: out = 16'(-297);
			4101: out = 16'(737);
			4102: out = 16'(-458);
			4103: out = 16'(-5836);
			4104: out = 16'(52);
			4105: out = 16'(1098);
			4106: out = 16'(-5380);
			4107: out = 16'(-3660);
			4108: out = 16'(4425);
			4109: out = 16'(4503);
			4110: out = 16'(-1109);
			4111: out = 16'(6058);
			4112: out = 16'(-3548);
			4113: out = 16'(-2434);
			4114: out = 16'(744);
			4115: out = 16'(1610);
			4116: out = 16'(-3319);
			4117: out = 16'(-425);
			4118: out = 16'(1958);
			4119: out = 16'(-2906);
			4120: out = 16'(-1563);
			4121: out = 16'(1243);
			4122: out = 16'(4902);
			4123: out = 16'(-1080);
			4124: out = 16'(-3220);
			4125: out = 16'(2821);
			4126: out = 16'(1600);
			4127: out = 16'(-9019);
			4128: out = 16'(1808);
			4129: out = 16'(10407);
			4130: out = 16'(-3432);
			4131: out = 16'(1632);
			4132: out = 16'(2084);
			4133: out = 16'(1028);
			4134: out = 16'(-14227);
			4135: out = 16'(6662);
			4136: out = 16'(3488);
			4137: out = 16'(-8645);
			4138: out = 16'(-1927);
			4139: out = 16'(6854);
			4140: out = 16'(1439);
			4141: out = 16'(-862);
			4142: out = 16'(5675);
			4143: out = 16'(-861);
			4144: out = 16'(-3906);
			4145: out = 16'(372);
			4146: out = 16'(-1562);
			4147: out = 16'(762);
			4148: out = 16'(-119);
			4149: out = 16'(-1358);
			4150: out = 16'(4083);
			4151: out = 16'(-793);
			4152: out = 16'(-3727);
			4153: out = 16'(604);
			4154: out = 16'(5301);
			4155: out = 16'(-2405);
			4156: out = 16'(-2492);
			4157: out = 16'(4335);
			4158: out = 16'(-3144);
			4159: out = 16'(-2680);
			4160: out = 16'(2197);
			4161: out = 16'(8317);
			4162: out = 16'(-2580);
			4163: out = 16'(-161);
			4164: out = 16'(-3547);
			4165: out = 16'(1187);
			4166: out = 16'(343);
			4167: out = 16'(-1524);
			4168: out = 16'(2254);
			4169: out = 16'(-386);
			4170: out = 16'(500);
			4171: out = 16'(1012);
			4172: out = 16'(2193);
			4173: out = 16'(-5466);
			4174: out = 16'(97);
			4175: out = 16'(126);
			4176: out = 16'(702);
			4177: out = 16'(-5805);
			4178: out = 16'(7925);
			4179: out = 16'(-3547);
			4180: out = 16'(976);
			4181: out = 16'(2459);
			4182: out = 16'(2887);
			4183: out = 16'(-5265);
			4184: out = 16'(-3323);
			4185: out = 16'(7394);
			4186: out = 16'(-5198);
			4187: out = 16'(4340);
			4188: out = 16'(2119);
			4189: out = 16'(1089);
			4190: out = 16'(-5283);
			4191: out = 16'(4500);
			4192: out = 16'(-405);
			4193: out = 16'(-1497);
			4194: out = 16'(1583);
			4195: out = 16'(729);
			4196: out = 16'(3719);
			4197: out = 16'(628);
			4198: out = 16'(-32);
			4199: out = 16'(-433);
			4200: out = 16'(-1153);
			4201: out = 16'(668);
			4202: out = 16'(1788);
			4203: out = 16'(-2617);
			4204: out = 16'(1058);
			4205: out = 16'(-5927);
			4206: out = 16'(5215);
			4207: out = 16'(-4268);
			4208: out = 16'(-4883);
			4209: out = 16'(-221);
			4210: out = 16'(-262);
			4211: out = 16'(628);
			4212: out = 16'(-1469);
			4213: out = 16'(-422);
			4214: out = 16'(-1509);
			4215: out = 16'(1602);
			4216: out = 16'(1720);
			4217: out = 16'(180);
			4218: out = 16'(-1413);
			4219: out = 16'(3907);
			4220: out = 16'(-2342);
			4221: out = 16'(752);
			4222: out = 16'(-1142);
			4223: out = 16'(-2952);
			4224: out = 16'(-6893);
			4225: out = 16'(7007);
			4226: out = 16'(-155);
			4227: out = 16'(906);
			4228: out = 16'(6319);
			4229: out = 16'(-1367);
			4230: out = 16'(-1681);
			4231: out = 16'(-2549);
			4232: out = 16'(-155);
			4233: out = 16'(-2151);
			4234: out = 16'(1718);
			4235: out = 16'(-2920);
			4236: out = 16'(4230);
			4237: out = 16'(1294);
			4238: out = 16'(-1333);
			4239: out = 16'(1637);
			4240: out = 16'(3436);
			4241: out = 16'(-118);
			4242: out = 16'(-4259);
			4243: out = 16'(2793);
			4244: out = 16'(-1046);
			4245: out = 16'(-341);
			4246: out = 16'(5905);
			4247: out = 16'(784);
			4248: out = 16'(-4737);
			4249: out = 16'(494);
			4250: out = 16'(-453);
			4251: out = 16'(-4234);
			4252: out = 16'(1861);
			4253: out = 16'(121);
			4254: out = 16'(969);
			4255: out = 16'(2029);
			4256: out = 16'(986);
			4257: out = 16'(-4457);
			4258: out = 16'(3803);
			4259: out = 16'(-4653);
			4260: out = 16'(2388);
			4261: out = 16'(115);
			4262: out = 16'(-837);
			4263: out = 16'(-120);
			4264: out = 16'(149);
			4265: out = 16'(4631);
			4266: out = 16'(-2769);
			4267: out = 16'(-5964);
			4268: out = 16'(-1389);
			4269: out = 16'(-148);
			4270: out = 16'(3554);
			4271: out = 16'(5707);
			4272: out = 16'(1392);
			4273: out = 16'(-2927);
			4274: out = 16'(2559);
			4275: out = 16'(265);
			4276: out = 16'(1897);
			4277: out = 16'(-1277);
			4278: out = 16'(1079);
			4279: out = 16'(3187);
			4280: out = 16'(-5598);
			4281: out = 16'(1993);
			4282: out = 16'(-2519);
			4283: out = 16'(-2171);
			4284: out = 16'(-419);
			4285: out = 16'(-1096);
			4286: out = 16'(2775);
			4287: out = 16'(-7686);
			4288: out = 16'(2686);
			4289: out = 16'(1261);
			4290: out = 16'(-1971);
			4291: out = 16'(-4267);
			4292: out = 16'(5274);
			4293: out = 16'(5066);
			4294: out = 16'(-8257);
			4295: out = 16'(6818);
			4296: out = 16'(-1997);
			4297: out = 16'(-1632);
			4298: out = 16'(2509);
			4299: out = 16'(1555);
			4300: out = 16'(-3997);
			4301: out = 16'(665);
			4302: out = 16'(931);
			4303: out = 16'(-889);
			4304: out = 16'(-299);
			4305: out = 16'(5539);
			4306: out = 16'(-4291);
			4307: out = 16'(-1195);
			4308: out = 16'(-1856);
			4309: out = 16'(1064);
			4310: out = 16'(-2006);
			4311: out = 16'(-1813);
			4312: out = 16'(4601);
			4313: out = 16'(280);
			4314: out = 16'(-1207);
			4315: out = 16'(-4666);
			4316: out = 16'(2101);
			4317: out = 16'(-964);
			4318: out = 16'(-5014);
			4319: out = 16'(-325);
			4320: out = 16'(2296);
			4321: out = 16'(-1855);
			4322: out = 16'(-3505);
			4323: out = 16'(4517);
			4324: out = 16'(-580);
			4325: out = 16'(-3735);
			4326: out = 16'(2660);
			4327: out = 16'(5365);
			4328: out = 16'(239);
			4329: out = 16'(-11401);
			4330: out = 16'(2786);
			4331: out = 16'(1843);
			4332: out = 16'(-5649);
			4333: out = 16'(21);
			4334: out = 16'(4749);
			4335: out = 16'(558);
			4336: out = 16'(-7118);
			4337: out = 16'(3333);
			4338: out = 16'(2254);
			4339: out = 16'(-3441);
			4340: out = 16'(-999);
			4341: out = 16'(113);
			4342: out = 16'(1400);
			4343: out = 16'(-9287);
			4344: out = 16'(4554);
			4345: out = 16'(5710);
			4346: out = 16'(-920);
			4347: out = 16'(-2114);
			4348: out = 16'(5511);
			4349: out = 16'(2736);
			4350: out = 16'(-3808);
			4351: out = 16'(425);
			4352: out = 16'(-1386);
			4353: out = 16'(-2560);
			4354: out = 16'(-1232);
			4355: out = 16'(2452);
			4356: out = 16'(4283);
			4357: out = 16'(1421);
			4358: out = 16'(-5966);
			4359: out = 16'(209);
			4360: out = 16'(749);
			4361: out = 16'(1215);
			4362: out = 16'(-1948);
			4363: out = 16'(6177);
			4364: out = 16'(6723);
			4365: out = 16'(587);
			4366: out = 16'(5472);
			4367: out = 16'(-2216);
			4368: out = 16'(-4597);
			4369: out = 16'(196);
			4370: out = 16'(163);
			4371: out = 16'(359);
			4372: out = 16'(-884);
			4373: out = 16'(2181);
			4374: out = 16'(-361);
			4375: out = 16'(1282);
			4376: out = 16'(-1374);
			4377: out = 16'(1565);
			4378: out = 16'(-4990);
			4379: out = 16'(-303);
			4380: out = 16'(-282);
			4381: out = 16'(-129);
			4382: out = 16'(-825);
			4383: out = 16'(4191);
			4384: out = 16'(-1314);
			4385: out = 16'(1982);
			4386: out = 16'(-928);
			4387: out = 16'(4404);
			4388: out = 16'(-4093);
			4389: out = 16'(409);
			4390: out = 16'(4592);
			4391: out = 16'(1741);
			4392: out = 16'(-343);
			4393: out = 16'(-3714);
			4394: out = 16'(1484);
			4395: out = 16'(-6371);
			4396: out = 16'(-92);
			4397: out = 16'(3195);
			4398: out = 16'(-4166);
			4399: out = 16'(-6849);
			4400: out = 16'(2361);
			4401: out = 16'(1243);
			4402: out = 16'(-460);
			4403: out = 16'(-6268);
			4404: out = 16'(6768);
			4405: out = 16'(-2780);
			4406: out = 16'(2423);
			4407: out = 16'(-1021);
			4408: out = 16'(-564);
			4409: out = 16'(-887);
			4410: out = 16'(-3640);
			4411: out = 16'(6122);
			4412: out = 16'(-1644);
			4413: out = 16'(-33);
			4414: out = 16'(-1338);
			4415: out = 16'(3194);
			4416: out = 16'(198);
			4417: out = 16'(-7621);
			4418: out = 16'(1594);
			4419: out = 16'(-3651);
			4420: out = 16'(2842);
			4421: out = 16'(2826);
			4422: out = 16'(3805);
			4423: out = 16'(1980);
			4424: out = 16'(-847);
			4425: out = 16'(3621);
			4426: out = 16'(-424);
			4427: out = 16'(563);
			4428: out = 16'(-132);
			4429: out = 16'(-855);
			4430: out = 16'(1491);
			4431: out = 16'(-533);
			4432: out = 16'(1838);
			4433: out = 16'(-134);
			4434: out = 16'(557);
			4435: out = 16'(-6491);
			4436: out = 16'(-1464);
			4437: out = 16'(2696);
			4438: out = 16'(-2110);
			4439: out = 16'(716);
			4440: out = 16'(-813);
			4441: out = 16'(5620);
			4442: out = 16'(-1698);
			4443: out = 16'(-2819);
			4444: out = 16'(1391);
			4445: out = 16'(-3493);
			4446: out = 16'(779);
			4447: out = 16'(-983);
			4448: out = 16'(1702);
			4449: out = 16'(-2952);
			4450: out = 16'(-816);
			4451: out = 16'(6366);
			4452: out = 16'(-8317);
			4453: out = 16'(114);
			4454: out = 16'(-4724);
			4455: out = 16'(4440);
			4456: out = 16'(1443);
			4457: out = 16'(734);
			4458: out = 16'(2427);
			4459: out = 16'(-1423);
			4460: out = 16'(2226);
			4461: out = 16'(456);
			4462: out = 16'(1412);
			4463: out = 16'(-4343);
			4464: out = 16'(-56);
			4465: out = 16'(7722);
			4466: out = 16'(-2362);
			4467: out = 16'(1291);
			4468: out = 16'(-2154);
			4469: out = 16'(-1679);
			4470: out = 16'(714);
			4471: out = 16'(1533);
			4472: out = 16'(-1396);
			4473: out = 16'(-7098);
			4474: out = 16'(5739);
			4475: out = 16'(1420);
			4476: out = 16'(1479);
			4477: out = 16'(-2212);
			4478: out = 16'(1650);
			4479: out = 16'(-3942);
			4480: out = 16'(-1503);
			4481: out = 16'(2786);
			4482: out = 16'(-768);
			4483: out = 16'(1906);
			4484: out = 16'(2243);
			4485: out = 16'(-3350);
			4486: out = 16'(-1281);
			4487: out = 16'(-2870);
			4488: out = 16'(5927);
			4489: out = 16'(-6747);
			4490: out = 16'(1053);
			4491: out = 16'(1747);
			4492: out = 16'(-3453);
			4493: out = 16'(-260);
			4494: out = 16'(-2752);
			4495: out = 16'(237);
			4496: out = 16'(136);
			4497: out = 16'(-60);
			4498: out = 16'(2384);
			4499: out = 16'(197);
			4500: out = 16'(1643);
			4501: out = 16'(420);
			4502: out = 16'(1804);
			4503: out = 16'(-4144);
			4504: out = 16'(-1833);
			4505: out = 16'(1405);
			4506: out = 16'(-1420);
			4507: out = 16'(6906);
			4508: out = 16'(-163);
			4509: out = 16'(3786);
			4510: out = 16'(-1924);
			4511: out = 16'(5486);
			4512: out = 16'(-2732);
			4513: out = 16'(-7209);
			4514: out = 16'(1974);
			4515: out = 16'(2793);
			4516: out = 16'(-2554);
			4517: out = 16'(-6612);
			4518: out = 16'(2343);
			4519: out = 16'(-6847);
			4520: out = 16'(-4021);
			4521: out = 16'(4875);
			4522: out = 16'(25);
			4523: out = 16'(196);
			4524: out = 16'(-3220);
			4525: out = 16'(1549);
			4526: out = 16'(2623);
			4527: out = 16'(62);
			4528: out = 16'(4003);
			4529: out = 16'(-2974);
			4530: out = 16'(-5625);
			4531: out = 16'(1471);
			4532: out = 16'(12);
			4533: out = 16'(878);
			4534: out = 16'(-2537);
			4535: out = 16'(2671);
			4536: out = 16'(-40);
			4537: out = 16'(-2228);
			4538: out = 16'(-1852);
			4539: out = 16'(5145);
			4540: out = 16'(-5438);
			4541: out = 16'(1202);
			4542: out = 16'(6005);
			4543: out = 16'(-520);
			4544: out = 16'(1277);
			4545: out = 16'(780);
			4546: out = 16'(-3641);
			4547: out = 16'(128);
			4548: out = 16'(-622);
			4549: out = 16'(1187);
			4550: out = 16'(959);
			4551: out = 16'(1231);
			4552: out = 16'(4986);
			4553: out = 16'(-1370);
			4554: out = 16'(287);
			4555: out = 16'(-3358);
			4556: out = 16'(1216);
			4557: out = 16'(-3473);
			4558: out = 16'(1672);
			4559: out = 16'(-2935);
			4560: out = 16'(452);
			4561: out = 16'(5699);
			4562: out = 16'(-61);
			4563: out = 16'(-2775);
			4564: out = 16'(388);
			4565: out = 16'(-1799);
			4566: out = 16'(1740);
			4567: out = 16'(701);
			4568: out = 16'(1915);
			4569: out = 16'(-5596);
			4570: out = 16'(-1106);
			4571: out = 16'(6666);
			4572: out = 16'(-3047);
			4573: out = 16'(-3408);
			4574: out = 16'(88);
			4575: out = 16'(1127);
			4576: out = 16'(-5744);
			4577: out = 16'(1938);
			4578: out = 16'(3043);
			4579: out = 16'(654);
			4580: out = 16'(974);
			4581: out = 16'(-207);
			4582: out = 16'(2097);
			4583: out = 16'(-6838);
			4584: out = 16'(-1758);
			4585: out = 16'(4531);
			4586: out = 16'(912);
			4587: out = 16'(-3060);
			4588: out = 16'(5508);
			4589: out = 16'(2445);
			4590: out = 16'(-2158);
			4591: out = 16'(1802);
			4592: out = 16'(4094);
			4593: out = 16'(-7959);
			4594: out = 16'(886);
			4595: out = 16'(-118);
			4596: out = 16'(97);
			4597: out = 16'(-4705);
			4598: out = 16'(1610);
			4599: out = 16'(6454);
			4600: out = 16'(-4217);
			4601: out = 16'(1014);
			4602: out = 16'(-1322);
			4603: out = 16'(2093);
			4604: out = 16'(-3297);
			4605: out = 16'(1693);
			4606: out = 16'(8769);
			4607: out = 16'(-1932);
			4608: out = 16'(1118);
			4609: out = 16'(373);
			4610: out = 16'(-851);
			4611: out = 16'(-256);
			4612: out = 16'(-4180);
			4613: out = 16'(5375);
			4614: out = 16'(-8297);
			4615: out = 16'(1324);
			4616: out = 16'(2786);
			4617: out = 16'(2235);
			4618: out = 16'(2714);
			4619: out = 16'(-515);
			4620: out = 16'(422);
			4621: out = 16'(-3206);
			4622: out = 16'(-5034);
			4623: out = 16'(3059);
			4624: out = 16'(862);
			4625: out = 16'(930);
			4626: out = 16'(748);
			4627: out = 16'(6439);
			4628: out = 16'(-782);
			4629: out = 16'(-897);
			4630: out = 16'(375);
			4631: out = 16'(2186);
			4632: out = 16'(-3670);
			4633: out = 16'(-6487);
			4634: out = 16'(4785);
			4635: out = 16'(-4065);
			4636: out = 16'(-2975);
			4637: out = 16'(-3320);
			4638: out = 16'(566);
			4639: out = 16'(-4452);
			4640: out = 16'(171);
			4641: out = 16'(5865);
			4642: out = 16'(659);
			4643: out = 16'(309);
			4644: out = 16'(1099);
			4645: out = 16'(3558);
			4646: out = 16'(254);
			4647: out = 16'(-4757);
			4648: out = 16'(2547);
			4649: out = 16'(133);
			4650: out = 16'(-134);
			4651: out = 16'(-829);
			4652: out = 16'(771);
			4653: out = 16'(689);
			4654: out = 16'(-2498);
			4655: out = 16'(5625);
			4656: out = 16'(2049);
			4657: out = 16'(-5176);
			4658: out = 16'(-190);
			4659: out = 16'(2321);
			4660: out = 16'(-381);
			4661: out = 16'(-5162);
			4662: out = 16'(5090);
			4663: out = 16'(-218);
			4664: out = 16'(-650);
			4665: out = 16'(805);
			4666: out = 16'(3027);
			4667: out = 16'(-667);
			4668: out = 16'(3570);
			4669: out = 16'(1390);
			4670: out = 16'(-415);
			4671: out = 16'(469);
			4672: out = 16'(-2354);
			4673: out = 16'(-4446);
			4674: out = 16'(-871);
			4675: out = 16'(-2827);
			4676: out = 16'(1040);
			4677: out = 16'(392);
			4678: out = 16'(-832);
			4679: out = 16'(321);
			4680: out = 16'(698);
			4681: out = 16'(-2544);
			4682: out = 16'(315);
			4683: out = 16'(2399);
			4684: out = 16'(-3021);
			4685: out = 16'(-430);
			4686: out = 16'(3472);
			4687: out = 16'(1771);
			4688: out = 16'(-1441);
			4689: out = 16'(-1286);
			4690: out = 16'(3186);
			4691: out = 16'(-7);
			4692: out = 16'(-5645);
			4693: out = 16'(3229);
			4694: out = 16'(-3609);
			4695: out = 16'(4614);
			4696: out = 16'(-4779);
			4697: out = 16'(1429);
			4698: out = 16'(-1307);
			4699: out = 16'(-1700);
			4700: out = 16'(666);
			4701: out = 16'(3106);
			4702: out = 16'(-4598);
			4703: out = 16'(-3197);
			4704: out = 16'(1471);
			4705: out = 16'(6364);
			4706: out = 16'(-4263);
			4707: out = 16'(-1574);
			4708: out = 16'(42);
			4709: out = 16'(2655);
			4710: out = 16'(-5662);
			4711: out = 16'(650);
			4712: out = 16'(5909);
			4713: out = 16'(-7901);
			4714: out = 16'(2197);
			4715: out = 16'(-427);
			4716: out = 16'(487);
			4717: out = 16'(-6015);
			4718: out = 16'(2739);
			4719: out = 16'(284);
			4720: out = 16'(-2242);
			4721: out = 16'(-1246);
			4722: out = 16'(-4339);
			4723: out = 16'(631);
			4724: out = 16'(2246);
			4725: out = 16'(-825);
			4726: out = 16'(827);
			4727: out = 16'(2679);
			4728: out = 16'(-1949);
			4729: out = 16'(-166);
			4730: out = 16'(2249);
			4731: out = 16'(-2169);
			4732: out = 16'(-3183);
			4733: out = 16'(917);
			4734: out = 16'(-269);
			4735: out = 16'(115);
			4736: out = 16'(-2265);
			4737: out = 16'(1724);
			4738: out = 16'(1056);
			4739: out = 16'(1121);
			4740: out = 16'(2746);
			4741: out = 16'(-4004);
			4742: out = 16'(2415);
			4743: out = 16'(-2963);
			4744: out = 16'(5716);
			4745: out = 16'(2259);
			4746: out = 16'(-1229);
			4747: out = 16'(501);
			4748: out = 16'(-496);
			4749: out = 16'(-3891);
			4750: out = 16'(-1357);
			4751: out = 16'(-2117);
			4752: out = 16'(-3644);
			4753: out = 16'(-3207);
			4754: out = 16'(3674);
			4755: out = 16'(-3910);
			4756: out = 16'(5257);
			4757: out = 16'(964);
			4758: out = 16'(-2554);
			4759: out = 16'(214);
			4760: out = 16'(-8658);
			4761: out = 16'(6578);
			4762: out = 16'(-5482);
			4763: out = 16'(3985);
			4764: out = 16'(3107);
			4765: out = 16'(3330);
			4766: out = 16'(-1689);
			4767: out = 16'(5508);
			4768: out = 16'(-3266);
			4769: out = 16'(-3086);
			4770: out = 16'(4341);
			4771: out = 16'(-4448);
			4772: out = 16'(-2353);
			4773: out = 16'(1963);
			4774: out = 16'(-520);
			4775: out = 16'(1822);
			4776: out = 16'(-3300);
			4777: out = 16'(6050);
			4778: out = 16'(-5816);
			4779: out = 16'(-3366);
			4780: out = 16'(3981);
			4781: out = 16'(161);
			4782: out = 16'(1624);
			4783: out = 16'(-1169);
			4784: out = 16'(1579);
			4785: out = 16'(-1657);
			4786: out = 16'(2713);
			4787: out = 16'(-588);
			4788: out = 16'(-3449);
			4789: out = 16'(4730);
			4790: out = 16'(-1244);
			4791: out = 16'(4197);
			4792: out = 16'(-889);
			4793: out = 16'(-2855);
			4794: out = 16'(-461);
			4795: out = 16'(-2833);
			4796: out = 16'(5239);
			4797: out = 16'(-3722);
			4798: out = 16'(10);
			4799: out = 16'(117);
			4800: out = 16'(2587);
			4801: out = 16'(-339);
			4802: out = 16'(359);
			4803: out = 16'(-342);
			4804: out = 16'(462);
			4805: out = 16'(-1327);
			4806: out = 16'(272);
			4807: out = 16'(-1528);
			4808: out = 16'(746);
			4809: out = 16'(-5596);
			4810: out = 16'(3513);
			4811: out = 16'(983);
			4812: out = 16'(-1847);
			4813: out = 16'(-1661);
			4814: out = 16'(1057);
			4815: out = 16'(174);
			4816: out = 16'(524);
			4817: out = 16'(3326);
			4818: out = 16'(-2799);
			4819: out = 16'(682);
			4820: out = 16'(-524);
			4821: out = 16'(2435);
			4822: out = 16'(428);
			4823: out = 16'(-740);
			4824: out = 16'(-845);
			4825: out = 16'(265);
			4826: out = 16'(2994);
			4827: out = 16'(-6573);
			4828: out = 16'(898);
			4829: out = 16'(3308);
			4830: out = 16'(-433);
			4831: out = 16'(-3347);
			4832: out = 16'(1980);
			4833: out = 16'(2284);
			4834: out = 16'(-1117);
			4835: out = 16'(630);
			4836: out = 16'(-592);
			4837: out = 16'(-2307);
			4838: out = 16'(-1221);
			4839: out = 16'(-694);
			4840: out = 16'(3961);
			4841: out = 16'(7722);
			4842: out = 16'(-4370);
			4843: out = 16'(4607);
			4844: out = 16'(367);
			4845: out = 16'(-47);
			4846: out = 16'(-9298);
			4847: out = 16'(5213);
			4848: out = 16'(704);
			4849: out = 16'(-1134);
			4850: out = 16'(601);
			4851: out = 16'(4260);
			4852: out = 16'(-4456);
			4853: out = 16'(73);
			4854: out = 16'(1843);
			4855: out = 16'(366);
			4856: out = 16'(-4926);
			4857: out = 16'(4894);
			4858: out = 16'(5071);
			4859: out = 16'(-2921);
			4860: out = 16'(233);
			4861: out = 16'(4299);
			4862: out = 16'(-3882);
			4863: out = 16'(-4637);
			4864: out = 16'(690);
			4865: out = 16'(-2609);
			4866: out = 16'(1916);
			4867: out = 16'(-3746);
			4868: out = 16'(3302);
			4869: out = 16'(-2228);
			4870: out = 16'(-3839);
			4871: out = 16'(2039);
			4872: out = 16'(2389);
			4873: out = 16'(-2228);
			4874: out = 16'(5019);
			4875: out = 16'(1577);
			4876: out = 16'(-3085);
			4877: out = 16'(518);
			4878: out = 16'(3042);
			4879: out = 16'(-3568);
			4880: out = 16'(2024);
			4881: out = 16'(6857);
			4882: out = 16'(-1630);
			4883: out = 16'(-2897);
			4884: out = 16'(1821);
			4885: out = 16'(-232);
			4886: out = 16'(-148);
			4887: out = 16'(-3371);
			4888: out = 16'(4310);
			4889: out = 16'(-4713);
			4890: out = 16'(4818);
			4891: out = 16'(2663);
			4892: out = 16'(-3712);
			4893: out = 16'(1955);
			4894: out = 16'(-5110);
			4895: out = 16'(-232);
			4896: out = 16'(4260);
			4897: out = 16'(201);
			4898: out = 16'(-3917);
			4899: out = 16'(4007);
			4900: out = 16'(4258);
			4901: out = 16'(-2534);
			4902: out = 16'(-1020);
			4903: out = 16'(-533);
			4904: out = 16'(68);
			4905: out = 16'(-7964);
			4906: out = 16'(2731);
			4907: out = 16'(5830);
			4908: out = 16'(-3894);
			4909: out = 16'(232);
			4910: out = 16'(3174);
			4911: out = 16'(-635);
			4912: out = 16'(-4863);
			4913: out = 16'(897);
			4914: out = 16'(3488);
			4915: out = 16'(-4243);
			4916: out = 16'(-3161);
			4917: out = 16'(4857);
			4918: out = 16'(-1929);
			4919: out = 16'(-4890);
			4920: out = 16'(1992);
			4921: out = 16'(4406);
			4922: out = 16'(-8857);
			4923: out = 16'(2861);
			4924: out = 16'(2288);
			4925: out = 16'(1026);
			4926: out = 16'(-3992);
			4927: out = 16'(1409);
			4928: out = 16'(1812);
			4929: out = 16'(-5669);
			4930: out = 16'(-386);
			4931: out = 16'(5855);
			4932: out = 16'(-1495);
			4933: out = 16'(257);
			4934: out = 16'(2802);
			4935: out = 16'(-432);
			4936: out = 16'(-3099);
			4937: out = 16'(-161);
			4938: out = 16'(1649);
			4939: out = 16'(-998);
			4940: out = 16'(3205);
			4941: out = 16'(-3462);
			4942: out = 16'(5825);
			4943: out = 16'(-4242);
			4944: out = 16'(-942);
			4945: out = 16'(4035);
			4946: out = 16'(-878);
			4947: out = 16'(-6166);
			4948: out = 16'(3042);
			4949: out = 16'(5064);
			4950: out = 16'(-8582);
			4951: out = 16'(5514);
			4952: out = 16'(2501);
			4953: out = 16'(-799);
			4954: out = 16'(-4328);
			4955: out = 16'(-1160);
			4956: out = 16'(427);
			4957: out = 16'(-5593);
			4958: out = 16'(5878);
			4959: out = 16'(462);
			4960: out = 16'(2765);
			4961: out = 16'(283);
			4962: out = 16'(-2234);
			4963: out = 16'(3257);
			4964: out = 16'(-1678);
			4965: out = 16'(-2506);
			4966: out = 16'(606);
			4967: out = 16'(-264);
			4968: out = 16'(1739);
			4969: out = 16'(-514);
			4970: out = 16'(2441);
			4971: out = 16'(-3259);
			4972: out = 16'(590);
			4973: out = 16'(2231);
			4974: out = 16'(-1717);
			4975: out = 16'(-978);
			4976: out = 16'(142);
			4977: out = 16'(270);
			4978: out = 16'(20);
			4979: out = 16'(413);
			4980: out = 16'(-1872);
			4981: out = 16'(1004);
			4982: out = 16'(555);
			4983: out = 16'(632);
			4984: out = 16'(2425);
			4985: out = 16'(-964);
			4986: out = 16'(-676);
			4987: out = 16'(-2891);
			4988: out = 16'(1909);
			4989: out = 16'(-1505);
			4990: out = 16'(-2565);
			4991: out = 16'(5624);
			4992: out = 16'(-393);
			4993: out = 16'(-528);
			4994: out = 16'(587);
			4995: out = 16'(881);
			4996: out = 16'(-5466);
			4997: out = 16'(-95);
			4998: out = 16'(7114);
			4999: out = 16'(-9984);
			5000: out = 16'(-844);
			5001: out = 16'(7092);
			5002: out = 16'(197);
			5003: out = 16'(-1876);
			5004: out = 16'(451);
			5005: out = 16'(707);
			5006: out = 16'(-3133);
			5007: out = 16'(1163);
			5008: out = 16'(889);
			5009: out = 16'(-3241);
			5010: out = 16'(1413);
			5011: out = 16'(3422);
			5012: out = 16'(-2239);
			5013: out = 16'(4);
			5014: out = 16'(-5748);
			5015: out = 16'(667);
			5016: out = 16'(5516);
			5017: out = 16'(580);
			5018: out = 16'(390);
			5019: out = 16'(1518);
			5020: out = 16'(1003);
			5021: out = 16'(-3212);
			5022: out = 16'(-66);
			5023: out = 16'(-4850);
			5024: out = 16'(-1546);
			5025: out = 16'(477);
			5026: out = 16'(-7);
			5027: out = 16'(-4998);
			5028: out = 16'(6101);
			5029: out = 16'(-1339);
			5030: out = 16'(49);
			5031: out = 16'(1044);
			5032: out = 16'(-3000);
			5033: out = 16'(-304);
			5034: out = 16'(480);
			5035: out = 16'(5840);
			5036: out = 16'(392);
			5037: out = 16'(-228);
			5038: out = 16'(3650);
			5039: out = 16'(-2156);
			5040: out = 16'(-2198);
			5041: out = 16'(3084);
			5042: out = 16'(-2131);
			5043: out = 16'(4083);
			5044: out = 16'(339);
			5045: out = 16'(-180);
			5046: out = 16'(285);
			5047: out = 16'(-1414);
			5048: out = 16'(-2051);
			5049: out = 16'(-7732);
			5050: out = 16'(4312);
			5051: out = 16'(-4638);
			5052: out = 16'(1403);
			5053: out = 16'(3679);
			5054: out = 16'(3062);
			5055: out = 16'(-4639);
			5056: out = 16'(4620);
			5057: out = 16'(-1583);
			5058: out = 16'(1693);
			5059: out = 16'(898);
			5060: out = 16'(969);
			5061: out = 16'(-1252);
			5062: out = 16'(99);
			5063: out = 16'(3482);
			5064: out = 16'(-4700);
			5065: out = 16'(1992);
			5066: out = 16'(-1197);
			5067: out = 16'(-237);
			5068: out = 16'(-1204);
			5069: out = 16'(2252);
			5070: out = 16'(-1870);
			5071: out = 16'(134);
			5072: out = 16'(1108);
			5073: out = 16'(682);
			5074: out = 16'(-1557);
			5075: out = 16'(3037);
			5076: out = 16'(-2489);
			5077: out = 16'(515);
			5078: out = 16'(3314);
			5079: out = 16'(193);
			5080: out = 16'(-695);
			5081: out = 16'(1664);
			5082: out = 16'(-2584);
			5083: out = 16'(5621);
			5084: out = 16'(-2603);
			5085: out = 16'(318);
			5086: out = 16'(-2507);
			5087: out = 16'(-304);
			5088: out = 16'(-1493);
			5089: out = 16'(-1321);
			5090: out = 16'(2471);
			5091: out = 16'(-224);
			5092: out = 16'(261);
			5093: out = 16'(809);
			5094: out = 16'(595);
			5095: out = 16'(-436);
			5096: out = 16'(-54);
			5097: out = 16'(1986);
			5098: out = 16'(-1632);
			5099: out = 16'(1880);
			5100: out = 16'(-2345);
			5101: out = 16'(-5338);
			5102: out = 16'(5169);
			5103: out = 16'(-5776);
			5104: out = 16'(-1130);
			5105: out = 16'(-256);
			5106: out = 16'(-1516);
			5107: out = 16'(-2248);
			5108: out = 16'(884);
			5109: out = 16'(3007);
			5110: out = 16'(-2935);
			5111: out = 16'(1646);
			5112: out = 16'(2562);
			5113: out = 16'(-3357);
			5114: out = 16'(-868);
			5115: out = 16'(4294);
			5116: out = 16'(2074);
			5117: out = 16'(-1298);
			5118: out = 16'(2443);
			5119: out = 16'(-607);
			5120: out = 16'(505);
			5121: out = 16'(1340);
			5122: out = 16'(-2104);
			5123: out = 16'(-788);
			5124: out = 16'(-1777);
			5125: out = 16'(-1260);
			5126: out = 16'(6209);
			5127: out = 16'(-5366);
			5128: out = 16'(-2735);
			5129: out = 16'(-267);
			5130: out = 16'(1465);
			5131: out = 16'(-6068);
			5132: out = 16'(1839);
			5133: out = 16'(-716);
			5134: out = 16'(403);
			5135: out = 16'(4305);
			5136: out = 16'(2288);
			5137: out = 16'(1649);
			5138: out = 16'(-1405);
			5139: out = 16'(96);
			5140: out = 16'(441);
			5141: out = 16'(-4166);
			5142: out = 16'(1746);
			5143: out = 16'(945);
			5144: out = 16'(-2059);
			5145: out = 16'(-1310);
			5146: out = 16'(-53);
			5147: out = 16'(2889);
			5148: out = 16'(-4742);
			5149: out = 16'(-942);
			5150: out = 16'(-222);
			5151: out = 16'(3984);
			5152: out = 16'(-2499);
			5153: out = 16'(2499);
			5154: out = 16'(3344);
			5155: out = 16'(414);
			5156: out = 16'(-603);
			5157: out = 16'(2982);
			5158: out = 16'(-1702);
			5159: out = 16'(-3818);
			5160: out = 16'(-4750);
			5161: out = 16'(4192);
			5162: out = 16'(-1813);
			5163: out = 16'(270);
			5164: out = 16'(917);
			5165: out = 16'(-2186);
			5166: out = 16'(-2195);
			5167: out = 16'(2429);
			5168: out = 16'(-827);
			5169: out = 16'(-893);
			5170: out = 16'(3102);
			5171: out = 16'(-2544);
			5172: out = 16'(258);
			5173: out = 16'(1229);
			5174: out = 16'(-1375);
			5175: out = 16'(1530);
			5176: out = 16'(1991);
			5177: out = 16'(662);
			5178: out = 16'(83);
			5179: out = 16'(-1934);
			5180: out = 16'(-1140);
			5181: out = 16'(-1596);
			5182: out = 16'(6339);
			5183: out = 16'(-5153);
			5184: out = 16'(-3394);
			5185: out = 16'(-1012);
			5186: out = 16'(-639);
			5187: out = 16'(-849);
			5188: out = 16'(2972);
			5189: out = 16'(2815);
			5190: out = 16'(-3177);
			5191: out = 16'(-283);
			5192: out = 16'(1826);
			5193: out = 16'(176);
			5194: out = 16'(1362);
			5195: out = 16'(-570);
			5196: out = 16'(5574);
			5197: out = 16'(-1349);
			5198: out = 16'(-532);
			5199: out = 16'(3712);
			5200: out = 16'(578);
			5201: out = 16'(-4996);
			5202: out = 16'(-2801);
			5203: out = 16'(5690);
			5204: out = 16'(-8095);
			5205: out = 16'(-3324);
			5206: out = 16'(4205);
			5207: out = 16'(3924);
			5208: out = 16'(-2063);
			5209: out = 16'(-4902);
			5210: out = 16'(4805);
			5211: out = 16'(-5133);
			5212: out = 16'(-1591);
			5213: out = 16'(6566);
			5214: out = 16'(795);
			5215: out = 16'(-3552);
			5216: out = 16'(2314);
			5217: out = 16'(577);
			5218: out = 16'(-1098);
			5219: out = 16'(-4849);
			5220: out = 16'(3091);
			5221: out = 16'(-3948);
			5222: out = 16'(718);
			5223: out = 16'(-2037);
			5224: out = 16'(638);
			5225: out = 16'(-1026);
			5226: out = 16'(495);
			5227: out = 16'(2069);
			5228: out = 16'(-524);
			5229: out = 16'(-212);
			5230: out = 16'(-6464);
			5231: out = 16'(6253);
			5232: out = 16'(97);
			5233: out = 16'(1733);
			5234: out = 16'(-220);
			5235: out = 16'(498);
			5236: out = 16'(-3665);
			5237: out = 16'(3154);
			5238: out = 16'(723);
			5239: out = 16'(-2509);
			5240: out = 16'(-706);
			5241: out = 16'(5173);
			5242: out = 16'(-669);
			5243: out = 16'(209);
			5244: out = 16'(-967);
			5245: out = 16'(1105);
			5246: out = 16'(1772);
			5247: out = 16'(1202);
			5248: out = 16'(690);
			5249: out = 16'(-4521);
			5250: out = 16'(3153);
			5251: out = 16'(-907);
			5252: out = 16'(3084);
			5253: out = 16'(-638);
			5254: out = 16'(1244);
			5255: out = 16'(-303);
			5256: out = 16'(1500);
			5257: out = 16'(224);
			5258: out = 16'(-913);
			5259: out = 16'(363);
			5260: out = 16'(-895);
			5261: out = 16'(-106);
			5262: out = 16'(1158);
			5263: out = 16'(-1019);
			5264: out = 16'(1116);
			5265: out = 16'(414);
			5266: out = 16'(1149);
			5267: out = 16'(-1133);
			5268: out = 16'(581);
			5269: out = 16'(-210);
			5270: out = 16'(-977);
			5271: out = 16'(2245);
			5272: out = 16'(-641);
			5273: out = 16'(905);
			5274: out = 16'(3637);
			5275: out = 16'(-498);
			5276: out = 16'(-1424);
			5277: out = 16'(674);
			5278: out = 16'(574);
			5279: out = 16'(-443);
			5280: out = 16'(1714);
			5281: out = 16'(-7);
			5282: out = 16'(92);
			5283: out = 16'(1884);
			5284: out = 16'(-575);
			5285: out = 16'(-1791);
			5286: out = 16'(-6035);
			5287: out = 16'(4048);
			5288: out = 16'(101);
			5289: out = 16'(-1937);
			5290: out = 16'(2921);
			5291: out = 16'(-1620);
			5292: out = 16'(223);
			5293: out = 16'(-163);
			5294: out = 16'(2001);
			5295: out = 16'(-5634);
			5296: out = 16'(-4752);
			5297: out = 16'(3812);
			5298: out = 16'(434);
			5299: out = 16'(708);
			5300: out = 16'(-19);
			5301: out = 16'(1098);
			5302: out = 16'(715);
			5303: out = 16'(1645);
			5304: out = 16'(549);
			5305: out = 16'(-3659);
			5306: out = 16'(-3076);
			5307: out = 16'(1012);
			5308: out = 16'(-3918);
			5309: out = 16'(28);
			5310: out = 16'(-1145);
			5311: out = 16'(294);
			5312: out = 16'(841);
			5313: out = 16'(884);
			5314: out = 16'(1552);
			5315: out = 16'(-148);
			5316: out = 16'(2756);
			5317: out = 16'(2147);
			5318: out = 16'(-650);
			5319: out = 16'(-268);
			5320: out = 16'(-1200);
			5321: out = 16'(2533);
			5322: out = 16'(-5532);
			5323: out = 16'(-579);
			5324: out = 16'(1882);
			5325: out = 16'(-3211);
			5326: out = 16'(-372);
			5327: out = 16'(4712);
			5328: out = 16'(-133);
			5329: out = 16'(-4168);
			5330: out = 16'(-396);
			5331: out = 16'(-408);
			5332: out = 16'(-847);
			5333: out = 16'(-247);
			5334: out = 16'(1544);
			5335: out = 16'(731);
			5336: out = 16'(386);
			5337: out = 16'(333);
			5338: out = 16'(3233);
			5339: out = 16'(-2617);
			5340: out = 16'(-720);
			5341: out = 16'(-611);
			5342: out = 16'(2410);
			5343: out = 16'(-5355);
			5344: out = 16'(213);
			5345: out = 16'(1295);
			5346: out = 16'(-1490);
			5347: out = 16'(-4852);
			5348: out = 16'(-2625);
			5349: out = 16'(3540);
			5350: out = 16'(-3677);
			5351: out = 16'(2058);
			5352: out = 16'(3820);
			5353: out = 16'(7);
			5354: out = 16'(413);
			5355: out = 16'(-3853);
			5356: out = 16'(1949);
			5357: out = 16'(-2798);
			5358: out = 16'(-3956);
			5359: out = 16'(5026);
			5360: out = 16'(66);
			5361: out = 16'(2237);
			5362: out = 16'(-1286);
			5363: out = 16'(877);
			5364: out = 16'(-3539);
			5365: out = 16'(377);
			5366: out = 16'(-836);
			5367: out = 16'(-4108);
			5368: out = 16'(1659);
			5369: out = 16'(-3773);
			5370: out = 16'(5025);
			5371: out = 16'(731);
			5372: out = 16'(2478);
			5373: out = 16'(3321);
			5374: out = 16'(-5118);
			5375: out = 16'(467);
			5376: out = 16'(1787);
			5377: out = 16'(1364);
			5378: out = 16'(1328);
			5379: out = 16'(-509);
			5380: out = 16'(1726);
			5381: out = 16'(-1144);
			5382: out = 16'(-720);
			5383: out = 16'(-1765);
			5384: out = 16'(-727);
			5385: out = 16'(-3701);
			5386: out = 16'(1588);
			5387: out = 16'(-355);
			5388: out = 16'(-1455);
			5389: out = 16'(3344);
			5390: out = 16'(-1317);
			5391: out = 16'(4787);
			5392: out = 16'(-2079);
			5393: out = 16'(-2034);
			5394: out = 16'(5528);
			5395: out = 16'(2713);
			5396: out = 16'(-5187);
			5397: out = 16'(251);
			5398: out = 16'(4007);
			5399: out = 16'(-617);
			5400: out = 16'(-2229);
			5401: out = 16'(4146);
			5402: out = 16'(-3433);
			5403: out = 16'(1062);
			5404: out = 16'(-1228);
			5405: out = 16'(64);
			5406: out = 16'(-2534);
			5407: out = 16'(-6052);
			5408: out = 16'(5834);
			5409: out = 16'(-5896);
			5410: out = 16'(191);
			5411: out = 16'(630);
			5412: out = 16'(7);
			5413: out = 16'(129);
			5414: out = 16'(320);
			5415: out = 16'(2805);
			5416: out = 16'(-1451);
			5417: out = 16'(-156);
			5418: out = 16'(913);
			5419: out = 16'(235);
			5420: out = 16'(-4068);
			5421: out = 16'(502);
			5422: out = 16'(1704);
			5423: out = 16'(-3636);
			5424: out = 16'(2779);
			5425: out = 16'(1681);
			5426: out = 16'(3056);
			5427: out = 16'(606);
			5428: out = 16'(-2215);
			5429: out = 16'(5071);
			5430: out = 16'(-5784);
			5431: out = 16'(3861);
			5432: out = 16'(1219);
			5433: out = 16'(3011);
			5434: out = 16'(-2995);
			5435: out = 16'(-99);
			5436: out = 16'(6375);
			5437: out = 16'(-642);
			5438: out = 16'(-769);
			5439: out = 16'(-1223);
			5440: out = 16'(1336);
			5441: out = 16'(-5424);
			5442: out = 16'(-3855);
			5443: out = 16'(1299);
			5444: out = 16'(2544);
			5445: out = 16'(433);
			5446: out = 16'(1572);
			5447: out = 16'(475);
			5448: out = 16'(-1417);
			5449: out = 16'(-4732);
			5450: out = 16'(5447);
			5451: out = 16'(493);
			5452: out = 16'(-2291);
			5453: out = 16'(-344);
			5454: out = 16'(1447);
			5455: out = 16'(498);
			5456: out = 16'(-2910);
			5457: out = 16'(2473);
			5458: out = 16'(-4114);
			5459: out = 16'(-648);
			5460: out = 16'(1947);
			5461: out = 16'(664);
			5462: out = 16'(-1652);
			5463: out = 16'(-2487);
			5464: out = 16'(3532);
			5465: out = 16'(-2533);
			5466: out = 16'(-47);
			5467: out = 16'(-907);
			5468: out = 16'(1711);
			5469: out = 16'(5652);
			5470: out = 16'(-3089);
			5471: out = 16'(235);
			5472: out = 16'(-669);
			5473: out = 16'(-431);
			5474: out = 16'(-2022);
			5475: out = 16'(2497);
			5476: out = 16'(41);
			5477: out = 16'(566);
			5478: out = 16'(50);
			5479: out = 16'(189);
			5480: out = 16'(-446);
			5481: out = 16'(555);
			5482: out = 16'(3025);
			5483: out = 16'(-506);
			5484: out = 16'(-2936);
			5485: out = 16'(2192);
			5486: out = 16'(-108);
			5487: out = 16'(506);
			5488: out = 16'(-1142);
			5489: out = 16'(812);
			5490: out = 16'(-114);
			5491: out = 16'(-5771);
			5492: out = 16'(2130);
			5493: out = 16'(2839);
			5494: out = 16'(664);
			5495: out = 16'(-1768);
			5496: out = 16'(5821);
			5497: out = 16'(-1415);
			5498: out = 16'(-7349);
			5499: out = 16'(3964);
			5500: out = 16'(601);
			5501: out = 16'(-2780);
			5502: out = 16'(1282);
			5503: out = 16'(-1210);
			5504: out = 16'(986);
			5505: out = 16'(-296);
			5506: out = 16'(4039);
			5507: out = 16'(681);
			5508: out = 16'(-2198);
			5509: out = 16'(2761);
			5510: out = 16'(708);
			5511: out = 16'(-4);
			5512: out = 16'(-4110);
			5513: out = 16'(2072);
			5514: out = 16'(-357);
			5515: out = 16'(-1242);
			5516: out = 16'(3625);
			5517: out = 16'(-2897);
			5518: out = 16'(4547);
			5519: out = 16'(-140);
			5520: out = 16'(109);
			5521: out = 16'(-302);
			5522: out = 16'(-391);
			5523: out = 16'(-202);
			5524: out = 16'(-281);
			5525: out = 16'(-215);
			5526: out = 16'(-3616);
			5527: out = 16'(2346);
			5528: out = 16'(1166);
			5529: out = 16'(-1051);
			5530: out = 16'(3236);
			5531: out = 16'(-1717);
			5532: out = 16'(3247);
			5533: out = 16'(-4365);
			5534: out = 16'(1790);
			5535: out = 16'(-1724);
			5536: out = 16'(3528);
			5537: out = 16'(673);
			5538: out = 16'(261);
			5539: out = 16'(584);
			5540: out = 16'(-3696);
			5541: out = 16'(-3810);
			5542: out = 16'(1762);
			5543: out = 16'(1252);
			5544: out = 16'(-2822);
			5545: out = 16'(2635);
			5546: out = 16'(810);
			5547: out = 16'(-434);
			5548: out = 16'(-2031);
			5549: out = 16'(3672);
			5550: out = 16'(-5348);
			5551: out = 16'(2746);
			5552: out = 16'(-4275);
			5553: out = 16'(3);
			5554: out = 16'(12);
			5555: out = 16'(4560);
			5556: out = 16'(1421);
			5557: out = 16'(-3790);
			5558: out = 16'(297);
			5559: out = 16'(-3749);
			5560: out = 16'(3899);
			5561: out = 16'(1729);
			5562: out = 16'(-3283);
			5563: out = 16'(1745);
			5564: out = 16'(806);
			5565: out = 16'(-682);
			5566: out = 16'(1213);
			5567: out = 16'(27);
			5568: out = 16'(-1233);
			5569: out = 16'(-2284);
			5570: out = 16'(2873);
			5571: out = 16'(-158);
			5572: out = 16'(483);
			5573: out = 16'(71);
			5574: out = 16'(1351);
			5575: out = 16'(-391);
			5576: out = 16'(400);
			5577: out = 16'(-375);
			5578: out = 16'(228);
			5579: out = 16'(218);
			5580: out = 16'(-274);
			5581: out = 16'(9);
			5582: out = 16'(-3932);
			5583: out = 16'(-1032);
			5584: out = 16'(1935);
			5585: out = 16'(-3731);
			5586: out = 16'(700);
			5587: out = 16'(2117);
			5588: out = 16'(861);
			5589: out = 16'(1898);
			5590: out = 16'(147);
			5591: out = 16'(-447);
			5592: out = 16'(-1497);
			5593: out = 16'(-66);
			5594: out = 16'(881);
			5595: out = 16'(598);
			5596: out = 16'(99);
			5597: out = 16'(-1147);
			5598: out = 16'(2168);
			5599: out = 16'(-5017);
			5600: out = 16'(1151);
			5601: out = 16'(-104);
			5602: out = 16'(-4932);
			5603: out = 16'(-328);
			5604: out = 16'(2050);
			5605: out = 16'(-1291);
			5606: out = 16'(1558);
			5607: out = 16'(1624);
			5608: out = 16'(319);
			5609: out = 16'(-2754);
			5610: out = 16'(3190);
			5611: out = 16'(-1508);
			5612: out = 16'(-324);
			5613: out = 16'(2471);
			5614: out = 16'(601);
			5615: out = 16'(-237);
			5616: out = 16'(2068);
			5617: out = 16'(3298);
			5618: out = 16'(-4544);
			5619: out = 16'(4535);
			5620: out = 16'(-926);
			5621: out = 16'(-852);
			5622: out = 16'(-1504);
			5623: out = 16'(946);
			5624: out = 16'(-2466);
			5625: out = 16'(293);
			5626: out = 16'(-3385);
			5627: out = 16'(-134);
			5628: out = 16'(491);
			5629: out = 16'(584);
			5630: out = 16'(611);
			5631: out = 16'(1314);
			5632: out = 16'(1447);
			5633: out = 16'(1117);
			5634: out = 16'(-74);
			5635: out = 16'(353);
			5636: out = 16'(-280);
			5637: out = 16'(59);
			5638: out = 16'(-83);
			5639: out = 16'(1414);
			5640: out = 16'(-774);
			5641: out = 16'(122);
			5642: out = 16'(-1715);
			5643: out = 16'(-164);
			5644: out = 16'(-4854);
			5645: out = 16'(1335);
			5646: out = 16'(2259);
			5647: out = 16'(21);
			5648: out = 16'(-1160);
			5649: out = 16'(-337);
			5650: out = 16'(3036);
			5651: out = 16'(-3240);
			5652: out = 16'(312);
			5653: out = 16'(953);
			5654: out = 16'(1568);
			5655: out = 16'(-3180);
			5656: out = 16'(1910);
			5657: out = 16'(47);
			5658: out = 16'(-3009);
			5659: out = 16'(-212);
			5660: out = 16'(2249);
			5661: out = 16'(-4606);
			5662: out = 16'(1485);
			5663: out = 16'(2107);
			5664: out = 16'(1521);
			5665: out = 16'(-732);
			5666: out = 16'(648);
			5667: out = 16'(-614);
			5668: out = 16'(2067);
			5669: out = 16'(814);
			5670: out = 16'(-1181);
			5671: out = 16'(4097);
			5672: out = 16'(-1350);
			5673: out = 16'(486);
			5674: out = 16'(-383);
			5675: out = 16'(-320);
			5676: out = 16'(-2534);
			5677: out = 16'(-197);
			5678: out = 16'(510);
			5679: out = 16'(-645);
			5680: out = 16'(430);
			5681: out = 16'(617);
			5682: out = 16'(-831);
			5683: out = 16'(-562);
			5684: out = 16'(1024);
			5685: out = 16'(407);
			5686: out = 16'(-1198);
			5687: out = 16'(2144);
			5688: out = 16'(309);
			5689: out = 16'(-1166);
			5690: out = 16'(736);
			5691: out = 16'(218);
			5692: out = 16'(-43);
			5693: out = 16'(-2718);
			5694: out = 16'(1390);
			5695: out = 16'(2750);
			5696: out = 16'(-5795);
			5697: out = 16'(1039);
			5698: out = 16'(-5122);
			5699: out = 16'(2111);
			5700: out = 16'(-2889);
			5701: out = 16'(-79);
			5702: out = 16'(-611);
			5703: out = 16'(-687);
			5704: out = 16'(1218);
			5705: out = 16'(1722);
			5706: out = 16'(338);
			5707: out = 16'(-4225);
			5708: out = 16'(2632);
			5709: out = 16'(2552);
			5710: out = 16'(-1557);
			5711: out = 16'(4116);
			5712: out = 16'(-1290);
			5713: out = 16'(-693);
			5714: out = 16'(-1946);
			5715: out = 16'(4440);
			5716: out = 16'(-2725);
			5717: out = 16'(-4129);
			5718: out = 16'(906);
			5719: out = 16'(35);
			5720: out = 16'(-70);
			5721: out = 16'(-3576);
			5722: out = 16'(3210);
			5723: out = 16'(2229);
			5724: out = 16'(1713);
			5725: out = 16'(-3176);
			5726: out = 16'(-203);
			5727: out = 16'(-111);
			5728: out = 16'(-815);
			5729: out = 16'(99);
			5730: out = 16'(4691);
			5731: out = 16'(-3248);
			5732: out = 16'(454);
			5733: out = 16'(629);
			5734: out = 16'(463);
			5735: out = 16'(-4482);
			5736: out = 16'(-1038);
			5737: out = 16'(975);
			5738: out = 16'(-131);
			5739: out = 16'(312);
			5740: out = 16'(2027);
			5741: out = 16'(3699);
			5742: out = 16'(-4757);
			5743: out = 16'(561);
			5744: out = 16'(2546);
			5745: out = 16'(-3812);
			5746: out = 16'(1180);
			5747: out = 16'(630);
			5748: out = 16'(2012);
			5749: out = 16'(-1404);
			5750: out = 16'(549);
			5751: out = 16'(1904);
			5752: out = 16'(-1710);
			5753: out = 16'(-12);
			5754: out = 16'(225);
			5755: out = 16'(-1925);
			5756: out = 16'(-427);
			5757: out = 16'(-2133);
			5758: out = 16'(1194);
			5759: out = 16'(-4606);
			5760: out = 16'(401);
			5761: out = 16'(-594);
			5762: out = 16'(-499);
			5763: out = 16'(-1056);
			5764: out = 16'(273);
			5765: out = 16'(4085);
			5766: out = 16'(-1379);
			5767: out = 16'(1861);
			5768: out = 16'(-170);
			5769: out = 16'(-1243);
			5770: out = 16'(-480);
			5771: out = 16'(136);
			5772: out = 16'(2021);
			5773: out = 16'(2015);
			5774: out = 16'(-3155);
			5775: out = 16'(139);
			5776: out = 16'(46);
			5777: out = 16'(-3432);
			5778: out = 16'(668);
			5779: out = 16'(2570);
			5780: out = 16'(-291);
			5781: out = 16'(-354);
			5782: out = 16'(540);
			5783: out = 16'(18);
			5784: out = 16'(-915);
			5785: out = 16'(264);
			5786: out = 16'(-217);
			5787: out = 16'(-2176);
			5788: out = 16'(-2178);
			5789: out = 16'(2678);
			5790: out = 16'(2386);
			5791: out = 16'(1256);
			5792: out = 16'(-199);
			5793: out = 16'(-219);
			5794: out = 16'(-2887);
			5795: out = 16'(-2738);
			5796: out = 16'(1031);
			5797: out = 16'(-175);
			5798: out = 16'(-1389);
			5799: out = 16'(1345);
			5800: out = 16'(4635);
			5801: out = 16'(-2605);
			5802: out = 16'(1424);
			5803: out = 16'(1825);
			5804: out = 16'(-5337);
			5805: out = 16'(-1604);
			5806: out = 16'(1421);
			5807: out = 16'(-488);
			5808: out = 16'(-268);
			5809: out = 16'(1637);
			5810: out = 16'(2249);
			5811: out = 16'(1265);
			5812: out = 16'(-2715);
			5813: out = 16'(288);
			5814: out = 16'(378);
			5815: out = 16'(632);
			5816: out = 16'(-876);
			5817: out = 16'(-377);
			5818: out = 16'(756);
			5819: out = 16'(-698);
			5820: out = 16'(-205);
			5821: out = 16'(-2073);
			5822: out = 16'(1220);
			5823: out = 16'(-1579);
			5824: out = 16'(2924);
			5825: out = 16'(1671);
			5826: out = 16'(661);
			5827: out = 16'(-2004);
			5828: out = 16'(2316);
			5829: out = 16'(4079);
			5830: out = 16'(-4959);
			5831: out = 16'(-2168);
			5832: out = 16'(-2649);
			5833: out = 16'(-1303);
			5834: out = 16'(2061);
			5835: out = 16'(612);
			5836: out = 16'(-822);
			5837: out = 16'(84);
			5838: out = 16'(-152);
			5839: out = 16'(175);
			5840: out = 16'(-134);
			5841: out = 16'(-1025);
			5842: out = 16'(-1320);
			5843: out = 16'(544);
			5844: out = 16'(1238);
			5845: out = 16'(-1685);
			5846: out = 16'(-621);
			5847: out = 16'(646);
			5848: out = 16'(14);
			5849: out = 16'(-1578);
			5850: out = 16'(1263);
			5851: out = 16'(-621);
			5852: out = 16'(4192);
			5853: out = 16'(1298);
			5854: out = 16'(-791);
			5855: out = 16'(29);
			5856: out = 16'(-1333);
			5857: out = 16'(320);
			5858: out = 16'(-3693);
			5859: out = 16'(771);
			5860: out = 16'(-6443);
			5861: out = 16'(3665);
			5862: out = 16'(3518);
			5863: out = 16'(1683);
			5864: out = 16'(598);
			5865: out = 16'(-1081);
			5866: out = 16'(-1376);
			5867: out = 16'(276);
			5868: out = 16'(-804);
			5869: out = 16'(3091);
			5870: out = 16'(-2074);
			5871: out = 16'(722);
			5872: out = 16'(2891);
			5873: out = 16'(-3301);
			5874: out = 16'(1004);
			5875: out = 16'(-4006);
			5876: out = 16'(-1424);
			5877: out = 16'(-859);
			5878: out = 16'(2635);
			5879: out = 16'(-241);
			5880: out = 16'(1552);
			5881: out = 16'(-587);
			5882: out = 16'(-1042);
			5883: out = 16'(83);
			5884: out = 16'(-2864);
			5885: out = 16'(-1771);
			5886: out = 16'(1842);
			5887: out = 16'(799);
			5888: out = 16'(1948);
			5889: out = 16'(5433);
			5890: out = 16'(1862);
			5891: out = 16'(-2434);
			5892: out = 16'(-2955);
			5893: out = 16'(-487);
			5894: out = 16'(-171);
			5895: out = 16'(-3538);
			5896: out = 16'(2922);
			5897: out = 16'(2986);
			5898: out = 16'(-1695);
			5899: out = 16'(1305);
			5900: out = 16'(273);
			5901: out = 16'(-33);
			5902: out = 16'(371);
			5903: out = 16'(-2425);
			5904: out = 16'(-874);
			5905: out = 16'(-2512);
			5906: out = 16'(4251);
			5907: out = 16'(1418);
			5908: out = 16'(1835);
			5909: out = 16'(3398);
			5910: out = 16'(-2342);
			5911: out = 16'(-723);
			5912: out = 16'(-1127);
			5913: out = 16'(-179);
			5914: out = 16'(1287);
			5915: out = 16'(-461);
			5916: out = 16'(-383);
			5917: out = 16'(-151);
			5918: out = 16'(1753);
			5919: out = 16'(-2385);
			5920: out = 16'(535);
			5921: out = 16'(-2797);
			5922: out = 16'(-2385);
			5923: out = 16'(1051);
			5924: out = 16'(881);
			5925: out = 16'(1089);
			5926: out = 16'(1479);
			5927: out = 16'(1407);
			5928: out = 16'(-1137);
			5929: out = 16'(2162);
			5930: out = 16'(-757);
			5931: out = 16'(-1241);
			5932: out = 16'(-1112);
			5933: out = 16'(-356);
			5934: out = 16'(-60);
			5935: out = 16'(2372);
			5936: out = 16'(-885);
			5937: out = 16'(-1215);
			5938: out = 16'(-3187);
			5939: out = 16'(4525);
			5940: out = 16'(-4645);
			5941: out = 16'(1786);
			5942: out = 16'(-138);
			5943: out = 16'(545);
			5944: out = 16'(2135);
			5945: out = 16'(-835);
			5946: out = 16'(2681);
			5947: out = 16'(-3884);
			5948: out = 16'(-344);
			5949: out = 16'(3071);
			5950: out = 16'(-3982);
			5951: out = 16'(-2586);
			5952: out = 16'(-36);
			5953: out = 16'(2168);
			5954: out = 16'(89);
			5955: out = 16'(-921);
			5956: out = 16'(-312);
			5957: out = 16'(-1385);
			5958: out = 16'(-293);
			5959: out = 16'(184);
			5960: out = 16'(411);
			5961: out = 16'(-2588);
			5962: out = 16'(991);
			5963: out = 16'(3389);
			5964: out = 16'(-710);
			5965: out = 16'(1858);
			5966: out = 16'(-8);
			5967: out = 16'(313);
			5968: out = 16'(430);
			5969: out = 16'(-3990);
			5970: out = 16'(1983);
			5971: out = 16'(-289);
			5972: out = 16'(-763);
			5973: out = 16'(2629);
			5974: out = 16'(1552);
			5975: out = 16'(-5842);
			5976: out = 16'(196);
			5977: out = 16'(-451);
			5978: out = 16'(-3379);
			5979: out = 16'(1839);
			5980: out = 16'(938);
			5981: out = 16'(1255);
			5982: out = 16'(118);
			5983: out = 16'(-142);
			5984: out = 16'(3817);
			5985: out = 16'(-299);
			5986: out = 16'(1138);
			5987: out = 16'(-42);
			5988: out = 16'(-263);
			5989: out = 16'(-863);
			5990: out = 16'(-780);
			5991: out = 16'(1586);
			5992: out = 16'(-1629);
			5993: out = 16'(234);
			5994: out = 16'(-758);
			5995: out = 16'(-1329);
			5996: out = 16'(-1744);
			5997: out = 16'(2467);
			5998: out = 16'(2494);
			5999: out = 16'(-4547);
			6000: out = 16'(677);
			6001: out = 16'(1321);
			6002: out = 16'(-23);
			6003: out = 16'(2406);
			6004: out = 16'(-1830);
			6005: out = 16'(1878);
			6006: out = 16'(-243);
			6007: out = 16'(405);
			6008: out = 16'(31);
			6009: out = 16'(664);
			6010: out = 16'(-5167);
			6011: out = 16'(738);
			6012: out = 16'(1495);
			6013: out = 16'(-375);
			6014: out = 16'(0);
			6015: out = 16'(-576);
			6016: out = 16'(3069);
			6017: out = 16'(312);
			6018: out = 16'(-2860);
			6019: out = 16'(4215);
			6020: out = 16'(-1082);
			6021: out = 16'(-2389);
			6022: out = 16'(-282);
			6023: out = 16'(589);
			6024: out = 16'(-1584);
			6025: out = 16'(-1166);
			6026: out = 16'(698);
			6027: out = 16'(1316);
			6028: out = 16'(-1713);
			6029: out = 16'(3710);
			6030: out = 16'(2952);
			6031: out = 16'(-1292);
			6032: out = 16'(-4527);
			6033: out = 16'(408);
			6034: out = 16'(-1121);
			6035: out = 16'(-1548);
			6036: out = 16'(1615);
			6037: out = 16'(-2240);
			6038: out = 16'(-1088);
			6039: out = 16'(686);
			6040: out = 16'(4274);
			6041: out = 16'(-662);
			6042: out = 16'(519);
			6043: out = 16'(-1543);
			6044: out = 16'(1504);
			6045: out = 16'(-18);
			6046: out = 16'(2736);
			6047: out = 16'(1286);
			6048: out = 16'(-3192);
			6049: out = 16'(1580);
			6050: out = 16'(1272);
			6051: out = 16'(-1461);
			6052: out = 16'(-1057);
			6053: out = 16'(1029);
			6054: out = 16'(135);
			6055: out = 16'(886);
			6056: out = 16'(353);
			6057: out = 16'(-599);
			6058: out = 16'(-44);
			6059: out = 16'(92);
			6060: out = 16'(-4836);
			6061: out = 16'(600);
			6062: out = 16'(2189);
			6063: out = 16'(-2421);
			6064: out = 16'(6107);
			6065: out = 16'(2263);
			6066: out = 16'(-1564);
			6067: out = 16'(-3925);
			6068: out = 16'(1364);
			6069: out = 16'(-1304);
			6070: out = 16'(-1659);
			6071: out = 16'(467);
			6072: out = 16'(358);
			6073: out = 16'(1266);
			6074: out = 16'(259);
			6075: out = 16'(359);
			6076: out = 16'(-1792);
			6077: out = 16'(-1348);
			6078: out = 16'(-2486);
			6079: out = 16'(563);
			6080: out = 16'(-786);
			6081: out = 16'(1431);
			6082: out = 16'(-965);
			6083: out = 16'(4397);
			6084: out = 16'(109);
			6085: out = 16'(1616);
			6086: out = 16'(-1786);
			6087: out = 16'(-1495);
			6088: out = 16'(-2099);
			6089: out = 16'(-229);
			6090: out = 16'(847);
			6091: out = 16'(-1);
			6092: out = 16'(4290);
			6093: out = 16'(-1316);
			6094: out = 16'(-32);
			6095: out = 16'(-2400);
			6096: out = 16'(7);
			6097: out = 16'(-186);
			6098: out = 16'(-2109);
			6099: out = 16'(577);
			6100: out = 16'(-782);
			6101: out = 16'(-285);
			6102: out = 16'(1015);
			6103: out = 16'(34);
			6104: out = 16'(-259);
			6105: out = 16'(-787);
			6106: out = 16'(643);
			6107: out = 16'(2652);
			6108: out = 16'(1677);
			6109: out = 16'(-4298);
			6110: out = 16'(-1898);
			6111: out = 16'(-516);
			6112: out = 16'(-1285);
			6113: out = 16'(-514);
			6114: out = 16'(1668);
			6115: out = 16'(-2386);
			6116: out = 16'(34);
			6117: out = 16'(-197);
			6118: out = 16'(2050);
			6119: out = 16'(-1839);
			6120: out = 16'(742);
			6121: out = 16'(-104);
			6122: out = 16'(967);
			6123: out = 16'(2410);
			6124: out = 16'(-1602);
			6125: out = 16'(171);
			6126: out = 16'(-401);
			6127: out = 16'(-1016);
			6128: out = 16'(-4311);
			6129: out = 16'(-1502);
			6130: out = 16'(2575);
			6131: out = 16'(-705);
			6132: out = 16'(3081);
			6133: out = 16'(1561);
			6134: out = 16'(-187);
			6135: out = 16'(-2399);
			6136: out = 16'(975);
			6137: out = 16'(-33);
			6138: out = 16'(-2963);
			6139: out = 16'(-2471);
			6140: out = 16'(1079);
			6141: out = 16'(2801);
			6142: out = 16'(-304);
			6143: out = 16'(2600);
			6144: out = 16'(2313);
			6145: out = 16'(-1660);
			6146: out = 16'(290);
			6147: out = 16'(-838);
			6148: out = 16'(2294);
			6149: out = 16'(-1904);
			6150: out = 16'(271);
			6151: out = 16'(4327);
			6152: out = 16'(-2125);
			6153: out = 16'(75);
			6154: out = 16'(-1808);
			6155: out = 16'(3019);
			6156: out = 16'(-3233);
			6157: out = 16'(-1104);
			6158: out = 16'(628);
			6159: out = 16'(-1723);
			6160: out = 16'(2297);
			6161: out = 16'(126);
			6162: out = 16'(-1270);
			6163: out = 16'(2073);
			6164: out = 16'(-3572);
			6165: out = 16'(1046);
			6166: out = 16'(947);
			6167: out = 16'(-3563);
			6168: out = 16'(570);
			6169: out = 16'(3076);
			6170: out = 16'(888);
			6171: out = 16'(-1776);
			6172: out = 16'(807);
			6173: out = 16'(-4348);
			6174: out = 16'(-957);
			6175: out = 16'(780);
			6176: out = 16'(1654);
			6177: out = 16'(-1135);
			6178: out = 16'(-1930);
			6179: out = 16'(3297);
			6180: out = 16'(189);
			6181: out = 16'(475);
			6182: out = 16'(-422);
			6183: out = 16'(-1158);
			6184: out = 16'(298);
			6185: out = 16'(-40);
			6186: out = 16'(3138);
			6187: out = 16'(-3154);
			6188: out = 16'(-2196);
			6189: out = 16'(-1175);
			6190: out = 16'(2322);
			6191: out = 16'(-1628);
			6192: out = 16'(-257);
			6193: out = 16'(4491);
			6194: out = 16'(-4383);
			6195: out = 16'(2890);
			6196: out = 16'(412);
			6197: out = 16'(-310);
			6198: out = 16'(336);
			6199: out = 16'(-17);
			6200: out = 16'(644);
			6201: out = 16'(-1351);
			6202: out = 16'(43);
			6203: out = 16'(2667);
			6204: out = 16'(201);
			6205: out = 16'(-1500);
			6206: out = 16'(860);
			6207: out = 16'(1288);
			6208: out = 16'(-2434);
			6209: out = 16'(919);
			6210: out = 16'(499);
			6211: out = 16'(-658);
			6212: out = 16'(208);
			6213: out = 16'(-601);
			6214: out = 16'(1492);
			6215: out = 16'(691);
			6216: out = 16'(-1147);
			6217: out = 16'(1503);
			6218: out = 16'(1211);
			6219: out = 16'(-848);
			6220: out = 16'(-2743);
			6221: out = 16'(1646);
			6222: out = 16'(1738);
			6223: out = 16'(-366);
			6224: out = 16'(722);
			6225: out = 16'(265);
			6226: out = 16'(-2714);
			6227: out = 16'(-3824);
			6228: out = 16'(3528);
			6229: out = 16'(-5697);
			6230: out = 16'(352);
			6231: out = 16'(1744);
			6232: out = 16'(-483);
			6233: out = 16'(-622);
			6234: out = 16'(-2314);
			6235: out = 16'(593);
			6236: out = 16'(1318);
			6237: out = 16'(-45);
			6238: out = 16'(-3010);
			6239: out = 16'(1723);
			6240: out = 16'(628);
			6241: out = 16'(1179);
			6242: out = 16'(5561);
			6243: out = 16'(-692);
			6244: out = 16'(-5802);
			6245: out = 16'(2310);
			6246: out = 16'(-852);
			6247: out = 16'(92);
			6248: out = 16'(-2104);
			6249: out = 16'(3140);
			6250: out = 16'(-4159);
			6251: out = 16'(1018);
			6252: out = 16'(1362);
			6253: out = 16'(-2900);
			6254: out = 16'(-459);
			6255: out = 16'(349);
			6256: out = 16'(2141);
			6257: out = 16'(-3306);
			6258: out = 16'(-61);
			6259: out = 16'(855);
			6260: out = 16'(1858);
			6261: out = 16'(-663);
			6262: out = 16'(-2763);
			6263: out = 16'(-962);
			6264: out = 16'(3516);
			6265: out = 16'(-1309);
			6266: out = 16'(1710);
			6267: out = 16'(654);
			6268: out = 16'(35);
			6269: out = 16'(-978);
			6270: out = 16'(458);
			6271: out = 16'(223);
			6272: out = 16'(-7625);
			6273: out = 16'(2174);
			6274: out = 16'(-397);
			6275: out = 16'(818);
			6276: out = 16'(-1087);
			6277: out = 16'(1827);
			6278: out = 16'(-637);
			6279: out = 16'(100);
			6280: out = 16'(2073);
			6281: out = 16'(895);
			6282: out = 16'(-1199);
			6283: out = 16'(-1258);
			6284: out = 16'(-386);
			6285: out = 16'(-2987);
			6286: out = 16'(1659);
			6287: out = 16'(506);
			6288: out = 16'(-719);
			6289: out = 16'(393);
			6290: out = 16'(-147);
			6291: out = 16'(391);
			6292: out = 16'(1350);
			6293: out = 16'(-3517);
			6294: out = 16'(-680);
			6295: out = 16'(-106);
			6296: out = 16'(-1223);
			6297: out = 16'(-1459);
			6298: out = 16'(2142);
			6299: out = 16'(378);
			6300: out = 16'(761);
			6301: out = 16'(1964);
			6302: out = 16'(182);
			6303: out = 16'(-3919);
			6304: out = 16'(-980);
			6305: out = 16'(810);
			6306: out = 16'(1209);
			6307: out = 16'(-504);
			6308: out = 16'(1201);
			6309: out = 16'(964);
			6310: out = 16'(2278);
			6311: out = 16'(-2782);
			6312: out = 16'(-2470);
			6313: out = 16'(316);
			6314: out = 16'(-2262);
			6315: out = 16'(51);
			6316: out = 16'(738);
			6317: out = 16'(-2474);
			6318: out = 16'(809);
			6319: out = 16'(3722);
			6320: out = 16'(2436);
			6321: out = 16'(-5254);
			6322: out = 16'(-830);
			6323: out = 16'(1729);
			6324: out = 16'(-1896);
			6325: out = 16'(2180);
			6326: out = 16'(1794);
			6327: out = 16'(3311);
			6328: out = 16'(-4808);
			6329: out = 16'(-688);
			6330: out = 16'(-2344);
			6331: out = 16'(-627);
			6332: out = 16'(-147);
			6333: out = 16'(-440);
			6334: out = 16'(-462);
			6335: out = 16'(-1513);
			6336: out = 16'(5814);
			6337: out = 16'(974);
			6338: out = 16'(643);
			6339: out = 16'(-290);
			6340: out = 16'(-3034);
			6341: out = 16'(-1391);
			6342: out = 16'(-224);
			6343: out = 16'(181);
			6344: out = 16'(-417);
			6345: out = 16'(-924);
			6346: out = 16'(3535);
			6347: out = 16'(667);
			6348: out = 16'(-443);
			6349: out = 16'(-2208);
			6350: out = 16'(142);
			6351: out = 16'(-541);
			6352: out = 16'(-2350);
			6353: out = 16'(410);
			6354: out = 16'(-2741);
			6355: out = 16'(3375);
			6356: out = 16'(2655);
			6357: out = 16'(354);
			6358: out = 16'(1310);
			6359: out = 16'(-194);
			6360: out = 16'(-726);
			6361: out = 16'(423);
			6362: out = 16'(837);
			6363: out = 16'(1410);
			6364: out = 16'(-228);
			6365: out = 16'(3124);
			6366: out = 16'(-96);
			6367: out = 16'(-3766);
			6368: out = 16'(-2292);
			6369: out = 16'(977);
			6370: out = 16'(-177);
			6371: out = 16'(427);
			6372: out = 16'(948);
			6373: out = 16'(-3235);
			6374: out = 16'(1700);
			6375: out = 16'(-75);
			6376: out = 16'(3655);
			6377: out = 16'(-2460);
			6378: out = 16'(-442);
			6379: out = 16'(359);
			6380: out = 16'(1989);
			6381: out = 16'(2144);
			6382: out = 16'(2230);
			6383: out = 16'(-3080);
			6384: out = 16'(-371);
			6385: out = 16'(1669);
			6386: out = 16'(-208);
			6387: out = 16'(1087);
			6388: out = 16'(-678);
			6389: out = 16'(-1408);
			6390: out = 16'(-18);
			6391: out = 16'(-303);
			6392: out = 16'(-1331);
			6393: out = 16'(-602);
			6394: out = 16'(-2307);
			6395: out = 16'(-253);
			6396: out = 16'(1903);
			6397: out = 16'(-105);
			6398: out = 16'(686);
			6399: out = 16'(3874);
			6400: out = 16'(58);
			6401: out = 16'(1171);
			6402: out = 16'(-254);
			6403: out = 16'(-4252);
			6404: out = 16'(-199);
			6405: out = 16'(1736);
			6406: out = 16'(-1686);
			6407: out = 16'(-2164);
			6408: out = 16'(-1315);
			6409: out = 16'(1109);
			6410: out = 16'(409);
			6411: out = 16'(1856);
			6412: out = 16'(-1183);
			6413: out = 16'(-3650);
			6414: out = 16'(1275);
			6415: out = 16'(-178);
			6416: out = 16'(1094);
			6417: out = 16'(-289);
			6418: out = 16'(-1114);
			6419: out = 16'(1019);
			6420: out = 16'(681);
			6421: out = 16'(161);
			6422: out = 16'(-3147);
			6423: out = 16'(-229);
			6424: out = 16'(1464);
			6425: out = 16'(-261);
			6426: out = 16'(3588);
			6427: out = 16'(-107);
			6428: out = 16'(-1553);
			6429: out = 16'(-1867);
			6430: out = 16'(-2229);
			6431: out = 16'(-2010);
			6432: out = 16'(-1853);
			6433: out = 16'(-99);
			6434: out = 16'(933);
			6435: out = 16'(2424);
			6436: out = 16'(1558);
			6437: out = 16'(3524);
			6438: out = 16'(-1204);
			6439: out = 16'(256);
			6440: out = 16'(-1306);
			6441: out = 16'(935);
			6442: out = 16'(-619);
			6443: out = 16'(833);
			6444: out = 16'(1116);
			6445: out = 16'(-1390);
			6446: out = 16'(-385);
			6447: out = 16'(-69);
			6448: out = 16'(-484);
			6449: out = 16'(-1241);
			6450: out = 16'(855);
			6451: out = 16'(584);
			6452: out = 16'(1388);
			6453: out = 16'(-3420);
			6454: out = 16'(4498);
			6455: out = 16'(-332);
			6456: out = 16'(898);
			6457: out = 16'(453);
			6458: out = 16'(677);
			6459: out = 16'(-1351);
			6460: out = 16'(-1843);
			6461: out = 16'(2355);
			6462: out = 16'(-1192);
			6463: out = 16'(1309);
			6464: out = 16'(-3011);
			6465: out = 16'(1823);
			6466: out = 16'(485);
			6467: out = 16'(56);
			6468: out = 16'(-4104);
			6469: out = 16'(2933);
			6470: out = 16'(-246);
			6471: out = 16'(-711);
			6472: out = 16'(2163);
			6473: out = 16'(1231);
			6474: out = 16'(-4956);
			6475: out = 16'(459);
			6476: out = 16'(2096);
			6477: out = 16'(704);
			6478: out = 16'(798);
			6479: out = 16'(-1107);
			6480: out = 16'(356);
			6481: out = 16'(245);
			6482: out = 16'(3455);
			6483: out = 16'(-715);
			6484: out = 16'(1066);
			6485: out = 16'(-837);
			6486: out = 16'(-73);
			6487: out = 16'(-1275);
			6488: out = 16'(-3375);
			6489: out = 16'(1874);
			6490: out = 16'(260);
			6491: out = 16'(2717);
			6492: out = 16'(-159);
			6493: out = 16'(1264);
			6494: out = 16'(-9);
			6495: out = 16'(-1251);
			6496: out = 16'(3286);
			6497: out = 16'(-2079);
			6498: out = 16'(-1468);
			6499: out = 16'(268);
			6500: out = 16'(1754);
			6501: out = 16'(-91);
			6502: out = 16'(-2675);
			6503: out = 16'(2476);
			6504: out = 16'(-856);
			6505: out = 16'(-1222);
			6506: out = 16'(542);
			6507: out = 16'(-4478);
			6508: out = 16'(443);
			6509: out = 16'(-917);
			6510: out = 16'(1873);
			6511: out = 16'(2090);
			6512: out = 16'(-1849);
			6513: out = 16'(1178);
			6514: out = 16'(3867);
			6515: out = 16'(3999);
			6516: out = 16'(-2548);
			6517: out = 16'(293);
			6518: out = 16'(-241);
			6519: out = 16'(-1456);
			6520: out = 16'(170);
			6521: out = 16'(2595);
			6522: out = 16'(-277);
			6523: out = 16'(-1977);
			6524: out = 16'(-674);
			6525: out = 16'(912);
			6526: out = 16'(354);
			6527: out = 16'(-3638);
			6528: out = 16'(1042);
			6529: out = 16'(-468);
			6530: out = 16'(-2426);
			6531: out = 16'(660);
			6532: out = 16'(695);
			6533: out = 16'(-411);
			6534: out = 16'(-397);
			6535: out = 16'(-942);
			6536: out = 16'(279);
			6537: out = 16'(-1379);
			6538: out = 16'(1612);
			6539: out = 16'(-313);
			6540: out = 16'(322);
			6541: out = 16'(-170);
			6542: out = 16'(2856);
			6543: out = 16'(856);
			6544: out = 16'(255);
			6545: out = 16'(1226);
			6546: out = 16'(-1960);
			6547: out = 16'(550);
			6548: out = 16'(-1652);
			6549: out = 16'(1184);
			6550: out = 16'(-2148);
			6551: out = 16'(1747);
			6552: out = 16'(-1043);
			6553: out = 16'(1560);
			6554: out = 16'(-4050);
			6555: out = 16'(1590);
			6556: out = 16'(370);
			6557: out = 16'(-1111);
			6558: out = 16'(381);
			6559: out = 16'(-413);
			6560: out = 16'(2898);
			6561: out = 16'(51);
			6562: out = 16'(-826);
			6563: out = 16'(-242);
			6564: out = 16'(-1910);
			6565: out = 16'(538);
			6566: out = 16'(229);
			6567: out = 16'(-1497);
			6568: out = 16'(684);
			6569: out = 16'(-1653);
			6570: out = 16'(2224);
			6571: out = 16'(280);
			6572: out = 16'(527);
			6573: out = 16'(-118);
			6574: out = 16'(848);
			6575: out = 16'(40);
			6576: out = 16'(-1713);
			6577: out = 16'(1502);
			6578: out = 16'(-2012);
			6579: out = 16'(-2420);
			6580: out = 16'(0);
			6581: out = 16'(2102);
			6582: out = 16'(-1274);
			6583: out = 16'(294);
			6584: out = 16'(-1884);
			6585: out = 16'(3064);
			6586: out = 16'(-2672);
			6587: out = 16'(154);
			6588: out = 16'(2531);
			6589: out = 16'(205);
			6590: out = 16'(285);
			6591: out = 16'(2724);
			6592: out = 16'(-172);
			6593: out = 16'(-457);
			6594: out = 16'(-2324);
			6595: out = 16'(-79);
			6596: out = 16'(-28);
			6597: out = 16'(-3470);
			6598: out = 16'(3628);
			6599: out = 16'(465);
			6600: out = 16'(2061);
			6601: out = 16'(365);
			6602: out = 16'(917);
			6603: out = 16'(-2744);
			6604: out = 16'(-1883);
			6605: out = 16'(289);
			6606: out = 16'(648);
			6607: out = 16'(-953);
			6608: out = 16'(-1726);
			6609: out = 16'(559);
			6610: out = 16'(913);
			6611: out = 16'(-1590);
			6612: out = 16'(1401);
			6613: out = 16'(-1098);
			6614: out = 16'(1996);
			6615: out = 16'(450);
			6616: out = 16'(1211);
			6617: out = 16'(-309);
			6618: out = 16'(-2064);
			6619: out = 16'(-370);
			6620: out = 16'(690);
			6621: out = 16'(-731);
			6622: out = 16'(-3178);
			6623: out = 16'(-284);
			6624: out = 16'(-1878);
			6625: out = 16'(1805);
			6626: out = 16'(412);
			6627: out = 16'(-357);
			6628: out = 16'(493);
			6629: out = 16'(2059);
			6630: out = 16'(1105);
			6631: out = 16'(-897);
			6632: out = 16'(-707);
			6633: out = 16'(172);
			6634: out = 16'(117);
			6635: out = 16'(-1060);
			6636: out = 16'(-5084);
			6637: out = 16'(-1713);
			6638: out = 16'(-120);
			6639: out = 16'(2013);
			6640: out = 16'(164);
			6641: out = 16'(796);
			6642: out = 16'(510);
			6643: out = 16'(318);
			6644: out = 16'(3278);
			6645: out = 16'(-272);
			6646: out = 16'(-1788);
			6647: out = 16'(164);
			6648: out = 16'(150);
			6649: out = 16'(236);
			6650: out = 16'(-1328);
			6651: out = 16'(-3471);
			6652: out = 16'(3393);
			6653: out = 16'(1640);
			6654: out = 16'(-116);
			6655: out = 16'(8);
			6656: out = 16'(426);
			6657: out = 16'(-2960);
			6658: out = 16'(-761);
			6659: out = 16'(1308);
			6660: out = 16'(-229);
			6661: out = 16'(2650);
			6662: out = 16'(-1264);
			6663: out = 16'(178);
			6664: out = 16'(-5035);
			6665: out = 16'(2632);
			6666: out = 16'(-419);
			6667: out = 16'(1152);
			6668: out = 16'(2468);
			6669: out = 16'(-1543);
			6670: out = 16'(477);
			6671: out = 16'(499);
			6672: out = 16'(1718);
			6673: out = 16'(-2296);
			6674: out = 16'(-1793);
			6675: out = 16'(-3365);
			6676: out = 16'(1768);
			6677: out = 16'(60);
			6678: out = 16'(591);
			6679: out = 16'(1171);
			6680: out = 16'(-486);
			6681: out = 16'(-903);
			6682: out = 16'(2786);
			6683: out = 16'(-1326);
			6684: out = 16'(2348);
			6685: out = 16'(-1966);
			6686: out = 16'(-262);
			6687: out = 16'(-394);
			6688: out = 16'(-808);
			6689: out = 16'(-960);
			6690: out = 16'(2729);
			6691: out = 16'(1125);
			6692: out = 16'(-2374);
			6693: out = 16'(-1131);
			6694: out = 16'(-386);
			6695: out = 16'(601);
			6696: out = 16'(-90);
			6697: out = 16'(-1727);
			6698: out = 16'(2371);
			6699: out = 16'(-74);
			6700: out = 16'(1879);
			6701: out = 16'(1402);
			6702: out = 16'(-306);
			6703: out = 16'(-1163);
			6704: out = 16'(-129);
			6705: out = 16'(3611);
			6706: out = 16'(294);
			6707: out = 16'(-1469);
			6708: out = 16'(12);
			6709: out = 16'(2374);
			6710: out = 16'(-215);
			6711: out = 16'(-309);
			6712: out = 16'(-3512);
			6713: out = 16'(-732);
			6714: out = 16'(-2672);
			6715: out = 16'(1158);
			6716: out = 16'(491);
			6717: out = 16'(3108);
			6718: out = 16'(-1746);
			6719: out = 16'(386);
			6720: out = 16'(-215);
			6721: out = 16'(-1609);
			6722: out = 16'(-3015);
			6723: out = 16'(-1670);
			6724: out = 16'(3403);
			6725: out = 16'(-866);
			6726: out = 16'(424);
			6727: out = 16'(-266);
			6728: out = 16'(2471);
			6729: out = 16'(-2956);
			6730: out = 16'(2804);
			6731: out = 16'(-201);
			6732: out = 16'(-1266);
			6733: out = 16'(526);
			6734: out = 16'(1480);
			6735: out = 16'(1723);
			6736: out = 16'(-4222);
			6737: out = 16'(-761);
			6738: out = 16'(721);
			6739: out = 16'(2689);
			6740: out = 16'(-1456);
			6741: out = 16'(202);
			6742: out = 16'(-3416);
			6743: out = 16'(1864);
			6744: out = 16'(-249);
			6745: out = 16'(195);
			6746: out = 16'(-161);
			6747: out = 16'(-310);
			6748: out = 16'(1281);
			6749: out = 16'(296);
			6750: out = 16'(1754);
			6751: out = 16'(-2429);
			6752: out = 16'(376);
			6753: out = 16'(163);
			6754: out = 16'(438);
			6755: out = 16'(939);
			6756: out = 16'(-174);
			6757: out = 16'(-14);
			6758: out = 16'(3451);
			6759: out = 16'(203);
			6760: out = 16'(1035);
			6761: out = 16'(-3147);
			6762: out = 16'(2530);
			6763: out = 16'(-1245);
			6764: out = 16'(58);
			6765: out = 16'(-1580);
			6766: out = 16'(14);
			6767: out = 16'(-1042);
			6768: out = 16'(-268);
			6769: out = 16'(1996);
			6770: out = 16'(-496);
			6771: out = 16'(221);
			6772: out = 16'(31);
			6773: out = 16'(3097);
			6774: out = 16'(-142);
			6775: out = 16'(1180);
			6776: out = 16'(-386);
			6777: out = 16'(3640);
			6778: out = 16'(-4784);
			6779: out = 16'(-800);
			6780: out = 16'(-1779);
			6781: out = 16'(-1062);
			6782: out = 16'(-171);
			6783: out = 16'(2129);
			6784: out = 16'(582);
			6785: out = 16'(-1171);
			6786: out = 16'(343);
			6787: out = 16'(488);
			6788: out = 16'(-472);
			6789: out = 16'(14);
			6790: out = 16'(126);
			6791: out = 16'(2422);
			6792: out = 16'(-189);
			6793: out = 16'(-97);
			6794: out = 16'(2635);
			6795: out = 16'(-1789);
			6796: out = 16'(-1292);
			6797: out = 16'(390);
			6798: out = 16'(-1644);
			6799: out = 16'(-2605);
			6800: out = 16'(1495);
			6801: out = 16'(2915);
			6802: out = 16'(667);
			6803: out = 16'(-4508);
			6804: out = 16'(2178);
			6805: out = 16'(548);
			6806: out = 16'(-2386);
			6807: out = 16'(3805);
			6808: out = 16'(-274);
			6809: out = 16'(-1150);
			6810: out = 16'(1800);
			6811: out = 16'(4542);
			6812: out = 16'(-1595);
			6813: out = 16'(-3856);
			6814: out = 16'(-1352);
			6815: out = 16'(1787);
			6816: out = 16'(410);
			6817: out = 16'(-747);
			6818: out = 16'(3159);
			6819: out = 16'(-1795);
			6820: out = 16'(-44);
			6821: out = 16'(123);
			6822: out = 16'(675);
			6823: out = 16'(-2641);
			6824: out = 16'(2089);
			6825: out = 16'(1314);
			6826: out = 16'(-39);
			6827: out = 16'(215);
			6828: out = 16'(504);
			6829: out = 16'(1077);
			6830: out = 16'(-1780);
			6831: out = 16'(-316);
			6832: out = 16'(-1377);
			6833: out = 16'(-247);
			6834: out = 16'(473);
			6835: out = 16'(1104);
			6836: out = 16'(569);
			6837: out = 16'(-260);
			6838: out = 16'(-2678);
			6839: out = 16'(1795);
			6840: out = 16'(-221);
			6841: out = 16'(-4681);
			6842: out = 16'(2042);
			6843: out = 16'(-4138);
			6844: out = 16'(3654);
			6845: out = 16'(-989);
			6846: out = 16'(589);
			6847: out = 16'(1805);
			6848: out = 16'(-2493);
			6849: out = 16'(488);
			6850: out = 16'(23);
			6851: out = 16'(-188);
			6852: out = 16'(-3278);
			6853: out = 16'(1963);
			6854: out = 16'(364);
			6855: out = 16'(133);
			6856: out = 16'(1612);
			6857: out = 16'(1858);
			6858: out = 16'(-5052);
			6859: out = 16'(1299);
			6860: out = 16'(-2513);
			6861: out = 16'(722);
			6862: out = 16'(-2232);
			6863: out = 16'(3183);
			6864: out = 16'(1498);
			6865: out = 16'(-57);
			6866: out = 16'(2203);
			6867: out = 16'(51);
			6868: out = 16'(-165);
			6869: out = 16'(-1393);
			6870: out = 16'(909);
			6871: out = 16'(-475);
			6872: out = 16'(-853);
			6873: out = 16'(-1819);
			6874: out = 16'(5028);
			6875: out = 16'(-4296);
			6876: out = 16'(-3322);
			6877: out = 16'(1393);
			6878: out = 16'(-103);
			6879: out = 16'(-955);
			6880: out = 16'(739);
			6881: out = 16'(752);
			6882: out = 16'(2199);
			6883: out = 16'(-1632);
			6884: out = 16'(2112);
			6885: out = 16'(371);
			6886: out = 16'(-3337);
			6887: out = 16'(39);
			6888: out = 16'(3383);
			6889: out = 16'(937);
			6890: out = 16'(-5852);
			6891: out = 16'(1278);
			6892: out = 16'(1309);
			6893: out = 16'(297);
			6894: out = 16'(44);
			6895: out = 16'(553);
			6896: out = 16'(-119);
			6897: out = 16'(-3459);
			6898: out = 16'(436);
			6899: out = 16'(-1618);
			6900: out = 16'(-1693);
			6901: out = 16'(1512);
			6902: out = 16'(390);
			6903: out = 16'(3431);
			6904: out = 16'(-2129);
			6905: out = 16'(1244);
			6906: out = 16'(292);
			6907: out = 16'(849);
			6908: out = 16'(-1367);
			6909: out = 16'(497);
			6910: out = 16'(-992);
			6911: out = 16'(-508);
			6912: out = 16'(3472);
			6913: out = 16'(-5229);
			6914: out = 16'(630);
			6915: out = 16'(843);
			6916: out = 16'(-1203);
			6917: out = 16'(-1811);
			6918: out = 16'(1467);
			6919: out = 16'(-1498);
			6920: out = 16'(1698);
			6921: out = 16'(1326);
			6922: out = 16'(449);
			6923: out = 16'(-2309);
			6924: out = 16'(1321);
			6925: out = 16'(135);
			6926: out = 16'(1703);
			6927: out = 16'(263);
			6928: out = 16'(-2877);
			6929: out = 16'(-422);
			6930: out = 16'(-3025);
			6931: out = 16'(4374);
			6932: out = 16'(-5472);
			6933: out = 16'(4209);
			6934: out = 16'(564);
			6935: out = 16'(-326);
			6936: out = 16'(886);
			6937: out = 16'(-3566);
			6938: out = 16'(-638);
			6939: out = 16'(-1306);
			6940: out = 16'(326);
			6941: out = 16'(647);
			6942: out = 16'(-1770);
			6943: out = 16'(-1420);
			6944: out = 16'(4262);
			6945: out = 16'(2999);
			6946: out = 16'(-791);
			6947: out = 16'(-177);
			6948: out = 16'(-355);
			6949: out = 16'(-3939);
			6950: out = 16'(4222);
			6951: out = 16'(-2274);
			6952: out = 16'(137);
			6953: out = 16'(-3185);
			6954: out = 16'(1497);
			6955: out = 16'(-4288);
			6956: out = 16'(30);
			6957: out = 16'(1312);
			6958: out = 16'(556);
			6959: out = 16'(-473);
			6960: out = 16'(453);
			6961: out = 16'(2643);
			6962: out = 16'(-3694);
			6963: out = 16'(-497);
			6964: out = 16'(3596);
			6965: out = 16'(-3017);
			6966: out = 16'(-599);
			6967: out = 16'(142);
			6968: out = 16'(1028);
			6969: out = 16'(-329);
			6970: out = 16'(-652);
			6971: out = 16'(1256);
			6972: out = 16'(-2408);
			6973: out = 16'(2538);
			6974: out = 16'(598);
			6975: out = 16'(2035);
			6976: out = 16'(-3079);
			6977: out = 16'(1823);
			6978: out = 16'(-876);
			6979: out = 16'(478);
			6980: out = 16'(-241);
			6981: out = 16'(-1650);
			6982: out = 16'(2245);
			6983: out = 16'(83);
			6984: out = 16'(-50);
			6985: out = 16'(2090);
			6986: out = 16'(-43);
			6987: out = 16'(-576);
			6988: out = 16'(1001);
			6989: out = 16'(894);
			6990: out = 16'(-2197);
			6991: out = 16'(-2300);
			6992: out = 16'(3600);
			6993: out = 16'(-3409);
			6994: out = 16'(372);
			6995: out = 16'(1769);
			6996: out = 16'(-847);
			6997: out = 16'(-20);
			6998: out = 16'(-1411);
			6999: out = 16'(1965);
			7000: out = 16'(-3345);
			7001: out = 16'(334);
			7002: out = 16'(474);
			7003: out = 16'(1461);
			7004: out = 16'(-2438);
			7005: out = 16'(-1255);
			7006: out = 16'(2677);
			7007: out = 16'(372);
			7008: out = 16'(-2586);
			7009: out = 16'(1271);
			7010: out = 16'(1749);
			7011: out = 16'(-4240);
			7012: out = 16'(512);
			7013: out = 16'(3466);
			7014: out = 16'(-2542);
			7015: out = 16'(-4831);
			7016: out = 16'(621);
			7017: out = 16'(403);
			7018: out = 16'(-1215);
			7019: out = 16'(246);
			7020: out = 16'(33);
			7021: out = 16'(-967);
			7022: out = 16'(308);
			7023: out = 16'(418);
			7024: out = 16'(857);
			7025: out = 16'(-702);
			7026: out = 16'(-59);
			7027: out = 16'(1377);
			7028: out = 16'(-1148);
			7029: out = 16'(-982);
			7030: out = 16'(-345);
			7031: out = 16'(603);
			7032: out = 16'(491);
			7033: out = 16'(-4959);
			7034: out = 16'(1710);
			7035: out = 16'(-850);
			7036: out = 16'(568);
			7037: out = 16'(-992);
			7038: out = 16'(3034);
			7039: out = 16'(-4909);
			7040: out = 16'(1898);
			7041: out = 16'(3084);
			7042: out = 16'(0);
			7043: out = 16'(-1145);
			7044: out = 16'(624);
			7045: out = 16'(1731);
			7046: out = 16'(-989);
			7047: out = 16'(-762);
			7048: out = 16'(-1392);
			7049: out = 16'(61);
			7050: out = 16'(-680);
			7051: out = 16'(4426);
			7052: out = 16'(-482);
			7053: out = 16'(-709);
			7054: out = 16'(-71);
			7055: out = 16'(1843);
			7056: out = 16'(-1141);
			7057: out = 16'(-216);
			7058: out = 16'(-1089);
			7059: out = 16'(-271);
			7060: out = 16'(-84);
			7061: out = 16'(1678);
			7062: out = 16'(-375);
			7063: out = 16'(-3412);
			7064: out = 16'(-399);
			7065: out = 16'(-290);
			7066: out = 16'(1354);
			7067: out = 16'(-3891);
			7068: out = 16'(1545);
			7069: out = 16'(1803);
			7070: out = 16'(-37);
			7071: out = 16'(-503);
			7072: out = 16'(2700);
			7073: out = 16'(-2229);
			7074: out = 16'(-2392);
			7075: out = 16'(1104);
			7076: out = 16'(-863);
			7077: out = 16'(-2188);
			7078: out = 16'(74);
			7079: out = 16'(2004);
			7080: out = 16'(5225);
			7081: out = 16'(-476);
			7082: out = 16'(-1433);
			7083: out = 16'(1281);
			7084: out = 16'(303);
			7085: out = 16'(-4130);
			7086: out = 16'(494);
			7087: out = 16'(480);
			7088: out = 16'(-5457);
			7089: out = 16'(928);
			7090: out = 16'(3971);
			7091: out = 16'(3965);
			7092: out = 16'(-5558);
			7093: out = 16'(3483);
			7094: out = 16'(-460);
			7095: out = 16'(-3736);
			7096: out = 16'(333);
			7097: out = 16'(1233);
			7098: out = 16'(1343);
			7099: out = 16'(-1029);
			7100: out = 16'(-300);
			7101: out = 16'(1671);
			7102: out = 16'(-4059);
			7103: out = 16'(-306);
			7104: out = 16'(321);
			7105: out = 16'(-385);
			7106: out = 16'(556);
			7107: out = 16'(1153);
			7108: out = 16'(3467);
			7109: out = 16'(-1017);
			7110: out = 16'(1730);
			7111: out = 16'(-2978);
			7112: out = 16'(538);
			7113: out = 16'(-109);
			7114: out = 16'(861);
			7115: out = 16'(234);
			7116: out = 16'(112);
			7117: out = 16'(1104);
			7118: out = 16'(-1005);
			7119: out = 16'(-900);
			7120: out = 16'(168);
			7121: out = 16'(1601);
			7122: out = 16'(-4355);
			7123: out = 16'(1707);
			7124: out = 16'(-1858);
			7125: out = 16'(423);
			7126: out = 16'(176);
			7127: out = 16'(810);
			7128: out = 16'(1199);
			7129: out = 16'(110);
			7130: out = 16'(-1538);
			7131: out = 16'(2175);
			7132: out = 16'(-3539);
			7133: out = 16'(271);
			7134: out = 16'(-207);
			7135: out = 16'(-79);
			7136: out = 16'(1860);
			7137: out = 16'(-477);
			7138: out = 16'(-528);
			7139: out = 16'(-796);
			7140: out = 16'(3206);
			7141: out = 16'(-2401);
			7142: out = 16'(2673);
			7143: out = 16'(-539);
			7144: out = 16'(-4302);
			7145: out = 16'(2919);
			7146: out = 16'(132);
			7147: out = 16'(-160);
			7148: out = 16'(-345);
			7149: out = 16'(-517);
			7150: out = 16'(2339);
			7151: out = 16'(-1591);
			7152: out = 16'(636);
			7153: out = 16'(370);
			7154: out = 16'(-155);
			7155: out = 16'(-3267);
			7156: out = 16'(3521);
			7157: out = 16'(-1658);
			7158: out = 16'(-2690);
			7159: out = 16'(3399);
			7160: out = 16'(1772);
			7161: out = 16'(497);
			7162: out = 16'(-588);
			7163: out = 16'(1636);
			7164: out = 16'(-1851);
			7165: out = 16'(-1343);
			7166: out = 16'(2729);
			7167: out = 16'(429);
			7168: out = 16'(-2664);
			7169: out = 16'(1278);
			7170: out = 16'(3655);
			7171: out = 16'(165);
			7172: out = 16'(-3148);
			7173: out = 16'(184);
			7174: out = 16'(-2030);
			7175: out = 16'(1355);
			7176: out = 16'(-696);
			7177: out = 16'(-138);
			7178: out = 16'(-143);
			7179: out = 16'(-1992);
			7180: out = 16'(1623);
			7181: out = 16'(-208);
			7182: out = 16'(-1664);
			7183: out = 16'(-113);
			7184: out = 16'(52);
			7185: out = 16'(1260);
			7186: out = 16'(1051);
			7187: out = 16'(-949);
			7188: out = 16'(485);
			7189: out = 16'(952);
			7190: out = 16'(560);
			7191: out = 16'(489);
			7192: out = 16'(-387);
			7193: out = 16'(-1468);
			7194: out = 16'(-216);
			7195: out = 16'(-1754);
			7196: out = 16'(147);
			7197: out = 16'(652);
			7198: out = 16'(-959);
			7199: out = 16'(1749);
			7200: out = 16'(126);
			7201: out = 16'(2013);
			7202: out = 16'(-204);
			7203: out = 16'(715);
			7204: out = 16'(-202);
			7205: out = 16'(-1043);
			7206: out = 16'(-817);
			7207: out = 16'(1754);
			7208: out = 16'(1742);
			7209: out = 16'(-2601);
			7210: out = 16'(332);
			7211: out = 16'(1214);
			7212: out = 16'(479);
			7213: out = 16'(-14);
			7214: out = 16'(-324);
			7215: out = 16'(1144);
			7216: out = 16'(-518);
			7217: out = 16'(1503);
			7218: out = 16'(-36);
			7219: out = 16'(-644);
			7220: out = 16'(-2168);
			7221: out = 16'(784);
			7222: out = 16'(145);
			7223: out = 16'(-1524);
			7224: out = 16'(703);
			7225: out = 16'(188);
			7226: out = 16'(2789);
			7227: out = 16'(-402);
			7228: out = 16'(160);
			7229: out = 16'(-2048);
			7230: out = 16'(-33);
			7231: out = 16'(-331);
			7232: out = 16'(1229);
			7233: out = 16'(-3912);
			7234: out = 16'(1073);
			7235: out = 16'(-431);
			7236: out = 16'(2230);
			7237: out = 16'(2477);
			7238: out = 16'(-3658);
			7239: out = 16'(-596);
			7240: out = 16'(1301);
			7241: out = 16'(1599);
			7242: out = 16'(-1853);
			7243: out = 16'(1927);
			7244: out = 16'(263);
			7245: out = 16'(92);
			7246: out = 16'(-317);
			7247: out = 16'(935);
			7248: out = 16'(-2679);
			7249: out = 16'(-1283);
			7250: out = 16'(-97);
			7251: out = 16'(400);
			7252: out = 16'(-2751);
			7253: out = 16'(911);
			7254: out = 16'(-145);
			7255: out = 16'(-232);
			7256: out = 16'(402);
			7257: out = 16'(-129);
			7258: out = 16'(577);
			7259: out = 16'(-1276);
			7260: out = 16'(1982);
			7261: out = 16'(-206);
			7262: out = 16'(-2241);
			7263: out = 16'(609);
			7264: out = 16'(63);
			7265: out = 16'(-2474);
			7266: out = 16'(1812);
			7267: out = 16'(1159);
			7268: out = 16'(217);
			7269: out = 16'(-1459);
			7270: out = 16'(1886);
			7271: out = 16'(-192);
			7272: out = 16'(-1248);
			7273: out = 16'(-232);
			7274: out = 16'(1869);
			7275: out = 16'(1335);
			7276: out = 16'(304);
			7277: out = 16'(1243);
			7278: out = 16'(387);
			7279: out = 16'(-1500);
			7280: out = 16'(-599);
			7281: out = 16'(2301);
			7282: out = 16'(-2186);
			7283: out = 16'(-3238);
			7284: out = 16'(-671);
			7285: out = 16'(3950);
			7286: out = 16'(2215);
			7287: out = 16'(-1789);
			7288: out = 16'(-2034);
			7289: out = 16'(-1668);
			7290: out = 16'(-1030);
			7291: out = 16'(1618);
			7292: out = 16'(833);
			7293: out = 16'(3038);
			7294: out = 16'(-688);
			7295: out = 16'(253);
			7296: out = 16'(2245);
			7297: out = 16'(-1265);
			7298: out = 16'(-4984);
			7299: out = 16'(255);
			7300: out = 16'(1852);
			7301: out = 16'(-3429);
			7302: out = 16'(1457);
			7303: out = 16'(358);
			7304: out = 16'(959);
			7305: out = 16'(-3791);
			7306: out = 16'(1623);
			7307: out = 16'(-1622);
			7308: out = 16'(229);
			7309: out = 16'(146);
			7310: out = 16'(1330);
			7311: out = 16'(1006);
			7312: out = 16'(-2723);
			7313: out = 16'(774);
			7314: out = 16'(-2018);
			7315: out = 16'(3643);
			7316: out = 16'(-3078);
			7317: out = 16'(1088);
			7318: out = 16'(1306);
			7319: out = 16'(101);
			7320: out = 16'(-221);
			7321: out = 16'(-125);
			7322: out = 16'(-857);
			7323: out = 16'(-645);
			7324: out = 16'(-569);
			7325: out = 16'(-569);
			7326: out = 16'(-15);
			7327: out = 16'(254);
			7328: out = 16'(1728);
			7329: out = 16'(368);
			7330: out = 16'(-329);
			7331: out = 16'(2293);
			7332: out = 16'(-535);
			7333: out = 16'(-1281);
			7334: out = 16'(1263);
			7335: out = 16'(368);
			7336: out = 16'(-1771);
			7337: out = 16'(1821);
			7338: out = 16'(-2769);
			7339: out = 16'(-2333);
			7340: out = 16'(-289);
			7341: out = 16'(-1331);
			7342: out = 16'(244);
			7343: out = 16'(1184);
			7344: out = 16'(-1663);
			7345: out = 16'(1226);
			7346: out = 16'(2078);
			7347: out = 16'(-705);
			7348: out = 16'(-1059);
			7349: out = 16'(-1753);
			7350: out = 16'(382);
			7351: out = 16'(-1926);
			7352: out = 16'(2133);
			7353: out = 16'(590);
			7354: out = 16'(536);
			7355: out = 16'(400);
			7356: out = 16'(274);
			7357: out = 16'(-215);
			7358: out = 16'(972);
			7359: out = 16'(-419);
			7360: out = 16'(-966);
			7361: out = 16'(1861);
			7362: out = 16'(-2373);
			7363: out = 16'(-1601);
			7364: out = 16'(332);
			7365: out = 16'(2808);
			7366: out = 16'(-4755);
			7367: out = 16'(478);
			7368: out = 16'(-2687);
			7369: out = 16'(745);
			7370: out = 16'(602);
			7371: out = 16'(1055);
			7372: out = 16'(-206);
			7373: out = 16'(266);
			7374: out = 16'(-258);
			7375: out = 16'(-1633);
			7376: out = 16'(925);
			7377: out = 16'(549);
			7378: out = 16'(-676);
			7379: out = 16'(77);
			7380: out = 16'(3484);
			7381: out = 16'(-2887);
			7382: out = 16'(-2377);
			7383: out = 16'(507);
			7384: out = 16'(2888);
			7385: out = 16'(-974);
			7386: out = 16'(380);
			7387: out = 16'(3174);
			7388: out = 16'(-2149);
			7389: out = 16'(237);
			7390: out = 16'(971);
			7391: out = 16'(-1094);
			7392: out = 16'(-39);
			7393: out = 16'(-2859);
			7394: out = 16'(3615);
			7395: out = 16'(571);
			7396: out = 16'(-1194);
			7397: out = 16'(2270);
			7398: out = 16'(-652);
			7399: out = 16'(-499);
			7400: out = 16'(-4234);
			7401: out = 16'(534);
			7402: out = 16'(1769);
			7403: out = 16'(-1464);
			7404: out = 16'(-539);
			7405: out = 16'(1089);
			7406: out = 16'(-689);
			7407: out = 16'(-1877);
			7408: out = 16'(-1398);
			7409: out = 16'(601);
			7410: out = 16'(-1208);
			7411: out = 16'(1140);
			7412: out = 16'(-803);
			7413: out = 16'(1785);
			7414: out = 16'(-1064);
			7415: out = 16'(-62);
			7416: out = 16'(1182);
			7417: out = 16'(-2966);
			7418: out = 16'(-774);
			7419: out = 16'(-917);
			7420: out = 16'(2824);
			7421: out = 16'(-1516);
			7422: out = 16'(1667);
			7423: out = 16'(-1518);
			7424: out = 16'(48);
			7425: out = 16'(-2065);
			7426: out = 16'(271);
			7427: out = 16'(1083);
			7428: out = 16'(-2549);
			7429: out = 16'(3032);
			7430: out = 16'(101);
			7431: out = 16'(-618);
			7432: out = 16'(2040);
			7433: out = 16'(-1005);
			7434: out = 16'(-430);
			7435: out = 16'(773);
			7436: out = 16'(-218);
			7437: out = 16'(286);
			7438: out = 16'(-636);
			7439: out = 16'(1763);
			7440: out = 16'(-1684);
			7441: out = 16'(-67);
			7442: out = 16'(466);
			7443: out = 16'(2088);
			7444: out = 16'(-1834);
			7445: out = 16'(-525);
			7446: out = 16'(1050);
			7447: out = 16'(159);
			7448: out = 16'(-353);
			7449: out = 16'(176);
			7450: out = 16'(51);
			7451: out = 16'(-56);
			7452: out = 16'(-1005);
			7453: out = 16'(811);
			7454: out = 16'(322);
			7455: out = 16'(-2950);
			7456: out = 16'(752);
			7457: out = 16'(726);
			7458: out = 16'(-1457);
			7459: out = 16'(428);
			7460: out = 16'(1261);
			7461: out = 16'(-390);
			7462: out = 16'(2585);
			7463: out = 16'(-3227);
			7464: out = 16'(258);
			7465: out = 16'(-1260);
			7466: out = 16'(-1188);
			7467: out = 16'(-1263);
			7468: out = 16'(364);
			7469: out = 16'(-1570);
			7470: out = 16'(317);
			7471: out = 16'(2435);
			7472: out = 16'(1734);
			7473: out = 16'(-1745);
			7474: out = 16'(1216);
			7475: out = 16'(-351);
			7476: out = 16'(321);
			7477: out = 16'(-714);
			7478: out = 16'(-1647);
			7479: out = 16'(2099);
			7480: out = 16'(-440);
			7481: out = 16'(2733);
			7482: out = 16'(-1202);
			7483: out = 16'(-411);
			7484: out = 16'(-2780);
			7485: out = 16'(-293);
			7486: out = 16'(651);
			7487: out = 16'(-757);
			7488: out = 16'(-835);
			7489: out = 16'(-135);
			7490: out = 16'(2096);
			7491: out = 16'(244);
			7492: out = 16'(-812);
			7493: out = 16'(-132);
			7494: out = 16'(2533);
			7495: out = 16'(-1244);
			7496: out = 16'(2980);
			7497: out = 16'(40);
			7498: out = 16'(-302);
			7499: out = 16'(370);
			7500: out = 16'(170);
			7501: out = 16'(-2337);
			7502: out = 16'(-1120);
			7503: out = 16'(1363);
			7504: out = 16'(-9);
			7505: out = 16'(1893);
			7506: out = 16'(-112);
			7507: out = 16'(313);
			7508: out = 16'(269);
			7509: out = 16'(1196);
			7510: out = 16'(106);
			7511: out = 16'(-445);
			7512: out = 16'(512);
			7513: out = 16'(-1041);
			7514: out = 16'(-1016);
			7515: out = 16'(2200);
			7516: out = 16'(-254);
			7517: out = 16'(-1365);
			7518: out = 16'(8);
			7519: out = 16'(-417);
			7520: out = 16'(759);
			7521: out = 16'(1610);
			7522: out = 16'(633);
			7523: out = 16'(-463);
			7524: out = 16'(-20);
			7525: out = 16'(-1804);
			7526: out = 16'(-75);
			7527: out = 16'(-141);
			7528: out = 16'(-4313);
			7529: out = 16'(2455);
			7530: out = 16'(344);
			7531: out = 16'(-1070);
			7532: out = 16'(1238);
			7533: out = 16'(2816);
			7534: out = 16'(49);
			7535: out = 16'(-1425);
			7536: out = 16'(1246);
			7537: out = 16'(251);
			7538: out = 16'(-2347);
			7539: out = 16'(381);
			7540: out = 16'(1764);
			7541: out = 16'(-537);
			7542: out = 16'(77);
			7543: out = 16'(-300);
			7544: out = 16'(1183);
			7545: out = 16'(-2513);
			7546: out = 16'(775);
			7547: out = 16'(234);
			7548: out = 16'(2004);
			7549: out = 16'(477);
			7550: out = 16'(365);
			7551: out = 16'(104);
			7552: out = 16'(372);
			7553: out = 16'(-116);
			7554: out = 16'(-1472);
			7555: out = 16'(-392);
			7556: out = 16'(185);
			7557: out = 16'(896);
			7558: out = 16'(-896);
			7559: out = 16'(3150);
			7560: out = 16'(-2181);
			7561: out = 16'(1710);
			7562: out = 16'(-21);
			7563: out = 16'(-1677);
			7564: out = 16'(675);
			7565: out = 16'(38);
			7566: out = 16'(-2198);
			7567: out = 16'(1837);
			7568: out = 16'(-875);
			7569: out = 16'(-1349);
			7570: out = 16'(730);
			7571: out = 16'(2099);
			7572: out = 16'(-408);
			7573: out = 16'(1303);
			7574: out = 16'(658);
			7575: out = 16'(-1879);
			7576: out = 16'(127);
			7577: out = 16'(-373);
			7578: out = 16'(981);
			7579: out = 16'(-750);
			7580: out = 16'(-1692);
			7581: out = 16'(-278);
			7582: out = 16'(3085);
			7583: out = 16'(348);
			7584: out = 16'(-1800);
			7585: out = 16'(-254);
			7586: out = 16'(777);
			7587: out = 16'(-1554);
			7588: out = 16'(-1636);
			7589: out = 16'(4030);
			7590: out = 16'(-414);
			7591: out = 16'(-186);
			7592: out = 16'(3974);
			7593: out = 16'(-245);
			7594: out = 16'(-2004);
			7595: out = 16'(-1650);
			7596: out = 16'(1178);
			7597: out = 16'(-127);
			7598: out = 16'(-3252);
			7599: out = 16'(2392);
			7600: out = 16'(-15);
			7601: out = 16'(-173);
			7602: out = 16'(-1123);
			7603: out = 16'(-1015);
			7604: out = 16'(-531);
			7605: out = 16'(-3444);
			7606: out = 16'(2798);
			7607: out = 16'(-66);
			7608: out = 16'(1097);
			7609: out = 16'(-140);
			7610: out = 16'(2040);
			7611: out = 16'(1934);
			7612: out = 16'(-2459);
			7613: out = 16'(-1798);
			7614: out = 16'(2735);
			7615: out = 16'(-1239);
			7616: out = 16'(1680);
			7617: out = 16'(-173);
			7618: out = 16'(231);
			7619: out = 16'(-229);
			7620: out = 16'(859);
			7621: out = 16'(-472);
			7622: out = 16'(-4235);
			7623: out = 16'(-48);
			7624: out = 16'(589);
			7625: out = 16'(904);
			7626: out = 16'(1766);
			7627: out = 16'(2151);
			7628: out = 16'(-1056);
			7629: out = 16'(2746);
			7630: out = 16'(-3124);
			7631: out = 16'(-1420);
			7632: out = 16'(-25);
			7633: out = 16'(-1838);
			7634: out = 16'(1874);
			7635: out = 16'(-634);
			7636: out = 16'(329);
			7637: out = 16'(516);
			7638: out = 16'(1623);
			7639: out = 16'(47);
			7640: out = 16'(-4317);
			7641: out = 16'(812);
			7642: out = 16'(-2755);
			7643: out = 16'(1908);
			7644: out = 16'(1250);
			7645: out = 16'(-836);
			7646: out = 16'(-647);
			7647: out = 16'(-294);
			7648: out = 16'(1800);
			7649: out = 16'(787);
			7650: out = 16'(-3208);
			7651: out = 16'(1927);
			7652: out = 16'(228);
			7653: out = 16'(994);
			7654: out = 16'(-294);
			7655: out = 16'(-731);
			7656: out = 16'(-271);
			7657: out = 16'(262);
			7658: out = 16'(-528);
			7659: out = 16'(-934);
			7660: out = 16'(923);
			7661: out = 16'(-966);
			7662: out = 16'(2637);
			7663: out = 16'(-30);
			7664: out = 16'(-706);
			7665: out = 16'(-525);
			7666: out = 16'(36);
			7667: out = 16'(899);
			7668: out = 16'(24);
			7669: out = 16'(2729);
			7670: out = 16'(-747);
			7671: out = 16'(-839);
			7672: out = 16'(-121);
			7673: out = 16'(397);
			7674: out = 16'(-166);
			7675: out = 16'(-1429);
			7676: out = 16'(2593);
			7677: out = 16'(233);
			7678: out = 16'(-241);
			7679: out = 16'(-1033);
			7680: out = 16'(-337);
			7681: out = 16'(-251);
			7682: out = 16'(-2136);
			7683: out = 16'(468);
			7684: out = 16'(-243);
			7685: out = 16'(-1572);
			7686: out = 16'(3189);
			7687: out = 16'(-86);
			7688: out = 16'(1838);
			7689: out = 16'(-1271);
			7690: out = 16'(-15);
			7691: out = 16'(-2082);
			7692: out = 16'(497);
			7693: out = 16'(829);
			7694: out = 16'(7);
			7695: out = 16'(6);
			7696: out = 16'(758);
			7697: out = 16'(1104);
			7698: out = 16'(104);
			7699: out = 16'(715);
			7700: out = 16'(-1104);
			7701: out = 16'(-309);
			7702: out = 16'(-73);
			7703: out = 16'(15);
			7704: out = 16'(-1191);
			7705: out = 16'(658);
			7706: out = 16'(473);
			7707: out = 16'(792);
			7708: out = 16'(-422);
			7709: out = 16'(-194);
			7710: out = 16'(261);
			7711: out = 16'(1611);
			7712: out = 16'(1125);
			7713: out = 16'(78);
			7714: out = 16'(-3120);
			7715: out = 16'(-634);
			7716: out = 16'(2137);
			7717: out = 16'(-2124);
			7718: out = 16'(286);
			7719: out = 16'(749);
			7720: out = 16'(-3972);
			7721: out = 16'(3137);
			7722: out = 16'(-1423);
			7723: out = 16'(-1096);
			7724: out = 16'(564);
			7725: out = 16'(1614);
			7726: out = 16'(505);
			7727: out = 16'(-496);
			7728: out = 16'(1106);
			7729: out = 16'(-21);
			7730: out = 16'(401);
			7731: out = 16'(343);
			7732: out = 16'(-103);
			7733: out = 16'(-2640);
			7734: out = 16'(-1276);
			7735: out = 16'(3495);
			7736: out = 16'(347);
			7737: out = 16'(-1127);
			7738: out = 16'(161);
			7739: out = 16'(1556);
			7740: out = 16'(190);
			7741: out = 16'(-3206);
			7742: out = 16'(1314);
			7743: out = 16'(-113);
			7744: out = 16'(138);
			7745: out = 16'(742);
			7746: out = 16'(1607);
			7747: out = 16'(-4312);
			7748: out = 16'(529);
			7749: out = 16'(1240);
			7750: out = 16'(-743);
			7751: out = 16'(359);
			7752: out = 16'(-1575);
			7753: out = 16'(198);
			7754: out = 16'(2912);
			7755: out = 16'(-368);
			7756: out = 16'(-2294);
			7757: out = 16'(-69);
			7758: out = 16'(-2135);
			7759: out = 16'(329);
			7760: out = 16'(-283);
			7761: out = 16'(574);
			7762: out = 16'(481);
			7763: out = 16'(-173);
			7764: out = 16'(-118);
			7765: out = 16'(-793);
			7766: out = 16'(337);
			7767: out = 16'(-78);
			7768: out = 16'(2458);
			7769: out = 16'(-1854);
			7770: out = 16'(888);
			7771: out = 16'(-879);
			7772: out = 16'(779);
			7773: out = 16'(187);
			7774: out = 16'(-902);
			7775: out = 16'(-298);
			7776: out = 16'(-25);
			7777: out = 16'(2220);
			7778: out = 16'(-941);
			7779: out = 16'(-251);
			7780: out = 16'(-788);
			7781: out = 16'(-389);
			7782: out = 16'(-2710);
			7783: out = 16'(-87);
			7784: out = 16'(1404);
			7785: out = 16'(-1551);
			7786: out = 16'(519);
			7787: out = 16'(2734);
			7788: out = 16'(-270);
			7789: out = 16'(1412);
			7790: out = 16'(-4232);
			7791: out = 16'(451);
			7792: out = 16'(-545);
			7793: out = 16'(-2318);
			7794: out = 16'(2805);
			7795: out = 16'(2588);
			7796: out = 16'(-1071);
			7797: out = 16'(-1703);
			7798: out = 16'(2623);
			7799: out = 16'(-3165);
			7800: out = 16'(-1107);
			7801: out = 16'(-297);
			7802: out = 16'(974);
			7803: out = 16'(196);
			7804: out = 16'(623);
			7805: out = 16'(-214);
			7806: out = 16'(560);
			7807: out = 16'(-961);
			7808: out = 16'(-30);
			7809: out = 16'(-1338);
			7810: out = 16'(619);
			7811: out = 16'(196);
			7812: out = 16'(2552);
			7813: out = 16'(3503);
			7814: out = 16'(-4118);
			7815: out = 16'(42);
			7816: out = 16'(2207);
			7817: out = 16'(-607);
			7818: out = 16'(-2805);
			7819: out = 16'(678);
			7820: out = 16'(250);
			7821: out = 16'(-1313);
			7822: out = 16'(3641);
			7823: out = 16'(-296);
			7824: out = 16'(-1747);
			7825: out = 16'(-450);
			7826: out = 16'(1840);
			7827: out = 16'(239);
			7828: out = 16'(-3099);
			7829: out = 16'(1363);
			7830: out = 16'(336);
			7831: out = 16'(196);
			7832: out = 16'(2346);
			7833: out = 16'(-228);
			7834: out = 16'(-3257);
			7835: out = 16'(-302);
			7836: out = 16'(1648);
			7837: out = 16'(-2293);
			7838: out = 16'(-2186);
			7839: out = 16'(1330);
			7840: out = 16'(5);
			7841: out = 16'(1610);
			7842: out = 16'(-688);
			7843: out = 16'(665);
			7844: out = 16'(321);
			7845: out = 16'(1070);
			7846: out = 16'(477);
			7847: out = 16'(346);
			7848: out = 16'(-590);
			7849: out = 16'(-1143);
			7850: out = 16'(2371);
			7851: out = 16'(121);
			7852: out = 16'(-1560);
			7853: out = 16'(864);
			7854: out = 16'(-14);
			7855: out = 16'(690);
			7856: out = 16'(-1700);
			7857: out = 16'(-542);
			7858: out = 16'(-2204);
			7859: out = 16'(-1054);
			7860: out = 16'(584);
			7861: out = 16'(-95);
			7862: out = 16'(3406);
			7863: out = 16'(-3);
			7864: out = 16'(-68);
			7865: out = 16'(-173);
			7866: out = 16'(-2377);
			7867: out = 16'(-2356);
			7868: out = 16'(991);
			7869: out = 16'(2307);
			7870: out = 16'(-2175);
			7871: out = 16'(3494);
			7872: out = 16'(466);
			7873: out = 16'(-91);
			7874: out = 16'(-399);
			7875: out = 16'(1470);
			7876: out = 16'(-3606);
			7877: out = 16'(-4776);
			7878: out = 16'(3013);
			7879: out = 16'(-172);
			7880: out = 16'(1013);
			7881: out = 16'(-51);
			7882: out = 16'(1958);
			7883: out = 16'(-857);
			7884: out = 16'(-3554);
			7885: out = 16'(300);
			7886: out = 16'(52);
			7887: out = 16'(-1276);
			7888: out = 16'(2316);
			7889: out = 16'(1020);
			7890: out = 16'(1386);
			7891: out = 16'(-1568);
			7892: out = 16'(-36);
			7893: out = 16'(27);
			7894: out = 16'(-1772);
			7895: out = 16'(90);
			7896: out = 16'(-509);
			7897: out = 16'(1233);
			7898: out = 16'(-734);
			7899: out = 16'(1978);
			7900: out = 16'(382);
			7901: out = 16'(-2780);
			7902: out = 16'(-388);
			7903: out = 16'(664);
			7904: out = 16'(300);
			7905: out = 16'(-303);
			7906: out = 16'(-151);
			7907: out = 16'(2501);
			7908: out = 16'(-871);
			7909: out = 16'(-1791);
			7910: out = 16'(-1360);
			7911: out = 16'(1957);
			7912: out = 16'(178);
			7913: out = 16'(1215);
			7914: out = 16'(-142);
			7915: out = 16'(-1502);
			7916: out = 16'(320);
			7917: out = 16'(223);
			7918: out = 16'(1757);
			7919: out = 16'(-3461);
			7920: out = 16'(-660);
			7921: out = 16'(1255);
			7922: out = 16'(748);
			7923: out = 16'(800);
			7924: out = 16'(-866);
			7925: out = 16'(337);
			7926: out = 16'(577);
			7927: out = 16'(2845);
			7928: out = 16'(-2917);
			7929: out = 16'(-1287);
			7930: out = 16'(969);
			7931: out = 16'(424);
			7932: out = 16'(1761);
			7933: out = 16'(236);
			7934: out = 16'(-259);
			7935: out = 16'(-819);
			7936: out = 16'(269);
			7937: out = 16'(644);
			7938: out = 16'(-4358);
			7939: out = 16'(-3293);
			7940: out = 16'(1978);
			7941: out = 16'(3097);
			7942: out = 16'(-1498);
			7943: out = 16'(-700);
			7944: out = 16'(390);
			7945: out = 16'(688);
			7946: out = 16'(-20);
			7947: out = 16'(-333);
			7948: out = 16'(-116);
			7949: out = 16'(1281);
			7950: out = 16'(-2538);
			7951: out = 16'(1893);
			7952: out = 16'(632);
			7953: out = 16'(-3589);
			7954: out = 16'(-484);
			7955: out = 16'(923);
			7956: out = 16'(-124);
			7957: out = 16'(320);
			7958: out = 16'(607);
			7959: out = 16'(-674);
			7960: out = 16'(1225);
			7961: out = 16'(248);
			7962: out = 16'(1579);
			7963: out = 16'(-141);
			7964: out = 16'(-2236);
			7965: out = 16'(67);
			7966: out = 16'(2114);
			7967: out = 16'(231);
			7968: out = 16'(-1464);
			7969: out = 16'(357);
			7970: out = 16'(1097);
			7971: out = 16'(320);
			7972: out = 16'(-231);
			7973: out = 16'(454);
			7974: out = 16'(-1372);
			7975: out = 16'(-1593);
			7976: out = 16'(424);
			7977: out = 16'(-94);
			7978: out = 16'(-1940);
			7979: out = 16'(2663);
			7980: out = 16'(-277);
			7981: out = 16'(882);
			7982: out = 16'(423);
			7983: out = 16'(-2655);
			7984: out = 16'(244);
			7985: out = 16'(-250);
			7986: out = 16'(-311);
			7987: out = 16'(-104);
			7988: out = 16'(-1907);
			7989: out = 16'(1645);
			7990: out = 16'(2333);
			7991: out = 16'(-772);
			7992: out = 16'(-156);
			7993: out = 16'(-3114);
			7994: out = 16'(1641);
			7995: out = 16'(-1378);
			7996: out = 16'(341);
			7997: out = 16'(-226);
			7998: out = 16'(2590);
			7999: out = 16'(222);
			8000: out = 16'(-419);
			8001: out = 16'(174);
			8002: out = 16'(-1749);
			8003: out = 16'(-134);
			8004: out = 16'(-163);
			8005: out = 16'(65);
			8006: out = 16'(185);
			8007: out = 16'(-1001);
			8008: out = 16'(1015);
			8009: out = 16'(782);
			8010: out = 16'(-844);
			8011: out = 16'(-2);
			8012: out = 16'(350);
			8013: out = 16'(-58);
			8014: out = 16'(1640);
			8015: out = 16'(-990);
			8016: out = 16'(-128);
			8017: out = 16'(1677);
			8018: out = 16'(-152);
			8019: out = 16'(1165);
			8020: out = 16'(-3521);
			8021: out = 16'(-47);
			8022: out = 16'(1707);
			8023: out = 16'(-1589);
			8024: out = 16'(53);
			8025: out = 16'(-162);
			8026: out = 16'(-415);
			8027: out = 16'(319);
			8028: out = 16'(2409);
			8029: out = 16'(-3054);
			8030: out = 16'(-2580);
			8031: out = 16'(3693);
			8032: out = 16'(-44);
			8033: out = 16'(-1317);
			8034: out = 16'(-491);
			8035: out = 16'(674);
			8036: out = 16'(1512);
			8037: out = 16'(-9);
			8038: out = 16'(2264);
			8039: out = 16'(-1554);
			8040: out = 16'(-916);
			8041: out = 16'(2161);
			8042: out = 16'(-1596);
			8043: out = 16'(93);
			8044: out = 16'(-2054);
			8045: out = 16'(1091);
			8046: out = 16'(2123);
			8047: out = 16'(-626);
			8048: out = 16'(-757);
			8049: out = 16'(-345);
			8050: out = 16'(-218);
			8051: out = 16'(-136);
			8052: out = 16'(171);
			8053: out = 16'(-2689);
			8054: out = 16'(153);
			8055: out = 16'(369);
			8056: out = 16'(771);
			8057: out = 16'(2668);
			8058: out = 16'(24);
			8059: out = 16'(-864);
			8060: out = 16'(-973);
			8061: out = 16'(114);
			8062: out = 16'(-632);
			8063: out = 16'(-635);
			8064: out = 16'(1214);
			8065: out = 16'(258);
			8066: out = 16'(1468);
			8067: out = 16'(590);
			8068: out = 16'(1440);
			8069: out = 16'(-1422);
			8070: out = 16'(-1913);
			8071: out = 16'(724);
			8072: out = 16'(-1387);
			8073: out = 16'(176);
			8074: out = 16'(600);
			8075: out = 16'(1050);
			8076: out = 16'(1960);
			8077: out = 16'(-183);
			8078: out = 16'(314);
			8079: out = 16'(-3180);
			8080: out = 16'(1977);
			8081: out = 16'(1383);
			8082: out = 16'(-1433);
			8083: out = 16'(-377);
			8084: out = 16'(1073);
			8085: out = 16'(-116);
			8086: out = 16'(274);
			8087: out = 16'(-883);
			8088: out = 16'(-569);
			8089: out = 16'(-183);
			8090: out = 16'(-427);
			8091: out = 16'(2040);
			8092: out = 16'(-2052);
			8093: out = 16'(-509);
			8094: out = 16'(414);
			8095: out = 16'(1987);
			8096: out = 16'(-1253);
			8097: out = 16'(22);
			8098: out = 16'(-1563);
			8099: out = 16'(580);
			8100: out = 16'(-15);
			8101: out = 16'(731);
			8102: out = 16'(-49);
			8103: out = 16'(-1740);
			8104: out = 16'(-670);
			8105: out = 16'(1016);
			8106: out = 16'(-296);
			8107: out = 16'(-3713);
			8108: out = 16'(3928);
			8109: out = 16'(339);
			8110: out = 16'(-64);
			8111: out = 16'(-198);
			8112: out = 16'(-1555);
			8113: out = 16'(1747);
			8114: out = 16'(-105);
			8115: out = 16'(-79);
			8116: out = 16'(-222);
			8117: out = 16'(-1847);
			8118: out = 16'(1858);
			8119: out = 16'(1249);
			8120: out = 16'(-766);
			8121: out = 16'(-1496);
			8122: out = 16'(-474);
			8123: out = 16'(248);
			8124: out = 16'(-705);
			8125: out = 16'(271);
			8126: out = 16'(-1877);
			8127: out = 16'(391);
			8128: out = 16'(391);
			8129: out = 16'(557);
			8130: out = 16'(-28);
			8131: out = 16'(-2532);
			8132: out = 16'(1374);
			8133: out = 16'(66);
			8134: out = 16'(-356);
			8135: out = 16'(1416);
			8136: out = 16'(2355);
			8137: out = 16'(-197);
			8138: out = 16'(-576);
			8139: out = 16'(-378);
			8140: out = 16'(-2288);
			8141: out = 16'(846);
			8142: out = 16'(-641);
			8143: out = 16'(-1120);
			8144: out = 16'(977);
			8145: out = 16'(-526);
			8146: out = 16'(2960);
			8147: out = 16'(1404);
			8148: out = 16'(-1164);
			8149: out = 16'(-844);
			8150: out = 16'(-87);
			8151: out = 16'(775);
			8152: out = 16'(66);
			8153: out = 16'(0);
			8154: out = 16'(928);
			8155: out = 16'(-391);
			8156: out = 16'(-268);
			8157: out = 16'(-1514);
			8158: out = 16'(339);
			8159: out = 16'(-861);
			8160: out = 16'(-324);
			8161: out = 16'(2555);
			8162: out = 16'(1231);
			8163: out = 16'(-419);
			8164: out = 16'(-292);
			8165: out = 16'(1903);
			8166: out = 16'(-2532);
			8167: out = 16'(-603);
			8168: out = 16'(119);
			8169: out = 16'(-143);
			8170: out = 16'(-1484);
			8171: out = 16'(1440);
			8172: out = 16'(270);
			8173: out = 16'(328);
			8174: out = 16'(273);
			8175: out = 16'(37);
			8176: out = 16'(270);
			8177: out = 16'(-111);
			8178: out = 16'(-321);
			8179: out = 16'(1286);
			8180: out = 16'(-1082);
			8181: out = 16'(-151);
			8182: out = 16'(497);
			8183: out = 16'(-2596);
			8184: out = 16'(-63);
			8185: out = 16'(821);
			8186: out = 16'(345);
			8187: out = 16'(-558);
			8188: out = 16'(335);
			8189: out = 16'(-702);
			8190: out = 16'(123);
			8191: out = 16'(1475);
			8192: out = 16'(-708);
			8193: out = 16'(-463);
			8194: out = 16'(-1855);
			8195: out = 16'(398);
			8196: out = 16'(2697);
			8197: out = 16'(-202);
			8198: out = 16'(325);
			8199: out = 16'(-475);
			8200: out = 16'(360);
			8201: out = 16'(-1877);
			8202: out = 16'(678);
			8203: out = 16'(266);
			8204: out = 16'(381);
			8205: out = 16'(1626);
			8206: out = 16'(-190);
			8207: out = 16'(-974);
			8208: out = 16'(-54);
			8209: out = 16'(737);
			8210: out = 16'(-742);
			8211: out = 16'(-59);
			8212: out = 16'(-415);
			8213: out = 16'(-1311);
			8214: out = 16'(2147);
			8215: out = 16'(370);
			8216: out = 16'(-1141);
			8217: out = 16'(-847);
			8218: out = 16'(-889);
			8219: out = 16'(-411);
			8220: out = 16'(2087);
			8221: out = 16'(-55);
			8222: out = 16'(-795);
			8223: out = 16'(981);
			8224: out = 16'(1374);
			8225: out = 16'(-263);
			8226: out = 16'(496);
			8227: out = 16'(-2222);
			8228: out = 16'(-311);
			8229: out = 16'(-303);
			8230: out = 16'(951);
			8231: out = 16'(-1124);
			8232: out = 16'(-743);
			8233: out = 16'(366);
			8234: out = 16'(395);
			8235: out = 16'(303);
			8236: out = 16'(-282);
			8237: out = 16'(-682);
			8238: out = 16'(375);
			8239: out = 16'(-77);
			8240: out = 16'(-738);
			8241: out = 16'(1787);
			8242: out = 16'(-1411);
			8243: out = 16'(-353);
			8244: out = 16'(48);
			8245: out = 16'(-215);
			8246: out = 16'(-401);
			8247: out = 16'(-178);
			8248: out = 16'(250);
			8249: out = 16'(-103);
			8250: out = 16'(-909);
			8251: out = 16'(-387);
			8252: out = 16'(2857);
			8253: out = 16'(882);
			8254: out = 16'(-2326);
			8255: out = 16'(773);
			8256: out = 16'(-1903);
			8257: out = 16'(-1577);
			8258: out = 16'(489);
			8259: out = 16'(86);
			8260: out = 16'(407);
			8261: out = 16'(1333);
			8262: out = 16'(531);
			8263: out = 16'(1361);
			8264: out = 16'(-8);
			8265: out = 16'(-128);
			8266: out = 16'(-635);
			8267: out = 16'(-1336);
			8268: out = 16'(336);
			8269: out = 16'(-1068);
			8270: out = 16'(1830);
			8271: out = 16'(-1055);
			8272: out = 16'(1563);
			8273: out = 16'(-229);
			8274: out = 16'(-360);
			8275: out = 16'(-93);
			8276: out = 16'(208);
			8277: out = 16'(-354);
			8278: out = 16'(343);
			8279: out = 16'(275);
			8280: out = 16'(18);
			8281: out = 16'(523);
			8282: out = 16'(659);
			8283: out = 16'(-163);
			8284: out = 16'(-2187);
			8285: out = 16'(-38);
			8286: out = 16'(-1068);
			8287: out = 16'(758);
			8288: out = 16'(-563);
			8289: out = 16'(-559);
			8290: out = 16'(-730);
			8291: out = 16'(-206);
			8292: out = 16'(-1773);
			8293: out = 16'(194);
			8294: out = 16'(-1239);
			8295: out = 16'(1757);
			8296: out = 16'(159);
			8297: out = 16'(1922);
			8298: out = 16'(83);
			8299: out = 16'(-1553);
			8300: out = 16'(1441);
			8301: out = 16'(-1033);
			8302: out = 16'(656);
			8303: out = 16'(-538);
			8304: out = 16'(66);
			8305: out = 16'(-1966);
			8306: out = 16'(-817);
			8307: out = 16'(-164);
			8308: out = 16'(-22);
			8309: out = 16'(-580);
			8310: out = 16'(-878);
			8311: out = 16'(892);
			8312: out = 16'(357);
			8313: out = 16'(1086);
			8314: out = 16'(2825);
			8315: out = 16'(415);
			8316: out = 16'(20);
			8317: out = 16'(-370);
			8318: out = 16'(-199);
			8319: out = 16'(-506);
			8320: out = 16'(522);
			8321: out = 16'(130);
			8322: out = 16'(206);
			8323: out = 16'(-189);
			8324: out = 16'(12);
			8325: out = 16'(1207);
			8326: out = 16'(-2765);
			8327: out = 16'(-117);
			8328: out = 16'(151);
			8329: out = 16'(-1859);
			8330: out = 16'(908);
			8331: out = 16'(5);
			8332: out = 16'(843);
			8333: out = 16'(-181);
			8334: out = 16'(381);
			8335: out = 16'(-510);
			8336: out = 16'(-881);
			8337: out = 16'(1808);
			8338: out = 16'(-685);
			8339: out = 16'(1769);
			8340: out = 16'(931);
			8341: out = 16'(4);
			8342: out = 16'(229);
			8343: out = 16'(-2594);
			8344: out = 16'(372);
			8345: out = 16'(-2205);
			8346: out = 16'(780);
			8347: out = 16'(-2276);
			8348: out = 16'(142);
			8349: out = 16'(1462);
			8350: out = 16'(-1130);
			8351: out = 16'(-50);
			8352: out = 16'(227);
			8353: out = 16'(563);
			8354: out = 16'(267);
			8355: out = 16'(858);
			8356: out = 16'(-252);
			8357: out = 16'(-122);
			8358: out = 16'(-93);
			8359: out = 16'(-202);
			8360: out = 16'(390);
			8361: out = 16'(-2348);
			8362: out = 16'(-897);
			8363: out = 16'(1750);
			8364: out = 16'(-3);
			8365: out = 16'(1462);
			8366: out = 16'(-746);
			8367: out = 16'(434);
			8368: out = 16'(-1708);
			8369: out = 16'(-331);
			8370: out = 16'(-102);
			8371: out = 16'(354);
			8372: out = 16'(679);
			8373: out = 16'(-869);
			8374: out = 16'(1443);
			8375: out = 16'(-2174);
			8376: out = 16'(-776);
			8377: out = 16'(1219);
			8378: out = 16'(-2405);
			8379: out = 16'(1980);
			8380: out = 16'(1130);
			8381: out = 16'(1226);
			8382: out = 16'(1359);
			8383: out = 16'(-249);
			8384: out = 16'(290);
			8385: out = 16'(-3131);
			8386: out = 16'(893);
			8387: out = 16'(-206);
			8388: out = 16'(79);
			8389: out = 16'(764);
			8390: out = 16'(554);
			8391: out = 16'(1199);
			8392: out = 16'(103);
			8393: out = 16'(-1432);
			8394: out = 16'(-857);
			8395: out = 16'(-2005);
			8396: out = 16'(-551);
			8397: out = 16'(868);
			8398: out = 16'(3486);
			8399: out = 16'(296);
			8400: out = 16'(-216);
			8401: out = 16'(-141);
			8402: out = 16'(-955);
			8403: out = 16'(-2367);
			8404: out = 16'(-759);
			8405: out = 16'(90);
			8406: out = 16'(-648);
			8407: out = 16'(1464);
			8408: out = 16'(-421);
			8409: out = 16'(2888);
			8410: out = 16'(-1044);
			8411: out = 16'(120);
			8412: out = 16'(-1160);
			8413: out = 16'(-2145);
			8414: out = 16'(574);
			8415: out = 16'(758);
			8416: out = 16'(841);
			8417: out = 16'(177);
			8418: out = 16'(623);
			8419: out = 16'(-259);
			8420: out = 16'(-278);
			8421: out = 16'(-3141);
			8422: out = 16'(-1313);
			8423: out = 16'(637);
			8424: out = 16'(1483);
			8425: out = 16'(358);
			8426: out = 16'(-2017);
			8427: out = 16'(-102);
			8428: out = 16'(123);
			8429: out = 16'(-553);
			8430: out = 16'(217);
			8431: out = 16'(79);
			8432: out = 16'(-1095);
			8433: out = 16'(2813);
			8434: out = 16'(343);
			8435: out = 16'(683);
			8436: out = 16'(284);
			8437: out = 16'(-873);
			8438: out = 16'(470);
			8439: out = 16'(576);
			8440: out = 16'(-1274);
			8441: out = 16'(49);
			8442: out = 16'(1342);
			8443: out = 16'(-187);
			8444: out = 16'(-12);
			8445: out = 16'(-533);
			8446: out = 16'(-2725);
			8447: out = 16'(1738);
			8448: out = 16'(1436);
			8449: out = 16'(-1628);
			8450: out = 16'(447);
			8451: out = 16'(288);
			8452: out = 16'(-1198);
			8453: out = 16'(-214);
			8454: out = 16'(837);
			8455: out = 16'(-538);
			8456: out = 16'(-517);
			8457: out = 16'(558);
			8458: out = 16'(1916);
			8459: out = 16'(153);
			8460: out = 16'(325);
			8461: out = 16'(-774);
			8462: out = 16'(-789);
			8463: out = 16'(-821);
			8464: out = 16'(891);
			8465: out = 16'(-898);
			8466: out = 16'(-164);
			8467: out = 16'(218);
			8468: out = 16'(1819);
			8469: out = 16'(-636);
			8470: out = 16'(3);
			8471: out = 16'(-616);
			8472: out = 16'(-1938);
			8473: out = 16'(-1278);
			8474: out = 16'(1378);
			8475: out = 16'(356);
			8476: out = 16'(853);
			8477: out = 16'(117);
			8478: out = 16'(-365);
			8479: out = 16'(-639);
			8480: out = 16'(-182);
			8481: out = 16'(2192);
			8482: out = 16'(-1641);
			8483: out = 16'(927);
			8484: out = 16'(-2004);
			8485: out = 16'(124);
			8486: out = 16'(-2288);
			8487: out = 16'(1033);
			8488: out = 16'(381);
			8489: out = 16'(-222);
			8490: out = 16'(274);
			8491: out = 16'(121);
			8492: out = 16'(-249);
			8493: out = 16'(-327);
			8494: out = 16'(816);
			8495: out = 16'(-123);
			8496: out = 16'(-833);
			8497: out = 16'(1336);
			8498: out = 16'(782);
			8499: out = 16'(-229);
			8500: out = 16'(193);
			8501: out = 16'(-409);
			8502: out = 16'(-543);
			8503: out = 16'(532);
			8504: out = 16'(76);
			8505: out = 16'(-1808);
			8506: out = 16'(64);
			8507: out = 16'(972);
			8508: out = 16'(246);
			8509: out = 16'(378);
			8510: out = 16'(333);
			8511: out = 16'(-1066);
			8512: out = 16'(-1177);
			8513: out = 16'(304);
			8514: out = 16'(407);
			8515: out = 16'(-106);
			8516: out = 16'(1758);
			8517: out = 16'(199);
			8518: out = 16'(119);
			8519: out = 16'(-1053);
			8520: out = 16'(-811);
			8521: out = 16'(-240);
			8522: out = 16'(-324);
			8523: out = 16'(-1078);
			8524: out = 16'(-1243);
			8525: out = 16'(2128);
			8526: out = 16'(-775);
			8527: out = 16'(1125);
			8528: out = 16'(-891);
			8529: out = 16'(-696);
			8530: out = 16'(172);
			8531: out = 16'(-1091);
			8532: out = 16'(1551);
			8533: out = 16'(-1889);
			8534: out = 16'(2922);
			8535: out = 16'(-1339);
			8536: out = 16'(-104);
			8537: out = 16'(-721);
			8538: out = 16'(874);
			8539: out = 16'(8);
			8540: out = 16'(-1491);
			8541: out = 16'(-114);
			8542: out = 16'(398);
			8543: out = 16'(531);
			8544: out = 16'(2131);
			8545: out = 16'(-298);
			8546: out = 16'(-514);
			8547: out = 16'(-338);
			8548: out = 16'(550);
			8549: out = 16'(706);
			8550: out = 16'(-2103);
			8551: out = 16'(488);
			8552: out = 16'(890);
			8553: out = 16'(525);
			8554: out = 16'(-729);
			8555: out = 16'(905);
			8556: out = 16'(-2478);
			8557: out = 16'(340);
			8558: out = 16'(1577);
			8559: out = 16'(1310);
			8560: out = 16'(145);
			8561: out = 16'(-595);
			8562: out = 16'(337);
			8563: out = 16'(-161);
			8564: out = 16'(-1957);
			8565: out = 16'(152);
			8566: out = 16'(451);
			8567: out = 16'(263);
			8568: out = 16'(230);
			8569: out = 16'(1207);
			8570: out = 16'(-2090);
			8571: out = 16'(236);
			8572: out = 16'(373);
			8573: out = 16'(-843);
			8574: out = 16'(359);
			8575: out = 16'(1629);
			8576: out = 16'(-179);
			8577: out = 16'(2535);
			8578: out = 16'(-1321);
			8579: out = 16'(-298);
			8580: out = 16'(-1216);
			8581: out = 16'(808);
			8582: out = 16'(380);
			8583: out = 16'(-750);
			8584: out = 16'(1229);
			8585: out = 16'(-807);
			8586: out = 16'(1815);
			8587: out = 16'(-875);
			8588: out = 16'(-316);
			8589: out = 16'(-2739);
			8590: out = 16'(-5);
			8591: out = 16'(131);
			8592: out = 16'(683);
			8593: out = 16'(1028);
			8594: out = 16'(894);
			8595: out = 16'(159);
			8596: out = 16'(-94);
			8597: out = 16'(-31);
			8598: out = 16'(307);
			8599: out = 16'(-798);
			8600: out = 16'(-674);
			8601: out = 16'(2371);
			8602: out = 16'(153);
			8603: out = 16'(529);
			8604: out = 16'(1309);
			8605: out = 16'(228);
			8606: out = 16'(-3174);
			8607: out = 16'(-325);
			8608: out = 16'(104);
			8609: out = 16'(-1765);
			8610: out = 16'(112);
			8611: out = 16'(357);
			8612: out = 16'(1415);
			8613: out = 16'(-1451);
			8614: out = 16'(2158);
			8615: out = 16'(144);
			8616: out = 16'(-915);
			8617: out = 16'(-144);
			8618: out = 16'(767);
			8619: out = 16'(254);
			8620: out = 16'(723);
			8621: out = 16'(12);
			8622: out = 16'(487);
			8623: out = 16'(-221);
			8624: out = 16'(-1886);
			8625: out = 16'(-91);
			8626: out = 16'(821);
			8627: out = 16'(-1099);
			8628: out = 16'(499);
			8629: out = 16'(303);
			8630: out = 16'(-1972);
			8631: out = 16'(2236);
			8632: out = 16'(-142);
			8633: out = 16'(286);
			8634: out = 16'(-148);
			8635: out = 16'(-225);
			8636: out = 16'(-276);
			8637: out = 16'(924);
			8638: out = 16'(346);
			8639: out = 16'(-172);
			8640: out = 16'(-1817);
			8641: out = 16'(-1373);
			8642: out = 16'(-144);
			8643: out = 16'(1741);
			8644: out = 16'(-3193);
			8645: out = 16'(2310);
			8646: out = 16'(-1230);
			8647: out = 16'(-107);
			8648: out = 16'(306);
			8649: out = 16'(452);
			8650: out = 16'(150);
			8651: out = 16'(-3387);
			8652: out = 16'(505);
			8653: out = 16'(1993);
			8654: out = 16'(1058);
			8655: out = 16'(-1382);
			8656: out = 16'(-333);
			8657: out = 16'(6);
			8658: out = 16'(-1893);
			8659: out = 16'(131);
			8660: out = 16'(2254);
			8661: out = 16'(-636);
			8662: out = 16'(4);
			8663: out = 16'(1058);
			8664: out = 16'(-232);
			8665: out = 16'(-2962);
			8666: out = 16'(279);
			8667: out = 16'(-6);
			8668: out = 16'(-324);
			8669: out = 16'(24);
			8670: out = 16'(414);
			8671: out = 16'(283);
			8672: out = 16'(534);
			8673: out = 16'(2888);
			8674: out = 16'(-1674);
			8675: out = 16'(-505);
			8676: out = 16'(-312);
			8677: out = 16'(-153);
			8678: out = 16'(1085);
			8679: out = 16'(-1969);
			8680: out = 16'(95);
			8681: out = 16'(-375);
			8682: out = 16'(1400);
			8683: out = 16'(-769);
			8684: out = 16'(-24);
			8685: out = 16'(-213);
			8686: out = 16'(-407);
			8687: out = 16'(968);
			8688: out = 16'(-208);
			8689: out = 16'(-8);
			8690: out = 16'(-779);
			8691: out = 16'(357);
			8692: out = 16'(-36);
			8693: out = 16'(-756);
			8694: out = 16'(346);
			8695: out = 16'(758);
			8696: out = 16'(-567);
			8697: out = 16'(691);
			8698: out = 16'(-200);
			8699: out = 16'(-638);
			8700: out = 16'(243);
			8701: out = 16'(-896);
			8702: out = 16'(419);
			8703: out = 16'(267);
			8704: out = 16'(-202);
			8705: out = 16'(205);
			8706: out = 16'(697);
			8707: out = 16'(-960);
			8708: out = 16'(-257);
			8709: out = 16'(322);
			8710: out = 16'(200);
			8711: out = 16'(-384);
			8712: out = 16'(982);
			8713: out = 16'(826);
			8714: out = 16'(-3212);
			8715: out = 16'(1986);
			8716: out = 16'(182);
			8717: out = 16'(-383);
			8718: out = 16'(-464);
			8719: out = 16'(904);
			8720: out = 16'(-2079);
			8721: out = 16'(594);
			8722: out = 16'(1110);
			8723: out = 16'(-683);
			8724: out = 16'(-698);
			8725: out = 16'(-66);
			8726: out = 16'(240);
			8727: out = 16'(-244);
			8728: out = 16'(-1437);
			8729: out = 16'(130);
			8730: out = 16'(864);
			8731: out = 16'(-450);
			8732: out = 16'(1899);
			8733: out = 16'(273);
			8734: out = 16'(-320);
			8735: out = 16'(-1610);
			8736: out = 16'(378);
			8737: out = 16'(1206);
			8738: out = 16'(290);
			8739: out = 16'(-139);
			8740: out = 16'(2107);
			8741: out = 16'(254);
			8742: out = 16'(-1507);
			8743: out = 16'(891);
			8744: out = 16'(160);
			8745: out = 16'(-1139);
			8746: out = 16'(-559);
			8747: out = 16'(2006);
			8748: out = 16'(-863);
			8749: out = 16'(-1040);
			8750: out = 16'(1675);
			8751: out = 16'(-923);
			8752: out = 16'(157);
			8753: out = 16'(162);
			8754: out = 16'(955);
			8755: out = 16'(-271);
			8756: out = 16'(-458);
			8757: out = 16'(-1165);
			8758: out = 16'(1297);
			8759: out = 16'(175);
			8760: out = 16'(313);
			8761: out = 16'(897);
			8762: out = 16'(-390);
			8763: out = 16'(-709);
			8764: out = 16'(1218);
			8765: out = 16'(2669);
			8766: out = 16'(-2873);
			8767: out = 16'(-334);
			8768: out = 16'(-817);
			8769: out = 16'(-2310);
			8770: out = 16'(134);
			8771: out = 16'(1489);
			8772: out = 16'(-896);
			8773: out = 16'(-1417);
			8774: out = 16'(-56);
			8775: out = 16'(-1157);
			8776: out = 16'(-518);
			8777: out = 16'(1892);
			8778: out = 16'(1000);
			8779: out = 16'(-638);
			8780: out = 16'(1600);
			8781: out = 16'(412);
			8782: out = 16'(1274);
			8783: out = 16'(-2226);
			8784: out = 16'(258);
			8785: out = 16'(-19);
			8786: out = 16'(-1094);
			8787: out = 16'(-41);
			8788: out = 16'(933);
			8789: out = 16'(-288);
			8790: out = 16'(-1499);
			8791: out = 16'(567);
			8792: out = 16'(-2324);
			8793: out = 16'(137);
			8794: out = 16'(621);
			8795: out = 16'(321);
			8796: out = 16'(810);
			8797: out = 16'(-107);
			8798: out = 16'(635);
			8799: out = 16'(1103);
			8800: out = 16'(353);
			8801: out = 16'(-1928);
			8802: out = 16'(-209);
			8803: out = 16'(604);
			8804: out = 16'(-2086);
			8805: out = 16'(1646);
			8806: out = 16'(295);
			8807: out = 16'(-92);
			8808: out = 16'(-261);
			8809: out = 16'(-235);
			8810: out = 16'(1169);
			8811: out = 16'(-1766);
			8812: out = 16'(755);
			8813: out = 16'(-712);
			8814: out = 16'(-610);
			8815: out = 16'(-545);
			8816: out = 16'(675);
			8817: out = 16'(2999);
			8818: out = 16'(-539);
			8819: out = 16'(-2686);
			8820: out = 16'(1572);
			8821: out = 16'(129);
			8822: out = 16'(-445);
			8823: out = 16'(718);
			8824: out = 16'(107);
			8825: out = 16'(-2773);
			8826: out = 16'(1670);
			8827: out = 16'(1450);
			8828: out = 16'(-836);
			8829: out = 16'(-301);
			8830: out = 16'(-39);
			8831: out = 16'(728);
			8832: out = 16'(-1710);
			8833: out = 16'(-74);
			8834: out = 16'(184);
			8835: out = 16'(1204);
			8836: out = 16'(-34);
			8837: out = 16'(1848);
			8838: out = 16'(-682);
			8839: out = 16'(-2246);
			8840: out = 16'(829);
			8841: out = 16'(26);
			8842: out = 16'(-93);
			8843: out = 16'(-1504);
			8844: out = 16'(562);
			8845: out = 16'(935);
			8846: out = 16'(-2740);
			8847: out = 16'(-481);
			8848: out = 16'(794);
			8849: out = 16'(-1044);
			8850: out = 16'(1255);
			8851: out = 16'(420);
			8852: out = 16'(1535);
			8853: out = 16'(-3201);
			8854: out = 16'(712);
			8855: out = 16'(1006);
			8856: out = 16'(306);
			8857: out = 16'(100);
			8858: out = 16'(135);
			8859: out = 16'(809);
			8860: out = 16'(-1721);
			8861: out = 16'(2475);
			8862: out = 16'(-107);
			8863: out = 16'(-1632);
			8864: out = 16'(97);
			8865: out = 16'(120);
			8866: out = 16'(168);
			8867: out = 16'(66);
			8868: out = 16'(260);
			8869: out = 16'(952);
			8870: out = 16'(-1126);
			8871: out = 16'(-642);
			8872: out = 16'(1175);
			8873: out = 16'(-177);
			8874: out = 16'(-980);
			8875: out = 16'(542);
			8876: out = 16'(375);
			8877: out = 16'(-468);
			8878: out = 16'(83);
			8879: out = 16'(663);
			8880: out = 16'(-454);
			8881: out = 16'(247);
			8882: out = 16'(570);
			8883: out = 16'(203);
			8884: out = 16'(-2162);
			8885: out = 16'(746);
			8886: out = 16'(286);
			8887: out = 16'(1208);
			8888: out = 16'(-496);
			8889: out = 16'(127);
			8890: out = 16'(-118);
			8891: out = 16'(-206);
			8892: out = 16'(-215);
			8893: out = 16'(-1600);
			8894: out = 16'(1033);
			8895: out = 16'(-2058);
			8896: out = 16'(-29);
			8897: out = 16'(860);
			8898: out = 16'(-654);
			8899: out = 16'(282);
			8900: out = 16'(1748);
			8901: out = 16'(-535);
			8902: out = 16'(-1142);
			8903: out = 16'(-1096);
			8904: out = 16'(866);
			8905: out = 16'(195);
			8906: out = 16'(-296);
			8907: out = 16'(381);
			8908: out = 16'(-229);
			8909: out = 16'(155);
			8910: out = 16'(1142);
			8911: out = 16'(1090);
			8912: out = 16'(-691);
			8913: out = 16'(-577);
			8914: out = 16'(611);
			8915: out = 16'(205);
			8916: out = 16'(-165);
			8917: out = 16'(1307);
			8918: out = 16'(-664);
			8919: out = 16'(-304);
			8920: out = 16'(-1738);
			8921: out = 16'(877);
			8922: out = 16'(696);
			8923: out = 16'(-2029);
			8924: out = 16'(1688);
			8925: out = 16'(-698);
			8926: out = 16'(123);
			8927: out = 16'(1645);
			8928: out = 16'(562);
			8929: out = 16'(-1859);
			8930: out = 16'(-987);
			8931: out = 16'(73);
			8932: out = 16'(-499);
			8933: out = 16'(-2110);
			8934: out = 16'(528);
			8935: out = 16'(924);
			8936: out = 16'(384);
			8937: out = 16'(281);
			8938: out = 16'(-66);
			8939: out = 16'(822);
			8940: out = 16'(-1657);
			8941: out = 16'(632);
			8942: out = 16'(587);
			8943: out = 16'(-2503);
			8944: out = 16'(729);
			8945: out = 16'(1013);
			8946: out = 16'(396);
			8947: out = 16'(-1592);
			8948: out = 16'(-7);
			8949: out = 16'(630);
			8950: out = 16'(-2152);
			8951: out = 16'(220);
			8952: out = 16'(-293);
			8953: out = 16'(-186);
			8954: out = 16'(-903);
			8955: out = 16'(1194);
			8956: out = 16'(445);
			8957: out = 16'(-818);
			8958: out = 16'(-2043);
			8959: out = 16'(871);
			8960: out = 16'(831);
			8961: out = 16'(-326);
			8962: out = 16'(-266);
			8963: out = 16'(144);
			8964: out = 16'(-1104);
			8965: out = 16'(328);
			8966: out = 16'(812);
			8967: out = 16'(511);
			8968: out = 16'(41);
			8969: out = 16'(-380);
			8970: out = 16'(23);
			8971: out = 16'(-1240);
			8972: out = 16'(270);
			8973: out = 16'(-460);
			8974: out = 16'(1164);
			8975: out = 16'(-577);
			8976: out = 16'(379);
			8977: out = 16'(1105);
			8978: out = 16'(-1053);
			8979: out = 16'(327);
			8980: out = 16'(1144);
			8981: out = 16'(-590);
			8982: out = 16'(-192);
			8983: out = 16'(316);
			8984: out = 16'(1090);
			8985: out = 16'(-338);
			8986: out = 16'(411);
			8987: out = 16'(-1403);
			8988: out = 16'(-1519);
			8989: out = 16'(220);
			8990: out = 16'(234);
			8991: out = 16'(-229);
			8992: out = 16'(-650);
			8993: out = 16'(658);
			8994: out = 16'(-101);
			8995: out = 16'(1117);
			8996: out = 16'(-88);
			8997: out = 16'(270);
			8998: out = 16'(-170);
			8999: out = 16'(-202);
			9000: out = 16'(1425);
			9001: out = 16'(525);
			9002: out = 16'(-445);
			9003: out = 16'(-1096);
			9004: out = 16'(81);
			9005: out = 16'(107);
			9006: out = 16'(-1550);
			9007: out = 16'(275);
			9008: out = 16'(-856);
			9009: out = 16'(322);
			9010: out = 16'(-49);
			9011: out = 16'(484);
			9012: out = 16'(-174);
			9013: out = 16'(-198);
			9014: out = 16'(399);
			9015: out = 16'(345);
			9016: out = 16'(30);
			9017: out = 16'(236);
			9018: out = 16'(12);
			9019: out = 16'(-529);
			9020: out = 16'(-505);
			9021: out = 16'(538);
			9022: out = 16'(184);
			9023: out = 16'(-230);
			9024: out = 16'(387);
			9025: out = 16'(-41);
			9026: out = 16'(144);
			9027: out = 16'(-642);
			9028: out = 16'(-404);
			9029: out = 16'(1434);
			9030: out = 16'(-1299);
			9031: out = 16'(351);
			9032: out = 16'(-40);
			9033: out = 16'(-128);
			9034: out = 16'(-99);
			9035: out = 16'(1760);
			9036: out = 16'(32);
			9037: out = 16'(-1214);
			9038: out = 16'(265);
			9039: out = 16'(274);
			9040: out = 16'(-188);
			9041: out = 16'(-1887);
			9042: out = 16'(371);
			9043: out = 16'(-1472);
			9044: out = 16'(742);
			9045: out = 16'(582);
			9046: out = 16'(1360);
			9047: out = 16'(-220);
			9048: out = 16'(-632);
			9049: out = 16'(-306);
			9050: out = 16'(234);
			9051: out = 16'(111);
			9052: out = 16'(-744);
			9053: out = 16'(14);
			9054: out = 16'(1114);
			9055: out = 16'(175);
			9056: out = 16'(1677);
			9057: out = 16'(-44);
			9058: out = 16'(-1699);
			9059: out = 16'(-292);
			9060: out = 16'(982);
			9061: out = 16'(-754);
			9062: out = 16'(-253);
			9063: out = 16'(387);
			9064: out = 16'(656);
			9065: out = 16'(-1115);
			9066: out = 16'(277);
			9067: out = 16'(-53);
			9068: out = 16'(-1996);
			9069: out = 16'(187);
			9070: out = 16'(629);
			9071: out = 16'(363);
			9072: out = 16'(-127);
			9073: out = 16'(916);
			9074: out = 16'(2239);
			9075: out = 16'(-1377);
			9076: out = 16'(-1088);
			9077: out = 16'(-126);
			9078: out = 16'(-798);
			9079: out = 16'(-1136);
			9080: out = 16'(-897);
			9081: out = 16'(2191);
			9082: out = 16'(-2251);
			9083: out = 16'(475);
			9084: out = 16'(1433);
			9085: out = 16'(-227);
			9086: out = 16'(-1526);
			9087: out = 16'(1116);
			9088: out = 16'(59);
			9089: out = 16'(-1066);
			9090: out = 16'(16);
			9091: out = 16'(186);
			9092: out = 16'(-879);
			9093: out = 16'(-204);
			9094: out = 16'(244);
			9095: out = 16'(-188);
			9096: out = 16'(-628);
			9097: out = 16'(-452);
			9098: out = 16'(-640);
			9099: out = 16'(564);
			9100: out = 16'(387);
			9101: out = 16'(231);
			9102: out = 16'(210);
			9103: out = 16'(-885);
			9104: out = 16'(-142);
			9105: out = 16'(581);
			9106: out = 16'(-194);
			9107: out = 16'(-545);
			9108: out = 16'(35);
			9109: out = 16'(832);
			9110: out = 16'(-1542);
			9111: out = 16'(1438);
			9112: out = 16'(-298);
			9113: out = 16'(510);
			9114: out = 16'(204);
			9115: out = 16'(-1762);
			9116: out = 16'(1438);
			9117: out = 16'(-1356);
			9118: out = 16'(673);
			9119: out = 16'(-261);
			9120: out = 16'(-156);
			9121: out = 16'(-603);
			9122: out = 16'(531);
			9123: out = 16'(479);
			9124: out = 16'(288);
			9125: out = 16'(-98);
			9126: out = 16'(590);
			9127: out = 16'(-759);
			9128: out = 16'(-25);
			9129: out = 16'(-957);
			9130: out = 16'(1904);
			9131: out = 16'(-1036);
			9132: out = 16'(-14);
			9133: out = 16'(-74);
			9134: out = 16'(-228);
			9135: out = 16'(-855);
			9136: out = 16'(211);
			9137: out = 16'(-1482);
			9138: out = 16'(54);
			9139: out = 16'(252);
			9140: out = 16'(944);
			9141: out = 16'(300);
			9142: out = 16'(-430);
			9143: out = 16'(690);
			9144: out = 16'(297);
			9145: out = 16'(229);
			9146: out = 16'(-162);
			9147: out = 16'(-347);
			9148: out = 16'(271);
			9149: out = 16'(35);
			9150: out = 16'(-124);
			9151: out = 16'(1574);
			9152: out = 16'(-2269);
			9153: out = 16'(8);
			9154: out = 16'(-50);
			9155: out = 16'(557);
			9156: out = 16'(-1859);
			9157: out = 16'(70);
			9158: out = 16'(788);
			9159: out = 16'(-1958);
			9160: out = 16'(1206);
			9161: out = 16'(2278);
			9162: out = 16'(-791);
			9163: out = 16'(574);
			9164: out = 16'(-125);
			9165: out = 16'(175);
			9166: out = 16'(-991);
			9167: out = 16'(-213);
			9168: out = 16'(-320);
			9169: out = 16'(-460);
			9170: out = 16'(37);
			9171: out = 16'(681);
			9172: out = 16'(221);
			9173: out = 16'(704);
			9174: out = 16'(-936);
			9175: out = 16'(85);
			9176: out = 16'(-1103);
			9177: out = 16'(-80);
			9178: out = 16'(853);
			9179: out = 16'(1718);
			9180: out = 16'(79);
			9181: out = 16'(692);
			9182: out = 16'(-1586);
			9183: out = 16'(-1018);
			9184: out = 16'(-341);
			9185: out = 16'(-33);
			9186: out = 16'(-3);
			9187: out = 16'(-32);
			9188: out = 16'(2191);
			9189: out = 16'(-922);
			9190: out = 16'(647);
			9191: out = 16'(131);
			9192: out = 16'(-1833);
			9193: out = 16'(-169);
			9194: out = 16'(-4);
			9195: out = 16'(777);
			9196: out = 16'(732);
			9197: out = 16'(-406);
			9198: out = 16'(1833);
			9199: out = 16'(-487);
			9200: out = 16'(171);
			9201: out = 16'(16);
			9202: out = 16'(-548);
			9203: out = 16'(-811);
			9204: out = 16'(1457);
			9205: out = 16'(-175);
			9206: out = 16'(-136);
			9207: out = 16'(-331);
			9208: out = 16'(-108);
			9209: out = 16'(-2194);
			9210: out = 16'(1039);
			9211: out = 16'(-1408);
			9212: out = 16'(538);
			9213: out = 16'(680);
			9214: out = 16'(-57);
			9215: out = 16'(-560);
			9216: out = 16'(183);
			9217: out = 16'(33);
			9218: out = 16'(936);
			9219: out = 16'(31);
			9220: out = 16'(-108);
			9221: out = 16'(-554);
			9222: out = 16'(60);
			9223: out = 16'(1964);
			9224: out = 16'(-1458);
			9225: out = 16'(-677);
			9226: out = 16'(-1856);
			9227: out = 16'(882);
			9228: out = 16'(609);
			9229: out = 16'(1119);
			9230: out = 16'(370);
			9231: out = 16'(790);
			9232: out = 16'(43);
			9233: out = 16'(633);
			9234: out = 16'(433);
			9235: out = 16'(-359);
			9236: out = 16'(-1150);
			9237: out = 16'(-145);
			9238: out = 16'(506);
			9239: out = 16'(-572);
			9240: out = 16'(312);
			9241: out = 16'(204);
			9242: out = 16'(-1114);
			9243: out = 16'(204);
			9244: out = 16'(-372);
			9245: out = 16'(0);
			9246: out = 16'(-397);
			9247: out = 16'(342);
			9248: out = 16'(239);
			9249: out = 16'(244);
			9250: out = 16'(1225);
			9251: out = 16'(-79);
			9252: out = 16'(-371);
			9253: out = 16'(-224);
			9254: out = 16'(-1110);
			9255: out = 16'(-715);
			9256: out = 16'(1017);
			9257: out = 16'(1503);
			9258: out = 16'(255);
			9259: out = 16'(-197);
			9260: out = 16'(102);
			9261: out = 16'(-381);
			9262: out = 16'(62);
			9263: out = 16'(-755);
			9264: out = 16'(-745);
			9265: out = 16'(65);
			9266: out = 16'(647);
			9267: out = 16'(-1115);
			9268: out = 16'(485);
			9269: out = 16'(-328);
			9270: out = 16'(-1083);
			9271: out = 16'(499);
			9272: out = 16'(99);
			9273: out = 16'(83);
			9274: out = 16'(211);
			9275: out = 16'(184);
			9276: out = 16'(-21);
			9277: out = 16'(-1559);
			9278: out = 16'(1064);
			9279: out = 16'(-1381);
			9280: out = 16'(314);
			9281: out = 16'(121);
			9282: out = 16'(194);
			9283: out = 16'(593);
			9284: out = 16'(-15);
			9285: out = 16'(-525);
			9286: out = 16'(96);
			9287: out = 16'(131);
			9288: out = 16'(867);
			9289: out = 16'(97);
			9290: out = 16'(1279);
			9291: out = 16'(-200);
			9292: out = 16'(419);
			9293: out = 16'(-1415);
			9294: out = 16'(1);
			9295: out = 16'(220);
			9296: out = 16'(-1423);
			9297: out = 16'(-175);
			9298: out = 16'(-310);
			9299: out = 16'(226);
			9300: out = 16'(-322);
			9301: out = 16'(-177);
			9302: out = 16'(-125);
			9303: out = 16'(258);
			9304: out = 16'(-1867);
			9305: out = 16'(266);
			9306: out = 16'(1292);
			9307: out = 16'(445);
			9308: out = 16'(873);
			9309: out = 16'(1200);
			9310: out = 16'(-1642);
			9311: out = 16'(254);
			9312: out = 16'(-571);
			9313: out = 16'(-128);
			9314: out = 16'(-152);
			9315: out = 16'(432);
			9316: out = 16'(-1169);
			9317: out = 16'(387);
			9318: out = 16'(1078);
			9319: out = 16'(-792);
			9320: out = 16'(-249);
			9321: out = 16'(-1038);
			9322: out = 16'(-816);
			9323: out = 16'(102);
			9324: out = 16'(-95);
			9325: out = 16'(-20);
			9326: out = 16'(-629);
			9327: out = 16'(87);
			9328: out = 16'(1155);
			9329: out = 16'(-212);
			9330: out = 16'(87);
			9331: out = 16'(-1470);
			9332: out = 16'(158);
			9333: out = 16'(-385);
			9334: out = 16'(1069);
			9335: out = 16'(9);
			9336: out = 16'(-1089);
			9337: out = 16'(384);
			9338: out = 16'(273);
			9339: out = 16'(-138);
			9340: out = 16'(-449);
			9341: out = 16'(-135);
			9342: out = 16'(-1200);
			9343: out = 16'(1513);
			9344: out = 16'(217);
			9345: out = 16'(-133);
			9346: out = 16'(-261);
			9347: out = 16'(680);
			9348: out = 16'(158);
			9349: out = 16'(-257);
			9350: out = 16'(742);
			9351: out = 16'(-965);
			9352: out = 16'(410);
			9353: out = 16'(-235);
			9354: out = 16'(29);
			9355: out = 16'(-1096);
			9356: out = 16'(-140);
			9357: out = 16'(45);
			9358: out = 16'(933);
			9359: out = 16'(-1752);
			9360: out = 16'(-9);
			9361: out = 16'(-894);
			9362: out = 16'(226);
			9363: out = 16'(653);
			9364: out = 16'(-29);
			9365: out = 16'(1389);
			9366: out = 16'(-1413);
			9367: out = 16'(1570);
			9368: out = 16'(-136);
			9369: out = 16'(-1617);
			9370: out = 16'(-12);
			9371: out = 16'(-180);
			9372: out = 16'(-342);
			9373: out = 16'(-16);
			9374: out = 16'(186);
			9375: out = 16'(-182);
			9376: out = 16'(282);
			9377: out = 16'(404);
			9378: out = 16'(-315);
			9379: out = 16'(-21);
			9380: out = 16'(153);
			9381: out = 16'(146);
			9382: out = 16'(668);
			9383: out = 16'(-1586);
			9384: out = 16'(-661);
			9385: out = 16'(538);
			9386: out = 16'(-149);
			9387: out = 16'(-39);
			9388: out = 16'(-178);
			9389: out = 16'(144);
			9390: out = 16'(279);
			9391: out = 16'(862);
			9392: out = 16'(-266);
			9393: out = 16'(-156);
			9394: out = 16'(-1419);
			9395: out = 16'(-63);
			9396: out = 16'(-517);
			9397: out = 16'(505);
			9398: out = 16'(-1326);
			9399: out = 16'(1313);
			9400: out = 16'(75);
			9401: out = 16'(-900);
			9402: out = 16'(354);
			9403: out = 16'(312);
			9404: out = 16'(-784);
			9405: out = 16'(288);
			9406: out = 16'(1834);
			9407: out = 16'(-95);
			9408: out = 16'(554);
			9409: out = 16'(-191);
			9410: out = 16'(619);
			9411: out = 16'(-1972);
			9412: out = 16'(-136);
			9413: out = 16'(729);
			9414: out = 16'(-1);
			9415: out = 16'(199);
			9416: out = 16'(166);
			9417: out = 16'(1392);
			9418: out = 16'(-1811);
			9419: out = 16'(944);
			9420: out = 16'(-296);
			9421: out = 16'(-1035);
			9422: out = 16'(429);
			9423: out = 16'(1113);
			9424: out = 16'(581);
			9425: out = 16'(-1547);
			9426: out = 16'(669);
			9427: out = 16'(-581);
			9428: out = 16'(-244);
			9429: out = 16'(135);
			9430: out = 16'(-1064);
			9431: out = 16'(-317);
			9432: out = 16'(-51);
			9433: out = 16'(617);
			9434: out = 16'(1591);
			9435: out = 16'(-367);
			9436: out = 16'(-1192);
			9437: out = 16'(-48);
			9438: out = 16'(-192);
			9439: out = 16'(-1231);
			9440: out = 16'(95);
			9441: out = 16'(-42);
			9442: out = 16'(-357);
			9443: out = 16'(-26);
			9444: out = 16'(941);
			9445: out = 16'(-1162);
			9446: out = 16'(-709);
			9447: out = 16'(1072);
			9448: out = 16'(-72);
			9449: out = 16'(18);
			9450: out = 16'(-165);
			9451: out = 16'(-611);
			9452: out = 16'(1309);
			9453: out = 16'(-190);
			9454: out = 16'(-230);
			9455: out = 16'(-666);
			9456: out = 16'(-444);
			9457: out = 16'(-219);
			9458: out = 16'(222);
			9459: out = 16'(848);
			9460: out = 16'(-2096);
			9461: out = 16'(800);
			9462: out = 16'(274);
			9463: out = 16'(-32);
			9464: out = 16'(218);
			9465: out = 16'(223);
			9466: out = 16'(-132);
			9467: out = 16'(-210);
			9468: out = 16'(1084);
			9469: out = 16'(553);
			9470: out = 16'(-1818);
			9471: out = 16'(-760);
			9472: out = 16'(178);
			9473: out = 16'(-124);
			9474: out = 16'(-582);
			9475: out = 16'(-107);
			9476: out = 16'(-77);
			9477: out = 16'(-46);
			9478: out = 16'(671);
			9479: out = 16'(-376);
			9480: out = 16'(-1040);
			9481: out = 16'(237);
			9482: out = 16'(-180);
			9483: out = 16'(754);
			9484: out = 16'(-392);
			9485: out = 16'(-351);
			9486: out = 16'(785);
			9487: out = 16'(1767);
			9488: out = 16'(-2523);
			9489: out = 16'(46);
			9490: out = 16'(-132);
			9491: out = 16'(-172);
			9492: out = 16'(-66);
			9493: out = 16'(861);
			9494: out = 16'(22);
			9495: out = 16'(-2239);
			9496: out = 16'(2230);
			9497: out = 16'(323);
			9498: out = 16'(-1894);
			9499: out = 16'(-2594);
			9500: out = 16'(279);
			9501: out = 16'(638);
			9502: out = 16'(-972);
			9503: out = 16'(454);
			9504: out = 16'(352);
			9505: out = 16'(-1043);
			9506: out = 16'(584);
			9507: out = 16'(-134);
			9508: out = 16'(-20);
			9509: out = 16'(-895);
			9510: out = 16'(218);
			9511: out = 16'(1411);
			9512: out = 16'(-546);
			9513: out = 16'(220);
			9514: out = 16'(-235);
			9515: out = 16'(-194);
			9516: out = 16'(-1580);
			9517: out = 16'(-433);
			9518: out = 16'(489);
			9519: out = 16'(-2166);
			9520: out = 16'(1547);
			9521: out = 16'(612);
			9522: out = 16'(-32);
			9523: out = 16'(-45);
			9524: out = 16'(2531);
			9525: out = 16'(-1064);
			9526: out = 16'(-375);
			9527: out = 16'(259);
			9528: out = 16'(399);
			9529: out = 16'(-1545);
			9530: out = 16'(53);
			9531: out = 16'(925);
			9532: out = 16'(-1577);
			9533: out = 16'(1166);
			9534: out = 16'(-1313);
			9535: out = 16'(346);
			9536: out = 16'(-355);
			9537: out = 16'(240);
			9538: out = 16'(124);
			9539: out = 16'(218);
			9540: out = 16'(-88);
			9541: out = 16'(-181);
			9542: out = 16'(1242);
			9543: out = 16'(-166);
			9544: out = 16'(36);
			9545: out = 16'(-586);
			9546: out = 16'(-76);
			9547: out = 16'(-1177);
			9548: out = 16'(242);
			9549: out = 16'(630);
			9550: out = 16'(-668);
			9551: out = 16'(-50);
			9552: out = 16'(491);
			9553: out = 16'(130);
			9554: out = 16'(-1827);
			9555: out = 16'(139);
			9556: out = 16'(-169);
			9557: out = 16'(-9);
			9558: out = 16'(452);
			9559: out = 16'(-190);
			9560: out = 16'(-335);
			9561: out = 16'(-164);
			9562: out = 16'(-528);
			9563: out = 16'(1845);
			9564: out = 16'(-1705);
			9565: out = 16'(33);
			9566: out = 16'(260);
			9567: out = 16'(-24);
			9568: out = 16'(104);
			9569: out = 16'(270);
			9570: out = 16'(279);
			9571: out = 16'(-217);
			9572: out = 16'(170);
			9573: out = 16'(973);
			9574: out = 16'(621);
			9575: out = 16'(-1712);
			9576: out = 16'(198);
			9577: out = 16'(528);
			9578: out = 16'(-661);
			9579: out = 16'(-212);
			9580: out = 16'(521);
			9581: out = 16'(-711);
			9582: out = 16'(50);
			9583: out = 16'(861);
			9584: out = 16'(197);
			9585: out = 16'(-548);
			9586: out = 16'(217);
			9587: out = 16'(-202);
			9588: out = 16'(779);
			9589: out = 16'(-1433);
			9590: out = 16'(-658);
			9591: out = 16'(1394);
			9592: out = 16'(172);
			9593: out = 16'(259);
			9594: out = 16'(828);
			9595: out = 16'(-1850);
			9596: out = 16'(-174);
			9597: out = 16'(103);
			9598: out = 16'(1497);
			9599: out = 16'(-2839);
			9600: out = 16'(1097);
			9601: out = 16'(1654);
			9602: out = 16'(97);
			9603: out = 16'(108);
			9604: out = 16'(-1389);
			9605: out = 16'(-525);
			9606: out = 16'(-2616);
			9607: out = 16'(1586);
			9608: out = 16'(245);
			9609: out = 16'(-1830);
			9610: out = 16'(477);
			9611: out = 16'(1372);
			9612: out = 16'(1142);
			9613: out = 16'(-1419);
			9614: out = 16'(-693);
			9615: out = 16'(208);
			9616: out = 16'(-1250);
			9617: out = 16'(467);
			9618: out = 16'(-61);
			9619: out = 16'(372);
			9620: out = 16'(-1541);
			9621: out = 16'(1629);
			9622: out = 16'(-689);
			9623: out = 16'(-1036);
			9624: out = 16'(-518);
			9625: out = 16'(1073);
			9626: out = 16'(1096);
			9627: out = 16'(-572);
			9628: out = 16'(1068);
			9629: out = 16'(1169);
			9630: out = 16'(-673);
			9631: out = 16'(420);
			9632: out = 16'(41);
			9633: out = 16'(-339);
			9634: out = 16'(-1191);
			9635: out = 16'(287);
			9636: out = 16'(1159);
			9637: out = 16'(-1016);
			9638: out = 16'(216);
			9639: out = 16'(-352);
			9640: out = 16'(1232);
			9641: out = 16'(111);
			9642: out = 16'(679);
			9643: out = 16'(141);
			9644: out = 16'(-1316);
			9645: out = 16'(-87);
			9646: out = 16'(191);
			9647: out = 16'(-256);
			9648: out = 16'(-863);
			9649: out = 16'(873);
			9650: out = 16'(436);
			9651: out = 16'(214);
			9652: out = 16'(-313);
			9653: out = 16'(662);
			9654: out = 16'(-101);
			9655: out = 16'(-976);
			9656: out = 16'(208);
			9657: out = 16'(114);
			9658: out = 16'(-38);
			9659: out = 16'(-519);
			9660: out = 16'(908);
			9661: out = 16'(-30);
			9662: out = 16'(-29);
			9663: out = 16'(165);
			9664: out = 16'(479);
			9665: out = 16'(-1026);
			9666: out = 16'(107);
			9667: out = 16'(-743);
			9668: out = 16'(1695);
			9669: out = 16'(-598);
			9670: out = 16'(1725);
			9671: out = 16'(256);
			9672: out = 16'(-379);
			9673: out = 16'(-44);
			9674: out = 16'(-212);
			9675: out = 16'(-1359);
			9676: out = 16'(-1446);
			9677: out = 16'(174);
			9678: out = 16'(1123);
			9679: out = 16'(-634);
			9680: out = 16'(241);
			9681: out = 16'(465);
			9682: out = 16'(-102);
			9683: out = 16'(187);
			9684: out = 16'(-232);
			9685: out = 16'(587);
			9686: out = 16'(-901);
			9687: out = 16'(709);
			9688: out = 16'(1547);
			9689: out = 16'(-389);
			9690: out = 16'(-154);
			9691: out = 16'(129);
			9692: out = 16'(-125);
			9693: out = 16'(-764);
			9694: out = 16'(-1092);
			9695: out = 16'(1286);
			9696: out = 16'(129);
			9697: out = 16'(128);
			9698: out = 16'(788);
			9699: out = 16'(197);
			9700: out = 16'(-2844);
			9701: out = 16'(138);
			9702: out = 16'(195);
			9703: out = 16'(602);
			9704: out = 16'(-2269);
			9705: out = 16'(213);
			9706: out = 16'(567);
			9707: out = 16'(661);
			9708: out = 16'(328);
			9709: out = 16'(-22);
			9710: out = 16'(-74);
			9711: out = 16'(-756);
			9712: out = 16'(1247);
			9713: out = 16'(-112);
			9714: out = 16'(-719);
			9715: out = 16'(-172);
			9716: out = 16'(1103);
			9717: out = 16'(-380);
			9718: out = 16'(-283);
			9719: out = 16'(-589);
			9720: out = 16'(814);
			9721: out = 16'(-408);
			9722: out = 16'(762);
			9723: out = 16'(455);
			9724: out = 16'(-1648);
			9725: out = 16'(1469);
			9726: out = 16'(626);
			9727: out = 16'(445);
			9728: out = 16'(-118);
			9729: out = 16'(-1388);
			9730: out = 16'(400);
			9731: out = 16'(-14);
			9732: out = 16'(-545);
			9733: out = 16'(440);
			9734: out = 16'(-1522);
			9735: out = 16'(-188);
			9736: out = 16'(415);
			9737: out = 16'(-15);
			9738: out = 16'(-1000);
			9739: out = 16'(-245);
			9740: out = 16'(672);
			9741: out = 16'(0);
			9742: out = 16'(571);
			9743: out = 16'(-356);
			9744: out = 16'(-160);
			9745: out = 16'(168);
			9746: out = 16'(1129);
			9747: out = 16'(123);
			9748: out = 16'(-54);
			9749: out = 16'(-70);
			9750: out = 16'(-52);
			9751: out = 16'(294);
			9752: out = 16'(593);
			9753: out = 16'(-547);
			9754: out = 16'(-1492);
			9755: out = 16'(490);
			9756: out = 16'(-163);
			9757: out = 16'(150);
			9758: out = 16'(1072);
			9759: out = 16'(-761);
			9760: out = 16'(2020);
			9761: out = 16'(-1133);
			9762: out = 16'(-2010);
			9763: out = 16'(-625);
			9764: out = 16'(421);
			9765: out = 16'(1186);
			9766: out = 16'(-657);
			9767: out = 16'(601);
			9768: out = 16'(-970);
			9769: out = 16'(1296);
			9770: out = 16'(946);
			9771: out = 16'(-873);
			9772: out = 16'(144);
			9773: out = 16'(-1664);
			9774: out = 16'(296);
			9775: out = 16'(1926);
			9776: out = 16'(-338);
			9777: out = 16'(74);
			9778: out = 16'(-264);
			9779: out = 16'(172);
			9780: out = 16'(-947);
			9781: out = 16'(-432);
			9782: out = 16'(-452);
			9783: out = 16'(25);
			9784: out = 16'(322);
			9785: out = 16'(-81);
			9786: out = 16'(1554);
			9787: out = 16'(-63);
			9788: out = 16'(254);
			9789: out = 16'(227);
			9790: out = 16'(-283);
			9791: out = 16'(-1568);
			9792: out = 16'(-496);
			9793: out = 16'(518);
			9794: out = 16'(366);
			9795: out = 16'(237);
			9796: out = 16'(-80);
			9797: out = 16'(-46);
			9798: out = 16'(129);
			9799: out = 16'(-153);
			9800: out = 16'(247);
			9801: out = 16'(-346);
			9802: out = 16'(851);
			9803: out = 16'(-188);
			9804: out = 16'(854);
			9805: out = 16'(315);
			9806: out = 16'(-533);
			9807: out = 16'(46);
			9808: out = 16'(-671);
			9809: out = 16'(-868);
			9810: out = 16'(97);
			9811: out = 16'(-1142);
			9812: out = 16'(534);
			9813: out = 16'(1160);
			9814: out = 16'(-193);
			9815: out = 16'(-51);
			9816: out = 16'(-110);
			9817: out = 16'(115);
			9818: out = 16'(-1727);
			9819: out = 16'(1177);
			9820: out = 16'(405);
			9821: out = 16'(-294);
			9822: out = 16'(-182);
			9823: out = 16'(574);
			9824: out = 16'(-237);
			9825: out = 16'(-1764);
			9826: out = 16'(1582);
			9827: out = 16'(369);
			9828: out = 16'(-378);
			9829: out = 16'(-435);
			9830: out = 16'(977);
			9831: out = 16'(323);
			9832: out = 16'(-78);
			9833: out = 16'(-452);
			9834: out = 16'(-59);
			9835: out = 16'(-1266);
			9836: out = 16'(281);
			9837: out = 16'(354);
			9838: out = 16'(-531);
			9839: out = 16'(-498);
			9840: out = 16'(144);
			9841: out = 16'(-264);
			9842: out = 16'(20);
			9843: out = 16'(-53);
			9844: out = 16'(-44);
			9845: out = 16'(1460);
			9846: out = 16'(168);
			9847: out = 16'(207);
			9848: out = 16'(77);
			9849: out = 16'(-793);
			9850: out = 16'(-1198);
			9851: out = 16'(186);
			9852: out = 16'(-609);
			9853: out = 16'(-629);
			9854: out = 16'(107);
			9855: out = 16'(474);
			9856: out = 16'(576);
			9857: out = 16'(849);
			9858: out = 16'(-740);
			9859: out = 16'(-1072);
			9860: out = 16'(-58);
			9861: out = 16'(-501);
			9862: out = 16'(147);
			9863: out = 16'(285);
			9864: out = 16'(569);
			9865: out = 16'(342);
			9866: out = 16'(499);
			9867: out = 16'(-724);
			9868: out = 16'(-1422);
			9869: out = 16'(541);
			9870: out = 16'(-1263);
			9871: out = 16'(283);
			9872: out = 16'(78);
			9873: out = 16'(-76);
			9874: out = 16'(328);
			9875: out = 16'(838);
			9876: out = 16'(728);
			9877: out = 16'(-1201);
			9878: out = 16'(-476);
			9879: out = 16'(-325);
			9880: out = 16'(158);
			9881: out = 16'(134);
			9882: out = 16'(100);
			9883: out = 16'(472);
			9884: out = 16'(-30);
			9885: out = 16'(1236);
			9886: out = 16'(-193);
			9887: out = 16'(-1230);
			9888: out = 16'(239);
			9889: out = 16'(-93);
			9890: out = 16'(1054);
			9891: out = 16'(206);
			9892: out = 16'(-149);
			9893: out = 16'(489);
			9894: out = 16'(768);
			9895: out = 16'(-1044);
			9896: out = 16'(-2170);
			9897: out = 16'(743);
			9898: out = 16'(-742);
			9899: out = 16'(448);
			9900: out = 16'(738);
			9901: out = 16'(-58);
			9902: out = 16'(-1351);
			9903: out = 16'(97);
			9904: out = 16'(1807);
			9905: out = 16'(-1319);
			9906: out = 16'(-516);
			9907: out = 16'(-398);
			9908: out = 16'(313);
			9909: out = 16'(-619);
			9910: out = 16'(1353);
			9911: out = 16'(190);
			9912: out = 16'(-902);
			9913: out = 16'(188);
			9914: out = 16'(1125);
			9915: out = 16'(70);
			9916: out = 16'(-721);
			9917: out = 16'(-117);
			9918: out = 16'(1006);
			9919: out = 16'(-391);
			9920: out = 16'(161);
			9921: out = 16'(-44);
			9922: out = 16'(124);
			9923: out = 16'(-225);
			9924: out = 16'(-472);
			9925: out = 16'(159);
			9926: out = 16'(-1035);
			9927: out = 16'(-125);
			9928: out = 16'(-466);
			9929: out = 16'(184);
			9930: out = 16'(-90);
			9931: out = 16'(-269);
			9932: out = 16'(360);
			9933: out = 16'(1166);
			9934: out = 16'(-227);
			9935: out = 16'(-640);
			9936: out = 16'(144);
			9937: out = 16'(-193);
			9938: out = 16'(-626);
			9939: out = 16'(245);
			9940: out = 16'(-506);
			9941: out = 16'(867);
			9942: out = 16'(70);
			9943: out = 16'(805);
			9944: out = 16'(-32);
			9945: out = 16'(-550);
			9946: out = 16'(-144);
			9947: out = 16'(-140);
			9948: out = 16'(-506);
			9949: out = 16'(-567);
			9950: out = 16'(1066);
			9951: out = 16'(-109);
			9952: out = 16'(-548);
			9953: out = 16'(1404);
			9954: out = 16'(-1534);
			9955: out = 16'(178);
			9956: out = 16'(-663);
			9957: out = 16'(-1729);
			9958: out = 16'(-554);
			9959: out = 16'(685);
			9960: out = 16'(521);
			9961: out = 16'(331);
			9962: out = 16'(219);
			9963: out = 16'(91);
			9964: out = 16'(29);
			9965: out = 16'(80);
			9966: out = 16'(-221);
			9967: out = 16'(163);
			9968: out = 16'(-935);
			9969: out = 16'(228);
			9970: out = 16'(256);
			9971: out = 16'(562);
			9972: out = 16'(-535);
			9973: out = 16'(53);
			9974: out = 16'(206);
			9975: out = 16'(-878);
			9976: out = 16'(679);
			9977: out = 16'(-535);
			9978: out = 16'(247);
			9979: out = 16'(-1524);
			9980: out = 16'(-177);
			9981: out = 16'(282);
			9982: out = 16'(-555);
			9983: out = 16'(-1464);
			9984: out = 16'(699);
			9985: out = 16'(-238);
			9986: out = 16'(207);
			9987: out = 16'(-1460);
			9988: out = 16'(712);
			9989: out = 16'(396);
			9990: out = 16'(291);
			9991: out = 16'(377);
			9992: out = 16'(-147);
			9993: out = 16'(-96);
			9994: out = 16'(-501);
			9995: out = 16'(527);
			9996: out = 16'(-166);
			9997: out = 16'(-1977);
			9998: out = 16'(-861);
			9999: out = 16'(726);
			10000: out = 16'(56);
			10001: out = 16'(-286);
			10002: out = 16'(549);
			10003: out = 16'(219);
			10004: out = 16'(252);
			10005: out = 16'(144);
			10006: out = 16'(-697);
			10007: out = 16'(-1119);
			10008: out = 16'(543);
			10009: out = 16'(258);
			10010: out = 16'(75);
			10011: out = 16'(841);
			10012: out = 16'(-1494);
			10013: out = 16'(-78);
			10014: out = 16'(-9);
			10015: out = 16'(543);
			10016: out = 16'(-1179);
			10017: out = 16'(-71);
			10018: out = 16'(152);
			10019: out = 16'(588);
			10020: out = 16'(-78);
			10021: out = 16'(443);
			10022: out = 16'(-512);
			10023: out = 16'(-44);
			10024: out = 16'(798);
			10025: out = 16'(-668);
			10026: out = 16'(702);
			10027: out = 16'(-1234);
			10028: out = 16'(568);
			10029: out = 16'(1769);
			10030: out = 16'(-259);
			10031: out = 16'(-115);
			10032: out = 16'(-427);
			10033: out = 16'(406);
			10034: out = 16'(-515);
			10035: out = 16'(132);
			10036: out = 16'(-417);
			10037: out = 16'(-1004);
			10038: out = 16'(778);
			10039: out = 16'(-6);
			10040: out = 16'(405);
			10041: out = 16'(-260);
			10042: out = 16'(-957);
			10043: out = 16'(1236);
			10044: out = 16'(-374);
			10045: out = 16'(26);
			10046: out = 16'(-1210);
			10047: out = 16'(-746);
			10048: out = 16'(716);
			10049: out = 16'(-35);
			10050: out = 16'(1293);
			10051: out = 16'(209);
			10052: out = 16'(-7);
			10053: out = 16'(-86);
			10054: out = 16'(1315);
			10055: out = 16'(-1501);
			10056: out = 16'(-538);
			10057: out = 16'(-243);
			10058: out = 16'(82);
			10059: out = 16'(-90);
			10060: out = 16'(-118);
			10061: out = 16'(832);
			10062: out = 16'(128);
			10063: out = 16'(-986);
			10064: out = 16'(1117);
			10065: out = 16'(-480);
			10066: out = 16'(127);
			10067: out = 16'(-196);
			10068: out = 16'(1210);
			10069: out = 16'(117);
			10070: out = 16'(-18);
			10071: out = 16'(69);
			10072: out = 16'(-171);
			10073: out = 16'(-51);
			10074: out = 16'(-1137);
			10075: out = 16'(-265);
			10076: out = 16'(198);
			10077: out = 16'(271);
			10078: out = 16'(1581);
			10079: out = 16'(10);
			10080: out = 16'(258);
			10081: out = 16'(-823);
			10082: out = 16'(-591);
			10083: out = 16'(-105);
			10084: out = 16'(-1917);
			10085: out = 16'(749);
			10086: out = 16'(-358);
			10087: out = 16'(968);
			10088: out = 16'(-921);
			10089: out = 16'(620);
			10090: out = 16'(-1193);
			10091: out = 16'(182);
			10092: out = 16'(79);
			10093: out = 16'(-60);
			10094: out = 16'(1157);
			10095: out = 16'(96);
			10096: out = 16'(134);
			10097: out = 16'(-176);
			10098: out = 16'(-946);
			10099: out = 16'(-137);
			10100: out = 16'(0);
			10101: out = 16'(-505);
			10102: out = 16'(-114);
			10103: out = 16'(172);
			10104: out = 16'(254);
			10105: out = 16'(941);
			10106: out = 16'(-83);
			10107: out = 16'(-335);
			10108: out = 16'(-854);
			10109: out = 16'(23);
			10110: out = 16'(462);
			10111: out = 16'(-449);
			10112: out = 16'(23);
			10113: out = 16'(759);
			10114: out = 16'(-431);
			10115: out = 16'(-130);
			10116: out = 16'(-195);
			10117: out = 16'(-222);
			10118: out = 16'(-34);
			10119: out = 16'(-100);
			10120: out = 16'(1289);
			10121: out = 16'(-699);
			10122: out = 16'(214);
			10123: out = 16'(-45);
			10124: out = 16'(209);
			10125: out = 16'(-555);
			10126: out = 16'(-669);
			10127: out = 16'(431);
			10128: out = 16'(-100);
			10129: out = 16'(481);
			10130: out = 16'(129);
			10131: out = 16'(207);
			10132: out = 16'(-1113);
			10133: out = 16'(-154);
			10134: out = 16'(445);
			10135: out = 16'(-116);
			10136: out = 16'(280);
			10137: out = 16'(-637);
			10138: out = 16'(1210);
			10139: out = 16'(365);
			10140: out = 16'(-338);
			10141: out = 16'(-1541);
			10142: out = 16'(87);
			10143: out = 16'(-1944);
			10144: out = 16'(87);
			10145: out = 16'(434);
			10146: out = 16'(-198);
			10147: out = 16'(254);
			10148: out = 16'(1575);
			10149: out = 16'(223);
			10150: out = 16'(10);
			10151: out = 16'(-1674);
			10152: out = 16'(10);
			10153: out = 16'(260);
			10154: out = 16'(-235);
			10155: out = 16'(1436);
			10156: out = 16'(88);
			10157: out = 16'(-1);
			10158: out = 16'(-1138);
			10159: out = 16'(1547);
			10160: out = 16'(-1806);
			10161: out = 16'(-68);
			10162: out = 16'(325);
			10163: out = 16'(-130);
			10164: out = 16'(-504);
			10165: out = 16'(1121);
			10166: out = 16'(-812);
			10167: out = 16'(-281);
			10168: out = 16'(-134);
			10169: out = 16'(412);
			10170: out = 16'(-819);
			10171: out = 16'(-93);
			10172: out = 16'(543);
			10173: out = 16'(-30);
			10174: out = 16'(265);
			10175: out = 16'(-835);
			10176: out = 16'(-74);
			10177: out = 16'(157);
			10178: out = 16'(134);
			10179: out = 16'(658);
			10180: out = 16'(105);
			10181: out = 16'(-114);
			10182: out = 16'(-662);
			10183: out = 16'(768);
			10184: out = 16'(-47);
			10185: out = 16'(-1052);
			10186: out = 16'(322);
			10187: out = 16'(721);
			10188: out = 16'(246);
			10189: out = 16'(157);
			10190: out = 16'(99);
			10191: out = 16'(-574);
			10192: out = 16'(-537);
			10193: out = 16'(-789);
			10194: out = 16'(942);
			10195: out = 16'(-444);
			10196: out = 16'(498);
			10197: out = 16'(1098);
			10198: out = 16'(302);
			10199: out = 16'(-1284);
			10200: out = 16'(-528);
			10201: out = 16'(-444);
			10202: out = 16'(-1047);
			10203: out = 16'(-281);
			10204: out = 16'(438);
			10205: out = 16'(1358);
			10206: out = 16'(-231);
			10207: out = 16'(92);
			10208: out = 16'(106);
			10209: out = 16'(-652);
			10210: out = 16'(-732);
			10211: out = 16'(430);
			10212: out = 16'(1374);
			10213: out = 16'(-888);
			10214: out = 16'(1441);
			10215: out = 16'(588);
			10216: out = 16'(-453);
			10217: out = 16'(-584);
			10218: out = 16'(14);
			10219: out = 16'(-418);
			10220: out = 16'(-1681);
			10221: out = 16'(82);
			10222: out = 16'(-38);
			10223: out = 16'(215);
			10224: out = 16'(670);
			10225: out = 16'(-675);
			10226: out = 16'(151);
			10227: out = 16'(-712);
			10228: out = 16'(97);
			10229: out = 16'(229);
			10230: out = 16'(499);
			10231: out = 16'(-829);
			10232: out = 16'(497);
			10233: out = 16'(1298);
			10234: out = 16'(-1497);
			10235: out = 16'(21);
			10236: out = 16'(150);
			10237: out = 16'(-167);
			10238: out = 16'(-272);
			10239: out = 16'(289);
			10240: out = 16'(1238);
			10241: out = 16'(-593);
			10242: out = 16'(-818);
			10243: out = 16'(382);
			10244: out = 16'(-524);
			10245: out = 16'(365);
			10246: out = 16'(-563);
			10247: out = 16'(490);
			10248: out = 16'(-1084);
			10249: out = 16'(992);
			10250: out = 16'(-142);
			10251: out = 16'(-155);
			10252: out = 16'(41);
			10253: out = 16'(-533);
			10254: out = 16'(-36);
			10255: out = 16'(0);
			10256: out = 16'(775);
			10257: out = 16'(150);
			10258: out = 16'(-213);
			10259: out = 16'(746);
			10260: out = 16'(-431);
			10261: out = 16'(-648);
			10262: out = 16'(-992);
			10263: out = 16'(-84);
			10264: out = 16'(810);
			10265: out = 16'(-192);
			10266: out = 16'(295);
			10267: out = 16'(409);
			10268: out = 16'(752);
			10269: out = 16'(-1313);
			10270: out = 16'(612);
			10271: out = 16'(-1119);
			10272: out = 16'(-757);
			10273: out = 16'(1184);
			10274: out = 16'(-481);
			10275: out = 16'(278);
			10276: out = 16'(-1159);
			10277: out = 16'(117);
			10278: out = 16'(-27);
			10279: out = 16'(188);
			10280: out = 16'(-510);
			10281: out = 16'(-441);
			10282: out = 16'(733);
			10283: out = 16'(498);
			10284: out = 16'(186);
			10285: out = 16'(71);
			10286: out = 16'(61);
			10287: out = 16'(-718);
			10288: out = 16'(523);
			10289: out = 16'(-26);
			10290: out = 16'(-1171);
			10291: out = 16'(-1412);
			10292: out = 16'(1171);
			10293: out = 16'(11);
			10294: out = 16'(499);
			10295: out = 16'(361);
			10296: out = 16'(-180);
			10297: out = 16'(-109);
			10298: out = 16'(256);
			10299: out = 16'(213);
			10300: out = 16'(-824);
			10301: out = 16'(-292);
			10302: out = 16'(96);
			10303: out = 16'(118);
			10304: out = 16'(-5);
			10305: out = 16'(-116);
			10306: out = 16'(222);
			10307: out = 16'(340);
			10308: out = 16'(-259);
			10309: out = 16'(-1547);
			10310: out = 16'(597);
			10311: out = 16'(-1145);
			10312: out = 16'(677);
			10313: out = 16'(-53);
			10314: out = 16'(-87);
			10315: out = 16'(342);
			10316: out = 16'(-258);
			10317: out = 16'(404);
			10318: out = 16'(-630);
			10319: out = 16'(-33);
			10320: out = 16'(-46);
			10321: out = 16'(235);
			10322: out = 16'(719);
			10323: out = 16'(422);
			10324: out = 16'(176);
			10325: out = 16'(-198);
			10326: out = 16'(-1766);
			10327: out = 16'(-914);
			10328: out = 16'(-204);
			10329: out = 16'(1103);
			10330: out = 16'(-1065);
			10331: out = 16'(-76);
			10332: out = 16'(426);
			10333: out = 16'(155);
			10334: out = 16'(921);
			10335: out = 16'(-335);
			10336: out = 16'(-1308);
			10337: out = 16'(234);
			10338: out = 16'(-431);
			10339: out = 16'(-410);
			10340: out = 16'(959);
			10341: out = 16'(0);
			10342: out = 16'(484);
			10343: out = 16'(483);
			10344: out = 16'(-404);
			10345: out = 16'(-743);
			10346: out = 16'(-120);
			10347: out = 16'(944);
			10348: out = 16'(-620);
			10349: out = 16'(149);
			10350: out = 16'(189);
			10351: out = 16'(902);
			10352: out = 16'(79);
			10353: out = 16'(13);
			10354: out = 16'(-269);
			10355: out = 16'(-132);
			10356: out = 16'(100);
			10357: out = 16'(675);
			10358: out = 16'(-277);
			10359: out = 16'(-2);
			10360: out = 16'(92);
			10361: out = 16'(-490);
			10362: out = 16'(692);
			10363: out = 16'(-1262);
			10364: out = 16'(185);
			10365: out = 16'(-737);
			10366: out = 16'(-67);
			10367: out = 16'(-287);
			10368: out = 16'(-75);
			10369: out = 16'(264);
			10370: out = 16'(-122);
			10371: out = 16'(-187);
			10372: out = 16'(279);
			10373: out = 16'(-124);
			10374: out = 16'(1089);
			10375: out = 16'(-69);
			10376: out = 16'(-111);
			10377: out = 16'(-48);
			10378: out = 16'(318);
			10379: out = 16'(-469);
			10380: out = 16'(-185);
			10381: out = 16'(-398);
			10382: out = 16'(-451);
			10383: out = 16'(450);
			10384: out = 16'(548);
			10385: out = 16'(-869);
			10386: out = 16'(-10);
			10387: out = 16'(-1062);
			10388: out = 16'(-1005);
			10389: out = 16'(308);
			10390: out = 16'(166);
			10391: out = 16'(41);
			10392: out = 16'(1100);
			10393: out = 16'(344);
			10394: out = 16'(-872);
			10395: out = 16'(194);
			10396: out = 16'(139);
			10397: out = 16'(250);
			10398: out = 16'(-141);
			10399: out = 16'(1181);
			10400: out = 16'(-1058);
			10401: out = 16'(-226);
			10402: out = 16'(1002);
			10403: out = 16'(-250);
			10404: out = 16'(-359);
			10405: out = 16'(-1551);
			10406: out = 16'(-417);
			10407: out = 16'(761);
			10408: out = 16'(-358);
			10409: out = 16'(459);
			10410: out = 16'(-995);
			10411: out = 16'(1336);
			10412: out = 16'(-321);
			10413: out = 16'(77);
			10414: out = 16'(356);
			10415: out = 16'(-216);
			10416: out = 16'(108);
			10417: out = 16'(-217);
			10418: out = 16'(-494);
			10419: out = 16'(161);
			10420: out = 16'(-737);
			10421: out = 16'(170);
			10422: out = 16'(-1039);
			10423: out = 16'(-186);
			10424: out = 16'(248);
			10425: out = 16'(-138);
			10426: out = 16'(-159);
			10427: out = 16'(516);
			10428: out = 16'(714);
			10429: out = 16'(-627);
			10430: out = 16'(657);
			10431: out = 16'(-76);
			10432: out = 16'(28);
			10433: out = 16'(300);
			10434: out = 16'(140);
			10435: out = 16'(-509);
			10436: out = 16'(-241);
			10437: out = 16'(-55);
			10438: out = 16'(-70);
			10439: out = 16'(1043);
			10440: out = 16'(-705);
			10441: out = 16'(-57);
			10442: out = 16'(503);
			10443: out = 16'(-806);
			10444: out = 16'(-258);
			10445: out = 16'(455);
			10446: out = 16'(90);
			10447: out = 16'(-744);
			10448: out = 16'(657);
			10449: out = 16'(-809);
			10450: out = 16'(-999);
			10451: out = 16'(563);
			10452: out = 16'(1080);
			10453: out = 16'(-748);
			10454: out = 16'(862);
			10455: out = 16'(-1240);
			10456: out = 16'(480);
			10457: out = 16'(-90);
			10458: out = 16'(-101);
			10459: out = 16'(-459);
			10460: out = 16'(160);
			10461: out = 16'(489);
			10462: out = 16'(578);
			10463: out = 16'(67);
			10464: out = 16'(-1288);
			10465: out = 16'(-172);
			10466: out = 16'(-129);
			10467: out = 16'(181);
			10468: out = 16'(-994);
			10469: out = 16'(1476);
			10470: out = 16'(489);
			10471: out = 16'(24);
			10472: out = 16'(-368);
			10473: out = 16'(843);
			10474: out = 16'(-952);
			10475: out = 16'(-698);
			10476: out = 16'(578);
			10477: out = 16'(-136);
			10478: out = 16'(-269);
			10479: out = 16'(204);
			10480: out = 16'(172);
			10481: out = 16'(-154);
			10482: out = 16'(-1114);
			10483: out = 16'(-154);
			10484: out = 16'(-67);
			10485: out = 16'(-91);
			10486: out = 16'(222);
			10487: out = 16'(1040);
			10488: out = 16'(273);
			10489: out = 16'(77);
			10490: out = 16'(-910);
			10491: out = 16'(683);
			10492: out = 16'(-926);
			10493: out = 16'(-749);
			10494: out = 16'(665);
			10495: out = 16'(103);
			10496: out = 16'(-431);
			10497: out = 16'(585);
			10498: out = 16'(192);
			10499: out = 16'(-687);
			10500: out = 16'(-770);
			10501: out = 16'(977);
			10502: out = 16'(-108);
			10503: out = 16'(-519);
			10504: out = 16'(218);
			10505: out = 16'(-585);
			10506: out = 16'(403);
			10507: out = 16'(-352);
			10508: out = 16'(168);
			10509: out = 16'(-166);
			10510: out = 16'(-691);
			10511: out = 16'(-168);
			10512: out = 16'(1083);
			10513: out = 16'(190);
			10514: out = 16'(-589);
			10515: out = 16'(591);
			10516: out = 16'(-86);
			10517: out = 16'(-861);
			10518: out = 16'(71);
			10519: out = 16'(836);
			10520: out = 16'(-225);
			10521: out = 16'(-757);
			10522: out = 16'(234);
			10523: out = 16'(-625);
			10524: out = 16'(354);
			10525: out = 16'(-447);
			10526: out = 16'(289);
			10527: out = 16'(-566);
			10528: out = 16'(-560);
			10529: out = 16'(1083);
			10530: out = 16'(97);
			10531: out = 16'(26);
			10532: out = 16'(660);
			10533: out = 16'(-910);
			10534: out = 16'(158);
			10535: out = 16'(-643);
			10536: out = 16'(-23);
			10537: out = 16'(163);
			10538: out = 16'(211);
			10539: out = 16'(152);
			10540: out = 16'(139);
			10541: out = 16'(374);
			10542: out = 16'(-992);
			10543: out = 16'(181);
			10544: out = 16'(-452);
			10545: out = 16'(-925);
			10546: out = 16'(468);
			10547: out = 16'(570);
			10548: out = 16'(-66);
			10549: out = 16'(-59);
			10550: out = 16'(-253);
			10551: out = 16'(-77);
			10552: out = 16'(-702);
			10553: out = 16'(-30);
			10554: out = 16'(-502);
			10555: out = 16'(10);
			10556: out = 16'(244);
			10557: out = 16'(1032);
			10558: out = 16'(15);
			10559: out = 16'(129);
			10560: out = 16'(64);
			10561: out = 16'(349);
			10562: out = 16'(373);
			10563: out = 16'(-1012);
			10564: out = 16'(805);
			10565: out = 16'(-436);
			10566: out = 16'(38);
			10567: out = 16'(-311);
			10568: out = 16'(-195);
			10569: out = 16'(383);
			10570: out = 16'(-427);
			10571: out = 16'(778);
			10572: out = 16'(-292);
			10573: out = 16'(-425);
			10574: out = 16'(67);
			10575: out = 16'(275);
			10576: out = 16'(828);
			10577: out = 16'(-565);
			10578: out = 16'(1057);
			10579: out = 16'(-82);
			10580: out = 16'(-145);
			10581: out = 16'(-143);
			10582: out = 16'(-1197);
			10583: out = 16'(-141);
			10584: out = 16'(-599);
			10585: out = 16'(351);
			10586: out = 16'(-98);
			10587: out = 16'(-344);
			10588: out = 16'(722);
			10589: out = 16'(-259);
			10590: out = 16'(82);
			10591: out = 16'(-601);
			10592: out = 16'(134);
			10593: out = 16'(-768);
			10594: out = 16'(9);
			10595: out = 16'(-165);
			10596: out = 16'(1239);
			10597: out = 16'(512);
			10598: out = 16'(93);
			10599: out = 16'(-93);
			10600: out = 16'(-1161);
			10601: out = 16'(78);
			10602: out = 16'(264);
			10603: out = 16'(-105);
			10604: out = 16'(-301);
			10605: out = 16'(-512);
			10606: out = 16'(147);
			10607: out = 16'(-404);
			10608: out = 16'(112);
			10609: out = 16'(97);
			10610: out = 16'(-1370);
			10611: out = 16'(1260);
			10612: out = 16'(-184);
			10613: out = 16'(734);
			10614: out = 16'(736);
			10615: out = 16'(-310);
			10616: out = 16'(387);
			10617: out = 16'(-205);
			10618: out = 16'(91);
			10619: out = 16'(-1118);
			10620: out = 16'(815);
			10621: out = 16'(-132);
			10622: out = 16'(-277);
			10623: out = 16'(-33);
			10624: out = 16'(-670);
			10625: out = 16'(648);
			10626: out = 16'(88);
			10627: out = 16'(-801);
			10628: out = 16'(-96);
			10629: out = 16'(514);
			10630: out = 16'(-212);
			10631: out = 16'(11);
			10632: out = 16'(-210);
			10633: out = 16'(488);
			10634: out = 16'(-194);
			10635: out = 16'(65);
			10636: out = 16'(227);
			10637: out = 16'(131);
			10638: out = 16'(-898);
			10639: out = 16'(156);
			10640: out = 16'(412);
			10641: out = 16'(-34);
			10642: out = 16'(-791);
			10643: out = 16'(-3);
			10644: out = 16'(251);
			10645: out = 16'(-1390);
			10646: out = 16'(783);
			10647: out = 16'(-65);
			10648: out = 16'(598);
			10649: out = 16'(-683);
			10650: out = 16'(285);
			10651: out = 16'(253);
			10652: out = 16'(-634);
			10653: out = 16'(-569);
			10654: out = 16'(808);
			10655: out = 16'(364);
			10656: out = 16'(-220);
			10657: out = 16'(394);
			10658: out = 16'(-54);
			10659: out = 16'(-722);
			10660: out = 16'(-14);
			10661: out = 16'(-161);
			10662: out = 16'(-691);
			10663: out = 16'(396);
			10664: out = 16'(4);
			10665: out = 16'(757);
			10666: out = 16'(388);
			10667: out = 16'(-53);
			10668: out = 16'(-187);
			10669: out = 16'(-215);
			10670: out = 16'(126);
			10671: out = 16'(1);
			10672: out = 16'(52);
			10673: out = 16'(-132);
			10674: out = 16'(-447);
			10675: out = 16'(735);
			10676: out = 16'(794);
			10677: out = 16'(-1210);
			10678: out = 16'(29);
			10679: out = 16'(217);
			10680: out = 16'(-385);
			10681: out = 16'(359);
			10682: out = 16'(591);
			10683: out = 16'(-238);
			10684: out = 16'(-879);
			10685: out = 16'(668);
			10686: out = 16'(-712);
			10687: out = 16'(-54);
			10688: out = 16'(110);
			10689: out = 16'(307);
			10690: out = 16'(146);
			10691: out = 16'(-38);
			10692: out = 16'(-62);
			10693: out = 16'(9);
			10694: out = 16'(-303);
			10695: out = 16'(112);
			10696: out = 16'(582);
			10697: out = 16'(-99);
			10698: out = 16'(55);
			10699: out = 16'(20);
			10700: out = 16'(-117);
			10701: out = 16'(-931);
			10702: out = 16'(-574);
			10703: out = 16'(117);
			10704: out = 16'(17);
			10705: out = 16'(-102);
			10706: out = 16'(852);
			10707: out = 16'(240);
			10708: out = 16'(24);
			10709: out = 16'(-560);
			10710: out = 16'(-114);
			10711: out = 16'(-950);
			10712: out = 16'(-341);
			10713: out = 16'(827);
			10714: out = 16'(-48);
			10715: out = 16'(13);
			10716: out = 16'(335);
			10717: out = 16'(-159);
			10718: out = 16'(-307);
			10719: out = 16'(-298);
			10720: out = 16'(-154);
			10721: out = 16'(371);
			10722: out = 16'(-149);
			10723: out = 16'(-101);
			10724: out = 16'(1210);
			10725: out = 16'(165);
			10726: out = 16'(-1483);
			10727: out = 16'(-189);
			10728: out = 16'(-793);
			10729: out = 16'(-939);
			10730: out = 16'(-100);
			10731: out = 16'(1135);
			10732: out = 16'(166);
			10733: out = 16'(-236);
			10734: out = 16'(1025);
			10735: out = 16'(166);
			10736: out = 16'(-614);
			10737: out = 16'(-818);
			10738: out = 16'(188);
			10739: out = 16'(-588);
			10740: out = 16'(-717);
			10741: out = 16'(1177);
			10742: out = 16'(45);
			10743: out = 16'(-324);
			10744: out = 16'(-433);
			10745: out = 16'(398);
			10746: out = 16'(-306);
			10747: out = 16'(-583);
			10748: out = 16'(477);
			10749: out = 16'(43);
			10750: out = 16'(-72);
			10751: out = 16'(272);
			10752: out = 16'(-90);
			10753: out = 16'(-61);
			10754: out = 16'(-408);
			10755: out = 16'(-56);
			10756: out = 16'(463);
			10757: out = 16'(-299);
			10758: out = 16'(-177);
			10759: out = 16'(897);
			10760: out = 16'(-14);
			10761: out = 16'(-645);
			10762: out = 16'(520);
			10763: out = 16'(-633);
			10764: out = 16'(-84);
			10765: out = 16'(252);
			10766: out = 16'(256);
			10767: out = 16'(78);
			10768: out = 16'(-779);
			10769: out = 16'(104);
			10770: out = 16'(87);
			10771: out = 16'(-595);
			10772: out = 16'(-1019);
			10773: out = 16'(277);
			10774: out = 16'(435);
			10775: out = 16'(146);
			10776: out = 16'(345);
			10777: out = 16'(-84);
			10778: out = 16'(-761);
			10779: out = 16'(-93);
			10780: out = 16'(369);
			10781: out = 16'(484);
			10782: out = 16'(-403);
			10783: out = 16'(708);
			10784: out = 16'(37);
			10785: out = 16'(-332);
			10786: out = 16'(427);
			10787: out = 16'(-26);
			10788: out = 16'(-71);
			10789: out = 16'(-1075);
			10790: out = 16'(300);
			10791: out = 16'(140);
			10792: out = 16'(-94);
			10793: out = 16'(-107);
			10794: out = 16'(96);
			10795: out = 16'(-44);
			10796: out = 16'(-728);
			10797: out = 16'(361);
			10798: out = 16'(-463);
			10799: out = 16'(381);
			10800: out = 16'(2);
			10801: out = 16'(-166);
			10802: out = 16'(-349);
			10803: out = 16'(-57);
			10804: out = 16'(52);
			10805: out = 16'(74);
			10806: out = 16'(-89);
			10807: out = 16'(-630);
			10808: out = 16'(398);
			10809: out = 16'(199);
			10810: out = 16'(-337);
			10811: out = 16'(515);
			10812: out = 16'(8);
			10813: out = 16'(-276);
			10814: out = 16'(459);
			10815: out = 16'(823);
			10816: out = 16'(109);
			10817: out = 16'(-508);
			10818: out = 16'(233);
			10819: out = 16'(-382);
			10820: out = 16'(87);
			10821: out = 16'(-126);
			10822: out = 16'(-448);
			10823: out = 16'(269);
			10824: out = 16'(-574);
			10825: out = 16'(297);
			10826: out = 16'(-156);
			10827: out = 16'(-696);
			10828: out = 16'(-183);
			10829: out = 16'(143);
			10830: out = 16'(271);
			10831: out = 16'(-302);
			10832: out = 16'(714);
			10833: out = 16'(162);
			10834: out = 16'(-887);
			10835: out = 16'(85);
			10836: out = 16'(202);
			10837: out = 16'(-851);
			10838: out = 16'(195);
			10839: out = 16'(-15);
			10840: out = 16'(310);
			10841: out = 16'(-57);
			10842: out = 16'(950);
			10843: out = 16'(-356);
			10844: out = 16'(142);
			10845: out = 16'(-918);
			10846: out = 16'(-101);
			10847: out = 16'(-172);
			10848: out = 16'(297);
			10849: out = 16'(468);
			10850: out = 16'(-443);
			10851: out = 16'(-61);
			10852: out = 16'(-90);
			10853: out = 16'(39);
			10854: out = 16'(-339);
			10855: out = 16'(-231);
			10856: out = 16'(-484);
			10857: out = 16'(289);
			10858: out = 16'(345);
			10859: out = 16'(499);
			10860: out = 16'(453);
			10861: out = 16'(238);
			10862: out = 16'(-587);
			10863: out = 16'(-917);
			10864: out = 16'(-496);
			10865: out = 16'(159);
			10866: out = 16'(287);
			10867: out = 16'(-344);
			10868: out = 16'(190);
			10869: out = 16'(630);
			10870: out = 16'(315);
			10871: out = 16'(-520);
			10872: out = 16'(-513);
			10873: out = 16'(-847);
			10874: out = 16'(-46);
			10875: out = 16'(400);
			10876: out = 16'(529);
			10877: out = 16'(77);
			10878: out = 16'(-1123);
			10879: out = 16'(347);
			10880: out = 16'(145);
			10881: out = 16'(-332);
			10882: out = 16'(121);
			10883: out = 16'(-67);
			10884: out = 16'(536);
			10885: out = 16'(345);
			10886: out = 16'(-10);
			10887: out = 16'(8);
			10888: out = 16'(-136);
			10889: out = 16'(-1106);
			10890: out = 16'(-402);
			10891: out = 16'(835);
			10892: out = 16'(-344);
			10893: out = 16'(659);
			10894: out = 16'(646);
			10895: out = 16'(-155);
			10896: out = 16'(-642);
			10897: out = 16'(-18);
			10898: out = 16'(126);
			10899: out = 16'(-118);
			10900: out = 16'(-10);
			10901: out = 16'(-217);
			10902: out = 16'(484);
			10903: out = 16'(-335);
			10904: out = 16'(109);
			10905: out = 16'(16);
			10906: out = 16'(-771);
			10907: out = 16'(-562);
			10908: out = 16'(-11);
			10909: out = 16'(390);
			10910: out = 16'(-4);
			10911: out = 16'(452);
			10912: out = 16'(190);
			10913: out = 16'(-897);
			10914: out = 16'(100);
			10915: out = 16'(-90);
			10916: out = 16'(-35);
			10917: out = 16'(-484);
			10918: out = 16'(-19);
			10919: out = 16'(787);
			10920: out = 16'(-76);
			10921: out = 16'(-307);
			10922: out = 16'(116);
			10923: out = 16'(-1035);
			10924: out = 16'(-184);
			10925: out = 16'(249);
			10926: out = 16'(560);
			10927: out = 16'(-162);
			10928: out = 16'(141);
			10929: out = 16'(380);
			10930: out = 16'(59);
			10931: out = 16'(-61);
			10932: out = 16'(-267);
			10933: out = 16'(594);
			10934: out = 16'(-154);
			10935: out = 16'(-295);
			10936: out = 16'(410);
			10937: out = 16'(-23);
			10938: out = 16'(-496);
			10939: out = 16'(301);
			10940: out = 16'(44);
			10941: out = 16'(-793);
			10942: out = 16'(-891);
			10943: out = 16'(866);
			10944: out = 16'(27);
			10945: out = 16'(-679);
			10946: out = 16'(334);
			10947: out = 16'(292);
			10948: out = 16'(-971);
			10949: out = 16'(600);
			10950: out = 16'(0);
			10951: out = 16'(320);
			10952: out = 16'(-548);
			10953: out = 16'(151);
			10954: out = 16'(556);
			10955: out = 16'(-738);
			10956: out = 16'(8);
			10957: out = 16'(58);
			10958: out = 16'(-273);
			10959: out = 16'(-143);
			10960: out = 16'(621);
			10961: out = 16'(206);
			10962: out = 16'(-7);
			10963: out = 16'(-278);
			10964: out = 16'(-32);
			10965: out = 16'(-269);
			10966: out = 16'(-327);
			10967: out = 16'(53);
			10968: out = 16'(211);
			10969: out = 16'(508);
			10970: out = 16'(-6);
			10971: out = 16'(562);
			10972: out = 16'(10);
			10973: out = 16'(-1097);
			10974: out = 16'(70);
			10975: out = 16'(69);
			10976: out = 16'(46);
			10977: out = 16'(154);
			10978: out = 16'(785);
			10979: out = 16'(193);
			10980: out = 16'(-366);
			10981: out = 16'(253);
			10982: out = 16'(-173);
			10983: out = 16'(-615);
			10984: out = 16'(-152);
			10985: out = 16'(-123);
			10986: out = 16'(851);
			10987: out = 16'(-373);
			10988: out = 16'(160);
			10989: out = 16'(481);
			10990: out = 16'(-462);
			10991: out = 16'(-1520);
			10992: out = 16'(341);
			10993: out = 16'(215);
			10994: out = 16'(-1298);
			10995: out = 16'(864);
			10996: out = 16'(314);
			10997: out = 16'(-294);
			10998: out = 16'(168);
			10999: out = 16'(360);
			11000: out = 16'(-512);
			11001: out = 16'(-453);
			11002: out = 16'(8);
			11003: out = 16'(492);
			11004: out = 16'(513);
			11005: out = 16'(108);
			11006: out = 16'(-114);
			11007: out = 16'(-136);
			11008: out = 16'(-871);
			11009: out = 16'(463);
			11010: out = 16'(37);
			11011: out = 16'(87);
			11012: out = 16'(-724);
			11013: out = 16'(-12);
			11014: out = 16'(233);
			11015: out = 16'(-266);
			11016: out = 16'(124);
			11017: out = 16'(93);
			11018: out = 16'(-825);
			11019: out = 16'(-154);
			11020: out = 16'(207);
			11021: out = 16'(584);
			11022: out = 16'(-808);
			11023: out = 16'(302);
			11024: out = 16'(128);
			11025: out = 16'(190);
			11026: out = 16'(-342);
			11027: out = 16'(175);
			11028: out = 16'(287);
			11029: out = 16'(-1143);
			11030: out = 16'(828);
			11031: out = 16'(20);
			11032: out = 16'(-338);
			11033: out = 16'(-99);
			11034: out = 16'(-510);
			11035: out = 16'(8);
			11036: out = 16'(-378);
			11037: out = 16'(-172);
			11038: out = 16'(729);
			11039: out = 16'(81);
			11040: out = 16'(-1030);
			11041: out = 16'(194);
			11042: out = 16'(465);
			11043: out = 16'(-113);
			11044: out = 16'(108);
			11045: out = 16'(-117);
			11046: out = 16'(-344);
			11047: out = 16'(83);
			11048: out = 16'(634);
			11049: out = 16'(273);
			11050: out = 16'(-753);
			11051: out = 16'(-153);
			11052: out = 16'(-211);
			11053: out = 16'(-26);
			11054: out = 16'(137);
			11055: out = 16'(-99);
			11056: out = 16'(288);
			11057: out = 16'(-615);
			11058: out = 16'(20);
			11059: out = 16'(-255);
			11060: out = 16'(510);
			11061: out = 16'(-50);
			11062: out = 16'(-344);
			11063: out = 16'(772);
			11064: out = 16'(-385);
			11065: out = 16'(185);
			11066: out = 16'(679);
			11067: out = 16'(58);
			11068: out = 16'(-431);
			11069: out = 16'(-657);
			11070: out = 16'(0);
			11071: out = 16'(-115);
			11072: out = 16'(-128);
			11073: out = 16'(-99);
			11074: out = 16'(-44);
			11075: out = 16'(-262);
			11076: out = 16'(71);
			11077: out = 16'(386);
			11078: out = 16'(-4);
			11079: out = 16'(-36);
			11080: out = 16'(183);
			11081: out = 16'(-147);
			11082: out = 16'(-454);
			11083: out = 16'(50);
			11084: out = 16'(-85);
			11085: out = 16'(-71);
			11086: out = 16'(92);
			11087: out = 16'(148);
			11088: out = 16'(145);
			11089: out = 16'(168);
			11090: out = 16'(-667);
			11091: out = 16'(-92);
			11092: out = 16'(-480);
			11093: out = 16'(-144);
			11094: out = 16'(28);
			11095: out = 16'(138);
			11096: out = 16'(282);
			11097: out = 16'(97);
			11098: out = 16'(360);
			11099: out = 16'(-437);
			11100: out = 16'(-34);
			11101: out = 16'(-258);
			11102: out = 16'(-230);
			11103: out = 16'(-270);
			11104: out = 16'(210);
			11105: out = 16'(120);
			11106: out = 16'(491);
			11107: out = 16'(-498);
			11108: out = 16'(-57);
			11109: out = 16'(66);
			11110: out = 16'(-695);
			11111: out = 16'(-542);
			11112: out = 16'(394);
			11113: out = 16'(156);
			11114: out = 16'(259);
			11115: out = 16'(44);
			11116: out = 16'(523);
			11117: out = 16'(-78);
			11118: out = 16'(-342);
			11119: out = 16'(-100);
			11120: out = 16'(-244);
			11121: out = 16'(-88);
			11122: out = 16'(5);
			11123: out = 16'(233);
			11124: out = 16'(110);
			11125: out = 16'(-138);
			11126: out = 16'(-17);
			11127: out = 16'(-404);
			11128: out = 16'(98);
			11129: out = 16'(-378);
			11130: out = 16'(50);
			11131: out = 16'(155);
			11132: out = 16'(-65);
			11133: out = 16'(650);
			11134: out = 16'(82);
			11135: out = 16'(-76);
			11136: out = 16'(-825);
			11137: out = 16'(-77);
			11138: out = 16'(406);
			11139: out = 16'(-223);
			11140: out = 16'(-132);
			11141: out = 16'(54);
			11142: out = 16'(-34);
			11143: out = 16'(202);
			11144: out = 16'(-314);
			11145: out = 16'(77);
			11146: out = 16'(-117);
			11147: out = 16'(-172);
			11148: out = 16'(673);
			11149: out = 16'(-189);
			11150: out = 16'(244);
			11151: out = 16'(-428);
			11152: out = 16'(57);
			11153: out = 16'(-262);
			11154: out = 16'(-264);
			11155: out = 16'(-160);
			11156: out = 16'(163);
			11157: out = 16'(14);
			11158: out = 16'(79);
			11159: out = 16'(137);
			11160: out = 16'(-95);
			11161: out = 16'(471);
			11162: out = 16'(-104);
			11163: out = 16'(-479);
			11164: out = 16'(-309);
			11165: out = 16'(441);
			11166: out = 16'(330);
			11167: out = 16'(6);
			11168: out = 16'(61);
			11169: out = 16'(-909);
			11170: out = 16'(43);
			11171: out = 16'(222);
			11172: out = 16'(-687);
			11173: out = 16'(58);
			11174: out = 16'(-71);
			11175: out = 16'(122);
			11176: out = 16'(430);
			11177: out = 16'(-88);
			11178: out = 16'(-236);
			11179: out = 16'(-878);
			11180: out = 16'(-450);
			11181: out = 16'(-374);
			11182: out = 16'(382);
			11183: out = 16'(890);
			11184: out = 16'(38);
			11185: out = 16'(-87);
			11186: out = 16'(-347);
			11187: out = 16'(-112);
			11188: out = 16'(634);
			11189: out = 16'(-660);
			11190: out = 16'(-72);
			11191: out = 16'(-148);
			11192: out = 16'(-204);
			11193: out = 16'(691);
			11194: out = 16'(0);
			11195: out = 16'(17);
			11196: out = 16'(-579);
			11197: out = 16'(-417);
			11198: out = 16'(205);
			11199: out = 16'(133);
			11200: out = 16'(43);
			11201: out = 16'(276);
			11202: out = 16'(70);
			11203: out = 16'(-40);
			11204: out = 16'(-480);
			11205: out = 16'(38);
			11206: out = 16'(-523);
			11207: out = 16'(28);
			11208: out = 16'(-121);
			11209: out = 16'(115);
			11210: out = 16'(109);
			11211: out = 16'(532);
			11212: out = 16'(9);
			11213: out = 16'(-104);
			11214: out = 16'(-349);
			11215: out = 16'(-125);
			11216: out = 16'(175);
			11217: out = 16'(75);
			11218: out = 16'(116);
			11219: out = 16'(-762);
			11220: out = 16'(448);
			11221: out = 16'(-861);
			11222: out = 16'(120);
			11223: out = 16'(338);
			11224: out = 16'(-178);
			11225: out = 16'(790);
			11226: out = 16'(-18);
			11227: out = 16'(-650);
			11228: out = 16'(176);
			11229: out = 16'(-548);
			11230: out = 16'(-85);
			11231: out = 16'(-372);
			11232: out = 16'(275);
			11233: out = 16'(465);
			11234: out = 16'(-101);
			11235: out = 16'(-96);
			11236: out = 16'(-562);
			11237: out = 16'(105);
			11238: out = 16'(-207);
			11239: out = 16'(-56);
			11240: out = 16'(404);
			11241: out = 16'(-184);
			11242: out = 16'(-74);
			11243: out = 16'(137);
			11244: out = 16'(577);
			11245: out = 16'(-510);
			11246: out = 16'(-599);
			11247: out = 16'(-19);
			11248: out = 16'(-307);
			11249: out = 16'(6);
			11250: out = 16'(87);
			11251: out = 16'(441);
			11252: out = 16'(104);
			11253: out = 16'(242);
			11254: out = 16'(-692);
			11255: out = 16'(-167);
			11256: out = 16'(-1204);
			11257: out = 16'(63);
			11258: out = 16'(467);
			11259: out = 16'(-380);
			11260: out = 16'(105);
			11261: out = 16'(795);
			11262: out = 16'(-161);
			11263: out = 16'(86);
			11264: out = 16'(-200);
			11265: out = 16'(-23);
			11266: out = 16'(72);
			11267: out = 16'(-53);
			11268: out = 16'(549);
			11269: out = 16'(43);
			11270: out = 16'(-11);
			11271: out = 16'(-636);
			11272: out = 16'(318);
			11273: out = 16'(-579);
			11274: out = 16'(-893);
			11275: out = 16'(503);
			11276: out = 16'(-49);
			11277: out = 16'(263);
			11278: out = 16'(147);
			11279: out = 16'(449);
			11280: out = 16'(-158);
			11281: out = 16'(78);
			11282: out = 16'(317);
			11283: out = 16'(-98);
			11284: out = 16'(-95);
			11285: out = 16'(-78);
			11286: out = 16'(-82);
			11287: out = 16'(0);
			11288: out = 16'(-277);
			11289: out = 16'(-204);
			11290: out = 16'(-171);
			11291: out = 16'(-290);
			11292: out = 16'(105);
			11293: out = 16'(487);
			11294: out = 16'(35);
			11295: out = 16'(-52);
			11296: out = 16'(329);
			11297: out = 16'(-625);
			11298: out = 16'(-24);
			11299: out = 16'(-342);
			11300: out = 16'(488);
			11301: out = 16'(73);
			11302: out = 16'(73);
			11303: out = 16'(-64);
			11304: out = 16'(13);
			11305: out = 16'(-608);
			11306: out = 16'(62);
			11307: out = 16'(-54);
			11308: out = 16'(-272);
			11309: out = 16'(-348);
			11310: out = 16'(642);
			11311: out = 16'(242);
			11312: out = 16'(197);
			11313: out = 16'(-468);
			11314: out = 16'(208);
			11315: out = 16'(-474);
			11316: out = 16'(59);
			11317: out = 16'(345);
			11318: out = 16'(-128);
			11319: out = 16'(97);
			11320: out = 16'(-363);
			11321: out = 16'(544);
			11322: out = 16'(28);
			11323: out = 16'(-232);
			11324: out = 16'(-146);
			11325: out = 16'(-194);
			11326: out = 16'(-467);
			11327: out = 16'(327);
			11328: out = 16'(593);
			11329: out = 16'(-65);
			11330: out = 16'(-609);
			11331: out = 16'(610);
			11332: out = 16'(-307);
			11333: out = 16'(95);
			11334: out = 16'(47);
			11335: out = 16'(258);
			11336: out = 16'(-532);
			11337: out = 16'(-59);
			11338: out = 16'(473);
			11339: out = 16'(-76);
			11340: out = 16'(-209);
			11341: out = 16'(-234);
			11342: out = 16'(104);
			11343: out = 16'(2);
			11344: out = 16'(-99);
			11345: out = 16'(587);
			11346: out = 16'(0);
			11347: out = 16'(-616);
			11348: out = 16'(-372);
			11349: out = 16'(426);
			11350: out = 16'(-34);
			11351: out = 16'(-265);
			11352: out = 16'(515);
			11353: out = 16'(-176);
			11354: out = 16'(-393);
			11355: out = 16'(-159);
			11356: out = 16'(326);
			11357: out = 16'(-192);
			11358: out = 16'(-554);
			11359: out = 16'(149);
			11360: out = 16'(93);
			11361: out = 16'(28);
			11362: out = 16'(123);
			11363: out = 16'(212);
			11364: out = 16'(-261);
			11365: out = 16'(-455);
			11366: out = 16'(62);
			11367: out = 16'(8);
			11368: out = 16'(312);
			11369: out = 16'(-98);
			11370: out = 16'(-33);
			11371: out = 16'(418);
			11372: out = 16'(-381);
			11373: out = 16'(13);
			11374: out = 16'(-552);
			11375: out = 16'(-582);
			11376: out = 16'(-218);
			11377: out = 16'(274);
			11378: out = 16'(566);
			11379: out = 16'(-127);
			11380: out = 16'(789);
			11381: out = 16'(-663);
			11382: out = 16'(213);
			11383: out = 16'(-382);
			11384: out = 16'(85);
			11385: out = 16'(-171);
			11386: out = 16'(53);
			11387: out = 16'(262);
			11388: out = 16'(300);
			11389: out = 16'(0);
			11390: out = 16'(-248);
			11391: out = 16'(-368);
			11392: out = 16'(-316);
			11393: out = 16'(-102);
			11394: out = 16'(-405);
			11395: out = 16'(237);
			11396: out = 16'(106);
			11397: out = 16'(117);
			11398: out = 16'(7);
			11399: out = 16'(-138);
			11400: out = 16'(-412);
			11401: out = 16'(167);
			11402: out = 16'(-46);
			11403: out = 16'(-60);
			11404: out = 16'(-320);
			11405: out = 16'(-22);
			11406: out = 16'(340);
			11407: out = 16'(-144);
			11408: out = 16'(-65);
			11409: out = 16'(-56);
			11410: out = 16'(-420);
			11411: out = 16'(55);
			11412: out = 16'(-43);
			11413: out = 16'(-94);
			11414: out = 16'(-242);
			11415: out = 16'(376);
			11416: out = 16'(-165);
			11417: out = 16'(-58);
			11418: out = 16'(39);
			11419: out = 16'(-10);
			11420: out = 16'(186);
			11421: out = 16'(-66);
			11422: out = 16'(-133);
			11423: out = 16'(12);
			11424: out = 16'(-255);
			11425: out = 16'(-50);
			11426: out = 16'(-16);
			11427: out = 16'(-40);
			11428: out = 16'(-59);
			11429: out = 16'(-143);
			11430: out = 16'(39);
			11431: out = 16'(-264);
			11432: out = 16'(-8);
			11433: out = 16'(-450);
			11434: out = 16'(-8);
			11435: out = 16'(89);
			11436: out = 16'(104);
			11437: out = 16'(-3);
			11438: out = 16'(299);
			11439: out = 16'(130);
			11440: out = 16'(28);
			11441: out = 16'(-46);
			11442: out = 16'(-62);
			11443: out = 16'(-343);
			11444: out = 16'(134);
			11445: out = 16'(72);
			11446: out = 16'(-149);
			11447: out = 16'(59);
			11448: out = 16'(-181);
			11449: out = 16'(-168);
			11450: out = 16'(-200);
			11451: out = 16'(-49);
			11452: out = 16'(-88);
			11453: out = 16'(-38);
			11454: out = 16'(-267);
			11455: out = 16'(-34);
			11456: out = 16'(448);
			11457: out = 16'(-236);
			11458: out = 16'(13);
			11459: out = 16'(0);
			11460: out = 16'(-93);
			11461: out = 16'(81);
			11462: out = 16'(-62);
			11463: out = 16'(17);
			11464: out = 16'(-83);
			11465: out = 16'(-90);
			11466: out = 16'(51);
			11467: out = 16'(431);
			11468: out = 16'(-132);
			11469: out = 16'(-274);
			11470: out = 16'(151);
			11471: out = 16'(-527);
			11472: out = 16'(-406);
			11473: out = 16'(50);
			11474: out = 16'(-40);
			11475: out = 16'(-322);
			11476: out = 16'(-82);
			11477: out = 16'(303);
			11478: out = 16'(-140);
			11479: out = 16'(469);
			11480: out = 16'(60);
			11481: out = 16'(-9);
			11482: out = 16'(-436);
			11483: out = 16'(33);
			11484: out = 16'(234);
			11485: out = 16'(33);
			11486: out = 16'(-551);
			11487: out = 16'(248);
			11488: out = 16'(198);
			11489: out = 16'(-260);
			11490: out = 16'(-179);
			11491: out = 16'(39);
			11492: out = 16'(-652);
			11493: out = 16'(-59);
			11494: out = 16'(333);
			11495: out = 16'(-29);
			11496: out = 16'(506);
			11497: out = 16'(52);
			11498: out = 16'(81);
			11499: out = 16'(-550);
			11500: out = 16'(-172);
			11501: out = 16'(-38);
			11502: out = 16'(171);
			11503: out = 16'(-145);
			11504: out = 16'(-154);
			11505: out = 16'(267);
			11506: out = 16'(220);
			11507: out = 16'(12);
			11508: out = 16'(-75);
			11509: out = 16'(-277);
			11510: out = 16'(-598);
			11511: out = 16'(-43);
			11512: out = 16'(597);
			11513: out = 16'(40);
			11514: out = 16'(-105);
			11515: out = 16'(102);
			11516: out = 16'(493);
			11517: out = 16'(-93);
			11518: out = 16'(-115);
			11519: out = 16'(-150);
			11520: out = 16'(-473);
			11521: out = 16'(-143);
			11522: out = 16'(147);
			11523: out = 16'(111);
			11524: out = 16'(-301);
			11525: out = 16'(-69);
			11526: out = 16'(153);
			11527: out = 16'(-293);
			11528: out = 16'(-126);
			11529: out = 16'(304);
			11530: out = 16'(54);
			11531: out = 16'(34);
			11532: out = 16'(27);
			11533: out = 16'(152);
			11534: out = 16'(-231);
			11535: out = 16'(-5);
			11536: out = 16'(-56);
			11537: out = 16'(-106);
			11538: out = 16'(-364);
			11539: out = 16'(89);
			11540: out = 16'(543);
			11541: out = 16'(-111);
			11542: out = 16'(-375);
			11543: out = 16'(358);
			11544: out = 16'(-124);
			11545: out = 16'(-160);
			11546: out = 16'(166);
			11547: out = 16'(63);
			11548: out = 16'(-465);
			11549: out = 16'(-300);
			11550: out = 16'(217);
			11551: out = 16'(-79);
			11552: out = 16'(-73);
			11553: out = 16'(-362);
			11554: out = 16'(495);
			11555: out = 16'(-2);
			11556: out = 16'(-442);
			11557: out = 16'(203);
			11558: out = 16'(383);
			11559: out = 16'(21);
			11560: out = 16'(-275);
			11561: out = 16'(504);
			11562: out = 16'(-463);
			11563: out = 16'(-89);
			11564: out = 16'(78);
			11565: out = 16'(419);
			11566: out = 16'(-22);
			11567: out = 16'(-68);
			11568: out = 16'(-8);
			11569: out = 16'(-237);
			11570: out = 16'(-150);
			11571: out = 16'(80);
			11572: out = 16'(188);
			11573: out = 16'(-228);
			11574: out = 16'(241);
			11575: out = 16'(275);
			11576: out = 16'(-419);
			11577: out = 16'(-522);
			11578: out = 16'(247);
			11579: out = 16'(-409);
			11580: out = 16'(72);
			11581: out = 16'(-72);
			11582: out = 16'(69);
			11583: out = 16'(193);
			11584: out = 16'(105);
			11585: out = 16'(351);
			11586: out = 16'(-29);
			11587: out = 16'(-282);
			11588: out = 16'(-73);
			11589: out = 16'(-111);
			11590: out = 16'(-76);
			11591: out = 16'(-639);
			11592: out = 16'(358);
			11593: out = 16'(307);
			11594: out = 16'(-403);
			11595: out = 16'(159);
			11596: out = 16'(-74);
			11597: out = 16'(6);
			11598: out = 16'(-74);
			11599: out = 16'(132);
			11600: out = 16'(-22);
			11601: out = 16'(58);
			11602: out = 16'(116);
			11603: out = 16'(-93);
			11604: out = 16'(-62);
			11605: out = 16'(-368);
			11606: out = 16'(34);
			11607: out = 16'(29);
			11608: out = 16'(-485);
			11609: out = 16'(-425);
			11610: out = 16'(161);
			11611: out = 16'(-25);
			11612: out = 16'(-11);
			11613: out = 16'(479);
			11614: out = 16'(15);
			11615: out = 16'(8);
			11616: out = 16'(-217);
			11617: out = 16'(165);
			11618: out = 16'(12);
			11619: out = 16'(-442);
			11620: out = 16'(388);
			11621: out = 16'(13);
			11622: out = 16'(-73);
			11623: out = 16'(-54);
			11624: out = 16'(327);
			11625: out = 16'(75);
			11626: out = 16'(-458);
			11627: out = 16'(-12);
			11628: out = 16'(-62);
			11629: out = 16'(-446);
			11630: out = 16'(219);
			11631: out = 16'(75);
			11632: out = 16'(-8);
			11633: out = 16'(-289);
			11634: out = 16'(447);
			11635: out = 16'(-126);
			11636: out = 16'(-210);
			11637: out = 16'(-30);
			11638: out = 16'(-682);
			11639: out = 16'(232);
			11640: out = 16'(-273);
			11641: out = 16'(151);
			11642: out = 16'(371);
			11643: out = 16'(-291);
			11644: out = 16'(-321);
			11645: out = 16'(271);
			11646: out = 16'(29);
			11647: out = 16'(-171);
			11648: out = 16'(-61);
			11649: out = 16'(-174);
			11650: out = 16'(44);
			11651: out = 16'(245);
			11652: out = 16'(-21);
			11653: out = 16'(-75);
			11654: out = 16'(-195);
			11655: out = 16'(-111);
			11656: out = 16'(68);
			11657: out = 16'(-6);
			11658: out = 16'(9);
			11659: out = 16'(-186);
			11660: out = 16'(107);
			11661: out = 16'(-156);
			11662: out = 16'(306);
			11663: out = 16'(122);
			11664: out = 16'(-43);
			11665: out = 16'(-192);
			11666: out = 16'(-110);
			11667: out = 16'(-256);
			11668: out = 16'(0);
			11669: out = 16'(197);
			11670: out = 16'(-70);
			11671: out = 16'(14);
			11672: out = 16'(-45);
			11673: out = 16'(-336);
			11674: out = 16'(190);
			11675: out = 16'(169);
			11676: out = 16'(-490);
			11677: out = 16'(-1);
			11678: out = 16'(-156);
			11679: out = 16'(321);
			11680: out = 16'(17);
			11681: out = 16'(-131);
			11682: out = 16'(-185);
			11683: out = 16'(41);
			11684: out = 16'(-20);
			11685: out = 16'(10);
			11686: out = 16'(-54);
			11687: out = 16'(-364);
			11688: out = 16'(71);
			11689: out = 16'(173);
			11690: out = 16'(88);
			11691: out = 16'(-265);
			11692: out = 16'(-1);
			11693: out = 16'(-21);
			11694: out = 16'(67);
			11695: out = 16'(-158);
			11696: out = 16'(-36);
			11697: out = 16'(14);
			11698: out = 16'(-35);
			11699: out = 16'(-31);
			11700: out = 16'(9);
			11701: out = 16'(-32);
			11702: out = 16'(46);
			11703: out = 16'(1);
			11704: out = 16'(-69);
			11705: out = 16'(-153);
			11706: out = 16'(-133);
			11707: out = 16'(-49);
			11708: out = 16'(-52);
			11709: out = 16'(-28);
			11710: out = 16'(-76);
			11711: out = 16'(68);
			11712: out = 16'(-38);
			11713: out = 16'(-86);
			11714: out = 16'(-94);
			11715: out = 16'(124);
			11716: out = 16'(-21);
			11717: out = 16'(20);
			11718: out = 16'(23);
			11719: out = 16'(-57);
			11720: out = 16'(-92);
			11721: out = 16'(-21);
			11722: out = 16'(18);
			11723: out = 16'(-116);
			11724: out = 16'(57);
			11725: out = 16'(-174);
			11726: out = 16'(-288);
			11727: out = 16'(39);
			11728: out = 16'(-312);
			11729: out = 16'(-17);
			11730: out = 16'(52);
			11731: out = 16'(84);
			11732: out = 16'(-67);
			11733: out = 16'(79);
			11734: out = 16'(5);
			11735: out = 16'(5);
			11736: out = 16'(-145);
			11737: out = 16'(-129);
			11738: out = 16'(115);
			11739: out = 16'(-331);
			11740: out = 16'(-78);
			11741: out = 16'(3);
			11742: out = 16'(122);
			11743: out = 16'(-269);
			11744: out = 16'(-22);
			11745: out = 16'(71);
			11746: out = 16'(-175);
			11747: out = 16'(-151);
			11748: out = 16'(255);
			11749: out = 16'(-82);
			11750: out = 16'(-78);
			11751: out = 16'(-116);
			11752: out = 16'(244);
			11753: out = 16'(-74);
			11754: out = 16'(-373);
			11755: out = 16'(-265);
			11756: out = 16'(17);
			11757: out = 16'(78);
			11758: out = 16'(-164);
			11759: out = 16'(349);
			11760: out = 16'(133);
			11761: out = 16'(-8);
			11762: out = 16'(4);
			11763: out = 16'(-228);
			11764: out = 16'(-264);
			11765: out = 16'(-431);
			11766: out = 16'(51);
			11767: out = 16'(306);
			11768: out = 16'(-249);
			11769: out = 16'(-93);
			11770: out = 16'(170);
			11771: out = 16'(-44);
			11772: out = 16'(-137);
			11773: out = 16'(13);
			11774: out = 16'(-21);
			11775: out = 16'(12);
			11776: out = 16'(-12);
			11777: out = 16'(-28);
			11778: out = 16'(-50);
			11779: out = 16'(-22);
			11780: out = 16'(431);
			11781: out = 16'(-226);
			11782: out = 16'(-425);
			11783: out = 16'(-237);
			11784: out = 16'(-24);
			11785: out = 16'(143);
			11786: out = 16'(-103);
			11787: out = 16'(288);
			11788: out = 16'(-163);
			11789: out = 16'(30);
			11790: out = 16'(-31);
			11791: out = 16'(-175);
			11792: out = 16'(-158);
			11793: out = 16'(-184);
			11794: out = 16'(43);
			11795: out = 16'(-21);
			11796: out = 16'(-70);
			11797: out = 16'(247);
			11798: out = 16'(-4);
			11799: out = 16'(291);
			11800: out = 16'(-361);
			11801: out = 16'(-24);
			11802: out = 16'(110);
			11803: out = 16'(22);
			11804: out = 16'(10);
			11805: out = 16'(-9);
			11806: out = 16'(-358);
			11807: out = 16'(-75);
			11808: out = 16'(81);
			11809: out = 16'(35);
			11810: out = 16'(-130);
			11811: out = 16'(-26);
			11812: out = 16'(59);
			11813: out = 16'(124);
			11814: out = 16'(0);
			11815: out = 16'(4);
			11816: out = 16'(-247);
			11817: out = 16'(-389);
			11818: out = 16'(190);
			11819: out = 16'(-51);
			11820: out = 16'(206);
			11821: out = 16'(-430);
			11822: out = 16'(257);
			11823: out = 16'(-213);
			11824: out = 16'(-66);
			11825: out = 16'(-176);
			11826: out = 16'(-54);
			11827: out = 16'(-313);
			11828: out = 16'(-225);
			11829: out = 16'(567);
			11830: out = 16'(58);
			11831: out = 16'(-257);
			11832: out = 16'(128);
			11833: out = 16'(-404);
			11834: out = 16'(14);
			11835: out = 16'(9);
			11836: out = 16'(200);
			11837: out = 16'(252);
			11838: out = 16'(-128);
			11839: out = 16'(66);
			11840: out = 16'(7);
			11841: out = 16'(-169);
			11842: out = 16'(-336);
			11843: out = 16'(-43);
			11844: out = 16'(-69);
			11845: out = 16'(-203);
			11846: out = 16'(26);
			11847: out = 16'(129);
			11848: out = 16'(48);
			11849: out = 16'(-60);
			11850: out = 16'(-31);
			11851: out = 16'(121);
			11852: out = 16'(-120);
			11853: out = 16'(-53);
			11854: out = 16'(176);
			11855: out = 16'(-102);
			11856: out = 16'(-146);
			11857: out = 16'(121);
			11858: out = 16'(203);
			11859: out = 16'(-309);
			11860: out = 16'(-368);
			11861: out = 16'(80);
			11862: out = 16'(-62);
			11863: out = 16'(-173);
			11864: out = 16'(238);
			11865: out = 16'(-140);
			11866: out = 16'(-92);
			11867: out = 16'(113);
			11868: out = 16'(-123);
			11869: out = 16'(67);
			11870: out = 16'(-354);
			11871: out = 16'(-11);
			11872: out = 16'(0);
			11873: out = 16'(-203);
			11874: out = 16'(-22);
			11875: out = 16'(82);
			11876: out = 16'(-36);
			11877: out = 16'(96);
			11878: out = 16'(-70);
			11879: out = 16'(43);
			11880: out = 16'(-101);
			11881: out = 16'(47);
			11882: out = 16'(-41);
			11883: out = 16'(-138);
			11884: out = 16'(7);
			11885: out = 16'(-165);
			11886: out = 16'(9);
			11887: out = 16'(-199);
			11888: out = 16'(16);
			11889: out = 16'(38);
			11890: out = 16'(-25);
			11891: out = 16'(-195);
			11892: out = 16'(-38);
			11893: out = 16'(29);
			11894: out = 16'(-61);
			11895: out = 16'(-47);
			11896: out = 16'(65);
			11897: out = 16'(-39);
			11898: out = 16'(-1);
			11899: out = 16'(46);
			11900: out = 16'(-74);
			11901: out = 16'(-245);
			11902: out = 16'(-95);
			11903: out = 16'(2);
			11904: out = 16'(135);
			11905: out = 16'(-67);
			11906: out = 16'(-61);
			11907: out = 16'(227);
			11908: out = 16'(-22);
			11909: out = 16'(-236);
			11910: out = 16'(-49);
			11911: out = 16'(-178);
			11912: out = 16'(-49);
			11913: out = 16'(6);
			11914: out = 16'(232);
			11915: out = 16'(-216);
			11916: out = 16'(-27);
			11917: out = 16'(75);
			11918: out = 16'(-205);
			11919: out = 16'(-28);
			11920: out = 16'(-120);
			11921: out = 16'(10);
			11922: out = 16'(-134);
			11923: out = 16'(-70);
			11924: out = 16'(-59);
			11925: out = 16'(71);
			11926: out = 16'(-255);
			11927: out = 16'(-57);
			11928: out = 16'(21);
			11929: out = 16'(-18);
			11930: out = 16'(-170);
			11931: out = 16'(119);
			11932: out = 16'(-39);
			11933: out = 16'(-78);
			11934: out = 16'(-16);
			11935: out = 16'(-41);
			11936: out = 16'(0);
			11937: out = 16'(-54);
			11938: out = 16'(162);
			11939: out = 16'(-26);
			11940: out = 16'(-62);
			11941: out = 16'(-162);
			11942: out = 16'(46);
			11943: out = 16'(-74);
			11944: out = 16'(-93);
			11945: out = 16'(18);
			11946: out = 16'(-8);
			11947: out = 16'(110);
			11948: out = 16'(-45);
			11949: out = 16'(-60);
			11950: out = 16'(-339);
			11951: out = 16'(-122);
			11952: out = 16'(6);
			11953: out = 16'(45);
			11954: out = 16'(217);
			11955: out = 16'(-112);
			11956: out = 16'(-149);
			11957: out = 16'(-14);
			11958: out = 16'(-41);
			11959: out = 16'(-127);
			11960: out = 16'(-121);
			11961: out = 16'(-90);
			11962: out = 16'(35);
			11963: out = 16'(49);
			11964: out = 16'(13);
			11965: out = 16'(-26);
			11966: out = 16'(92);
			11967: out = 16'(-16);
			11968: out = 16'(28);
			11969: out = 16'(-21);
			11970: out = 16'(-130);
			11971: out = 16'(9);
			11972: out = 16'(-9);
			11973: out = 16'(-65);
			11974: out = 16'(-45);
			11975: out = 16'(0);
			11976: out = 16'(-127);
			11977: out = 16'(-13);
			11978: out = 16'(-47);
			11979: out = 16'(-277);
			11980: out = 16'(122);
			11981: out = 16'(-23);
			11982: out = 16'(24);
			11983: out = 16'(-164);
			11984: out = 16'(-26);
			11985: out = 16'(6);
			11986: out = 16'(-65);
			11987: out = 16'(113);
			11988: out = 16'(-206);
			11989: out = 16'(12);
			11990: out = 16'(-122);
			11991: out = 16'(0);
			11992: out = 16'(-21);
			11993: out = 16'(31);
			11994: out = 16'(-8);
			11995: out = 16'(-52);
			11996: out = 16'(-39);
			11997: out = 16'(19);
			11998: out = 16'(20);
			11999: out = 16'(-48);
			12000: out = 16'(-110);
			12001: out = 16'(-160);
			12002: out = 16'(-47);
			12003: out = 16'(-19);
			12004: out = 16'(10);
			12005: out = 16'(-4);
			12006: out = 16'(-41);
			12007: out = 16'(20);
			12008: out = 16'(3);
			12009: out = 16'(-64);
			12010: out = 16'(-204);
			12011: out = 16'(-254);
			12012: out = 16'(-124);
			12013: out = 16'(40);
			12014: out = 16'(151);
			12015: out = 16'(170);
			12016: out = 16'(-14);
			12017: out = 16'(-12);
			12018: out = 16'(-68);
			12019: out = 16'(-223);
			12020: out = 16'(-188);
			12021: out = 16'(0);
			default: out = 0;
		endcase
	end
endmodule
