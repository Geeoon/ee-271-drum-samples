module open_hihat_lookup(index, out);
	input logic unsigned [9:0] index;
	output logic signed [23:0] out;
	always_comb begin
		case(index)
			0: out = 0;
			1: out = 0;
			2: out = 144;
			3: out = -244;
			4: out = 210;
			5: out = -326;
			6: out = 291;
			7: out = -431;
			8: out = 426;
			9: out = -582;
			10: out = 595;
			11: out = -770;
			12: out = 775;
			13: out = 2225;
			14: out = 8523;
			15: out = -12479;
			16: out = -680;
			17: out = 15705;
			18: out = 19528;
			19: out = -8997;
			20: out = -24513;
			21: out = -8816;
			22: out = 14127;
			23: out = 10488;
			24: out = -7222;
			25: out = 5310;
			26: out = 525;
			27: out = 9793;
			28: out = 16446;
			29: out = -11450;
			30: out = -24617;
			31: out = -14226;
			32: out = 11029;
			33: out = 21315;
			34: out = 13754;
			35: out = -1002;
			36: out = -14513;
			37: out = -15604;
			38: out = -10052;
			39: out = -2247;
			40: out = -7655;
			41: out = -1525;
			42: out = 14399;
			43: out = -2166;
			44: out = -7438;
			45: out = -5980;
			46: out = 9843;
			47: out = 1921;
			48: out = -7514;
			49: out = -15508;
			50: out = 3217;
			51: out = 2884;
			52: out = -4116;
			53: out = -7837;
			54: out = -3803;
			55: out = 2082;
			56: out = 3581;
			57: out = 8398;
			58: out = 3869;
			59: out = -2238;
			60: out = -14156;
			61: out = -3734;
			62: out = -3344;
			63: out = -8963;
			64: out = -13716;
			65: out = -1865;
			66: out = 4451;
			67: out = -10806;
			68: out = -11132;
			69: out = -1465;
			70: out = 13966;
			71: out = -322;
			72: out = -4441;
			73: out = -7656;
			74: out = 989;
			75: out = -15859;
			76: out = -16318;
			77: out = -5347;
			78: out = 1880;
			79: out = -711;
			80: out = -4714;
			81: out = 2012;
			82: out = -2613;
			83: out = 516;
			84: out = 898;
			85: out = -2792;
			86: out = -16034;
			87: out = -16758;
			88: out = 3404;
			89: out = 1942;
			90: out = -830;
			91: out = -3404;
			92: out = 3352;
			93: out = 3873;
			94: out = 180;
			95: out = -6063;
			96: out = -3418;
			97: out = 4549;
			98: out = 9586;
			99: out = 2310;
			100: out = -12889;
			101: out = -17433;
			102: out = 5404;
			103: out = -6684;
			104: out = 4873;
			105: out = 13640;
			106: out = 1862;
			107: out = -6222;
			108: out = -3071;
			109: out = 13889;
			110: out = 9816;
			111: out = 11853;
			112: out = 9156;
			113: out = -5694;
			114: out = 4412;
			115: out = 18913;
			116: out = 25125;
			117: out = 8904;
			118: out = -2777;
			119: out = -9424;
			120: out = -17429;
			121: out = -1126;
			122: out = 9318;
			123: out = 5356;
			124: out = 4691;
			125: out = -6199;
			126: out = -8445;
			127: out = 15252;
			128: out = 4042;
			129: out = 605;
			130: out = 7391;
			131: out = -427;
			132: out = -5393;
			133: out = -7677;
			134: out = 17073;
			135: out = -8940;
			136: out = 70;
			137: out = 30142;
			138: out = 9691;
			139: out = -463;
			140: out = -8951;
			141: out = 914;
			142: out = 6989;
			143: out = 19954;
			144: out = 18295;
			145: out = -25077;
			146: out = -25669;
			147: out = -9276;
			148: out = -4335;
			149: out = 23088;
			150: out = 24511;
			151: out = 7871;
			152: out = -3027;
			153: out = -8884;
			154: out = -3329;
			155: out = -937;
			156: out = 16170;
			157: out = 4183;
			158: out = -12559;
			159: out = 29156;
			160: out = 14447;
			161: out = -5428;
			162: out = -10567;
			163: out = -27476;
			164: out = -20155;
			165: out = 4551;
			166: out = 28189;
			167: out = 20665;
			168: out = 710;
			169: out = -25496;
			170: out = -3945;
			171: out = 4306;
			172: out = -38;
			173: out = 1855;
			174: out = -6485;
			175: out = -9121;
			176: out = 4186;
			177: out = -28043;
			178: out = -9423;
			179: out = 27601;
			180: out = 7281;
			181: out = -12089;
			182: out = -30632;
			183: out = -16910;
			184: out = -19716;
			185: out = 767;
			186: out = 11660;
			187: out = 2517;
			188: out = -17731;
			189: out = -22795;
			190: out = -3766;
			191: out = -9942;
			192: out = -16072;
			193: out = -15642;
			194: out = 21450;
			195: out = 9725;
			196: out = 3013;
			197: out = 8726;
			198: out = 1227;
			199: out = -735;
			200: out = 1801;
			201: out = 26909;
			202: out = -14386;
			203: out = -26776;
			204: out = 7567;
			205: out = -6406;
			206: out = 5432;
			207: out = 14426;
			208: out = -6729;
			209: out = 5168;
			210: out = 8558;
			211: out = 2483;
			212: out = 577;
			213: out = 4785;
			214: out = 5339;
			215: out = -26464;
			216: out = -6227;
			217: out = -3436;
			218: out = -22900;
			219: out = 17014;
			220: out = 29435;
			221: out = 24575;
			222: out = -25104;
			223: out = -916;
			224: out = 8913;
			225: out = 2105;
			226: out = -8870;
			227: out = 12388;
			228: out = 24668;
			229: out = -15352;
			230: out = -5715;
			231: out = 2493;
			232: out = 10903;
			233: out = -9974;
			234: out = -2345;
			235: out = 7696;
			236: out = -4099;
			237: out = 10804;
			238: out = 8176;
			239: out = -3903;
			240: out = -28925;
			241: out = -18916;
			242: out = 2904;
			243: out = 25549;
			244: out = -16457;
			245: out = -19152;
			246: out = 8231;
			247: out = 13630;
			248: out = -7727;
			249: out = -14540;
			250: out = 31144;
			251: out = 10536;
			252: out = -10172;
			253: out = -29000;
			254: out = 15084;
			255: out = 21370;
			256: out = 18398;
			257: out = 10134;
			258: out = 4793;
			259: out = -2425;
			260: out = -8283;
			261: out = -7034;
			262: out = -11250;
			263: out = -5365;
			264: out = 15586;
			265: out = 10436;
			266: out = -1688;
			267: out = -16002;
			268: out = 12797;
			269: out = 1491;
			270: out = -7961;
			271: out = -15199;
			272: out = -7303;
			273: out = -17277;
			274: out = -28429;
			275: out = -13195;
			276: out = 7744;
			277: out = 24222;
			278: out = 28636;
			279: out = -2442;
			280: out = -12778;
			281: out = -1744;
			282: out = 11195;
			283: out = 11400;
			284: out = 1551;
			285: out = -5807;
			286: out = -1834;
			287: out = 5933;
			288: out = 8020;
			289: out = 2548;
			290: out = 1612;
			291: out = -1438;
			292: out = -12665;
			293: out = 680;
			294: out = 3908;
			295: out = 8012;
			296: out = -1501;
			297: out = 10553;
			298: out = -110;
			299: out = -20801;
			300: out = -24511;
			301: out = 9990;
			302: out = 31660;
			303: out = 28480;
			304: out = -5456;
			305: out = -20292;
			306: out = 1251;
			307: out = 16254;
			308: out = 11607;
			309: out = -882;
			310: out = 16100;
			311: out = 1696;
			312: out = 2132;
			313: out = 10329;
			314: out = 814;
			315: out = 3094;
			316: out = -1479;
			317: out = -18869;
			318: out = -30363;
			319: out = -17791;
			320: out = 9800;
			321: out = 11683;
			322: out = -10460;
			323: out = -23467;
			324: out = 16486;
			325: out = 7515;
			326: out = 10595;
			327: out = 15255;
			328: out = -3931;
			329: out = 5384;
			330: out = 13391;
			331: out = -441;
			332: out = 74;
			333: out = -2414;
			334: out = -301;
			335: out = 535;
			336: out = 10295;
			337: out = 13318;
			338: out = -1987;
			339: out = 19133;
			340: out = 11521;
			341: out = -8440;
			342: out = -1089;
			343: out = 10783;
			344: out = 21437;
			345: out = 9430;
			346: out = 12457;
			347: out = -14140;
			348: out = -29852;
			349: out = 14208;
			350: out = 30989;
			351: out = 8516;
			352: out = -27513;
			353: out = -30619;
			354: out = -19290;
			355: out = 3587;
			356: out = 8790;
			357: out = -13125;
			358: out = -28179;
			359: out = -5512;
			360: out = -12426;
			361: out = -2886;
			362: out = 2329;
			363: out = 13718;
			364: out = -15958;
			365: out = -25508;
			366: out = 1140;
			367: out = 10107;
			368: out = 8038;
			369: out = -676;
			370: out = 17528;
			371: out = -5959;
			372: out = -14820;
			373: out = 1228;
			374: out = -342;
			375: out = 5179;
			376: out = 6424;
			377: out = 12914;
			378: out = -18260;
			379: out = -28963;
			380: out = -13523;
			381: out = -1997;
			382: out = -8211;
			383: out = -13616;
			384: out = 25268;
			385: out = 10036;
			386: out = 6384;
			387: out = 9415;
			388: out = -15338;
			389: out = -29123;
			390: out = -25929;
			391: out = -2572;
			392: out = 21207;
			393: out = 20546;
			394: out = 4843;
			395: out = 27847;
			396: out = 16454;
			397: out = 2193;
			398: out = 10016;
			399: out = -12599;
			400: out = -9599;
			401: out = 16756;
			402: out = 691;
			403: out = 4241;
			404: out = 1759;
			405: out = 1351;
			406: out = -19313;
			407: out = -13640;
			408: out = 9228;
			409: out = -7440;
			410: out = -20140;
			411: out = -24074;
			412: out = 6351;
			413: out = 718;
			414: out = 5326;
			415: out = 5142;
			416: out = -24674;
			417: out = -26792;
			418: out = -10385;
			419: out = 4770;
			420: out = 21353;
			421: out = 11539;
			422: out = -10002;
			423: out = 987;
			424: out = -3217;
			425: out = -7694;
			426: out = -10762;
			427: out = 22736;
			428: out = 28842;
			429: out = 15259;
			430: out = 17858;
			431: out = -9939;
			432: out = -26367;
			433: out = -14277;
			434: out = 9383;
			435: out = 14263;
			436: out = 684;
			437: out = 15442;
			438: out = -6092;
			439: out = -10985;
			440: out = 10265;
			441: out = 13200;
			442: out = 13688;
			443: out = 7534;
			444: out = -7898;
			445: out = -5707;
			446: out = -8890;
			447: out = -31477;
			448: out = -6829;
			449: out = 6396;
			450: out = 7874;
			451: out = -29730;
			452: out = 6221;
			453: out = 26803;
			454: out = 1090;
			455: out = 784;
			456: out = -19207;
			457: out = -27963;
			458: out = -1534;
			459: out = 4957;
			460: out = 12328;
			461: out = 27737;
			462: out = 1566;
			463: out = -14958;
			464: out = -18359;
			465: out = 32135;
			466: out = -4186;
			467: out = -15110;
			468: out = 19903;
			469: out = -4798;
			470: out = -501;
			471: out = 5630;
			472: out = 5124;
			473: out = -2186;
			474: out = -9046;
			475: out = -9337;
			476: out = 1451;
			477: out = 18998;
			478: out = 24772;
			479: out = -6887;
			480: out = -807;
			481: out = 7367;
			482: out = 20737;
			483: out = -4222;
			484: out = 12310;
			485: out = 20488;
			486: out = -20799;
			487: out = -13354;
			488: out = 1725;
			489: out = 15313;
			490: out = 2161;
			491: out = -3956;
			492: out = -2630;
			493: out = 7291;
			494: out = 6009;
			495: out = 328;
			496: out = -4205;
			497: out = -27652;
			498: out = -14286;
			499: out = 4322;
			500: out = 4279;
			501: out = -17221;
			502: out = -13784;
			503: out = 19195;
			504: out = -17281;
			505: out = 2751;
			506: out = 14033;
			507: out = -24144;
			508: out = 6235;
			509: out = 11164;
			510: out = -2916;
			511: out = -18196;
			512: out = -3291;
			513: out = 15009;
			514: out = -2280;
			515: out = 10420;
			516: out = -7193;
			517: out = -26994;
			518: out = 14819;
			519: out = 29025;
			520: out = 23886;
			521: out = 676;
			522: out = -1587;
			523: out = -856;
			524: out = 870;
			525: out = -32767;
			526: out = -6603;
			527: out = 24881;
			528: out = 26057;
			529: out = -18212;
			530: out = -25551;
			531: out = -1431;
			532: out = 1512;
			533: out = -6699;
			534: out = -4488;
			535: out = 32320;
			536: out = 4963;
			537: out = 2350;
			538: out = 2803;
			539: out = 18451;
			540: out = 913;
			541: out = -10027;
			542: out = -14204;
			543: out = 19579;
			544: out = -1094;
			545: out = -31866;
			546: out = 23344;
			547: out = 5734;
			548: out = -12028;
			549: out = -9436;
			550: out = -11056;
			551: out = 12692;
			552: out = 21427;
			553: out = -27972;
			554: out = -25484;
			555: out = -14198;
			556: out = 5095;
			557: out = 6931;
			558: out = 8742;
			559: out = 6672;
			560: out = 32173;
			561: out = -11679;
			562: out = -24912;
			563: out = 4891;
			564: out = 28374;
			565: out = 18292;
			566: out = -5551;
			567: out = -7059;
			568: out = -15415;
			569: out = -19;
			570: out = 28535;
			571: out = -10310;
			572: out = -5522;
			573: out = 6873;
			574: out = 15833;
			575: out = -7707;
			576: out = -12471;
			577: out = 2987;
			578: out = 14848;
			579: out = -10177;
			580: out = -26122;
			581: out = 25978;
			582: out = 13056;
			583: out = -3502;
			584: out = -23193;
			585: out = 8850;
			586: out = 1565;
			587: out = -8747;
			588: out = 14769;
			589: out = -16881;
			590: out = -4594;
			591: out = 29742;
			592: out = -7209;
			593: out = -4575;
			594: out = 966;
			595: out = -11136;
			596: out = 20223;
			597: out = 8794;
			598: out = -27572;
			599: out = -25407;
			600: out = -4583;
			601: out = 15726;
			602: out = -7488;
			603: out = 28861;
			604: out = 14177;
			605: out = -16438;
			606: out = -11901;
			607: out = -9185;
			608: out = -7334;
			609: out = -8663;
			610: out = -7996;
			611: out = 2000;
			612: out = 12918;
			613: out = 2343;
			614: out = 1868;
			615: out = 9211;
			616: out = 29059;
			617: out = 5021;
			618: out = -3438;
			619: out = -3869;
			620: out = 9338;
			621: out = 725;
			622: out = -8267;
			623: out = -10886;
			624: out = 3394;
			625: out = 13501;
			626: out = 13553;
			627: out = -13051;
			628: out = -7337;
			629: out = -8458;
			630: out = -28594;
			631: out = -22572;
			632: out = -9398;
			633: out = 7134;
			634: out = -3187;
			635: out = 890;
			636: out = 2267;
			637: out = 14302;
			638: out = -22220;
			639: out = -7116;
			640: out = 22873;
			641: out = 20975;
			642: out = -12832;
			643: out = -31058;
			644: out = -3467;
			645: out = -26485;
			646: out = -2706;
			647: out = 23595;
			648: out = -148;
			649: out = 7301;
			650: out = 4530;
			651: out = 2525;
			652: out = 951;
			653: out = 16158;
			654: out = 19032;
			655: out = -15773;
			656: out = -8225;
			657: out = 16371;
			658: out = 30830;
			659: out = 12095;
			660: out = -6423;
			661: out = -12431;
			662: out = -8870;
			663: out = 11425;
			664: out = 1917;
			665: out = -29622;
			666: out = -28832;
			667: out = -17281;
			668: out = 6747;
			669: out = 25683;
			670: out = 10067;
			671: out = 4749;
			672: out = 15440;
			673: out = 4817;
			674: out = -3343;
			675: out = -9128;
			676: out = 13573;
			677: out = -8104;
			678: out = -20900;
			679: out = -24267;
			680: out = 18141;
			681: out = 21532;
			682: out = 14778;
			683: out = 7944;
			684: out = 4901;
			685: out = -9741;
			686: out = -28078;
			687: out = -3464;
			688: out = 11765;
			689: out = 11988;
			690: out = -18456;
			691: out = -4141;
			692: out = 11811;
			693: out = 28429;
			694: out = -13184;
			695: out = 9061;
			696: out = 14070;
			697: out = -26107;
			698: out = -30612;
			699: out = -19332;
			700: out = 14921;
			701: out = 6610;
			702: out = -2169;
			703: out = -14753;
			704: out = -17025;
			705: out = 15884;
			706: out = 32766;
			707: out = 21870;
			708: out = -20857;
			709: out = -28447;
			710: out = -9582;
			711: out = 10695;
			712: out = 29888;
			713: out = 18731;
			714: out = -8585;
			715: out = -30301;
			716: out = -17411;
			717: out = 8842;
			718: out = 17602;
			719: out = -13389;
			720: out = -31351;
			721: out = -25810;
			722: out = -14221;
			723: out = 16407;
			724: out = 28195;
			725: out = 21412;
			726: out = 7142;
			727: out = -2117;
			728: out = -4414;
			729: out = -10600;
			730: out = -8999;
			731: out = -2979;
			732: out = 12041;
			733: out = -14872;
			734: out = -10715;
			735: out = 3918;
			736: out = 2804;
			737: out = 4328;
			738: out = -85;
			739: out = -9518;
			740: out = 16826;
			741: out = 10035;
			742: out = -8730;
			743: out = -21937;
			744: out = -1995;
			745: out = 17038;
			746: out = 11836;
			747: out = 11040;
			748: out = -172;
			749: out = 6400;
			750: out = 29042;
			751: out = 23889;
			752: out = -1553;
			753: out = -30159;
			754: out = -9279;
			755: out = 18104;
			756: out = 29449;
			757: out = 12010;
			758: out = 1619;
			759: out = -7860;
			760: out = -1254;
			761: out = -23944;
			762: out = 4225;
			763: out = 21889;
			764: out = -12404;
			765: out = -11976;
			766: out = 523;
			767: out = 25210;
			768: out = -2375;
			769: out = 468;
			770: out = 1188;
			771: out = 4834;
			772: out = -7274;
			773: out = -5895;
			774: out = 171;
			775: out = 9939;
			776: out = -14352;
			777: out = -30620;
			778: out = -13222;
			779: out = 2397;
			780: out = 13059;
			781: out = 15995;
			782: out = 22998;
			783: out = 16452;
			784: out = -1908;
			785: out = -29083;
			786: out = -15061;
			787: out = 11520;
			788: out = 25263;
			789: out = -2075;
			790: out = -18880;
			791: out = -24879;
			792: out = -2490;
			793: out = 7678;
			794: out = 25883;
			795: out = 24957;
			796: out = -21087;
			797: out = -31682;
			798: out = -25198;
			799: out = 3652;
			800: out = 30659;
			801: out = 13225;
			802: out = -10582;
			803: out = -9782;
			804: out = 12929;
			805: out = 13786;
			806: out = -30279;
			807: out = -1209;
			808: out = 2612;
			809: out = -3004;
			810: out = 273;
			811: out = -2093;
			812: out = 356;
			813: out = 6041;
			814: out = -7086;
			815: out = -9659;
			816: out = -4177;
			817: out = -25201;
			818: out = -522;
			819: out = 12045;
			820: out = 7376;
			821: out = -24788;
			822: out = -11099;
			823: out = 23165;
			824: out = 13273;
			825: out = 13605;
			826: out = 70;
			827: out = -14296;
			828: out = -4246;
			829: out = -4900;
			830: out = -9606;
			831: out = 3968;
			832: out = 3368;
			833: out = 12534;
			834: out = 25200;
			835: out = -2348;
			836: out = -1412;
			837: out = 9716;
			838: out = 13930;
			839: out = 6078;
			840: out = -7941;
			841: out = -18186;
			842: out = 8804;
			843: out = 11727;
			844: out = 2332;
			845: out = -3198;
			846: out = 2663;
			847: out = 11881;
			848: out = 11594;
			849: out = 14470;
			850: out = 571;
			851: out = -16427;
			852: out = -31725;
			853: out = -11871;
			854: out = 15242;
			855: out = 28713;
			856: out = -19816;
			857: out = -2702;
			858: out = 18466;
			859: out = -7732;
			860: out = -6235;
			861: out = -9005;
			862: out = -1727;
			863: out = -24475;
			864: out = -4099;
			865: out = 13398;
			866: out = -318;
			867: out = 6034;
			868: out = -4754;
			869: out = -15788;
			870: out = 1638;
			871: out = 14775;
			872: out = 11471;
			873: out = -20031;
			874: out = -4725;
			875: out = -345;
			876: out = -3431;
			877: out = 13925;
			878: out = 2118;
			879: out = -7804;
			880: out = -4929;
			881: out = 11444;
			882: out = 18714;
			883: out = 8527;
			884: out = -24123;
			885: out = -25594;
			886: out = -10450;
			887: out = -401;
			888: out = 20163;
			889: out = 8064;
			890: out = -15047;
			891: out = 16525;
			892: out = 2125;
			893: out = -2752;
			894: out = 1682;
			895: out = 17652;
			896: out = -1192;
			897: out = -29392;
			898: out = 1963;
			899: out = 2245;
			900: out = 4874;
			901: out = 8720;
			902: out = 19615;
			903: out = 18692;
			904: out = 8776;
			905: out = -4821;
			906: out = -18849;
			907: out = -27288;
			908: out = -27683;
			909: out = 15575;
			910: out = 31027;
			911: out = 18767;
			912: out = -15844;
			913: out = -16895;
			914: out = -3784;
			915: out = 6795;
			916: out = 21236;
			917: out = 20385;
			918: out = 11600;
			919: out = -5819;
			920: out = -20626;
			921: out = -23421;
			922: out = -2444;
			923: out = -26980;
			924: out = -10957;
			925: out = 14713;
			926: out = 28209;
			927: out = 798;
			928: out = -25393;
			929: out = -29028;
			930: out = -360;
			931: out = 21998;
			932: out = 17964;
			933: out = -4700;
			934: out = 8155;
			935: out = 12525;
			936: out = -5523;
			937: out = 4054;
			938: out = -7721;
			939: out = -10278;
			940: out = -3556;
			941: out = 16794;
			942: out = 17645;
			943: out = 3995;
			944: out = -28510;
			945: out = -6770;
			946: out = 23204;
			947: out = -20380;
			948: out = 19292;
			949: out = 18930;
			950: out = -5893;
			951: out = -8511;
			952: out = -12510;
			953: out = -6821;
			954: out = 3591;
			955: out = 5429;
			956: out = -686;
			957: out = -8229;
			958: out = 344;
			959: out = 2646;
			960: out = -1942;
			961: out = -13941;
			962: out = -1798;
			963: out = 12312;
			964: out = 16958;
			965: out = 9906;
			966: out = -3514;
			967: out = -11655;
			968: out = -8239;
			969: out = -2488;
			970: out = 9323;
			971: out = 19357;
			972: out = -27104;
			973: out = -3015;
			974: out = 21782;
			975: out = 12335;
			976: out = 5882;
			977: out = 72;
			978: out = 1472;
			979: out = 1079;
			980: out = -9722;
			981: out = -17789;
			982: out = -6902;
			983: out = 8620;
			984: out = 18748;
			985: out = 14213;
			986: out = 2011;
			987: out = -2208;
			988: out = 3163;
			989: out = 8114;
			990: out = 11581;
			991: out = 421;
			992: out = -11210;
			993: out = 6519;
			994: out = 6876;
			995: out = 2504;
			996: out = -12784;
			997: out = 7867;
			998: out = 2778;
			999: out = -8611;
			1000: out = -3384;
			1001: out = -389;
			1002: out = 1324;
			1003: out = -101;
			1004: out = -20597;
			1005: out = -15147;
			1006: out = 3643;
			1007: out = -8797;
			1008: out = 4142;
			1009: out = 9596;
			1010: out = 13231;
			1011: out = -21918;
			1012: out = -29415;
			1013: out = -28555;
			1014: out = 10717;
			1015: out = 19022;
			1016: out = 20647;
			1017: out = 24290;
			1018: out = 183;
			1019: out = -13283;
			1020: out = -14210;
			1021: out = 986;
			1022: out = 17654;
			1023: out = 20124;
			1024: out = 10004;
			1025: out = -6079;
			1026: out = -8557;
			1027: out = -4860;
			1028: out = -7222;
			1029: out = -7663;
			1030: out = -572;
			1031: out = 12388;
			1032: out = 13437;
			1033: out = 8299;
			1034: out = -7020;
			1035: out = -30747;
			1036: out = -11660;
			1037: out = 784;
			1038: out = -5436;
			1039: out = 6460;
			1040: out = -5348;
			1041: out = -10324;
			1042: out = 24214;
			1043: out = -18723;
			1044: out = -9815;
			1045: out = 30651;
			1046: out = 13972;
			1047: out = -10710;
			1048: out = -31509;
			1049: out = -1760;
			1050: out = -3436;
			1051: out = 5909;
			1052: out = 4775;
			1053: out = 22582;
			1054: out = -8528;
			1055: out = -23954;
			1056: out = -5904;
			1057: out = 18178;
			1058: out = 13217;
			1059: out = -8517;
			1060: out = -23802;
			1061: out = -2992;
			1062: out = 18359;
			1063: out = 4593;
			1064: out = -530;
			1065: out = -6677;
			1066: out = 2806;
			1067: out = -16778;
			1068: out = 14737;
			1069: out = 21056;
			1070: out = -13028;
			1071: out = -5340;
			1072: out = -14229;
			1073: out = -18503;
			1074: out = 23109;
			1075: out = 14754;
			1076: out = 4204;
			1077: out = 313;
			1078: out = 3038;
			1079: out = 4467;
			1080: out = 4505;
			1081: out = 9168;
			1082: out = 6073;
			1083: out = 224;
			1084: out = -6542;
			1085: out = -1769;
			1086: out = 5383;
			1087: out = 12703;
			1088: out = 18136;
			1089: out = 4201;
			1090: out = -13795;
			1091: out = -25586;
			1092: out = -13637;
			1093: out = -4708;
			1094: out = -6385;
			1095: out = -8880;
			1096: out = -14312;
			1097: out = -11444;
			1098: out = -7679;
			1099: out = 10958;
			1100: out = -847;
			1101: out = -17311;
			1102: out = -8924;
			1103: out = 1357;
			1104: out = 9010;
			1105: out = 5819;
			1106: out = 2039;
			1107: out = 5536;
			1108: out = 12095;
			1109: out = -3292;
			1110: out = 3041;
			1111: out = -5541;
			1112: out = -13980;
			1113: out = 25055;
			1114: out = 25433;
			1115: out = 5237;
			1116: out = -15425;
			1117: out = -32184;
			1118: out = -10292;
			1119: out = 28857;
			1120: out = -2914;
			1121: out = -14528;
			1122: out = -8058;
			1123: out = 24364;
			1124: out = 8984;
			1125: out = -2205;
			1126: out = -172;
			1127: out = -8343;
			1128: out = 14196;
			1129: out = 24769;
			1130: out = 12058;
			1131: out = -20221;
			1132: out = -19114;
			1133: out = 16058;
			1134: out = -533;
			1135: out = -7649;
			1136: out = -7798;
			1137: out = 31439;
			1138: out = 9253;
			1139: out = 14510;
			1140: out = 20352;
			1141: out = 391;
			1142: out = -18096;
			1143: out = -25313;
			1144: out = -12930;
			1145: out = 8995;
			1146: out = 16120;
			1147: out = 5163;
			1148: out = -24592;
			1149: out = -19099;
			1150: out = 3793;
			1151: out = 10588;
			1152: out = 18046;
			1153: out = 1484;
			1154: out = -18270;
			1155: out = -15604;
			1156: out = 4874;
			1157: out = 17383;
			1158: out = -1763;
			1159: out = 5872;
			1160: out = -181;
			1161: out = 813;
			1162: out = -16952;
			1163: out = 13117;
			1164: out = 21946;
			1165: out = 3713;
			1166: out = -21866;
			1167: out = -10994;
			1168: out = 22324;
			1169: out = 12468;
			1170: out = 7652;
			1171: out = -9949;
			1172: out = -20009;
			1173: out = -13735;
			1174: out = -1910;
			1175: out = 3615;
			1176: out = 19388;
			1177: out = 4936;
			1178: out = -13007;
			1179: out = -31775;
			1180: out = 1981;
			1181: out = 11512;
			1182: out = 1524;
			1183: out = -15171;
			1184: out = -7643;
			1185: out = -8627;
			1186: out = -31427;
			1187: out = 14595;
			1188: out = 17710;
			1189: out = -5731;
			1190: out = -27924;
			1191: out = -23495;
			1192: out = 7770;
			1193: out = 31477;
			1194: out = 24627;
			1195: out = 19709;
			1196: out = 8267;
			1197: out = -14754;
			1198: out = -17245;
			1199: out = -2568;
			1200: out = 18802;
			1201: out = -21638;
			1202: out = -28887;
			1203: out = -17875;
			1204: out = 17446;
			1205: out = 5347;
			1206: out = 1117;
			1207: out = 1726;
			1208: out = 20988;
			1209: out = 5991;
			1210: out = -11400;
			1211: out = -20459;
			1212: out = 11212;
			1213: out = 8845;
			1214: out = -29776;
			1215: out = -6479;
			1216: out = 8298;
			1217: out = 27911;
			1218: out = 27454;
			1219: out = 12920;
			1220: out = -11131;
			1221: out = -19244;
			1222: out = -32431;
			1223: out = -10933;
			1224: out = 4944;
			1225: out = 13880;
			1226: out = -17025;
			1227: out = -8446;
			1228: out = 25905;
			1229: out = 24244;
			1230: out = 14604;
			1231: out = -4104;
			1232: out = -26644;
			1233: out = -5513;
			1234: out = 228;
			1235: out = -7847;
			1236: out = -4637;
			1237: out = 17892;
			1238: out = 19084;
			1239: out = -28911;
			1240: out = -25741;
			1241: out = -9260;
			1242: out = 20575;
			1243: out = -11396;
			1244: out = 17658;
			1245: out = 18716;
			1246: out = -25851;
			1247: out = -12655;
			1248: out = -3815;
			1249: out = 8385;
			1250: out = 27039;
			1251: out = 25787;
			1252: out = 13834;
			1253: out = 2469;
			1254: out = -1034;
			1255: out = 9006;
			1256: out = 15756;
			1257: out = 2234;
			1258: out = -8860;
			1259: out = -18817;
			1260: out = -26547;
			1261: out = 11673;
			1262: out = 24358;
			1263: out = 16082;
			1264: out = -12169;
			1265: out = -14340;
			1266: out = -8890;
			1267: out = 2633;
			1268: out = -22301;
			1269: out = -2765;
			1270: out = 25361;
			1271: out = -3731;
			1272: out = 456;
			1273: out = 1149;
			1274: out = 9529;
			1275: out = 12143;
			1276: out = 9708;
			1277: out = -1102;
			1278: out = 9955;
			1279: out = -16560;
			1280: out = -18977;
			1281: out = 3082;
			1282: out = -7854;
			1283: out = -17264;
			1284: out = -15235;
			1285: out = 27427;
			1286: out = 16766;
			1287: out = 11416;
			1288: out = 9123;
			1289: out = -13646;
			1290: out = -22063;
			1291: out = -17851;
			1292: out = -11038;
			1293: out = 8708;
			1294: out = 12065;
			1295: out = -2280;
			1296: out = -9469;
			1297: out = -25192;
			1298: out = -24651;
			1299: out = 5455;
			1300: out = 10682;
			1301: out = -4814;
			1302: out = -30104;
			1303: out = 3184;
			1304: out = 6527;
			1305: out = 3310;
			1306: out = 6217;
			1307: out = 24151;
			1308: out = 18229;
			1309: out = -12181;
			1310: out = 24617;
			1311: out = -5420;
			1312: out = -25509;
			1313: out = -7067;
			1314: out = 5553;
			1315: out = 3068;
			1316: out = -11001;
			1317: out = -18369;
			1318: out = -6181;
			1319: out = 9838;
			1320: out = 11488;
			1321: out = -157;
			1322: out = 2278;
			1323: out = 16550;
			1324: out = -26102;
			1325: out = -11325;
			1326: out = 7613;
			1327: out = 7619;
			1328: out = 1909;
			1329: out = -10052;
			1330: out = -13469;
			1331: out = 6076;
			1332: out = 24865;
			1333: out = 19704;
			1334: out = -22339;
			1335: out = 9392;
			1336: out = 17402;
			1337: out = 13272;
			1338: out = 23961;
			1339: out = 16749;
			1340: out = 3079;
			1341: out = -27170;
			1342: out = 11552;
			1343: out = 20438;
			1344: out = 11222;
			1345: out = -6450;
			1346: out = -11746;
			1347: out = -7852;
			1348: out = 11203;
			1349: out = -9183;
			1350: out = 3147;
			1351: out = 16333;
			1352: out = 8750;
			1353: out = -17285;
			1354: out = -21714;
			1355: out = 9698;
			1356: out = 22023;
			1357: out = 12626;
			1358: out = -6182;
			1359: out = -9780;
			1360: out = 8340;
			1361: out = 14536;
			1362: out = -7540;
			1363: out = -3572;
			1364: out = 0;
			1365: out = 14090;
			1366: out = 27600;
			1367: out = 12151;
			1368: out = -11556;
			1369: out = -27295;
			1370: out = 7182;
			1371: out = 14531;
			1372: out = -2160;
			1373: out = -11426;
			1374: out = -20966;
			1375: out = -12905;
			1376: out = -5740;
			1377: out = 1841;
			1378: out = -11350;
			1379: out = -17452;
			1380: out = -935;
			1381: out = 14901;
			1382: out = 13622;
			1383: out = 28;
			1384: out = -21060;
			1385: out = -14379;
			1386: out = 2677;
			1387: out = -3134;
			1388: out = 1955;
			1389: out = 3823;
			1390: out = 5633;
			1391: out = 1527;
			1392: out = -9653;
			1393: out = -17253;
			1394: out = -7149;
			1395: out = 10699;
			1396: out = 16246;
			1397: out = 2846;
			1398: out = 3897;
			1399: out = -17660;
			1400: out = -25230;
			1401: out = 13714;
			1402: out = -601;
			1403: out = -3502;
			1404: out = 4166;
			1405: out = 17997;
			1406: out = 3745;
			1407: out = -16967;
			1408: out = -17731;
			1409: out = -21859;
			1410: out = -12471;
			1411: out = -1858;
			1412: out = 3550;
			1413: out = 1042;
			1414: out = 3212;
			1415: out = 20739;
			1416: out = -5161;
			1417: out = -6668;
			1418: out = 14398;
			1419: out = 10317;
			1420: out = 16080;
			1421: out = 6293;
			1422: out = -3333;
			1423: out = -16638;
			1424: out = 1292;
			1425: out = 22392;
			1426: out = 14117;
			1427: out = -6282;
			1428: out = -14510;
			1429: out = 6959;
			1430: out = 6581;
			1431: out = -4410;
			1432: out = -21649;
			1433: out = -20116;
			1434: out = 13126;
			1435: out = 28653;
			1436: out = -1742;
			1437: out = 19867;
			1438: out = 10166;
			1439: out = -1641;
			1440: out = -538;
			1441: out = -6091;
			1442: out = -10871;
			1443: out = -4733;
			1444: out = -19150;
			1445: out = -5953;
			1446: out = 16724;
			1447: out = 13492;
			1448: out = 21162;
			1449: out = 13141;
			1450: out = -7112;
			1451: out = 9484;
			1452: out = 5161;
			1453: out = -5542;
			1454: out = 9860;
			1455: out = -5206;
			1456: out = -9890;
			1457: out = -3183;
			1458: out = 20594;
			1459: out = 16218;
			1460: out = 855;
			1461: out = 2413;
			1462: out = -6839;
			1463: out = 800;
			1464: out = 17570;
			1465: out = 2736;
			1466: out = -4422;
			1467: out = -10195;
			1468: out = -4324;
			1469: out = -8436;
			1470: out = 2810;
			1471: out = 20190;
			1472: out = 8311;
			1473: out = -13298;
			1474: out = -30052;
			1475: out = -4535;
			1476: out = -4925;
			1477: out = 3387;
			1478: out = 10901;
			1479: out = 3261;
			1480: out = -2984;
			1481: out = -5857;
			1482: out = -15454;
			1483: out = 12551;
			1484: out = 12265;
			1485: out = -12679;
			1486: out = 14104;
			1487: out = 5030;
			1488: out = -8754;
			1489: out = -26825;
			1490: out = -20745;
			1491: out = -8942;
			1492: out = 2330;
			1493: out = -16475;
			1494: out = -7640;
			1495: out = 5092;
			1496: out = 4887;
			1497: out = 6385;
			1498: out = -7546;
			1499: out = -28644;
			1500: out = -6384;
			1501: out = -6639;
			1502: out = -3375;
			1503: out = 4818;
			1504: out = 18476;
			1505: out = 15830;
			1506: out = 4969;
			1507: out = -17277;
			1508: out = -8015;
			1509: out = 261;
			1510: out = -13761;
			1511: out = -24581;
			1512: out = -18963;
			1513: out = 7341;
			1514: out = 5858;
			1515: out = 17627;
			1516: out = 12998;
			1517: out = 1454;
			1518: out = -7423;
			1519: out = -4595;
			1520: out = 3354;
			1521: out = 17670;
			1522: out = 2431;
			1523: out = -15187;
			1524: out = -23322;
			1525: out = 2932;
			1526: out = 20500;
			1527: out = 18428;
			1528: out = 5712;
			1529: out = -14238;
			1530: out = -18939;
			1531: out = 5185;
			1532: out = -2071;
			1533: out = 4921;
			1534: out = 8111;
			1535: out = 13389;
			1536: out = -6747;
			1537: out = -6132;
			1538: out = 23476;
			1539: out = 29148;
			1540: out = 18313;
			1541: out = -3409;
			1542: out = 9984;
			1543: out = -11240;
			1544: out = -12305;
			1545: out = 6842;
			1546: out = 490;
			1547: out = 1294;
			1548: out = 1943;
			1549: out = 2330;
			1550: out = -4725;
			1551: out = -4957;
			1552: out = 6542;
			1553: out = -11802;
			1554: out = -3264;
			1555: out = 12376;
			1556: out = 11792;
			1557: out = 9624;
			1558: out = -1906;
			1559: out = -11393;
			1560: out = -11872;
			1561: out = 3525;
			1562: out = 17034;
			1563: out = 15294;
			1564: out = 4853;
			1565: out = -3039;
			1566: out = 799;
			1567: out = 6044;
			1568: out = 6177;
			1569: out = -1317;
			1570: out = 1336;
			1571: out = -8160;
			1572: out = -4158;
			1573: out = 749;
			1574: out = 8052;
			1575: out = -15040;
			1576: out = -28945;
			1577: out = -7239;
			1578: out = 5093;
			1579: out = 1735;
			1580: out = -10018;
			1581: out = -8845;
			1582: out = 10654;
			1583: out = 22174;
			1584: out = -512;
			1585: out = 2252;
			1586: out = 1953;
			1587: out = 4901;
			1588: out = -10507;
			1589: out = -10785;
			1590: out = -2112;
			1591: out = 16409;
			1592: out = 7317;
			1593: out = -5189;
			1594: out = -17275;
			1595: out = 7087;
			1596: out = 1003;
			1597: out = -5618;
			1598: out = 7000;
			1599: out = -3103;
			1600: out = -3576;
			1601: out = -3878;
			1602: out = 11070;
			1603: out = -3034;
			1604: out = -14400;
			1605: out = -19766;
			1606: out = 6125;
			1607: out = 9111;
			1608: out = -4465;
			1609: out = -27716;
			1610: out = -17193;
			1611: out = -192;
			1612: out = 6550;
			1613: out = -22261;
			1614: out = -12114;
			1615: out = 22639;
			1616: out = 11030;
			1617: out = 5251;
			1618: out = -3590;
			1619: out = 10916;
			1620: out = -12802;
			1621: out = 627;
			1622: out = 23350;
			1623: out = 16380;
			1624: out = 18119;
			1625: out = 8895;
			1626: out = 852;
			1627: out = -18186;
			1628: out = -2277;
			1629: out = 20502;
			1630: out = 370;
			1631: out = -6369;
			1632: out = -9468;
			1633: out = 7674;
			1634: out = -10648;
			1635: out = -6085;
			1636: out = 1509;
			1637: out = 10953;
			1638: out = 3990;
			1639: out = 4125;
			1640: out = 7673;
			1641: out = 2943;
			1642: out = -13506;
			1643: out = -22976;
			1644: out = 6476;
			1645: out = 18199;
			1646: out = 16348;
			1647: out = -2427;
			1648: out = 16828;
			1649: out = 8279;
			1650: out = -4004;
			1651: out = -13294;
			1652: out = -7630;
			1653: out = 4363;
			1654: out = 12837;
			1655: out = -14400;
			1656: out = -25080;
			1657: out = -15872;
			1658: out = 20214;
			1659: out = 5376;
			1660: out = -9192;
			1661: out = -16258;
			1662: out = 1200;
			1663: out = -2258;
			1664: out = -11255;
			1665: out = 8490;
			1666: out = -10069;
			1667: out = -1898;
			1668: out = 20469;
			1669: out = 19719;
			1670: out = 16362;
			1671: out = 4539;
			1672: out = -21803;
			1673: out = -12410;
			1674: out = -4171;
			1675: out = 36;
			1676: out = -18225;
			1677: out = -8327;
			1678: out = 7209;
			1679: out = 19893;
			1680: out = 1000;
			1681: out = 750;
			1682: out = 11735;
			1683: out = 17955;
			1684: out = -7691;
			1685: out = -30107;
			1686: out = -15466;
			1687: out = -1158;
			1688: out = 9521;
			1689: out = 4042;
			1690: out = -9727;
			1691: out = -14890;
			1692: out = -8553;
			1693: out = 666;
			1694: out = -7019;
			1695: out = -13971;
			1696: out = -14483;
			1697: out = -29;
			1698: out = -2565;
			1699: out = -5031;
			1700: out = 3076;
			1701: out = 2664;
			1702: out = 7439;
			1703: out = 13838;
			1704: out = 21950;
			1705: out = 17339;
			1706: out = 7259;
			1707: out = 360;
			1708: out = -23585;
			1709: out = -17260;
			1710: out = 6744;
			1711: out = 7658;
			1712: out = 6533;
			1713: out = 255;
			1714: out = 4724;
			1715: out = 1787;
			1716: out = 13959;
			1717: out = 17924;
			1718: out = 3169;
			1719: out = -19665;
			1720: out = -19812;
			1721: out = 19960;
			1722: out = -10613;
			1723: out = -2491;
			1724: out = 10793;
			1725: out = 10368;
			1726: out = 9732;
			1727: out = 14209;
			1728: out = 20276;
			1729: out = 5143;
			1730: out = -6643;
			1731: out = -12762;
			1732: out = -18702;
			1733: out = 5126;
			1734: out = 11181;
			1735: out = -6298;
			1736: out = 342;
			1737: out = 4270;
			1738: out = 9810;
			1739: out = -4114;
			1740: out = 5817;
			1741: out = -6679;
			1742: out = -32324;
			1743: out = -2081;
			1744: out = 1106;
			1745: out = -7922;
			1746: out = -7927;
			1747: out = -3554;
			1748: out = 7954;
			1749: out = 14364;
			1750: out = -15086;
			1751: out = -28440;
			1752: out = -22749;
			1753: out = 9637;
			1754: out = 3579;
			1755: out = 6581;
			1756: out = 15651;
			1757: out = -24713;
			1758: out = -15267;
			1759: out = 14481;
			1760: out = 28386;
			1761: out = 23867;
			1762: out = 209;
			1763: out = -28075;
			1764: out = -20168;
			1765: out = -7763;
			1766: out = 2801;
			1767: out = -5824;
			1768: out = 8702;
			1769: out = 13140;
			1770: out = 13698;
			1771: out = -18028;
			1772: out = -9273;
			1773: out = 4687;
			1774: out = 9230;
			1775: out = -2391;
			1776: out = -9490;
			1777: out = -10319;
			1778: out = 12641;
			1779: out = -5693;
			1780: out = -21634;
			1781: out = -11296;
			1782: out = 13076;
			1783: out = 28486;
			1784: out = 25285;
			1785: out = 3168;
			1786: out = 2898;
			1787: out = 7036;
			1788: out = 6440;
			1789: out = -15977;
			1790: out = -16328;
			1791: out = 5604;
			1792: out = -532;
			1793: out = 13310;
			1794: out = 10661;
			1795: out = 3124;
			1796: out = -5569;
			1797: out = 4282;
			1798: out = 15543;
			1799: out = 14560;
			1800: out = 2619;
			1801: out = -6943;
			1802: out = -8834;
			1803: out = 8993;
			1804: out = 10592;
			1805: out = 924;
			1806: out = -17713;
			1807: out = -7991;
			1808: out = 10873;
			1809: out = 24745;
			1810: out = -11287;
			1811: out = -19761;
			1812: out = -8966;
			1813: out = 5858;
			1814: out = 158;
			1815: out = 613;
			1816: out = 17137;
			1817: out = -2097;
			1818: out = -2107;
			1819: out = 649;
			1820: out = -10177;
			1821: out = 6340;
			1822: out = 8221;
			1823: out = -12138;
			1824: out = -2672;
			1825: out = -17432;
			1826: out = -26013;
			1827: out = 13473;
			1828: out = -1429;
			1829: out = -12879;
			1830: out = -18034;
			1831: out = -2673;
			1832: out = -8572;
			1833: out = -17438;
			1834: out = -5471;
			1835: out = 1519;
			1836: out = 10880;
			1837: out = 17874;
			1838: out = -11418;
			1839: out = -8825;
			1840: out = 7290;
			1841: out = 23659;
			1842: out = 5759;
			1843: out = 2180;
			1844: out = 14553;
			1845: out = 164;
			1846: out = -12324;
			1847: out = -18532;
			1848: out = 15907;
			1849: out = 1217;
			1850: out = 3105;
			1851: out = 11856;
			1852: out = 18352;
			1853: out = 11899;
			1854: out = 533;
			1855: out = -12558;
			1856: out = -4118;
			1857: out = -2568;
			1858: out = -10398;
			1859: out = 21959;
			1860: out = 5704;
			1861: out = -16518;
			1862: out = -27539;
			1863: out = -15440;
			1864: out = 5521;
			1865: out = 18125;
			1866: out = 7825;
			1867: out = 6908;
			1868: out = 1097;
			1869: out = -14384;
			1870: out = -7076;
			1871: out = 4177;
			1872: out = 10752;
			1873: out = -10576;
			1874: out = -2621;
			1875: out = 15701;
			1876: out = 25178;
			1877: out = 15829;
			1878: out = -5294;
			1879: out = -19604;
			1880: out = -3456;
			1881: out = 17895;
			1882: out = 22521;
			1883: out = 7186;
			1884: out = -17870;
			1885: out = -31277;
			1886: out = -22687;
			1887: out = 14493;
			1888: out = 13389;
			1889: out = 4107;
			1890: out = -3457;
			1891: out = 11574;
			1892: out = 6504;
			1893: out = -8096;
			1894: out = -939;
			1895: out = -5763;
			1896: out = 637;
			1897: out = 18040;
			1898: out = -3502;
			1899: out = 1173;
			1900: out = 7934;
			1901: out = -10575;
			1902: out = -16836;
			1903: out = -5231;
			1904: out = 23162;
			1905: out = -22563;
			1906: out = -25185;
			1907: out = -3325;
			1908: out = 18141;
			1909: out = 16866;
			1910: out = -1034;
			1911: out = -24902;
			1912: out = -21631;
			1913: out = -1988;
			1914: out = 10871;
			1915: out = -14332;
			1916: out = -6805;
			1917: out = 2285;
			1918: out = 9802;
			1919: out = 12708;
			1920: out = 1606;
			1921: out = -6107;
			1922: out = 20635;
			1923: out = 3251;
			1924: out = -1581;
			1925: out = 2221;
			1926: out = 1952;
			1927: out = 3144;
			1928: out = 3321;
			1929: out = -240;
			1930: out = 9036;
			1931: out = 15727;
			1932: out = 16750;
			1933: out = 6038;
			1934: out = 4609;
			1935: out = 5332;
			1936: out = -2318;
			1937: out = 1220;
			1938: out = -7784;
			1939: out = -20454;
			1940: out = 9271;
			1941: out = 7542;
			1942: out = -6844;
			1943: out = -26783;
			1944: out = -9968;
			1945: out = 6685;
			1946: out = 6545;
			1947: out = 15079;
			1948: out = -10785;
			1949: out = -26648;
			1950: out = -11852;
			1951: out = 8287;
			1952: out = 12515;
			1953: out = 674;
			1954: out = -5269;
			1955: out = -157;
			1956: out = 7089;
			1957: out = -7581;
			1958: out = 4953;
			1959: out = 5582;
			1960: out = 7278;
			1961: out = -26147;
			1962: out = -9488;
			1963: out = 3046;
			1964: out = 895;
			1965: out = -18084;
			1966: out = -12102;
			1967: out = 7218;
			1968: out = 9144;
			1969: out = -7232;
			1970: out = -11197;
			1971: out = 22103;
			1972: out = 894;
			1973: out = -2030;
			1974: out = -2469;
			1975: out = 6027;
			1976: out = 3637;
			1977: out = -1678;
			1978: out = -11731;
			1979: out = 11339;
			1980: out = 15496;
			1981: out = 5928;
			1982: out = -4295;
			1983: out = -15257;
			1984: out = -7057;
			1985: out = 15379;
			1986: out = 8835;
			1987: out = -972;
			1988: out = -5316;
			1989: out = 22764;
			1990: out = 15504;
			1991: out = 2759;
			1992: out = -15510;
			1993: out = -8918;
			1994: out = -1289;
			1995: out = 6197;
			1996: out = 1050;
			1997: out = -1834;
			1998: out = -7815;
			1999: out = -5788;
			2000: out = -11891;
			2001: out = -4480;
			2002: out = 3112;
			2003: out = 24126;
			2004: out = -11401;
			2005: out = -22799;
			2006: out = 639;
			2007: out = 20810;
			2008: out = 12050;
			2009: out = -4269;
			2010: out = 21001;
			2011: out = 2984;
			2012: out = 2731;
			2013: out = 7710;
			2014: out = 8110;
			2015: out = 6888;
			2016: out = 7109;
			2017: out = -35;
			2018: out = 12780;
			2019: out = 10722;
			2020: out = -2561;
			2021: out = -20361;
			2022: out = -15827;
			2023: out = -4421;
			2024: out = -27315;
			2025: out = -1998;
			2026: out = 5461;
			2027: out = 2616;
			2028: out = -13546;
			2029: out = -174;
			2030: out = 13741;
			2031: out = 1435;
			2032: out = 2993;
			2033: out = -11359;
			2034: out = -29237;
			2035: out = -2410;
			2036: out = -2477;
			2037: out = -6203;
			2038: out = 1026;
			2039: out = 7728;
			2040: out = 10049;
			2041: out = 5599;
			2042: out = 1495;
			2043: out = -252;
			2044: out = -475;
			2045: out = -1969;
			2046: out = -11409;
			2047: out = -9086;
			2048: out = 3916;
			2049: out = -10883;
			2050: out = -2219;
			2051: out = 5844;
			2052: out = 14925;
			2053: out = -9375;
			2054: out = -12387;
			2055: out = 1282;
			2056: out = -2970;
			2057: out = 4935;
			2058: out = -1278;
			2059: out = -26683;
			2060: out = 937;
			2061: out = 14218;
			2062: out = 10379;
			2063: out = -746;
			2064: out = -2006;
			2065: out = 3003;
			2066: out = -287;
			2067: out = 15283;
			2068: out = 7107;
			2069: out = -5283;
			2070: out = -15961;
			2071: out = 7836;
			2072: out = 21596;
			2073: out = 7404;
			2074: out = 17182;
			2075: out = 11831;
			2076: out = 5185;
			2077: out = -8789;
			2078: out = -11825;
			2079: out = -14195;
			2080: out = -16039;
			2081: out = -6066;
			2082: out = -912;
			2083: out = 555;
			2084: out = 2341;
			2085: out = 4830;
			2086: out = 1942;
			2087: out = -9310;
			2088: out = -316;
			2089: out = 3253;
			2090: out = 3160;
			2091: out = -19751;
			2092: out = -5022;
			2093: out = 6342;
			2094: out = 8969;
			2095: out = 12297;
			2096: out = 11883;
			2097: out = 8578;
			2098: out = 10658;
			2099: out = -5499;
			2100: out = -8600;
			2101: out = 1105;
			2102: out = 1505;
			2103: out = -5217;
			2104: out = -6399;
			2105: out = 21019;
			2106: out = 18097;
			2107: out = 11606;
			2108: out = -2339;
			2109: out = 114;
			2110: out = -1290;
			2111: out = 133;
			2112: out = -11069;
			2113: out = -4335;
			2114: out = -7388;
			2115: out = -12300;
			2116: out = -32246;
			2117: out = -8703;
			2118: out = 15904;
			2119: out = -10482;
			2120: out = 213;
			2121: out = 2148;
			2122: out = 2228;
			2123: out = 8641;
			2124: out = 246;
			2125: out = -6279;
			2126: out = 5027;
			2127: out = 689;
			2128: out = 3076;
			2129: out = 7100;
			2130: out = 1865;
			2131: out = 7478;
			2132: out = 11189;
			2133: out = 8869;
			2134: out = -7091;
			2135: out = -11525;
			2136: out = -1575;
			2137: out = -3672;
			2138: out = 1377;
			2139: out = -1536;
			2140: out = -8157;
			2141: out = -1152;
			2142: out = 3248;
			2143: out = -659;
			2144: out = 9965;
			2145: out = -9246;
			2146: out = -20726;
			2147: out = -15005;
			2148: out = 7415;
			2149: out = 10117;
			2150: out = 2483;
			2151: out = 24142;
			2152: out = 9355;
			2153: out = -5767;
			2154: out = -12563;
			2155: out = -878;
			2156: out = 16862;
			2157: out = 22456;
			2158: out = 16232;
			2159: out = -6380;
			2160: out = -14668;
			2161: out = 935;
			2162: out = 6557;
			2163: out = -2013;
			2164: out = -13360;
			2165: out = 12950;
			2166: out = 12154;
			2167: out = -1008;
			2168: out = -30867;
			2169: out = -17496;
			2170: out = -9729;
			2171: out = -304;
			2172: out = 3604;
			2173: out = 18656;
			2174: out = 13956;
			2175: out = -11985;
			2176: out = -15132;
			2177: out = -17217;
			2178: out = -5443;
			2179: out = -684;
			2180: out = 20757;
			2181: out = 11546;
			2182: out = -17211;
			2183: out = -15518;
			2184: out = 2749;
			2185: out = 18763;
			2186: out = 4095;
			2187: out = -1385;
			2188: out = -2090;
			2189: out = 11153;
			2190: out = -4758;
			2191: out = -4040;
			2192: out = -4489;
			2193: out = -6320;
			2194: out = -1131;
			2195: out = 3142;
			2196: out = -1304;
			2197: out = 4928;
			2198: out = -2677;
			2199: out = -6997;
			2200: out = -9144;
			2201: out = -830;
			2202: out = 293;
			2203: out = 748;
			2204: out = -12295;
			2205: out = 5267;
			2206: out = 14067;
			2207: out = -8733;
			2208: out = -18355;
			2209: out = -10115;
			2210: out = 15519;
			2211: out = -4179;
			2212: out = -8791;
			2213: out = -8473;
			2214: out = 22765;
			2215: out = 220;
			2216: out = 2558;
			2217: out = 10138;
			2218: out = 12888;
			2219: out = -4094;
			2220: out = -7713;
			2221: out = 21849;
			2222: out = 9439;
			2223: out = -984;
			2224: out = -12950;
			2225: out = -3466;
			2226: out = -538;
			2227: out = 3708;
			2228: out = 2596;
			2229: out = 3806;
			2230: out = -10662;
			2231: out = -27040;
			2232: out = 3828;
			2233: out = 4514;
			2234: out = -3436;
			2235: out = -23144;
			2236: out = 6203;
			2237: out = 13181;
			2238: out = 8555;
			2239: out = 15294;
			2240: out = 19421;
			2241: out = 16367;
			2242: out = -1535;
			2243: out = 931;
			2244: out = -1545;
			2245: out = -2206;
			2246: out = -5615;
			2247: out = -2422;
			2248: out = 2853;
			2249: out = 10643;
			2250: out = -6552;
			2251: out = -12294;
			2252: out = -7625;
			2253: out = 5195;
			2254: out = 6013;
			2255: out = -3668;
			2256: out = -21376;
			2257: out = -4031;
			2258: out = 6652;
			2259: out = 7809;
			2260: out = -5846;
			2261: out = -3092;
			2262: out = 3936;
			2263: out = 9264;
			2264: out = 3963;
			2265: out = -5483;
			2266: out = -15054;
			2267: out = -10879;
			2268: out = -11589;
			2269: out = -4262;
			2270: out = 6956;
			2271: out = 16613;
			2272: out = 13797;
			2273: out = 6170;
			2274: out = 4345;
			2275: out = 1029;
			2276: out = -340;
			2277: out = -1681;
			2278: out = -1071;
			2279: out = 9595;
			2280: out = 15505;
			2281: out = -19024;
			2282: out = -3806;
			2283: out = 1197;
			2284: out = 331;
			2285: out = -3248;
			2286: out = 7339;
			2287: out = 3806;
			2288: out = -28590;
			2289: out = -28417;
			2290: out = -10865;
			2291: out = 19644;
			2292: out = 4047;
			2293: out = 4298;
			2294: out = 1186;
			2295: out = 2091;
			2296: out = 296;
			2297: out = 6763;
			2298: out = 11910;
			2299: out = 10847;
			2300: out = -1474;
			2301: out = -10148;
			2302: out = 1471;
			2303: out = -984;
			2304: out = 4771;
			2305: out = 11639;
			2306: out = -2208;
			2307: out = -5258;
			2308: out = -2067;
			2309: out = 12636;
			2310: out = -6349;
			2311: out = -9830;
			2312: out = 1665;
			2313: out = -3042;
			2314: out = 2001;
			2315: out = 4461;
			2316: out = 9779;
			2317: out = 253;
			2318: out = -3715;
			2319: out = -4827;
			2320: out = 6094;
			2321: out = 3102;
			2322: out = 197;
			2323: out = -4662;
			2324: out = 3337;
			2325: out = -7260;
			2326: out = -23226;
			2327: out = -147;
			2328: out = 7699;
			2329: out = 13904;
			2330: out = 20622;
			2331: out = -1425;
			2332: out = -9841;
			2333: out = -6409;
			2334: out = 9526;
			2335: out = 4686;
			2336: out = -5377;
			2337: out = -19790;
			2338: out = 8705;
			2339: out = 10527;
			2340: out = -1225;
			2341: out = -1391;
			2342: out = 425;
			2343: out = -3111;
			2344: out = -20612;
			2345: out = -18118;
			2346: out = -12078;
			2347: out = -2422;
			2348: out = 1557;
			2349: out = -823;
			2350: out = -511;
			2351: out = 8331;
			2352: out = 10331;
			2353: out = 8454;
			2354: out = 2170;
			2355: out = 1274;
			2356: out = 3249;
			2357: out = 3186;
			2358: out = -5209;
			2359: out = 15771;
			2360: out = 21039;
			2361: out = 18121;
			2362: out = -9719;
			2363: out = 518;
			2364: out = 3134;
			2365: out = -936;
			2366: out = -14939;
			2367: out = -3557;
			2368: out = 10598;
			2369: out = -8806;
			2370: out = -4189;
			2371: out = -2302;
			2372: out = 3785;
			2373: out = -9864;
			2374: out = -5708;
			2375: out = 2772;
			2376: out = 13144;
			2377: out = 4484;
			2378: out = -1495;
			2379: out = -4235;
			2380: out = -5030;
			2381: out = -7461;
			2382: out = -10012;
			2383: out = -17674;
			2384: out = 5287;
			2385: out = 14316;
			2386: out = 4896;
			2387: out = -349;
			2388: out = -9452;
			2389: out = -3808;
			2390: out = 18447;
			2391: out = 11714;
			2392: out = 5310;
			2393: out = -25;
			2394: out = -14055;
			2395: out = -16894;
			2396: out = -12402;
			2397: out = 505;
			2398: out = 17;
			2399: out = 3630;
			2400: out = 4857;
			2401: out = -10741;
			2402: out = -21335;
			2403: out = -19744;
			2404: out = 2599;
			2405: out = 10887;
			2406: out = 14761;
			2407: out = 8569;
			2408: out = 2747;
			2409: out = -8000;
			2410: out = -9302;
			2411: out = -2725;
			2412: out = 6912;
			2413: out = 6097;
			2414: out = 1764;
			2415: out = 1995;
			2416: out = 10752;
			2417: out = 10727;
			2418: out = -7580;
			2419: out = 4211;
			2420: out = 11116;
			2421: out = 13726;
			2422: out = -9644;
			2423: out = -5452;
			2424: out = -1394;
			2425: out = -3953;
			2426: out = -1536;
			2427: out = -4157;
			2428: out = -3821;
			2429: out = 17908;
			2430: out = 5332;
			2431: out = -11203;
			2432: out = -23402;
			2433: out = 1887;
			2434: out = 14765;
			2435: out = 9399;
			2436: out = 2449;
			2437: out = -12077;
			2438: out = -9613;
			2439: out = 5999;
			2440: out = 12542;
			2441: out = 8976;
			2442: out = 5093;
			2443: out = 8133;
			2444: out = 16004;
			2445: out = 9777;
			2446: out = -10831;
			2447: out = -13606;
			2448: out = -5467;
			2449: out = 9777;
			2450: out = 13598;
			2451: out = 5786;
			2452: out = -4988;
			2453: out = -6585;
			2454: out = -12938;
			2455: out = -6186;
			2456: out = 3012;
			2457: out = 13603;
			2458: out = 1124;
			2459: out = -10356;
			2460: out = -13446;
			2461: out = -19725;
			2462: out = -10535;
			2463: out = 1445;
			2464: out = 6143;
			2465: out = 5599;
			2466: out = 6984;
			2467: out = 11507;
			2468: out = -2203;
			2469: out = -1989;
			2470: out = -1269;
			2471: out = -14093;
			2472: out = 975;
			2473: out = 6823;
			2474: out = 2535;
			2475: out = 6531;
			2476: out = 2907;
			2477: out = -2312;
			2478: out = -10075;
			2479: out = -14126;
			2480: out = -13020;
			2481: out = -3405;
			2482: out = 10495;
			2483: out = 16786;
			2484: out = 8863;
			2485: out = -14746;
			2486: out = -10083;
			2487: out = -1337;
			2488: out = 3575;
			2489: out = 4163;
			2490: out = -1939;
			2491: out = -11618;
			2492: out = -29733;
			2493: out = -6003;
			2494: out = 3988;
			2495: out = -834;
			2496: out = 13823;
			2497: out = 12849;
			2498: out = 11051;
			2499: out = 6146;
			2500: out = 5801;
			2501: out = 2117;
			2502: out = -2128;
			2503: out = 701;
			2504: out = 393;
			2505: out = 4163;
			2506: out = 9801;
			2507: out = 1880;
			2508: out = -10491;
			2509: out = -16321;
			2510: out = 8280;
			2511: out = 15212;
			2512: out = 10892;
			2513: out = -1328;
			2514: out = -19551;
			2515: out = -23594;
			2516: out = -10333;
			2517: out = 4114;
			2518: out = 16207;
			2519: out = 11236;
			2520: out = -12795;
			2521: out = 6676;
			2522: out = 5814;
			2523: out = -998;
			2524: out = -6513;
			2525: out = 5419;
			2526: out = 10408;
			2527: out = -1285;
			2528: out = 4978;
			2529: out = 2721;
			2530: out = 920;
			2531: out = 93;
			2532: out = 3642;
			2533: out = 7238;
			2534: out = 6263;
			2535: out = 9756;
			2536: out = -4348;
			2537: out = -16072;
			2538: out = 10341;
			2539: out = 3821;
			2540: out = -4492;
			2541: out = -15918;
			2542: out = -2456;
			2543: out = 5730;
			2544: out = 7177;
			2545: out = -19555;
			2546: out = -8361;
			2547: out = -2156;
			2548: out = -1782;
			2549: out = -7746;
			2550: out = -6150;
			2551: out = -3347;
			2552: out = 8023;
			2553: out = -12117;
			2554: out = -9891;
			2555: out = 15106;
			2556: out = 13445;
			2557: out = 6299;
			2558: out = -5127;
			2559: out = 3047;
			2560: out = 676;
			2561: out = 1453;
			2562: out = -4178;
			2563: out = 8056;
			2564: out = 3011;
			2565: out = -856;
			2566: out = -9211;
			2567: out = 7649;
			2568: out = 6053;
			2569: out = -8502;
			2570: out = -9398;
			2571: out = -2896;
			2572: out = 1878;
			2573: out = -17937;
			2574: out = -4805;
			2575: out = 1611;
			2576: out = 6239;
			2577: out = 2886;
			2578: out = 8860;
			2579: out = 5989;
			2580: out = -13009;
			2581: out = 4409;
			2582: out = 13635;
			2583: out = 9138;
			2584: out = 11609;
			2585: out = -10863;
			2586: out = -17986;
			2587: out = 10823;
			2588: out = 11217;
			2589: out = 11346;
			2590: out = 4933;
			2591: out = -2355;
			2592: out = -2752;
			2593: out = 2016;
			2594: out = 3439;
			2595: out = 2505;
			2596: out = -4095;
			2597: out = -8048;
			2598: out = -1016;
			2599: out = 4447;
			2600: out = -268;
			2601: out = -23826;
			2602: out = -6082;
			2603: out = 3866;
			2604: out = 7514;
			2605: out = -18391;
			2606: out = -4681;
			2607: out = 4847;
			2608: out = 1807;
			2609: out = 1608;
			2610: out = 6864;
			2611: out = 10901;
			2612: out = 5361;
			2613: out = -2401;
			2614: out = -2618;
			2615: out = 4660;
			2616: out = 6681;
			2617: out = -2769;
			2618: out = -10661;
			2619: out = 2237;
			2620: out = 12459;
			2621: out = 7340;
			2622: out = -15121;
			2623: out = -15659;
			2624: out = -238;
			2625: out = 17221;
			2626: out = -7058;
			2627: out = -3245;
			2628: out = -8114;
			2629: out = -8185;
			2630: out = -4704;
			2631: out = 7028;
			2632: out = 10268;
			2633: out = 5626;
			2634: out = -2907;
			2635: out = -3842;
			2636: out = -2014;
			2637: out = 6756;
			2638: out = -6415;
			2639: out = -19021;
			2640: out = -9472;
			2641: out = 8762;
			2642: out = 11609;
			2643: out = -7472;
			2644: out = 5084;
			2645: out = -3664;
			2646: out = -6100;
			2647: out = 1809;
			2648: out = 7039;
			2649: out = 4288;
			2650: out = -3702;
			2651: out = 2007;
			2652: out = 804;
			2653: out = 568;
			2654: out = 3479;
			2655: out = 2380;
			2656: out = 1693;
			2657: out = 776;
			2658: out = -16533;
			2659: out = -12261;
			2660: out = -1416;
			2661: out = -811;
			2662: out = 3941;
			2663: out = 4133;
			2664: out = 7370;
			2665: out = -496;
			2666: out = 11767;
			2667: out = 14729;
			2668: out = -648;
			2669: out = -2368;
			2670: out = -2101;
			2671: out = 2479;
			2672: out = 8091;
			2673: out = 3986;
			2674: out = -1173;
			2675: out = 760;
			2676: out = 1536;
			2677: out = 5844;
			2678: out = 6750;
			2679: out = -8937;
			2680: out = -8978;
			2681: out = -5734;
			2682: out = -5323;
			2683: out = -3341;
			2684: out = -4657;
			2685: out = -4789;
			2686: out = 10982;
			2687: out = 4686;
			2688: out = -3887;
			2689: out = -10765;
			2690: out = 8213;
			2691: out = 8457;
			2692: out = -4634;
			2693: out = 192;
			2694: out = -6364;
			2695: out = -4504;
			2696: out = -3539;
			2697: out = 17916;
			2698: out = 12952;
			2699: out = -416;
			2700: out = -12207;
			2701: out = -4519;
			2702: out = 4472;
			2703: out = 5124;
			2704: out = -4176;
			2705: out = -4589;
			2706: out = 1967;
			2707: out = 3913;
			2708: out = 2612;
			2709: out = 2224;
			2710: out = 7304;
			2711: out = -4391;
			2712: out = -10488;
			2713: out = -11758;
			2714: out = -488;
			2715: out = 2231;
			2716: out = 4795;
			2717: out = 6823;
			2718: out = -6805;
			2719: out = -11752;
			2720: out = -7617;
			2721: out = 10017;
			2722: out = 7574;
			2723: out = 4198;
			2724: out = 186;
			2725: out = 14008;
			2726: out = 4463;
			2727: out = -9431;
			2728: out = -9047;
			2729: out = 1255;
			2730: out = 6891;
			2731: out = -3629;
			2732: out = 16302;
			2733: out = 92;
			2734: out = -17668;
			2735: out = -11929;
			2736: out = -10967;
			2737: out = -1580;
			2738: out = 7797;
			2739: out = 2946;
			2740: out = -3297;
			2741: out = -7222;
			2742: out = 2943;
			2743: out = -1393;
			2744: out = 2873;
			2745: out = 10761;
			2746: out = 8689;
			2747: out = 5818;
			2748: out = 205;
			2749: out = -9802;
			2750: out = -449;
			2751: out = 2495;
			2752: out = -2102;
			2753: out = 9281;
			2754: out = 10418;
			2755: out = 7788;
			2756: out = -8083;
			2757: out = -1394;
			2758: out = -4910;
			2759: out = -11656;
			2760: out = -6052;
			2761: out = -1094;
			2762: out = 2213;
			2763: out = 6309;
			2764: out = -6480;
			2765: out = -8252;
			2766: out = -2750;
			2767: out = -2881;
			2768: out = -10897;
			2769: out = -12457;
			2770: out = 9474;
			2771: out = -2406;
			2772: out = -4095;
			2773: out = -1727;
			2774: out = 6107;
			2775: out = 2453;
			2776: out = -4168;
			2777: out = -8389;
			2778: out = 2281;
			2779: out = 11848;
			2780: out = 11203;
			2781: out = -3885;
			2782: out = -9200;
			2783: out = -1961;
			2784: out = 10349;
			2785: out = 19087;
			2786: out = 10845;
			2787: out = -2233;
			2788: out = -6117;
			2789: out = 1669;
			2790: out = 8536;
			2791: out = 6016;
			2792: out = -1555;
			2793: out = -1139;
			2794: out = 4945;
			2795: out = -806;
			2796: out = -2201;
			2797: out = -1008;
			2798: out = 10327;
			2799: out = -10097;
			2800: out = -15289;
			2801: out = -10220;
			2802: out = 21215;
			2803: out = 5404;
			2804: out = -4757;
			2805: out = -4371;
			2806: out = 5208;
			2807: out = 3298;
			2808: out = -3080;
			2809: out = 1384;
			2810: out = 833;
			2811: out = 1022;
			2812: out = -991;
			2813: out = 608;
			2814: out = 2993;
			2815: out = 6254;
			2816: out = 6034;
			2817: out = 2446;
			2818: out = -9312;
			2819: out = -25541;
			2820: out = -2611;
			2821: out = 2209;
			2822: out = 594;
			2823: out = 1203;
			2824: out = -1819;
			2825: out = -6930;
			2826: out = -12818;
			2827: out = -7425;
			2828: out = 1375;
			2829: out = 9523;
			2830: out = 9120;
			2831: out = 2589;
			2832: out = -5694;
			2833: out = -6990;
			2834: out = -7591;
			2835: out = -758;
			2836: out = 2702;
			2837: out = 7010;
			2838: out = 2881;
			2839: out = 6699;
			2840: out = 8691;
			2841: out = 7720;
			2842: out = -7960;
			2843: out = -14123;
			2844: out = 1485;
			2845: out = 12338;
			2846: out = 8805;
			2847: out = -4332;
			2848: out = -12063;
			2849: out = -3491;
			2850: out = 5286;
			2851: out = -3208;
			2852: out = -9082;
			2853: out = -14792;
			2854: out = -11928;
			2855: out = 236;
			2856: out = 2307;
			2857: out = -496;
			2858: out = -3953;
			2859: out = 1240;
			2860: out = 2660;
			2861: out = 1771;
			2862: out = -8913;
			2863: out = 2658;
			2864: out = 8205;
			2865: out = -1753;
			2866: out = -300;
			2867: out = 9688;
			2868: out = 22088;
			2869: out = 10009;
			2870: out = 6139;
			2871: out = -2701;
			2872: out = -6762;
			2873: out = 2796;
			2874: out = 12411;
			2875: out = 11574;
			2876: out = 2710;
			2877: out = -6883;
			2878: out = -10326;
			2879: out = -9702;
			2880: out = 4490;
			2881: out = 4545;
			2882: out = -942;
			2883: out = 1425;
			2884: out = -4086;
			2885: out = -5118;
			2886: out = 4077;
			2887: out = -17462;
			2888: out = -7428;
			2889: out = 11424;
			2890: out = 6049;
			2891: out = -979;
			2892: out = -3362;
			2893: out = 14256;
			2894: out = -10991;
			2895: out = -8865;
			2896: out = -3316;
			2897: out = 8478;
			2898: out = -8430;
			2899: out = -8115;
			2900: out = 11561;
			2901: out = 2460;
			2902: out = -1372;
			2903: out = -5071;
			2904: out = -4657;
			2905: out = 5859;
			2906: out = 6031;
			2907: out = -9667;
			2908: out = 1695;
			2909: out = -3545;
			2910: out = -8427;
			2911: out = -10549;
			2912: out = -2255;
			2913: out = 5003;
			2914: out = 6956;
			2915: out = -999;
			2916: out = -3905;
			2917: out = 616;
			2918: out = 12139;
			2919: out = 7518;
			2920: out = 1358;
			2921: out = -871;
			2922: out = -1088;
			2923: out = 12302;
			2924: out = 18396;
			2925: out = -1536;
			2926: out = 8270;
			2927: out = 11206;
			2928: out = 11184;
			2929: out = -6874;
			2930: out = -9408;
			2931: out = -7524;
			2932: out = -1987;
			2933: out = -3898;
			2934: out = -2261;
			2935: out = -294;
			2936: out = 7915;
			2937: out = 3619;
			2938: out = -1565;
			2939: out = -10988;
			2940: out = 859;
			2941: out = -4262;
			2942: out = -16210;
			2943: out = -2427;
			2944: out = 9630;
			2945: out = 10898;
			2946: out = -4021;
			2947: out = -13771;
			2948: out = -8290;
			2949: out = 10782;
			2950: out = 14693;
			2951: out = 6375;
			2952: out = -9539;
			2953: out = -12372;
			2954: out = -13593;
			2955: out = 3411;
			2956: out = 17399;
			2957: out = 14252;
			2958: out = 4109;
			2959: out = -2665;
			2960: out = 5152;
			2961: out = -5803;
			2962: out = -4045;
			2963: out = 181;
			2964: out = 1401;
			2965: out = -4639;
			2966: out = -9072;
			2967: out = -7697;
			2968: out = -4513;
			2969: out = -1635;
			2970: out = -705;
			2971: out = -7880;
			2972: out = 294;
			2973: out = 4510;
			2974: out = -1410;
			2975: out = -12073;
			2976: out = -15417;
			2977: out = -6890;
			2978: out = 653;
			2979: out = 8034;
			2980: out = 9099;
			2981: out = 11445;
			2982: out = -5393;
			2983: out = -3663;
			2984: out = 2022;
			2985: out = 933;
			2986: out = -6355;
			2987: out = -3762;
			2988: out = 12654;
			2989: out = 4993;
			2990: out = 738;
			2991: out = -5260;
			2992: out = 2520;
			2993: out = -2780;
			2994: out = 721;
			2995: out = 6721;
			2996: out = -4783;
			2997: out = -11388;
			2998: out = -10024;
			2999: out = -3648;
			3000: out = 9958;
			3001: out = 10781;
			3002: out = 627;
			3003: out = 865;
			3004: out = -137;
			3005: out = 1019;
			3006: out = 1840;
			3007: out = 2632;
			3008: out = 5578;
			3009: out = 9920;
			3010: out = 9408;
			3011: out = 5919;
			3012: out = 1045;
			3013: out = -1734;
			3014: out = 3612;
			3015: out = 9663;
			3016: out = 11547;
			3017: out = 4630;
			3018: out = -187;
			3019: out = -3316;
			3020: out = -2251;
			3021: out = -2142;
			3022: out = 1569;
			3023: out = 4443;
			3024: out = 1474;
			3025: out = -3260;
			3026: out = -6053;
			3027: out = -7578;
			3028: out = -1439;
			3029: out = -9144;
			3030: out = -24554;
			3031: out = 1081;
			3032: out = 5058;
			3033: out = 4639;
			3034: out = -910;
			3035: out = 2705;
			3036: out = -718;
			3037: out = -6191;
			3038: out = 5147;
			3039: out = 4828;
			3040: out = 2285;
			3041: out = -5467;
			3042: out = 4811;
			3043: out = 4692;
			3044: out = -439;
			3045: out = -6272;
			3046: out = -208;
			3047: out = 3497;
			3048: out = -4282;
			3049: out = 2903;
			3050: out = 4995;
			3051: out = 3322;
			3052: out = -11483;
			3053: out = -12215;
			3054: out = -3004;
			3055: out = 13244;
			3056: out = -2468;
			3057: out = -9347;
			3058: out = -5901;
			3059: out = 12632;
			3060: out = 12425;
			3061: out = 1632;
			3062: out = -16558;
			3063: out = -13744;
			3064: out = -8203;
			3065: out = -513;
			3066: out = 9187;
			3067: out = 3932;
			3068: out = -3079;
			3069: out = -4927;
			3070: out = 8560;
			3071: out = 10762;
			3072: out = 2584;
			3073: out = 3215;
			3074: out = -10198;
			3075: out = -4284;
			3076: out = 16467;
			3077: out = 14870;
			3078: out = 4819;
			3079: out = -9180;
			3080: out = -2097;
			3081: out = -11158;
			3082: out = -8812;
			3083: out = 1458;
			3084: out = -5334;
			3085: out = -7346;
			3086: out = -6020;
			3087: out = 3355;
			3088: out = 2836;
			3089: out = 4591;
			3090: out = 7265;
			3091: out = 12260;
			3092: out = 9646;
			3093: out = 3723;
			3094: out = -6718;
			3095: out = -2489;
			3096: out = -1404;
			3097: out = -3394;
			3098: out = 253;
			3099: out = 6655;
			3100: out = 7228;
			3101: out = -10158;
			3102: out = -3623;
			3103: out = 2707;
			3104: out = 6744;
			3105: out = 9994;
			3106: out = 1972;
			3107: out = -8569;
			3108: out = -12022;
			3109: out = -9438;
			3110: out = -1984;
			3111: out = 3024;
			3112: out = 5428;
			3113: out = 2849;
			3114: out = 1985;
			3115: out = 6468;
			3116: out = -2858;
			3117: out = -12555;
			3118: out = -17745;
			3119: out = 5726;
			3120: out = 9984;
			3121: out = 5356;
			3122: out = -8488;
			3123: out = -5302;
			3124: out = -5047;
			3125: out = -3687;
			3126: out = -1532;
			3127: out = 9946;
			3128: out = 12607;
			3129: out = -1318;
			3130: out = -4481;
			3131: out = -4649;
			3132: out = 1692;
			3133: out = -11497;
			3134: out = 2658;
			3135: out = 11957;
			3136: out = 7686;
			3137: out = -1639;
			3138: out = -15702;
			3139: out = -24029;
			3140: out = -1375;
			3141: out = 3223;
			3142: out = 8162;
			3143: out = 16235;
			3144: out = 4246;
			3145: out = -3891;
			3146: out = -5007;
			3147: out = 16509;
			3148: out = 6541;
			3149: out = -4134;
			3150: out = -3532;
			3151: out = -11576;
			3152: out = -491;
			3153: out = 9088;
			3154: out = -13212;
			3155: out = -11985;
			3156: out = -1266;
			3157: out = 17505;
			3158: out = 8382;
			3159: out = 8315;
			3160: out = 4755;
			3161: out = -11324;
			3162: out = -14510;
			3163: out = -11077;
			3164: out = -3605;
			3165: out = 3018;
			3166: out = 5798;
			3167: out = 4906;
			3168: out = 1934;
			3169: out = -550;
			3170: out = -2326;
			3171: out = -2495;
			3172: out = 5336;
			3173: out = 6536;
			3174: out = 1651;
			3175: out = -5043;
			3176: out = -12380;
			3177: out = -8186;
			3178: out = 7430;
			3179: out = 787;
			3180: out = 5905;
			3181: out = 9354;
			3182: out = 6503;
			3183: out = -1705;
			3184: out = -9656;
			3185: out = -11373;
			3186: out = -10555;
			3187: out = 610;
			3188: out = 9686;
			3189: out = 6194;
			3190: out = 5713;
			3191: out = 3026;
			3192: out = 2628;
			3193: out = -10976;
			3194: out = -6114;
			3195: out = 997;
			3196: out = -6766;
			3197: out = 431;
			3198: out = 1005;
			3199: out = -2069;
			3200: out = -9193;
			3201: out = -4641;
			3202: out = 7793;
			3203: out = 20019;
			3204: out = 11599;
			3205: out = -2096;
			3206: out = -14047;
			3207: out = -10056;
			3208: out = -1938;
			3209: out = 3605;
			3210: out = -1963;
			3211: out = 7998;
			3212: out = 10395;
			3213: out = 6530;
			3214: out = 2485;
			3215: out = -7823;
			3216: out = -12908;
			3217: out = -458;
			3218: out = -4778;
			3219: out = -990;
			3220: out = 3255;
			3221: out = 3475;
			3222: out = 73;
			3223: out = -1855;
			3224: out = -3017;
			3225: out = 13288;
			3226: out = 14886;
			3227: out = 6162;
			3228: out = -3284;
			3229: out = -8189;
			3230: out = -11961;
			3231: out = -20674;
			3232: out = -7519;
			3233: out = 4053;
			3234: out = 10071;
			3235: out = 10700;
			3236: out = 5601;
			3237: out = 2642;
			3238: out = 4133;
			3239: out = 3238;
			3240: out = -703;
			3241: out = -5318;
			3242: out = -4754;
			3243: out = -881;
			3244: out = 3259;
			3245: out = 6266;
			3246: out = -13930;
			3247: out = -16974;
			3248: out = -4789;
			3249: out = 3873;
			3250: out = 9996;
			3251: out = 3651;
			3252: out = -10980;
			3253: out = -7831;
			3254: out = -4088;
			3255: out = 2631;
			3256: out = 8719;
			3257: out = 11886;
			3258: out = 9247;
			3259: out = 5016;
			3260: out = -6025;
			3261: out = -4812;
			3262: out = 1499;
			3263: out = 6556;
			3264: out = 50;
			3265: out = -3707;
			3266: out = -1179;
			3267: out = 3628;
			3268: out = -1422;
			3269: out = -5747;
			3270: out = 14693;
			3271: out = 6043;
			3272: out = 2750;
			3273: out = -431;
			3274: out = -7413;
			3275: out = -11408;
			3276: out = -8720;
			3277: out = -5396;
			3278: out = 6300;
			3279: out = 8826;
			3280: out = 6126;
			3281: out = -1467;
			3282: out = 3588;
			3283: out = 5262;
			3284: out = -11075;
			3285: out = -15577;
			3286: out = -12059;
			3287: out = 2862;
			3288: out = -1067;
			3289: out = 4733;
			3290: out = 4266;
			3291: out = 2059;
			3292: out = -8261;
			3293: out = -5258;
			3294: out = 6371;
			3295: out = 9636;
			3296: out = 4320;
			3297: out = -2904;
			3298: out = 2962;
			3299: out = -6232;
			3300: out = -6728;
			3301: out = -4437;
			3302: out = 14629;
			3303: out = 2932;
			3304: out = -7690;
			3305: out = -3406;
			3306: out = -1566;
			3307: out = -921;
			3308: out = -5222;
			3309: out = -3493;
			3310: out = -1407;
			3311: out = 5461;
			3312: out = 9536;
			3313: out = 5943;
			3314: out = -4946;
			3315: out = -12582;
			3316: out = -642;
			3317: out = 6027;
			3318: out = 7001;
			3319: out = 1576;
			3320: out = 8699;
			3321: out = 9399;
			3322: out = 4671;
			3323: out = 2642;
			3324: out = -6253;
			3325: out = -7553;
			3326: out = -1470;
			3327: out = 6879;
			3328: out = 741;
			3329: out = -9752;
			3330: out = 1502;
			3331: out = 1828;
			3332: out = 3348;
			3333: out = 1913;
			3334: out = -6259;
			3335: out = -11025;
			3336: out = -7083;
			3337: out = 7148;
			3338: out = 4771;
			3339: out = -843;
			3340: out = -2274;
			3341: out = -3741;
			3342: out = -315;
			3343: out = 2071;
			3344: out = 9950;
			3345: out = -3439;
			3346: out = -6806;
			3347: out = 4711;
			3348: out = 4037;
			3349: out = 8487;
			3350: out = 8928;
			3351: out = 3903;
			3352: out = 2816;
			3353: out = 1722;
			3354: out = 416;
			3355: out = -1910;
			3356: out = -754;
			3357: out = -324;
			3358: out = -7946;
			3359: out = -2089;
			3360: out = 3131;
			3361: out = 4496;
			3362: out = 941;
			3363: out = -4313;
			3364: out = -9565;
			3365: out = -16680;
			3366: out = -6648;
			3367: out = 3398;
			3368: out = 7664;
			3369: out = 2149;
			3370: out = -1340;
			3371: out = -2709;
			3372: out = 1684;
			3373: out = -2466;
			3374: out = 497;
			3375: out = 7570;
			3376: out = 9617;
			3377: out = 5189;
			3378: out = 373;
			3379: out = 5795;
			3380: out = -2674;
			3381: out = -5306;
			3382: out = -4712;
			3383: out = -5971;
			3384: out = -6884;
			3385: out = -6066;
			3386: out = 920;
			3387: out = 560;
			3388: out = 1358;
			3389: out = -411;
			3390: out = 9853;
			3391: out = -3953;
			3392: out = -13763;
			3393: out = -4658;
			3394: out = -828;
			3395: out = 2533;
			3396: out = 1211;
			3397: out = -856;
			3398: out = 950;
			3399: out = 4313;
			3400: out = 5225;
			3401: out = 2387;
			3402: out = 801;
			3403: out = 2936;
			3404: out = 11451;
			3405: out = 6952;
			3406: out = -981;
			3407: out = -5630;
			3408: out = -3899;
			3409: out = 4206;
			3410: out = 11553;
			3411: out = 9007;
			3412: out = 6201;
			3413: out = 1421;
			3414: out = 1293;
			3415: out = -10863;
			3416: out = -7774;
			3417: out = 621;
			3418: out = -2307;
			3419: out = -4023;
			3420: out = -1894;
			3421: out = 7999;
			3422: out = 531;
			3423: out = -4700;
			3424: out = -9685;
			3425: out = -4347;
			3426: out = -1380;
			3427: out = 3320;
			3428: out = 3217;
			3429: out = 9813;
			3430: out = 4648;
			3431: out = -1536;
			3432: out = -6388;
			3433: out = -410;
			3434: out = 2451;
			3435: out = 842;
			3436: out = 5825;
			3437: out = 10229;
			3438: out = 9114;
			3439: out = -295;
			3440: out = -11690;
			3441: out = -12893;
			3442: out = -195;
			3443: out = 8235;
			3444: out = 9435;
			3445: out = 2935;
			3446: out = -2931;
			3447: out = -7488;
			3448: out = -6377;
			3449: out = -1973;
			3450: out = -8833;
			3451: out = -5142;
			3452: out = 596;
			3453: out = 421;
			3454: out = -2729;
			3455: out = -4461;
			3456: out = -1281;
			3457: out = -5975;
			3458: out = -3022;
			3459: out = 1344;
			3460: out = 5104;
			3461: out = 1908;
			3462: out = -1202;
			3463: out = -1571;
			3464: out = -7364;
			3465: out = -1106;
			3466: out = 5712;
			3467: out = 6072;
			3468: out = 2867;
			3469: out = 2031;
			3470: out = 5272;
			3471: out = -3053;
			3472: out = -1504;
			3473: out = 834;
			3474: out = 3866;
			3475: out = -2530;
			3476: out = -4881;
			3477: out = -2658;
			3478: out = -3613;
			3479: out = -1018;
			3480: out = 950;
			3481: out = 4122;
			3482: out = -4653;
			3483: out = -7268;
			3484: out = -2470;
			3485: out = 5160;
			3486: out = 6833;
			3487: out = 2010;
			3488: out = -5519;
			3489: out = -1017;
			3490: out = 5867;
			3491: out = 9453;
			3492: out = 7819;
			3493: out = 2846;
			3494: out = 559;
			3495: out = 2496;
			3496: out = 6931;
			3497: out = 7996;
			3498: out = 5121;
			3499: out = -6043;
			3500: out = -2999;
			3501: out = 1088;
			3502: out = -220;
			3503: out = 1824;
			3504: out = 2929;
			3505: out = 3501;
			3506: out = -6529;
			3507: out = -4292;
			3508: out = -1319;
			3509: out = -171;
			3510: out = -5960;
			3511: out = -11255;
			3512: out = -13315;
			3513: out = -10802;
			3514: out = -305;
			3515: out = 7289;
			3516: out = 5206;
			3517: out = 4186;
			3518: out = 16;
			3519: out = 406;
			3520: out = -503;
			3521: out = 12917;
			3522: out = 11198;
			3523: out = -6601;
			3524: out = 423;
			3525: out = 4648;
			3526: out = 8201;
			3527: out = -7427;
			3528: out = 603;
			3529: out = 4170;
			3530: out = 5252;
			3531: out = -10199;
			3532: out = -10272;
			3533: out = -5846;
			3534: out = -7874;
			3535: out = -8694;
			3536: out = -6841;
			3537: out = -1082;
			3538: out = -1778;
			3539: out = -2108;
			3540: out = -3485;
			3541: out = -5580;
			3542: out = -1766;
			3543: out = 1075;
			3544: out = 1402;
			3545: out = -6021;
			3546: out = -2860;
			3547: out = 3529;
			3548: out = 3741;
			3549: out = 2818;
			3550: out = 3068;
			3551: out = 8574;
			3552: out = 983;
			3553: out = 4881;
			3554: out = 4355;
			3555: out = -2874;
			3556: out = -9765;
			3557: out = -9664;
			3558: out = -2466;
			3559: out = 6328;
			3560: out = 7805;
			3561: out = 4144;
			3562: out = -2998;
			3563: out = 3014;
			3564: out = 5751;
			3565: out = 4014;
			3566: out = -2336;
			3567: out = -2858;
			3568: out = -1958;
			3569: out = -4756;
			3570: out = 1148;
			3571: out = 2247;
			3572: out = -290;
			3573: out = 5434;
			3574: out = 2042;
			3575: out = 3784;
			3576: out = 11159;
			3577: out = 5275;
			3578: out = -7565;
			3579: out = -19441;
			3580: out = -822;
			3581: out = 9421;
			3582: out = 12589;
			3583: out = 3422;
			3584: out = 5421;
			3585: out = 2797;
			3586: out = 2555;
			3587: out = 3784;
			3588: out = 1963;
			3589: out = -5914;
			3590: out = -16389;
			3591: out = -10417;
			3592: out = -3693;
			3593: out = -2767;
			3594: out = -4627;
			3595: out = -7101;
			3596: out = -946;
			3597: out = 7162;
			3598: out = 14308;
			3599: out = 1791;
			3600: out = -15250;
			3601: out = -12621;
			3602: out = -3259;
			3603: out = 4409;
			3604: out = 736;
			3605: out = 1659;
			3606: out = 4567;
			3607: out = 10838;
			3608: out = 7463;
			3609: out = 6306;
			3610: out = -609;
			3611: out = -7151;
			3612: out = -5906;
			3613: out = 1536;
			3614: out = 7264;
			3615: out = -614;
			3616: out = 410;
			3617: out = -2294;
			3618: out = -5390;
			3619: out = -1946;
			3620: out = 8546;
			3621: out = 13634;
			3622: out = -4970;
			3623: out = -8150;
			3624: out = -10802;
			3625: out = -7886;
			3626: out = -11853;
			3627: out = -5085;
			3628: out = 3734;
			3629: out = 9376;
			3630: out = 6932;
			3631: out = 3078;
			3632: out = -322;
			3633: out = -3388;
			3634: out = -6212;
			3635: out = -5317;
			3636: out = 4041;
			3637: out = 1305;
			3638: out = -616;
			3639: out = 1321;
			3640: out = 7871;
			3641: out = 9393;
			3642: out = 6030;
			3643: out = 10529;
			3644: out = -7785;
			3645: out = -10056;
			3646: out = 1992;
			3647: out = 1047;
			3648: out = -5045;
			3649: out = -11722;
			3650: out = -1977;
			3651: out = -615;
			3652: out = 4179;
			3653: out = 5367;
			3654: out = -212;
			3655: out = -4630;
			3656: out = -4545;
			3657: out = 125;
			3658: out = -2706;
			3659: out = -4806;
			3660: out = -3340;
			3661: out = -2217;
			3662: out = 2760;
			3663: out = 5889;
			3664: out = 6197;
			3665: out = 2017;
			3666: out = -3401;
			3667: out = -8701;
			3668: out = 49;
			3669: out = -3745;
			3670: out = -6505;
			3671: out = -821;
			3672: out = 4399;
			3673: out = 6517;
			3674: out = 3248;
			3675: out = 6945;
			3676: out = 161;
			3677: out = -8117;
			3678: out = -19006;
			3679: out = -4895;
			3680: out = 6576;
			3681: out = 9595;
			3682: out = -5506;
			3683: out = -5154;
			3684: out = -1374;
			3685: out = -1717;
			3686: out = 1270;
			3687: out = 699;
			3688: out = 225;
			3689: out = -171;
			3690: out = 1155;
			3691: out = 590;
			3692: out = -1038;
			3693: out = 332;
			3694: out = 5380;
			3695: out = 10947;
			3696: out = 14405;
			3697: out = 6689;
			3698: out = -2437;
			3699: out = -4920;
			3700: out = -310;
			3701: out = 7445;
			3702: out = 8610;
			3703: out = 655;
			3704: out = -4137;
			3705: out = -1954;
			3706: out = 4863;
			3707: out = 6893;
			3708: out = 2618;
			3709: out = -3219;
			3710: out = -3466;
			3711: out = 199;
			3712: out = 1465;
			3713: out = -2829;
			3714: out = -5468;
			3715: out = -3262;
			3716: out = 1556;
			3717: out = -5349;
			3718: out = 3598;
			3719: out = 8736;
			3720: out = 9217;
			3721: out = -2582;
			3722: out = -4422;
			3723: out = 2449;
			3724: out = 10886;
			3725: out = 11674;
			3726: out = 2383;
			3727: out = -11589;
			3728: out = -8618;
			3729: out = -3466;
			3730: out = 1594;
			3731: out = 236;
			3732: out = 959;
			3733: out = -2956;
			3734: out = -8951;
			3735: out = 6579;
			3736: out = 3266;
			3737: out = -4351;
			3738: out = -5525;
			3739: out = -2130;
			3740: out = 2262;
			3741: out = 1226;
			3742: out = -956;
			3743: out = -3512;
			3744: out = -4429;
			3745: out = -13974;
			3746: out = -2749;
			3747: out = 228;
			3748: out = 141;
			3749: out = -863;
			3750: out = 7024;
			3751: out = 7168;
			3752: out = -7458;
			3753: out = -13094;
			3754: out = -9699;
			3755: out = 2149;
			3756: out = 8506;
			3757: out = 4172;
			3758: out = -4941;
			3759: out = -8705;
			3760: out = -1073;
			3761: out = 6859;
			3762: out = 7236;
			3763: out = 1354;
			3764: out = -3692;
			3765: out = -6935;
			3766: out = -11150;
			3767: out = -5431;
			3768: out = -1766;
			3769: out = 693;
			3770: out = 444;
			3771: out = 4389;
			3772: out = 6959;
			3773: out = 4768;
			3774: out = 5741;
			3775: out = 2800;
			3776: out = -658;
			3777: out = -6561;
			3778: out = -2282;
			3779: out = 3443;
			3780: out = 6028;
			3781: out = 2596;
			3782: out = 445;
			3783: out = 384;
			3784: out = 1280;
			3785: out = 552;
			3786: out = 860;
			3787: out = 3912;
			3788: out = -1831;
			3789: out = -3955;
			3790: out = -3591;
			3791: out = 877;
			3792: out = 4005;
			3793: out = 9796;
			3794: out = 16127;
			3795: out = 2419;
			3796: out = -7520;
			3797: out = -12187;
			3798: out = 671;
			3799: out = 532;
			3800: out = 835;
			3801: out = -359;
			3802: out = 5470;
			3803: out = 3425;
			3804: out = -188;
			3805: out = -7580;
			3806: out = 3504;
			3807: out = 5973;
			3808: out = -4742;
			3809: out = -317;
			3810: out = -218;
			3811: out = 245;
			3812: out = -10535;
			3813: out = -977;
			3814: out = 1279;
			3815: out = -4540;
			3816: out = 7946;
			3817: out = 8461;
			3818: out = 4150;
			3819: out = -8823;
			3820: out = -6426;
			3821: out = -9113;
			3822: out = -17293;
			3823: out = -3196;
			3824: out = 334;
			3825: out = 741;
			3826: out = 3212;
			3827: out = 687;
			3828: out = -57;
			3829: out = 592;
			3830: out = 10763;
			3831: out = 7023;
			3832: out = 1351;
			3833: out = 2968;
			3834: out = -3414;
			3835: out = -8166;
			3836: out = -10519;
			3837: out = -4039;
			3838: out = 4066;
			3839: out = 8513;
			3840: out = 1806;
			3841: out = 3430;
			3842: out = -276;
			3843: out = -4477;
			3844: out = -5481;
			3845: out = -3911;
			3846: out = -1408;
			3847: out = 3167;
			3848: out = 289;
			3849: out = 1530;
			3850: out = 3790;
			3851: out = -910;
			3852: out = -781;
			3853: out = 4301;
			3854: out = 11925;
			3855: out = 8233;
			3856: out = -2151;
			3857: out = -13506;
			3858: out = -7551;
			3859: out = 61;
			3860: out = 6291;
			3861: out = 3934;
			3862: out = -477;
			3863: out = -4304;
			3864: out = -2127;
			3865: out = -7970;
			3866: out = 2726;
			3867: out = 5195;
			3868: out = -6345;
			3869: out = -7451;
			3870: out = -4911;
			3871: out = 3012;
			3872: out = 1717;
			3873: out = 6626;
			3874: out = 6119;
			3875: out = 3796;
			3876: out = -3934;
			3877: out = -6943;
			3878: out = -7109;
			3879: out = 6731;
			3880: out = -3189;
			3881: out = -6979;
			3882: out = 1112;
			3883: out = 12259;
			3884: out = 9267;
			3885: out = -318;
			3886: out = 9296;
			3887: out = 3426;
			3888: out = 1729;
			3889: out = -1495;
			3890: out = -1815;
			3891: out = -7796;
			3892: out = -8583;
			3893: out = 8683;
			3894: out = 6777;
			3895: out = 955;
			3896: out = -5518;
			3897: out = 2786;
			3898: out = 7223;
			3899: out = 5137;
			3900: out = -9379;
			3901: out = -8780;
			3902: out = -4151;
			3903: out = 1013;
			3904: out = -165;
			3905: out = -133;
			3906: out = 2115;
			3907: out = 5512;
			3908: out = 13143;
			3909: out = 14074;
			3910: out = 6240;
			3911: out = -3168;
			3912: out = -12152;
			3913: out = -12424;
			3914: out = -2516;
			3915: out = 3389;
			3916: out = 2208;
			3917: out = -3456;
			3918: out = 3876;
			3919: out = 4751;
			3920: out = 3117;
			3921: out = -2121;
			3922: out = -948;
			3923: out = 213;
			3924: out = 872;
			3925: out = 1922;
			3926: out = 1921;
			3927: out = 1616;
			3928: out = -802;
			3929: out = 2532;
			3930: out = 861;
			3931: out = -3611;
			3932: out = 3826;
			3933: out = 1712;
			3934: out = -3355;
			3935: out = -8528;
			3936: out = -10234;
			3937: out = -7791;
			3938: out = -3754;
			3939: out = -764;
			3940: out = -199;
			3941: out = 1404;
			3942: out = 5822;
			3943: out = 2482;
			3944: out = -1009;
			3945: out = -3915;
			3946: out = -13469;
			3947: out = -8161;
			3948: out = 1554;
			3949: out = 10202;
			3950: out = -2786;
			3951: out = -7730;
			3952: out = -3352;
			3953: out = 3993;
			3954: out = 1476;
			3955: out = -5184;
			3956: out = -5603;
			3957: out = -8654;
			3958: out = -4311;
			3959: out = -362;
			3960: out = 5817;
			3961: out = -518;
			3962: out = -3122;
			3963: out = 662;
			3964: out = 7396;
			3965: out = 5459;
			3966: out = -1331;
			3967: out = -514;
			3968: out = -3303;
			3969: out = -2523;
			3970: out = 1825;
			3971: out = 873;
			3972: out = 3007;
			3973: out = 3634;
			3974: out = 3435;
			3975: out = -3021;
			3976: out = -2402;
			3977: out = 7415;
			3978: out = 14261;
			3979: out = 12419;
			3980: out = 3167;
			3981: out = -7298;
			3982: out = -6128;
			3983: out = -588;
			3984: out = 942;
			3985: out = 8264;
			3986: out = 7372;
			3987: out = 2830;
			3988: out = -12587;
			3989: out = -6534;
			3990: out = -2170;
			3991: out = -2999;
			3992: out = 2715;
			3993: out = 7452;
			3994: out = 10355;
			3995: out = 1218;
			3996: out = 3819;
			3997: out = -1043;
			3998: out = -8817;
			3999: out = -6792;
			4000: out = 1925;
			4001: out = 10641;
			4002: out = 10766;
			4003: out = 6772;
			4004: out = 2024;
			4005: out = 1976;
			4006: out = -3821;
			4007: out = -645;
			4008: out = 2109;
			4009: out = 2836;
			4010: out = -1001;
			4011: out = -3655;
			4012: out = -4825;
			4013: out = -197;
			4014: out = -283;
			4015: out = -704;
			4016: out = -2679;
			4017: out = 2365;
			4018: out = -1062;
			4019: out = -9737;
			4020: out = -8596;
			4021: out = -3813;
			4022: out = 1343;
			4023: out = -2630;
			4024: out = 1800;
			4025: out = 2147;
			4026: out = 1590;
			4027: out = -6387;
			4028: out = -8689;
			4029: out = -8776;
			4030: out = -3186;
			4031: out = -3780;
			4032: out = 2102;
			4033: out = 6779;
			4034: out = 806;
			4035: out = -6047;
			4036: out = -5858;
			4037: out = 9365;
			4038: out = 2392;
			4039: out = 427;
			4040: out = -1997;
			4041: out = -740;
			4042: out = -6323;
			4043: out = -8146;
			4044: out = -1685;
			4045: out = -903;
			4046: out = 2857;
			4047: out = 4232;
			4048: out = -5582;
			4049: out = -5194;
			4050: out = -1298;
			4051: out = 3092;
			4052: out = 4068;
			4053: out = 3088;
			4054: out = 1345;
			4055: out = 140;
			4056: out = 3648;
			4057: out = 7195;
			4058: out = 6433;
			4059: out = 7349;
			4060: out = 6160;
			4061: out = 6730;
			4062: out = 1305;
			4063: out = 7150;
			4064: out = 4245;
			4065: out = -8007;
			4066: out = -10544;
			4067: out = -7393;
			4068: out = 149;
			4069: out = 2736;
			4070: out = 5305;
			4071: out = 3976;
			4072: out = -1012;
			4073: out = 7726;
			4074: out = 4396;
			4075: out = -982;
			4076: out = 1970;
			4077: out = 2898;
			4078: out = -855;
			4079: out = -12118;
			4080: out = -9782;
			4081: out = -5761;
			4082: out = 1497;
			4083: out = 2496;
			4084: out = 7051;
			4085: out = 6472;
			4086: out = 3708;
			4087: out = -4177;
			4088: out = -7604;
			4089: out = -7523;
			4090: out = -1579;
			4091: out = 1220;
			4092: out = 8196;
			4093: out = 15305;
			4094: out = 5808;
			4095: out = -2685;
			4096: out = -9434;
			4097: out = -5228;
			4098: out = -3798;
			4099: out = 314;
			4100: out = 1762;
			4101: out = 3688;
			4102: out = -790;
			4103: out = -7117;
			4104: out = -19619;
			4105: out = -5971;
			4106: out = 6784;
			4107: out = 11039;
			4108: out = 2637;
			4109: out = -1981;
			4110: out = -4849;
			4111: out = -4930;
			4112: out = -5111;
			4113: out = 52;
			4114: out = 5950;
			4115: out = 4170;
			4116: out = -1672;
			4117: out = -4956;
			4118: out = 988;
			4119: out = 7805;
			4120: out = 5266;
			4121: out = -7346;
			4122: out = 1402;
			4123: out = -2195;
			4124: out = -1985;
			4125: out = -499;
			4126: out = 4009;
			4127: out = 3415;
			4128: out = 2148;
			4129: out = -2177;
			4130: out = 3941;
			4131: out = 7259;
			4132: out = 2639;
			4133: out = -1555;
			4134: out = -4893;
			4135: out = -4871;
			4136: out = 5962;
			4137: out = 2686;
			4138: out = -2101;
			4139: out = -5783;
			4140: out = 5027;
			4141: out = 4502;
			4142: out = -3016;
			4143: out = 2287;
			4144: out = 4879;
			4145: out = 6632;
			4146: out = -1179;
			4147: out = 337;
			4148: out = -5203;
			4149: out = -7139;
			4150: out = 4147;
			4151: out = 7907;
			4152: out = 5668;
			4153: out = -1012;
			4154: out = -152;
			4155: out = 402;
			4156: out = -282;
			4157: out = -4426;
			4158: out = -5933;
			4159: out = -5841;
			4160: out = -6097;
			4161: out = -3247;
			4162: out = -5081;
			4163: out = -5739;
			4164: out = 2988;
			4165: out = 2371;
			4166: out = -3736;
			4167: out = -13801;
			4168: out = -8177;
			4169: out = -2683;
			4170: out = 374;
			4171: out = -2389;
			4172: out = -1069;
			4173: out = 625;
			4174: out = -263;
			4175: out = 7969;
			4176: out = 2387;
			4177: out = -6016;
			4178: out = -12990;
			4179: out = 1306;
			4180: out = 8679;
			4181: out = -380;
			4182: out = 5261;
			4183: out = -2121;
			4184: out = -5765;
			4185: out = -6;
			4186: out = -829;
			4187: out = 812;
			4188: out = 6935;
			4189: out = 2286;
			4190: out = 2492;
			4191: out = 656;
			4192: out = 7168;
			4193: out = -10748;
			4194: out = -14401;
			4195: out = -4133;
			4196: out = 8556;
			4197: out = 5471;
			4198: out = -751;
			4199: out = 4551;
			4200: out = 2750;
			4201: out = -766;
			4202: out = -8183;
			4203: out = 993;
			4204: out = 6590;
			4205: out = 11720;
			4206: out = 6393;
			4207: out = 12020;
			4208: out = 4435;
			4209: out = -6032;
			4210: out = 3457;
			4211: out = 8414;
			4212: out = 10451;
			4213: out = 3854;
			4214: out = 1490;
			4215: out = -4952;
			4216: out = -7469;
			4217: out = 1296;
			4218: out = 7031;
			4219: out = 4613;
			4220: out = -6173;
			4221: out = -2732;
			4222: out = 1369;
			4223: out = 1959;
			4224: out = 14;
			4225: out = -6476;
			4226: out = -6526;
			4227: out = 378;
			4228: out = 7923;
			4229: out = 5477;
			4230: out = -1276;
			4231: out = -7099;
			4232: out = 229;
			4233: out = 5978;
			4234: out = 4336;
			4235: out = -6927;
			4236: out = -6782;
			4237: out = 1524;
			4238: out = -2758;
			4239: out = -3237;
			4240: out = -3889;
			4241: out = 1103;
			4242: out = 349;
			4243: out = 595;
			4244: out = -2373;
			4245: out = -10081;
			4246: out = -9726;
			4247: out = -5209;
			4248: out = 1136;
			4249: out = -5499;
			4250: out = -3427;
			4251: out = 1506;
			4252: out = -2904;
			4253: out = -3007;
			4254: out = -3685;
			4255: out = -1845;
			4256: out = 708;
			4257: out = 1986;
			4258: out = 647;
			4259: out = 927;
			4260: out = -374;
			4261: out = 1758;
			4262: out = 4864;
			4263: out = 5871;
			4264: out = 2982;
			4265: out = -321;
			4266: out = 1493;
			4267: out = 1053;
			4268: out = 870;
			4269: out = -311;
			4270: out = 5829;
			4271: out = 5763;
			4272: out = 2920;
			4273: out = -1616;
			4274: out = -5988;
			4275: out = -10339;
			4276: out = -12074;
			4277: out = 4748;
			4278: out = 9773;
			4279: out = 6057;
			4280: out = 375;
			4281: out = -5747;
			4282: out = -3272;
			4283: out = 3990;
			4284: out = 3598;
			4285: out = -1813;
			4286: out = -5886;
			4287: out = 5358;
			4288: out = 2265;
			4289: out = 2093;
			4290: out = 382;
			4291: out = 6512;
			4292: out = 3120;
			4293: out = -133;
			4294: out = -4627;
			4295: out = 4761;
			4296: out = 5532;
			4297: out = -539;
			4298: out = 1049;
			4299: out = 1202;
			4300: out = 827;
			4301: out = -4783;
			4302: out = -1447;
			4303: out = 353;
			4304: out = 714;
			4305: out = 4274;
			4306: out = -2851;
			4307: out = -9246;
			4308: out = -4575;
			4309: out = -603;
			4310: out = 5087;
			4311: out = 5150;
			4312: out = 1648;
			4313: out = -2751;
			4314: out = -1289;
			4315: out = 2469;
			4316: out = 1580;
			4317: out = -7439;
			4318: out = -16070;
			4319: out = -6577;
			4320: out = 2632;
			4321: out = 6416;
			4322: out = 1886;
			4323: out = 279;
			4324: out = 3050;
			4325: out = 6686;
			4326: out = -7407;
			4327: out = -7005;
			4328: out = -2304;
			4329: out = 4474;
			4330: out = 2251;
			4331: out = -3441;
			4332: out = -9335;
			4333: out = -5138;
			4334: out = 139;
			4335: out = 5770;
			4336: out = 6971;
			4337: out = -2128;
			4338: out = -7648;
			4339: out = -6136;
			4340: out = -973;
			4341: out = 1504;
			4342: out = 2694;
			4343: out = 8431;
			4344: out = -5871;
			4345: out = -4480;
			4346: out = 1863;
			4347: out = 6613;
			4348: out = 2226;
			4349: out = 1428;
			4350: out = 7131;
			4351: out = 5480;
			4352: out = 2113;
			4353: out = -2506;
			4354: out = 330;
			4355: out = -1563;
			4356: out = -1387;
			4357: out = -140;
			4358: out = 5204;
			4359: out = 7034;
			4360: out = 3226;
			4361: out = -9981;
			4362: out = -12367;
			4363: out = -8535;
			4364: out = -157;
			4365: out = 11402;
			4366: out = 8103;
			4367: out = -2710;
			4368: out = -7544;
			4369: out = -11513;
			4370: out = -6070;
			4371: out = 23;
			4372: out = 6148;
			4373: out = -2577;
			4374: out = -9587;
			4375: out = 2295;
			4376: out = 420;
			4377: out = -650;
			4378: out = -3855;
			4379: out = 1120;
			4380: out = 768;
			4381: out = 3858;
			4382: out = 14273;
			4383: out = 7224;
			4384: out = -73;
			4385: out = -7054;
			4386: out = -1480;
			4387: out = -5224;
			4388: out = -5060;
			4389: out = 9436;
			4390: out = 5767;
			4391: out = 4960;
			4392: out = 1922;
			4393: out = -3718;
			4394: out = -9363;
			4395: out = -6189;
			4396: out = 8912;
			4397: out = 7887;
			4398: out = 4014;
			4399: out = -3452;
			4400: out = -9030;
			4401: out = -8701;
			4402: out = -354;
			4403: out = 9096;
			4404: out = 9380;
			4405: out = 3729;
			4406: out = -2086;
			4407: out = -294;
			4408: out = 1345;
			4409: out = 1793;
			4410: out = 1023;
			4411: out = -599;
			4412: out = 1054;
			4413: out = 3508;
			4414: out = 6262;
			4415: out = -238;
			4416: out = -6272;
			4417: out = -7372;
			4418: out = 6280;
			4419: out = 10626;
			4420: out = 5648;
			4421: out = 1467;
			4422: out = -5937;
			4423: out = -7744;
			4424: out = -3925;
			4425: out = -1660;
			4426: out = 445;
			4427: out = 765;
			4428: out = 2230;
			4429: out = -1530;
			4430: out = -2466;
			4431: out = 760;
			4432: out = 739;
			4433: out = 321;
			4434: out = -95;
			4435: out = 1873;
			4436: out = 466;
			4437: out = -2236;
			4438: out = -4163;
			4439: out = -6713;
			4440: out = -3474;
			4441: out = 1228;
			4442: out = 5233;
			4443: out = -1430;
			4444: out = -7879;
			4445: out = -9407;
			4446: out = 209;
			4447: out = 4508;
			4448: out = 2819;
			4449: out = -4790;
			4450: out = -4453;
			4451: out = -3139;
			4452: out = -2455;
			4453: out = -2417;
			4454: out = -2897;
			4455: out = -2864;
			4456: out = 3217;
			4457: out = 1050;
			4458: out = 2560;
			4459: out = 2749;
			4460: out = -407;
			4461: out = -10399;
			4462: out = -11529;
			4463: out = 8967;
			4464: out = 12164;
			4465: out = 6946;
			4466: out = -5234;
			4467: out = -6688;
			4468: out = -3430;
			4469: out = 2795;
			4470: out = 1919;
			4471: out = 1535;
			4472: out = -415;
			4473: out = 555;
			4474: out = 2014;
			4475: out = 2255;
			4476: out = 1550;
			4477: out = 4980;
			4478: out = 3431;
			4479: out = 2015;
			4480: out = -1924;
			4481: out = 4868;
			4482: out = 547;
			4483: out = -1271;
			4484: out = -597;
			4485: out = 5393;
			4486: out = 4291;
			4487: out = 985;
			4488: out = 2623;
			4489: out = 6024;
			4490: out = 5134;
			4491: out = -835;
			4492: out = -12655;
			4493: out = -12546;
			4494: out = -1010;
			4495: out = 6810;
			4496: out = 4785;
			4497: out = -1237;
			4498: out = 558;
			4499: out = -4292;
			4500: out = 282;
			4501: out = 5177;
			4502: out = -2596;
			4503: out = -1499;
			4504: out = -422;
			4505: out = -1758;
			4506: out = 410;
			4507: out = -143;
			4508: out = -1097;
			4509: out = 6333;
			4510: out = 3551;
			4511: out = 1036;
			4512: out = -1817;
			4513: out = 9037;
			4514: out = 5456;
			4515: out = -4968;
			4516: out = -751;
			4517: out = -5004;
			4518: out = -3191;
			4519: out = 2029;
			4520: out = -789;
			4521: out = -3227;
			4522: out = -3352;
			4523: out = 297;
			4524: out = 2425;
			4525: out = 4222;
			4526: out = 6807;
			4527: out = -7116;
			4528: out = -12007;
			4529: out = -9779;
			4530: out = -1838;
			4531: out = -320;
			4532: out = 3736;
			4533: out = 13353;
			4534: out = -21;
			4535: out = -237;
			4536: out = 2273;
			4537: out = -278;
			4538: out = -1067;
			4539: out = -892;
			4540: out = 2475;
			4541: out = -3547;
			4542: out = -673;
			4543: out = 3591;
			4544: out = -651;
			4545: out = 3076;
			4546: out = 3922;
			4547: out = 2520;
			4548: out = -3932;
			4549: out = -6445;
			4550: out = -5715;
			4551: out = -2862;
			4552: out = 51;
			4553: out = 1180;
			4554: out = -509;
			4555: out = 5951;
			4556: out = 2951;
			4557: out = -1152;
			4558: out = 293;
			4559: out = -1462;
			4560: out = 86;
			4561: out = 4605;
			4562: out = -624;
			4563: out = 327;
			4564: out = -1594;
			4565: out = -9744;
			4566: out = -6211;
			4567: out = 3747;
			4568: out = 11632;
			4569: out = 10714;
			4570: out = 587;
			4571: out = -8287;
			4572: out = -7671;
			4573: out = -2562;
			4574: out = -1630;
			4575: out = -5210;
			4576: out = 287;
			4577: out = 6432;
			4578: out = 9209;
			4579: out = 2465;
			4580: out = -2138;
			4581: out = -4114;
			4582: out = -1337;
			4583: out = -2952;
			4584: out = -6675;
			4585: out = -9989;
			4586: out = -2749;
			4587: out = -5461;
			4588: out = -1197;
			4589: out = 4449;
			4590: out = 7060;
			4591: out = 7035;
			4592: out = 5365;
			4593: out = 3026;
			4594: out = 1259;
			4595: out = -1013;
			4596: out = -3563;
			4597: out = -7262;
			4598: out = -3982;
			4599: out = 2493;
			4600: out = 5845;
			4601: out = 9828;
			4602: out = 6334;
			4603: out = 288;
			4604: out = -7258;
			4605: out = -6071;
			4606: out = -2172;
			4607: out = 2295;
			4608: out = -4182;
			4609: out = -1068;
			4610: out = 6060;
			4611: out = 451;
			4612: out = 387;
			4613: out = -22;
			4614: out = 4810;
			4615: out = -208;
			4616: out = 182;
			4617: out = -1275;
			4618: out = -1882;
			4619: out = -9458;
			4620: out = -6636;
			4621: out = 8615;
			4622: out = 6663;
			4623: out = 5569;
			4624: out = 2078;
			4625: out = 3424;
			4626: out = 80;
			4627: out = -1199;
			4628: out = -1967;
			4629: out = 2419;
			4630: out = 1390;
			4631: out = -710;
			4632: out = 877;
			4633: out = 496;
			4634: out = 697;
			4635: out = -1;
			4636: out = -553;
			4637: out = -1583;
			4638: out = -2848;
			4639: out = -9227;
			4640: out = -3179;
			4641: out = 418;
			4642: out = 170;
			4643: out = -3300;
			4644: out = -2736;
			4645: out = 2300;
			4646: out = 12333;
			4647: out = 3353;
			4648: out = -3649;
			4649: out = -4912;
			4650: out = -4730;
			4651: out = -1340;
			4652: out = 1125;
			4653: out = 1979;
			4654: out = -549;
			4655: out = -1785;
			4656: out = 21;
			4657: out = -13;
			4658: out = 2370;
			4659: out = 3059;
			4660: out = 4236;
			4661: out = -423;
			4662: out = -4315;
			4663: out = -9291;
			4664: out = 944;
			4665: out = -3895;
			4666: out = -3879;
			4667: out = 3999;
			4668: out = 9067;
			4669: out = 758;
			4670: out = -14078;
			4671: out = -12405;
			4672: out = -4645;
			4673: out = 3598;
			4674: out = 4116;
			4675: out = -2352;
			4676: out = -3122;
			4677: out = 2756;
			4678: out = 3971;
			4679: out = 2704;
			4680: out = 1237;
			4681: out = 4746;
			4682: out = 6619;
			4683: out = 4393;
			4684: out = -1282;
			4685: out = 1374;
			4686: out = 710;
			4687: out = 1037;
			4688: out = 1001;
			4689: out = 1364;
			4690: out = 5093;
			4691: out = 7842;
			4692: out = -1367;
			4693: out = -6407;
			4694: out = -8422;
			4695: out = -3173;
			4696: out = -777;
			4697: out = 2375;
			4698: out = 3194;
			4699: out = 6153;
			4700: out = 1724;
			4701: out = -1916;
			4702: out = -2634;
			4703: out = 7;
			4704: out = 250;
			4705: out = -2332;
			4706: out = 1229;
			4707: out = -3844;
			4708: out = -3434;
			4709: out = 1380;
			4710: out = 8584;
			4711: out = 5784;
			4712: out = -450;
			4713: out = 845;
			4714: out = -1420;
			4715: out = -1765;
			4716: out = -575;
			4717: out = -3976;
			4718: out = -1844;
			4719: out = 405;
			4720: out = -1497;
			4721: out = -1392;
			4722: out = 4755;
			4723: out = 13882;
			4724: out = -345;
			4725: out = -9978;
			4726: out = -15497;
			4727: out = -9879;
			4728: out = -3241;
			4729: out = 3036;
			4730: out = 5622;
			4731: out = -8623;
			4732: out = -6694;
			4733: out = 2897;
			4734: out = 2080;
			4735: out = 3127;
			4736: out = 170;
			4737: out = 3239;
			4738: out = -11001;
			4739: out = 0;
			4740: out = 9768;
			4741: out = 3864;
			4742: out = 40;
			4743: out = 1245;
			4744: out = 8917;
			4745: out = 8999;
			4746: out = 4672;
			4747: out = -4097;
			4748: out = -10645;
			4749: out = -9491;
			4750: out = -5812;
			4751: out = -4899;
			4752: out = 63;
			4753: out = 367;
			4754: out = 1890;
			4755: out = 3989;
			4756: out = 1815;
			4757: out = -4386;
			4758: out = -10184;
			4759: out = 5967;
			4760: out = 4814;
			4761: out = -2204;
			4762: out = -10287;
			4763: out = -5383;
			4764: out = 2432;
			4765: out = 6309;
			4766: out = 6030;
			4767: out = -93;
			4768: out = -3514;
			4769: out = 247;
			4770: out = 3284;
			4771: out = 3146;
			4772: out = -1330;
			4773: out = -483;
			4774: out = -4216;
			4775: out = -1294;
			4776: out = 10576;
			4777: out = 10704;
			4778: out = 9563;
			4779: out = 4066;
			4780: out = 4178;
			4781: out = -7963;
			4782: out = -14393;
			4783: out = -9194;
			4784: out = -3429;
			4785: out = -1072;
			4786: out = -2586;
			4787: out = 1003;
			4788: out = 2947;
			4789: out = 3536;
			4790: out = -2066;
			4791: out = 4716;
			4792: out = 2911;
			4793: out = -485;
			4794: out = -271;
			4795: out = 191;
			4796: out = 606;
			4797: out = 126;
			4798: out = 3919;
			4799: out = 8213;
			4800: out = 10583;
			4801: out = 3362;
			4802: out = 1253;
			4803: out = -4303;
			4804: out = -9852;
			4805: out = -5770;
			4806: out = 183;
			4807: out = 1941;
			4808: out = -4577;
			4809: out = -5134;
			4810: out = 82;
			4811: out = 6778;
			4812: out = 2127;
			4813: out = -5718;
			4814: out = -10249;
			4815: out = -430;
			4816: out = 1745;
			4817: out = 520;
			4818: out = -4051;
			4819: out = -5787;
			4820: out = -1596;
			4821: out = 5892;
			4822: out = 11842;
			4823: out = 3055;
			4824: out = -3346;
			4825: out = -709;
			4826: out = -7595;
			4827: out = -3005;
			4828: out = 2705;
			4829: out = 8832;
			4830: out = 2178;
			4831: out = -2033;
			4832: out = -1900;
			4833: out = 6545;
			4834: out = 5771;
			4835: out = 1200;
			4836: out = -117;
			4837: out = -2116;
			4838: out = -1329;
			4839: out = -2375;
			4840: out = -877;
			4841: out = -6612;
			4842: out = -8983;
			4843: out = -3523;
			4844: out = 3183;
			4845: out = 4072;
			4846: out = -985;
			4847: out = -642;
			4848: out = -4279;
			4849: out = -6181;
			4850: out = -5504;
			4851: out = 37;
			4852: out = 4981;
			4853: out = 5527;
			4854: out = 4331;
			4855: out = -3307;
			4856: out = -6170;
			4857: out = 718;
			4858: out = 6240;
			4859: out = 6377;
			4860: out = 602;
			4861: out = -1536;
			4862: out = -4026;
			4863: out = -1722;
			4864: out = 3182;
			4865: out = 909;
			4866: out = -1285;
			4867: out = -2340;
			4868: out = 32;
			4869: out = 47;
			4870: out = 624;
			4871: out = 2128;
			4872: out = -550;
			4873: out = -1895;
			4874: out = -656;
			4875: out = 580;
			4876: out = 4671;
			4877: out = 5783;
			4878: out = 4694;
			4879: out = -7052;
			4880: out = -7901;
			4881: out = 678;
			4882: out = 10881;
			4883: out = 7803;
			4884: out = -385;
			4885: out = -5578;
			4886: out = -2647;
			4887: out = 5824;
			4888: out = 10504;
			4889: out = 3562;
			4890: out = 2254;
			4891: out = 943;
			4892: out = 71;
			4893: out = -478;
			4894: out = -586;
			4895: out = -1592;
			4896: out = -8703;
			4897: out = -5314;
			4898: out = 791;
			4899: out = 7674;
			4900: out = 138;
			4901: out = -2495;
			4902: out = -3880;
			4903: out = 2513;
			4904: out = -7447;
			4905: out = -10476;
			4906: out = -4746;
			4907: out = 6773;
			4908: out = 5515;
			4909: out = -1689;
			4910: out = -4139;
			4911: out = 501;
			4912: out = 6394;
			4913: out = 5549;
			4914: out = 4334;
			4915: out = -3741;
			4916: out = -9105;
			4917: out = -7146;
			4918: out = -2429;
			4919: out = 2819;
			4920: out = 5317;
			4921: out = -4570;
			4922: out = -6855;
			4923: out = -4253;
			4924: out = 606;
			4925: out = 2945;
			4926: out = 2094;
			4927: out = -771;
			4928: out = -2996;
			4929: out = -3088;
			4930: out = -1912;
			4931: out = -2473;
			4932: out = -375;
			4933: out = -41;
			4934: out = 0;
			4935: out = -2224;
			4936: out = -228;
			4937: out = 900;
			4938: out = -1128;
			4939: out = 60;
			4940: out = 945;
			4941: out = 1571;
			4942: out = 4370;
			4943: out = 2265;
			4944: out = 1368;
			4945: out = 4345;
			4946: out = 849;
			4947: out = -1235;
			4948: out = -384;
			4949: out = 4151;
			4950: out = 7719;
			4951: out = 7084;
			4952: out = 3669;
			4953: out = -7763;
			4954: out = -8455;
			4955: out = 800;
			4956: out = 2505;
			4957: out = 7138;
			4958: out = 5172;
			4959: out = -798;
			4960: out = -3297;
			4961: out = -3605;
			4962: out = -1801;
			4963: out = 3391;
			4964: out = 4067;
			4965: out = 2343;
			4966: out = -1960;
			4967: out = 432;
			4968: out = 729;
			4969: out = 1108;
			4970: out = 3373;
			4971: out = 3773;
			4972: out = 2791;
			4973: out = 1589;
			4974: out = 336;
			4975: out = 2320;
			4976: out = 3668;
			4977: out = -2782;
			4978: out = -5679;
			4979: out = -3211;
			4980: out = 8173;
			4981: out = 1518;
			4982: out = 1847;
			4983: out = 92;
			4984: out = -2030;
			4985: out = -12363;
			4986: out = -12990;
			4987: out = 1230;
			4988: out = -1077;
			4989: out = -1008;
			4990: out = -2634;
			4991: out = 3513;
			4992: out = -1149;
			4993: out = -2757;
			4994: out = -2510;
			4995: out = 3261;
			4996: out = 2051;
			4997: out = -1615;
			4998: out = -5840;
			4999: out = -2;
			5000: out = 3070;
			5001: out = -1263;
			5002: out = 1126;
			5003: out = -372;
			5004: out = -426;
			5005: out = -4203;
			5006: out = 4559;
			5007: out = 5995;
			5008: out = -1484;
			5009: out = -3353;
			5010: out = -6852;
			5011: out = -5613;
			5012: out = -402;
			5013: out = -208;
			5014: out = -3991;
			5015: out = -7603;
			5016: out = -1525;
			5017: out = 1537;
			5018: out = 1048;
			5019: out = 5256;
			5020: out = -8600;
			5021: out = -9640;
			5022: out = 3100;
			5023: out = 3153;
			5024: out = 6125;
			5025: out = 5139;
			5026: out = 2350;
			5027: out = 323;
			5028: out = 285;
			5029: out = 2411;
			5030: out = -3634;
			5031: out = 1874;
			5032: out = 5826;
			5033: out = 589;
			5034: out = -2395;
			5035: out = -1138;
			5036: out = 5596;
			5037: out = -4728;
			5038: out = -2794;
			5039: out = -480;
			5040: out = 3534;
			5041: out = 945;
			5042: out = 3440;
			5043: out = 6401;
			5044: out = 1467;
			5045: out = -2764;
			5046: out = -4737;
			5047: out = -1095;
			5048: out = 774;
			5049: out = 4231;
			5050: out = 6179;
			5051: out = 55;
			5052: out = -1134;
			5053: out = -1968;
			5054: out = -1331;
			5055: out = 659;
			5056: out = 3233;
			5057: out = 3508;
			5058: out = 8790;
			5059: out = -1943;
			5060: out = -6622;
			5061: out = 2728;
			5062: out = 6391;
			5063: out = 5547;
			5064: out = -485;
			5065: out = 6921;
			5066: out = 1205;
			5067: out = -2253;
			5068: out = -7195;
			5069: out = -1404;
			5070: out = -3056;
			5071: out = -4822;
			5072: out = -1371;
			5073: out = 2667;
			5074: out = 708;
			5075: out = -7959;
			5076: out = -7565;
			5077: out = -3213;
			5078: out = 3176;
			5079: out = 3250;
			5080: out = 53;
			5081: out = -3943;
			5082: out = -1855;
			5083: out = -5422;
			5084: out = -714;
			5085: out = 3731;
			5086: out = 5704;
			5087: out = 2195;
			5088: out = -891;
			5089: out = -2807;
			5090: out = 208;
			5091: out = -163;
			5092: out = -383;
			5093: out = -1003;
			5094: out = 7261;
			5095: out = 6681;
			5096: out = -4561;
			5097: out = -3944;
			5098: out = -4765;
			5099: out = -2060;
			5100: out = -6976;
			5101: out = 3905;
			5102: out = 5204;
			5103: out = 300;
			5104: out = -204;
			5105: out = 2929;
			5106: out = 4248;
			5107: out = -6548;
			5108: out = -1428;
			5109: out = 2723;
			5110: out = 5532;
			5111: out = 3043;
			5112: out = -1923;
			5113: out = -6392;
			5114: out = 448;
			5115: out = -2339;
			5116: out = 781;
			5117: out = 2305;
			5118: out = 3598;
			5119: out = -1552;
			5120: out = -4549;
			5121: out = -10206;
			5122: out = 1680;
			5123: out = 1646;
			5124: out = -3259;
			5125: out = -16611;
			5126: out = -2776;
			5127: out = 8668;
			5128: out = 314;
			5129: out = -2323;
			5130: out = 2250;
			5131: out = 12205;
			5132: out = 1116;
			5133: out = -5835;
			5134: out = -8303;
			5135: out = 6210;
			5136: out = 1527;
			5137: out = -1732;
			5138: out = -6779;
			5139: out = 5032;
			5140: out = 1965;
			5141: out = -187;
			5142: out = 1056;
			5143: out = -398;
			5144: out = 560;
			5145: out = 919;
			5146: out = 2537;
			5147: out = -3070;
			5148: out = -4869;
			5149: out = 185;
			5150: out = 4039;
			5151: out = 3523;
			5152: out = 544;
			5153: out = 1093;
			5154: out = 1562;
			5155: out = 2871;
			5156: out = 6864;
			5157: out = -6076;
			5158: out = -4430;
			5159: out = 3245;
			5160: out = 3409;
			5161: out = 370;
			5162: out = 115;
			5163: out = 7813;
			5164: out = 629;
			5165: out = -1697;
			5166: out = -2710;
			5167: out = -1842;
			5168: out = 1284;
			5169: out = 3608;
			5170: out = 5269;
			5171: out = -4527;
			5172: out = -4003;
			5173: out = 1125;
			5174: out = 5244;
			5175: out = -2753;
			5176: out = -6793;
			5177: out = 1081;
			5178: out = -5046;
			5179: out = -2839;
			5180: out = -1644;
			5181: out = -2288;
			5182: out = 122;
			5183: out = 3335;
			5184: out = 3308;
			5185: out = 5916;
			5186: out = 2374;
			5187: out = -1802;
			5188: out = -9384;
			5189: out = -4741;
			5190: out = -698;
			5191: out = 2405;
			5192: out = -445;
			5193: out = 3329;
			5194: out = 4658;
			5195: out = -197;
			5196: out = -5568;
			5197: out = -5112;
			5198: out = 277;
			5199: out = 5246;
			5200: out = 1608;
			5201: out = -4719;
			5202: out = -11623;
			5203: out = 876;
			5204: out = 6737;
			5205: out = 2178;
			5206: out = -8103;
			5207: out = -8090;
			5208: out = 1218;
			5209: out = 11869;
			5210: out = 2282;
			5211: out = -6794;
			5212: out = -9162;
			5213: out = -577;
			5214: out = 1166;
			5215: out = -314;
			5216: out = 2893;
			5217: out = -730;
			5218: out = -671;
			5219: out = -125;
			5220: out = 998;
			5221: out = 802;
			5222: out = 2606;
			5223: out = 6575;
			5224: out = 4188;
			5225: out = -352;
			5226: out = -4343;
			5227: out = 4318;
			5228: out = 3881;
			5229: out = 2273;
			5230: out = 1940;
			5231: out = 630;
			5232: out = 582;
			5233: out = 275;
			5234: out = -5618;
			5235: out = -550;
			5236: out = 4591;
			5237: out = -441;
			5238: out = 6461;
			5239: out = 2439;
			5240: out = -2679;
			5241: out = -13168;
			5242: out = 57;
			5243: out = 8816;
			5244: out = 1215;
			5245: out = -653;
			5246: out = -4654;
			5247: out = -3143;
			5248: out = 4724;
			5249: out = 6487;
			5250: out = 4695;
			5251: out = 90;
			5252: out = 1152;
			5253: out = -3020;
			5254: out = -7857;
			5255: out = -9304;
			5256: out = -2214;
			5257: out = 3062;
			5258: out = 1119;
			5259: out = -5797;
			5260: out = -5724;
			5261: out = 1945;
			5262: out = 1579;
			5263: out = 6679;
			5264: out = 3351;
			5265: out = -2797;
			5266: out = -13546;
			5267: out = -11139;
			5268: out = -1490;
			5269: out = 3295;
			5270: out = 7186;
			5271: out = 5590;
			5272: out = 43;
			5273: out = -1511;
			5274: out = -1930;
			5275: out = 200;
			5276: out = -5353;
			5277: out = 4293;
			5278: out = 4860;
			5279: out = -151;
			5280: out = -3622;
			5281: out = 4120;
			5282: out = 9977;
			5283: out = -479;
			5284: out = -5456;
			5285: out = -6325;
			5286: out = 1311;
			5287: out = -709;
			5288: out = 1661;
			5289: out = 500;
			5290: out = -7828;
			5291: out = -2323;
			5292: out = 101;
			5293: out = -867;
			5294: out = 4929;
			5295: out = 8276;
			5296: out = 5395;
			5297: out = -11448;
			5298: out = -11149;
			5299: out = -3883;
			5300: out = 7945;
			5301: out = -1175;
			5302: out = 347;
			5303: out = 2820;
			5304: out = 10455;
			5305: out = 1892;
			5306: out = 1275;
			5307: out = 4831;
			5308: out = 788;
			5309: out = -3541;
			5310: out = -7457;
			5311: out = -3573;
			5312: out = -613;
			5313: out = 7484;
			5314: out = 12102;
			5315: out = 7110;
			5316: out = -653;
			5317: out = -4931;
			5318: out = -201;
			5319: out = -1542;
			5320: out = -3595;
			5321: out = -6778;
			5322: out = 2751;
			5323: out = -769;
			5324: out = -5336;
			5325: out = -8682;
			5326: out = -2114;
			5327: out = 2959;
			5328: out = 4774;
			5329: out = 3993;
			5330: out = 2148;
			5331: out = -1029;
			5332: out = -6965;
			5333: out = -648;
			5334: out = 991;
			5335: out = -1036;
			5336: out = -8245;
			5337: out = -3880;
			5338: out = 3979;
			5339: out = 8499;
			5340: out = 2174;
			5341: out = -4099;
			5342: out = -6627;
			5343: out = -9189;
			5344: out = -619;
			5345: out = 2996;
			5346: out = -2764;
			5347: out = 212;
			5348: out = -529;
			5349: out = -1171;
			5350: out = -4104;
			5351: out = -635;
			5352: out = 2111;
			5353: out = 2183;
			5354: out = -1123;
			5355: out = 86;
			5356: out = 3203;
			5357: out = -9388;
			5358: out = 4973;
			5359: out = 9050;
			5360: out = 1115;
			5361: out = 1022;
			5362: out = 1619;
			5363: out = 5334;
			5364: out = 7781;
			5365: out = 2070;
			5366: out = -2813;
			5367: out = -210;
			5368: out = -1810;
			5369: out = 7440;
			5370: out = 11254;
			5371: out = -4273;
			5372: out = -1356;
			5373: out = 431;
			5374: out = 3145;
			5375: out = 2060;
			5376: out = 3277;
			5377: out = 188;
			5378: out = -7195;
			5379: out = -10581;
			5380: out = -4665;
			5381: out = 5406;
			5382: out = 3147;
			5383: out = -1147;
			5384: out = -4155;
			5385: out = 884;
			5386: out = 3191;
			5387: out = 293;
			5388: out = -8383;
			5389: out = 981;
			5390: out = 119;
			5391: out = 1175;
			5392: out = 6474;
			5393: out = 9798;
			5394: out = 8961;
			5395: out = 2737;
			5396: out = 3717;
			5397: out = -4188;
			5398: out = -7820;
			5399: out = -4874;
			5400: out = -267;
			5401: out = -2907;
			5402: out = -8810;
			5403: out = -1298;
			5404: out = 6260;
			5405: out = 9250;
			5406: out = 701;
			5407: out = -5526;
			5408: out = -11651;
			5409: out = -11055;
			5410: out = -6610;
			5411: out = -582;
			5412: out = 1472;
			5413: out = 1527;
			5414: out = -1504;
			5415: out = 351;
			5416: out = 3782;
			5417: out = -9140;
			5418: out = -2881;
			5419: out = 4012;
			5420: out = 1355;
			5421: out = 5418;
			5422: out = 2069;
			5423: out = -1417;
			5424: out = -5393;
			5425: out = 1200;
			5426: out = 5559;
			5427: out = 3639;
			5428: out = 1600;
			5429: out = 4158;
			5430: out = 8250;
			5431: out = -6587;
			5432: out = -2459;
			5433: out = -2764;
			5434: out = -15177;
			5435: out = 3693;
			5436: out = 7847;
			5437: out = 4176;
			5438: out = -1583;
			5439: out = -548;
			5440: out = 80;
			5441: out = -4667;
			5442: out = -727;
			5443: out = 2527;
			5444: out = 5802;
			5445: out = -259;
			5446: out = 1124;
			5447: out = 884;
			5448: out = 2446;
			5449: out = -2264;
			5450: out = 1832;
			5451: out = 6950;
			5452: out = 5994;
			5453: out = 2076;
			5454: out = -1008;
			5455: out = -42;
			5456: out = 4839;
			5457: out = 4051;
			5458: out = -1375;
			5459: out = -1802;
			5460: out = -2299;
			5461: out = 2960;
			5462: out = 6972;
			5463: out = 6806;
			5464: out = 36;
			5465: out = -6620;
			5466: out = -11591;
			5467: out = -6647;
			5468: out = -134;
			5469: out = 6427;
			5470: out = -4828;
			5471: out = -3456;
			5472: out = 1242;
			5473: out = 10557;
			5474: out = -2981;
			5475: out = -7800;
			5476: out = -3023;
			5477: out = 479;
			5478: out = -6743;
			5479: out = -11970;
			5480: out = 5363;
			5481: out = 10142;
			5482: out = 10496;
			5483: out = 2604;
			5484: out = -275;
			5485: out = -1572;
			5486: out = 652;
			5487: out = -3492;
			5488: out = -346;
			5489: out = -686;
			5490: out = -455;
			5491: out = -3740;
			5492: out = -1561;
			5493: out = -60;
			5494: out = -562;
			5495: out = -4962;
			5496: out = -7645;
			5497: out = -7164;
			5498: out = -7844;
			5499: out = -3547;
			5500: out = -887;
			5501: out = -4316;
			5502: out = -4386;
			5503: out = -4493;
			5504: out = -1959;
			5505: out = -4430;
			5506: out = 3588;
			5507: out = 7250;
			5508: out = -218;
			5509: out = -477;
			5510: out = -3623;
			5511: out = -3229;
			5512: out = 8240;
			5513: out = 9981;
			5514: out = 6561;
			5515: out = 362;
			5516: out = 3374;
			5517: out = 9060;
			5518: out = 12111;
			5519: out = -6099;
			5520: out = -6133;
			5521: out = -6364;
			5522: out = -9652;
			5523: out = -1590;
			5524: out = 4474;
			5525: out = 5502;
			5526: out = -2549;
			5527: out = -1762;
			5528: out = -592;
			5529: out = -7368;
			5530: out = 7295;
			5531: out = 489;
			5532: out = -10874;
			5533: out = -8229;
			5534: out = 3549;
			5535: out = 9733;
			5536: out = -431;
			5537: out = 7163;
			5538: out = 3280;
			5539: out = 646;
			5540: out = 55;
			5541: out = -58;
			5542: out = 2606;
			5543: out = 11788;
			5544: out = -4187;
			5545: out = -2119;
			5546: out = 2012;
			5547: out = -1264;
			5548: out = -923;
			5549: out = 2437;
			5550: out = 6119;
			5551: out = 10236;
			5552: out = 1994;
			5553: out = -7478;
			5554: out = -7520;
			5555: out = -1598;
			5556: out = -3272;
			5557: out = -17774;
			5558: out = 1337;
			5559: out = 5489;
			5560: out = 6680;
			5561: out = -982;
			5562: out = 4529;
			5563: out = 4437;
			5564: out = 1955;
			5565: out = -13842;
			5566: out = -9559;
			5567: out = 3621;
			5568: out = 10626;
			5569: out = 10387;
			5570: out = 4476;
			5571: out = -459;
			5572: out = -4501;
			5573: out = 658;
			5574: out = 6619;
			5575: out = 5938;
			5576: out = 3485;
			5577: out = -654;
			5578: out = -1934;
			5579: out = -14371;
			5580: out = -6064;
			5581: out = 3529;
			5582: out = -1361;
			5583: out = 2696;
			5584: out = -4694;
			5585: out = -15962;
			5586: out = -579;
			5587: out = 980;
			5588: out = 839;
			5589: out = -3681;
			5590: out = 1393;
			5591: out = -4535;
			5592: out = -13773;
			5593: out = 1376;
			5594: out = 5063;
			5595: out = 5614;
			5596: out = 5002;
			5597: out = -2869;
			5598: out = -5129;
			5599: out = -2484;
			5600: out = 9523;
			5601: out = -72;
			5602: out = -6377;
			5603: out = 6697;
			5604: out = 764;
			5605: out = 3378;
			5606: out = 4296;
			5607: out = 3384;
			5608: out = 1008;
			5609: out = -2361;
			5610: out = -12506;
			5611: out = -1629;
			5612: out = 2174;
			5613: out = 3749;
			5614: out = -6573;
			5615: out = 2384;
			5616: out = 6830;
			5617: out = 5288;
			5618: out = -10714;
			5619: out = -9066;
			5620: out = 3957;
			5621: out = 5415;
			5622: out = -139;
			5623: out = -9100;
			5624: out = -7585;
			5625: out = -9743;
			5626: out = -773;
			5627: out = 6461;
			5628: out = 11698;
			5629: out = -590;
			5630: out = -6106;
			5631: out = 5250;
			5632: out = -4239;
			5633: out = 2316;
			5634: out = 6624;
			5635: out = -1302;
			5636: out = -7258;
			5637: out = -5060;
			5638: out = 8390;
			5639: out = 6291;
			5640: out = 8881;
			5641: out = 5549;
			5642: out = -11073;
			5643: out = -6666;
			5644: out = -173;
			5645: out = 399;
			5646: out = 3938;
			5647: out = -1386;
			5648: out = -4593;
			5649: out = -1062;
			5650: out = 7797;
			5651: out = 10308;
			5652: out = 3802;
			5653: out = -992;
			5654: out = -7042;
			5655: out = -5634;
			5656: out = 6264;
			5657: out = 7713;
			5658: out = 5828;
			5659: out = 962;
			5660: out = -390;
			5661: out = -3608;
			5662: out = -2011;
			5663: out = 7650;
			5664: out = 6745;
			5665: out = 2531;
			5666: out = -4450;
			5667: out = -5973;
			5668: out = -4704;
			5669: out = -2838;
			5670: out = -12771;
			5671: out = 1175;
			5672: out = 3948;
			5673: out = -551;
			5674: out = 3829;
			5675: out = 2849;
			5676: out = 1551;
			5677: out = 2133;
			5678: out = -6531;
			5679: out = -11534;
			5680: out = -11338;
			5681: out = 4526;
			5682: out = 3708;
			5683: out = 148;
			5684: out = 449;
			5685: out = 1681;
			5686: out = 2068;
			5687: out = 1194;
			5688: out = 816;
			5689: out = 3396;
			5690: out = 3690;
			5691: out = -1335;
			5692: out = -2073;
			5693: out = 1799;
			5694: out = 8518;
			5695: out = 2243;
			5696: out = 3369;
			5697: out = 408;
			5698: out = -5315;
			5699: out = -4793;
			5700: out = -2183;
			5701: out = 771;
			5702: out = 2516;
			5703: out = 3278;
			5704: out = -866;
			5705: out = -13372;
			5706: out = 2052;
			5707: out = 9254;
			5708: out = 9345;
			5709: out = -9106;
			5710: out = -5068;
			5711: out = -2389;
			5712: out = -6579;
			5713: out = -5988;
			5714: out = -3197;
			5715: out = 1310;
			5716: out = -193;
			5717: out = 2232;
			5718: out = 4612;
			5719: out = 6837;
			5720: out = 2000;
			5721: out = -7067;
			5722: out = -14682;
			5723: out = 1676;
			5724: out = 228;
			5725: out = 1706;
			5726: out = 1835;
			5727: out = 4777;
			5728: out = -1197;
			5729: out = -5809;
			5730: out = -3016;
			5731: out = 7134;
			5732: out = 9203;
			5733: out = -778;
			5734: out = 2499;
			5735: out = -4572;
			5736: out = -7623;
			5737: out = 6980;
			5738: out = 3096;
			5739: out = 1860;
			5740: out = 1237;
			5741: out = 10331;
			5742: out = 4075;
			5743: out = -3102;
			5744: out = 1497;
			5745: out = 2402;
			5746: out = 4125;
			5747: out = 3779;
			5748: out = -1750;
			5749: out = -583;
			5750: out = 1879;
			5751: out = -526;
			5752: out = -1699;
			5753: out = -1797;
			5754: out = 891;
			5755: out = 203;
			5756: out = -299;
			5757: out = -2634;
			5758: out = -6302;
			5759: out = -1033;
			5760: out = 656;
			5761: out = -2597;
			5762: out = 3699;
			5763: out = 2390;
			5764: out = 998;
			5765: out = -3711;
			5766: out = -2777;
			5767: out = -3068;
			5768: out = -231;
			5769: out = -4251;
			5770: out = 6281;
			5771: out = 9551;
			5772: out = -624;
			5773: out = -4109;
			5774: out = -3261;
			5775: out = 1371;
			5776: out = -2071;
			5777: out = -3049;
			5778: out = -1066;
			5779: out = 5407;
			5780: out = 4283;
			5781: out = 434;
			5782: out = -3056;
			5783: out = 354;
			5784: out = 4539;
			5785: out = 4597;
			5786: out = 411;
			5787: out = -5746;
			5788: out = -427;
			5789: out = 8799;
			5790: out = 162;
			5791: out = -1395;
			5792: out = -1212;
			5793: out = 4582;
			5794: out = 562;
			5795: out = -3455;
			5796: out = -7799;
			5797: out = -4171;
			5798: out = -1316;
			5799: out = 2793;
			5800: out = 4754;
			5801: out = 1826;
			5802: out = -4292;
			5803: out = -8969;
			5804: out = 5027;
			5805: out = -3470;
			5806: out = -6529;
			5807: out = -1423;
			5808: out = 3737;
			5809: out = -179;
			5810: out = -8629;
			5811: out = -6012;
			5812: out = -5691;
			5813: out = -1045;
			5814: out = 2451;
			5815: out = 8040;
			5816: out = 7284;
			5817: out = 3827;
			5818: out = -2879;
			5819: out = -847;
			5820: out = -1877;
			5821: out = -9715;
			5822: out = 6620;
			5823: out = 3586;
			5824: out = -681;
			5825: out = 6384;
			5826: out = 8798;
			5827: out = 5517;
			5828: out = -6763;
			5829: out = 185;
			5830: out = -2752;
			5831: out = -4508;
			5832: out = -9663;
			5833: out = 1688;
			5834: out = 4899;
			5835: out = -161;
			5836: out = -4061;
			5837: out = -163;
			5838: out = 6598;
			5839: out = 501;
			5840: out = 5769;
			5841: out = 504;
			5842: out = -7406;
			5843: out = -9365;
			5844: out = -2151;
			5845: out = 5311;
			5846: out = 3959;
			5847: out = 3156;
			5848: out = 686;
			5849: out = 603;
			5850: out = 7908;
			5851: out = 6258;
			5852: out = -1681;
			5853: out = -14516;
			5854: out = -9411;
			5855: out = -1954;
			5856: out = 1461;
			5857: out = 8489;
			5858: out = 3559;
			5859: out = -281;
			5860: out = 1145;
			5861: out = 3768;
			5862: out = 1246;
			5863: out = -6309;
			5864: out = -5306;
			5865: out = -4050;
			5866: out = 1939;
			5867: out = 6124;
			5868: out = 8705;
			5869: out = 4434;
			5870: out = -722;
			5871: out = -5065;
			5872: out = -681;
			5873: out = 3952;
			5874: out = 5632;
			5875: out = -1257;
			5876: out = -2718;
			5877: out = 375;
			5878: out = -2399;
			5879: out = -1095;
			5880: out = 2082;
			5881: out = 7873;
			5882: out = 1992;
			5883: out = -5015;
			5884: out = -9945;
			5885: out = 191;
			5886: out = 2337;
			5887: out = 1868;
			5888: out = -144;
			5889: out = -5592;
			5890: out = -6810;
			5891: out = -3312;
			5892: out = 5384;
			5893: out = 3972;
			5894: out = -166;
			5895: out = -4043;
			5896: out = -4735;
			5897: out = -5069;
			5898: out = -4139;
			5899: out = -2368;
			5900: out = 3838;
			5901: out = 4183;
			5902: out = -5680;
			5903: out = -254;
			5904: out = -743;
			5905: out = -1531;
			5906: out = 954;
			5907: out = 1802;
			5908: out = 2026;
			5909: out = 675;
			5910: out = 3563;
			5911: out = 2423;
			5912: out = 832;
			5913: out = -378;
			5914: out = 4191;
			5915: out = 3831;
			5916: out = -5135;
			5917: out = 677;
			5918: out = -2202;
			5919: out = -4174;
			5920: out = 5532;
			5921: out = 1335;
			5922: out = 616;
			5923: out = 4823;
			5924: out = 1701;
			5925: out = 1456;
			5926: out = 271;
			5927: out = 984;
			5928: out = -7315;
			5929: out = -8181;
			5930: out = 2491;
			5931: out = -7206;
			5932: out = -917;
			5933: out = 6390;
			5934: out = 10872;
			5935: out = 3623;
			5936: out = -1836;
			5937: out = -4197;
			5938: out = 708;
			5939: out = -3182;
			5940: out = -6793;
			5941: out = 224;
			5942: out = 4032;
			5943: out = 6159;
			5944: out = 3280;
			5945: out = 1674;
			5946: out = -425;
			5947: out = 1230;
			5948: out = 5509;
			5949: out = 2001;
			5950: out = -530;
			5951: out = 530;
			5952: out = -5588;
			5953: out = -1784;
			5954: out = 510;
			5955: out = -2368;
			5956: out = -2062;
			5957: out = 2815;
			5958: out = 9422;
			5959: out = -1211;
			5960: out = -2018;
			5961: out = -3286;
			5962: out = -5122;
			5963: out = -1309;
			5964: out = 2309;
			5965: out = 3461;
			5966: out = 8613;
			5967: out = 5501;
			5968: out = 2840;
			5969: out = -459;
			5970: out = 1092;
			5971: out = -4414;
			5972: out = -10733;
			5973: out = -3058;
			5974: out = 871;
			5975: out = 2144;
			5976: out = 251;
			5977: out = -310;
			5978: out = 311;
			5979: out = 581;
			5980: out = 4512;
			5981: out = -3374;
			5982: out = -7385;
			5983: out = -3928;
			5984: out = 1630;
			5985: out = -1652;
			5986: out = -9157;
			5987: out = -6845;
			5988: out = 2936;
			5989: out = 9109;
			5990: out = -186;
			5991: out = 4707;
			5992: out = -251;
			5993: out = -2197;
			5994: out = -7042;
			5995: out = 2106;
			5996: out = 3499;
			5997: out = -2408;
			5998: out = 7;
			5999: out = 4408;
			6000: out = 6806;
			6001: out = 4427;
			6002: out = -2634;
			6003: out = -4417;
			6004: out = 241;
			6005: out = 1619;
			6006: out = -3480;
			6007: out = -9843;
			6008: out = -4673;
			6009: out = 1068;
			6010: out = 5556;
			6011: out = 3594;
			6012: out = 8132;
			6013: out = 3955;
			6014: out = -770;
			6015: out = -987;
			6016: out = -4411;
			6017: out = -4902;
			6018: out = -3901;
			6019: out = 1427;
			6020: out = -666;
			6021: out = -2951;
			6022: out = -242;
			6023: out = 5277;
			6024: out = 5709;
			6025: out = -83;
			6026: out = 3517;
			6027: out = 1230;
			6028: out = -2345;
			6029: out = -9050;
			6030: out = -8050;
			6031: out = -3275;
			6032: out = 3551;
			6033: out = 3130;
			6034: out = 2308;
			6035: out = 277;
			6036: out = 3209;
			6037: out = -4130;
			6038: out = -5413;
			6039: out = -2348;
			6040: out = -70;
			6041: out = -2394;
			6042: out = -3303;
			6043: out = 8622;
			6044: out = -2834;
			6045: out = -1009;
			6046: out = 7111;
			6047: out = -2676;
			6048: out = -3152;
			6049: out = -480;
			6050: out = 10069;
			6051: out = -2072;
			6052: out = -3822;
			6053: out = 1471;
			6054: out = -3426;
			6055: out = -422;
			6056: out = 2737;
			6057: out = 8986;
			6058: out = 32;
			6059: out = -4871;
			6060: out = -7309;
			6061: out = 7312;
			6062: out = -857;
			6063: out = -5590;
			6064: out = 1399;
			6065: out = 4788;
			6066: out = 1963;
			6067: out = -5970;
			6068: out = 519;
			6069: out = 2267;
			6070: out = 2145;
			6071: out = -11547;
			6072: out = 4167;
			6073: out = 3619;
			6074: out = 163;
			6075: out = -4432;
			6076: out = 4540;
			6077: out = 7964;
			6078: out = 2592;
			6079: out = -3614;
			6080: out = -2990;
			6081: out = 865;
			6082: out = -5930;
			6083: out = -6261;
			6084: out = -3156;
			6085: out = 3997;
			6086: out = 5680;
			6087: out = 1881;
			6088: out = -2842;
			6089: out = 5913;
			6090: out = 5240;
			6091: out = 1868;
			6092: out = -6928;
			6093: out = -6472;
			6094: out = -4781;
			6095: out = 335;
			6096: out = 144;
			6097: out = 3872;
			6098: out = 3817;
			6099: out = 4317;
			6100: out = -5349;
			6101: out = -193;
			6102: out = 6396;
			6103: out = -4866;
			6104: out = -1649;
			6105: out = -1160;
			6106: out = -84;
			6107: out = -4748;
			6108: out = -2647;
			6109: out = 1151;
			6110: out = 5891;
			6111: out = 2193;
			6112: out = 1518;
			6113: out = 4280;
			6114: out = -44;
			6115: out = -1462;
			6116: out = -2410;
			6117: out = -2046;
			6118: out = -309;
			6119: out = 3473;
			6120: out = 7682;
			6121: out = -1613;
			6122: out = -1007;
			6123: out = -713;
			6124: out = -8241;
			6125: out = -5370;
			6126: out = -503;
			6127: out = 5667;
			6128: out = 3064;
			6129: out = 2740;
			6130: out = 698;
			6131: out = 339;
			6132: out = -358;
			6133: out = 2610;
			6134: out = 3987;
			6135: out = -1065;
			6136: out = -6981;
			6137: out = -7078;
			6138: out = 1870;
			6139: out = 5567;
			6140: out = 2953;
			6141: out = -3402;
			6142: out = 6664;
			6143: out = 6473;
			6144: out = 4215;
			6145: out = -2976;
			6146: out = 3840;
			6147: out = 3531;
			6148: out = -1896;
			6149: out = -3500;
			6150: out = -5185;
			6151: out = -4457;
			6152: out = -10098;
			6153: out = 7176;
			6154: out = 3858;
			6155: out = -7439;
			6156: out = -1082;
			6157: out = 1746;
			6158: out = 3875;
			6159: out = -407;
			6160: out = -2750;
			6161: out = -5624;
			6162: out = -5159;
			6163: out = -799;
			6164: out = 2660;
			6165: out = 4408;
			6166: out = 2706;
			6167: out = 4474;
			6168: out = 1137;
			6169: out = -1285;
			6170: out = -754;
			6171: out = 4086;
			6172: out = 2842;
			6173: out = -4781;
			6174: out = -13117;
			6175: out = -8621;
			6176: out = 2781;
			6177: out = -55;
			6178: out = -1259;
			6179: out = -4206;
			6180: out = 1176;
			6181: out = -6297;
			6182: out = 713;
			6183: out = 6540;
			6184: out = 731;
			6185: out = -2471;
			6186: out = -2590;
			6187: out = 2775;
			6188: out = 2654;
			6189: out = 5736;
			6190: out = 6288;
			6191: out = 1600;
			6192: out = -889;
			6193: out = -3552;
			6194: out = -4460;
			6195: out = 1144;
			6196: out = 5811;
			6197: out = 6547;
			6198: out = -650;
			6199: out = 290;
			6200: out = 666;
			6201: out = 259;
			6202: out = 2283;
			6203: out = -79;
			6204: out = -2678;
			6205: out = -220;
			6206: out = -1422;
			6207: out = -1536;
			6208: out = -2117;
			6209: out = 5114;
			6210: out = 1933;
			6211: out = -2184;
			6212: out = -66;
			6213: out = -2155;
			6214: out = -2200;
			6215: out = -2156;
			6216: out = 1500;
			6217: out = -82;
			6218: out = -591;
			6219: out = 4276;
			6220: out = 3079;
			6221: out = 2865;
			6222: out = 1808;
			6223: out = 1678;
			6224: out = -592;
			6225: out = -1112;
			6226: out = 1360;
			6227: out = 144;
			6228: out = -1756;
			6229: out = -3117;
			6230: out = 163;
			6231: out = 2187;
			6232: out = 2352;
			6233: out = -576;
			6234: out = -394;
			6235: out = -20;
			6236: out = -288;
			6237: out = -8415;
			6238: out = -8064;
			6239: out = -2046;
			6240: out = 8566;
			6241: out = 36;
			6242: out = -4291;
			6243: out = -3609;
			6244: out = 5428;
			6245: out = 4939;
			6246: out = 760;
			6247: out = -3037;
			6248: out = -8339;
			6249: out = -5220;
			6250: out = 1806;
			6251: out = -173;
			6252: out = 4568;
			6253: out = 6306;
			6254: out = 4965;
			6255: out = 817;
			6256: out = -3156;
			6257: out = -4755;
			6258: out = -673;
			6259: out = 1008;
			6260: out = 326;
			6261: out = -4315;
			6262: out = 6847;
			6263: out = 3659;
			6264: out = -5338;
			6265: out = -3776;
			6266: out = -7415;
			6267: out = -3854;
			6268: out = 932;
			6269: out = 8185;
			6270: out = 2043;
			6271: out = -6585;
			6272: out = -7316;
			6273: out = -2613;
			6274: out = 902;
			6275: out = -1511;
			6276: out = 234;
			6277: out = -97;
			6278: out = 469;
			6279: out = -209;
			6280: out = 1419;
			6281: out = 1788;
			6282: out = 422;
			6283: out = 2267;
			6284: out = -2120;
			6285: out = -4641;
			6286: out = 4586;
			6287: out = 6491;
			6288: out = 6318;
			6289: out = 331;
			6290: out = 1887;
			6291: out = -3692;
			6292: out = -7133;
			6293: out = -8811;
			6294: out = -2294;
			6295: out = 622;
			6296: out = 445;
			6297: out = 3050;
			6298: out = 2691;
			6299: out = 165;
			6300: out = 2841;
			6301: out = -9541;
			6302: out = -9098;
			6303: out = 1473;
			6304: out = 1784;
			6305: out = -1773;
			6306: out = -3980;
			6307: out = 7410;
			6308: out = 5642;
			6309: out = 4323;
			6310: out = -309;
			6311: out = -1947;
			6312: out = -1516;
			6313: out = 2287;
			6314: out = 2712;
			6315: out = 3532;
			6316: out = 801;
			6317: out = -270;
			6318: out = -9704;
			6319: out = 1168;
			6320: out = 9404;
			6321: out = -897;
			6322: out = 8087;
			6323: out = 5875;
			6324: out = 287;
			6325: out = -6081;
			6326: out = -4002;
			6327: out = -1128;
			6328: out = -6453;
			6329: out = 2481;
			6330: out = 3693;
			6331: out = 2291;
			6332: out = 1422;
			6333: out = 4007;
			6334: out = 4611;
			6335: out = 1152;
			6336: out = -2212;
			6337: out = -1729;
			6338: out = 2418;
			6339: out = 3991;
			6340: out = 2391;
			6341: out = 385;
			6342: out = 4197;
			6343: out = -3068;
			6344: out = -4776;
			6345: out = -4218;
			6346: out = 5820;
			6347: out = 1836;
			6348: out = -346;
			6349: out = 1235;
			6350: out = 885;
			6351: out = -4660;
			6352: out = -10936;
			6353: out = -1309;
			6354: out = -56;
			6355: out = 884;
			6356: out = -556;
			6357: out = -3515;
			6358: out = -6753;
			6359: out = -6576;
			6360: out = -662;
			6361: out = 1469;
			6362: out = 1779;
			6363: out = 1691;
			6364: out = -1901;
			6365: out = -4793;
			6366: out = -5104;
			6367: out = 7231;
			6368: out = 3982;
			6369: out = 1845;
			6370: out = 212;
			6371: out = -404;
			6372: out = -2965;
			6373: out = -2882;
			6374: out = -481;
			6375: out = 6287;
			6376: out = 7431;
			6377: out = 3891;
			6378: out = -7700;
			6379: out = -9065;
			6380: out = -5053;
			6381: out = 314;
			6382: out = -3339;
			6383: out = -1952;
			6384: out = 5006;
			6385: out = 6925;
			6386: out = 1312;
			6387: out = -5686;
			6388: out = -2267;
			6389: out = -371;
			6390: out = -1498;
			6391: out = -8736;
			6392: out = 3350;
			6393: out = 6151;
			6394: out = 5258;
			6395: out = -6947;
			6396: out = -1005;
			6397: out = 1326;
			6398: out = 1060;
			6399: out = 732;
			6400: out = 2626;
			6401: out = 3923;
			6402: out = -450;
			6403: out = 2541;
			6404: out = -669;
			6405: out = -6787;
			6406: out = -634;
			6407: out = 2490;
			6408: out = 3069;
			6409: out = -5271;
			6410: out = -270;
			6411: out = 2264;
			6412: out = 4866;
			6413: out = -7462;
			6414: out = 1395;
			6415: out = 7781;
			6416: out = -169;
			6417: out = 1264;
			6418: out = 170;
			6419: out = 1294;
			6420: out = 349;
			6421: out = 2972;
			6422: out = 3174;
			6423: out = -481;
			6424: out = 196;
			6425: out = -2159;
			6426: out = -4514;
			6427: out = 1235;
			6428: out = 5559;
			6429: out = 8171;
			6430: out = 4077;
			6431: out = 4416;
			6432: out = -3953;
			6433: out = -12021;
			6434: out = -763;
			6435: out = -151;
			6436: out = -64;
			6437: out = 559;
			6438: out = 93;
			6439: out = 2664;
			6440: out = 5029;
			6441: out = -640;
			6442: out = -2533;
			6443: out = -5588;
			6444: out = -7188;
			6445: out = -2295;
			6446: out = 3893;
			6447: out = 5787;
			6448: out = -1789;
			6449: out = -3008;
			6450: out = -2698;
			6451: out = -2884;
			6452: out = 5749;
			6453: out = 3768;
			6454: out = -1231;
			6455: out = 1223;
			6456: out = -1869;
			6457: out = -4218;
			6458: out = -6359;
			6459: out = -464;
			6460: out = 1388;
			6461: out = 566;
			6462: out = 1371;
			6463: out = -1415;
			6464: out = -863;
			6465: out = 918;
			6466: out = 4260;
			6467: out = -2130;
			6468: out = -7933;
			6469: out = 4084;
			6470: out = 727;
			6471: out = -660;
			6472: out = -2750;
			6473: out = 4314;
			6474: out = 2561;
			6475: out = -196;
			6476: out = 3823;
			6477: out = -6051;
			6478: out = -6574;
			6479: out = 5047;
			6480: out = -7809;
			6481: out = 1278;
			6482: out = 7378;
			6483: out = 266;
			6484: out = -5539;
			6485: out = -8532;
			6486: out = -5396;
			6487: out = -7343;
			6488: out = -4715;
			6489: out = -2075;
			6490: out = 489;
			6491: out = 3983;
			6492: out = 6935;
			6493: out = 7676;
			6494: out = -4747;
			6495: out = -3825;
			6496: out = 1235;
			6497: out = 3205;
			6498: out = 2089;
			6499: out = 140;
			6500: out = 1411;
			6501: out = 6721;
			6502: out = 5599;
			6503: out = 656;
			6504: out = 1211;
			6505: out = -5403;
			6506: out = -759;
			6507: out = 6074;
			6508: out = 7682;
			6509: out = 1037;
			6510: out = -2496;
			6511: out = 2592;
			6512: out = 1316;
			6513: out = -3775;
			6514: out = -9182;
			6515: out = -1833;
			6516: out = 6137;
			6517: out = 9115;
			6518: out = 2184;
			6519: out = -1369;
			6520: out = -2669;
			6521: out = 243;
			6522: out = -1572;
			6523: out = -563;
			6524: out = 803;
			6525: out = 4860;
			6526: out = 4351;
			6527: out = 2840;
			6528: out = -789;
			6529: out = -3510;
			6530: out = -2756;
			6531: out = -490;
			6532: out = -636;
			6533: out = 3102;
			6534: out = 5224;
			6535: out = 6320;
			6536: out = -3324;
			6537: out = -1911;
			6538: out = -980;
			6539: out = 1866;
			6540: out = -4009;
			6541: out = 672;
			6542: out = 5413;
			6543: out = -1334;
			6544: out = -4144;
			6545: out = -3336;
			6546: out = 1709;
			6547: out = 4191;
			6548: out = -984;
			6549: out = -8673;
			6550: out = -2240;
			6551: out = -3167;
			6552: out = 790;
			6553: out = 5872;
			6554: out = -320;
			6555: out = -748;
			6556: out = 148;
			6557: out = -7905;
			6558: out = -711;
			6559: out = 3458;
			6560: out = 2561;
			6561: out = 2702;
			6562: out = 1061;
			6563: out = -584;
			6564: out = -6756;
			6565: out = -4493;
			6566: out = -2498;
			6567: out = 1418;
			6568: out = -85;
			6569: out = 4722;
			6570: out = 4538;
			6571: out = -4195;
			6572: out = -9494;
			6573: out = -6716;
			6574: out = 1406;
			6575: out = 2870;
			6576: out = -4017;
			6577: out = -9945;
			6578: out = -876;
			6579: out = 2901;
			6580: out = 5076;
			6581: out = 1617;
			6582: out = -640;
			6583: out = -2856;
			6584: out = -935;
			6585: out = 4175;
			6586: out = 1172;
			6587: out = -472;
			6588: out = 262;
			6589: out = 909;
			6590: out = 856;
			6591: out = 1539;
			6592: out = 4773;
			6593: out = 5398;
			6594: out = 2364;
			6595: out = -3457;
			6596: out = 1799;
			6597: out = 321;
			6598: out = 673;
			6599: out = 2966;
			6600: out = 658;
			6601: out = -1870;
			6602: out = -2376;
			6603: out = 915;
			6604: out = 4102;
			6605: out = 3886;
			6606: out = -1773;
			6607: out = -2980;
			6608: out = -5201;
			6609: out = -6380;
			6610: out = -6372;
			6611: out = -3166;
			6612: out = 814;
			6613: out = 3257;
			6614: out = 4570;
			6615: out = 4605;
			6616: out = 3954;
			6617: out = -2692;
			6618: out = -845;
			6619: out = 1073;
			6620: out = 1573;
			6621: out = 771;
			6622: out = 1486;
			6623: out = 2148;
			6624: out = 1682;
			6625: out = -1040;
			6626: out = -1212;
			6627: out = 2499;
			6628: out = 860;
			6629: out = -575;
			6630: out = -3278;
			6631: out = -10118;
			6632: out = -4235;
			6633: out = 3809;
			6634: out = 8076;
			6635: out = 1716;
			6636: out = -2573;
			6637: out = -2993;
			6638: out = 461;
			6639: out = 1811;
			6640: out = -1638;
			6641: out = -10718;
			6642: out = 1090;
			6643: out = 1789;
			6644: out = -89;
			6645: out = 1017;
			6646: out = 1894;
			6647: out = 2952;
			6648: out = 3799;
			6649: out = 261;
			6650: out = 637;
			6651: out = 2331;
			6652: out = 7286;
			6653: out = -2218;
			6654: out = -9213;
			6655: out = -10569;
			6656: out = 639;
			6657: out = 2056;
			6658: out = -122;
			6659: out = 3669;
			6660: out = 644;
			6661: out = -92;
			6662: out = -700;
			6663: out = -7083;
			6664: out = -8204;
			6665: out = -5159;
			6666: out = 1170;
			6667: out = 2357;
			6668: out = 2458;
			6669: out = 389;
			6670: out = -1369;
			6671: out = -6562;
			6672: out = -7220;
			6673: out = 699;
			6674: out = 6614;
			6675: out = 6378;
			6676: out = -308;
			6677: out = -2999;
			6678: out = -4080;
			6679: out = -587;
			6680: out = 1581;
			6681: out = 6281;
			6682: out = 5534;
			6683: out = 2535;
			6684: out = -2963;
			6685: out = -1556;
			6686: out = 611;
			6687: out = -1203;
			6688: out = -9;
			6689: out = 184;
			6690: out = 139;
			6691: out = -10299;
			6692: out = -6514;
			6693: out = 772;
			6694: out = 5443;
			6695: out = 3814;
			6696: out = 927;
			6697: out = -1297;
			6698: out = -7540;
			6699: out = -3698;
			6700: out = 882;
			6701: out = 1114;
			6702: out = 5057;
			6703: out = 6544;
			6704: out = 7383;
			6705: out = 4533;
			6706: out = 3135;
			6707: out = 71;
			6708: out = -1569;
			6709: out = -6663;
			6710: out = -3997;
			6711: out = 1568;
			6712: out = 5747;
			6713: out = 1811;
			6714: out = -1854;
			6715: out = -548;
			6716: out = -1947;
			6717: out = -729;
			6718: out = 2090;
			6719: out = 8633;
			6720: out = 8319;
			6721: out = 2949;
			6722: out = -6891;
			6723: out = -4845;
			6724: out = -1395;
			6725: out = 3098;
			6726: out = -110;
			6727: out = 4504;
			6728: out = 4626;
			6729: out = 984;
			6730: out = 634;
			6731: out = 215;
			6732: out = -399;
			6733: out = -6410;
			6734: out = -685;
			6735: out = 3187;
			6736: out = 1658;
			6737: out = 4440;
			6738: out = 3261;
			6739: out = 1583;
			6740: out = -7779;
			6741: out = -1097;
			6742: out = 2026;
			6743: out = 1895;
			6744: out = -5609;
			6745: out = -2566;
			6746: out = 733;
			6747: out = -10326;
			6748: out = -3508;
			6749: out = 3406;
			6750: out = 6432;
			6751: out = 1692;
			6752: out = -6709;
			6753: out = -11665;
			6754: out = -5813;
			6755: out = -110;
			6756: out = 1458;
			6757: out = -1924;
			6758: out = -1477;
			6759: out = 1837;
			6760: out = 5158;
			6761: out = 2203;
			6762: out = 970;
			6763: out = -142;
			6764: out = 1074;
			6765: out = 1688;
			6766: out = -764;
			6767: out = -3447;
			6768: out = 824;
			6769: out = -3720;
			6770: out = -6465;
			6771: out = -7855;
			6772: out = 3774;
			6773: out = 6096;
			6774: out = 5360;
			6775: out = 2411;
			6776: out = -2009;
			6777: out = -5632;
			6778: out = -4551;
			6779: out = -216;
			6780: out = 6821;
			6781: out = 7131;
			6782: out = -1788;
			6783: out = -3884;
			6784: out = -426;
			6785: out = 6624;
			6786: out = 125;
			6787: out = 270;
			6788: out = -112;
			6789: out = 869;
			6790: out = -435;
			6791: out = -3045;
			6792: out = -6580;
			6793: out = 4562;
			6794: out = 2371;
			6795: out = 407;
			6796: out = -123;
			6797: out = 3441;
			6798: out = 1229;
			6799: out = -3733;
			6800: out = 1882;
			6801: out = 1139;
			6802: out = 966;
			6803: out = 869;
			6804: out = 1520;
			6805: out = 1383;
			6806: out = 288;
			6807: out = -2285;
			6808: out = -3114;
			6809: out = -697;
			6810: out = 4664;
			6811: out = 1052;
			6812: out = -1822;
			6813: out = -3276;
			6814: out = 433;
			6815: out = 1670;
			6816: out = 3958;
			6817: out = 8384;
			6818: out = -452;
			6819: out = -1485;
			6820: out = 1395;
			6821: out = 1699;
			6822: out = 942;
			6823: out = -2362;
			6824: out = -5277;
			6825: out = -623;
			6826: out = 1988;
			6827: out = 2247;
			6828: out = 5931;
			6829: out = -132;
			6830: out = -4747;
			6831: out = -6972;
			6832: out = 3327;
			6833: out = 2896;
			6834: out = -2395;
			6835: out = 484;
			6836: out = -2340;
			6837: out = 544;
			6838: out = 4850;
			6839: out = 1668;
			6840: out = -3646;
			6841: out = -6600;
			6842: out = 1789;
			6843: out = 97;
			6844: out = 98;
			6845: out = 1650;
			6846: out = -330;
			6847: out = 322;
			6848: out = -297;
			6849: out = -6181;
			6850: out = -2227;
			6851: out = 3307;
			6852: out = 7442;
			6853: out = 2223;
			6854: out = -780;
			6855: out = -1414;
			6856: out = 2980;
			6857: out = -1125;
			6858: out = -4906;
			6859: out = -6688;
			6860: out = -492;
			6861: out = 2097;
			6862: out = 1490;
			6863: out = -900;
			6864: out = -3180;
			6865: out = -2007;
			6866: out = 1138;
			6867: out = -1701;
			6868: out = -1451;
			6869: out = -242;
			6870: out = 1697;
			6871: out = 2708;
			6872: out = 3608;
			6873: out = 4279;
			6874: out = 1482;
			6875: out = 984;
			6876: out = -197;
			6877: out = -60;
			6878: out = -3512;
			6879: out = -745;
			6880: out = 3859;
			6881: out = 28;
			6882: out = -1860;
			6883: out = -2325;
			6884: out = -51;
			6885: out = 966;
			6886: out = -3806;
			6887: out = -11092;
			6888: out = 923;
			6889: out = 843;
			6890: out = 318;
			6891: out = -3888;
			6892: out = 2444;
			6893: out = 2186;
			6894: out = 158;
			6895: out = -4402;
			6896: out = 2204;
			6897: out = 5458;
			6898: out = -854;
			6899: out = 1157;
			6900: out = -498;
			6901: out = -1531;
			6902: out = -8896;
			6903: out = -1338;
			6904: out = 6253;
			6905: out = 8906;
			6906: out = 2543;
			6907: out = -175;
			6908: out = 738;
			6909: out = -3256;
			6910: out = -522;
			6911: out = -523;
			6912: out = 622;
			6913: out = -4533;
			6914: out = 606;
			6915: out = 5396;
			6916: out = 4647;
			6917: out = -3508;
			6918: out = -6334;
			6919: out = -931;
			6920: out = 3644;
			6921: out = 705;
			6922: out = -5235;
			6923: out = -1961;
			6924: out = -938;
			6925: out = -57;
			6926: out = -2612;
			6927: out = 3863;
			6928: out = 5627;
			6929: out = 5963;
			6930: out = 3496;
			6931: out = 1440;
			6932: out = -456;
			6933: out = -1198;
			6934: out = -1142;
			6935: out = -1241;
			6936: out = -1022;
			6937: out = -2256;
			6938: out = 3957;
			6939: out = 2526;
			6940: out = -6015;
			6941: out = 3150;
			6942: out = 4630;
			6943: out = 3416;
			6944: out = -10734;
			6945: out = -1755;
			6946: out = -1711;
			6947: out = -8179;
			6948: out = 476;
			6949: out = 525;
			6950: out = 687;
			6951: out = 6197;
			6952: out = 319;
			6953: out = -70;
			6954: out = 2344;
			6955: out = 348;
			6956: out = -3438;
			6957: out = -5141;
			6958: out = 2268;
			6959: out = 621;
			6960: out = 1574;
			6961: out = 2321;
			6962: out = 3667;
			6963: out = 1876;
			6964: out = 983;
			6965: out = 4513;
			6966: out = -2026;
			6967: out = -3799;
			6968: out = -2868;
			6969: out = -8503;
			6970: out = -4724;
			6971: out = 1853;
			6972: out = 5097;
			6973: out = 6478;
			6974: out = 1433;
			6975: out = -4216;
			6976: out = -7761;
			6977: out = -2556;
			6978: out = 1515;
			6979: out = -439;
			6980: out = -3870;
			6981: out = -3478;
			6982: out = 1181;
			6983: out = 1868;
			6984: out = 4455;
			6985: out = 4884;
			6986: out = 3388;
			6987: out = 792;
			6988: out = -1144;
			6989: out = -1366;
			6990: out = -9885;
			6991: out = -2393;
			6992: out = 3399;
			6993: out = 5029;
			6994: out = -3459;
			6995: out = -3060;
			6996: out = 2930;
			6997: out = 10964;
			6998: out = 2136;
			6999: out = -6536;
			7000: out = -8021;
			7001: out = -3393;
			7002: out = 163;
			7003: out = 168;
			7004: out = -4072;
			7005: out = 722;
			7006: out = 3880;
			7007: out = 2820;
			7008: out = 1938;
			7009: out = 1265;
			7010: out = -21;
			7011: out = -331;
			7012: out = -5993;
			7013: out = -5817;
			7014: out = 129;
			7015: out = 8718;
			7016: out = 7214;
			7017: out = 2259;
			7018: out = -956;
			7019: out = 2269;
			7020: out = 3056;
			7021: out = 1260;
			7022: out = -2772;
			7023: out = 1714;
			7024: out = 4750;
			7025: out = -969;
			7026: out = -8461;
			7027: out = -6354;
			7028: out = 6727;
			7029: out = 6435;
			7030: out = 4312;
			7031: out = -1612;
			7032: out = -3020;
			7033: out = -4102;
			7034: out = -2531;
			7035: out = -1100;
			7036: out = -4978;
			7037: out = -1663;
			7038: out = 2984;
			7039: out = 5505;
			7040: out = 498;
			7041: out = 932;
			7042: out = 5978;
			7043: out = -8358;
			7044: out = -11402;
			7045: out = -8963;
			7046: out = 2205;
			7047: out = 2741;
			7048: out = 2938;
			7049: out = 1590;
			7050: out = 5720;
			7051: out = 2684;
			7052: out = 758;
			7053: out = 5423;
			7054: out = -3112;
			7055: out = -4898;
			7056: out = -1757;
			7057: out = 331;
			7058: out = 638;
			7059: out = 377;
			7060: out = 3261;
			7061: out = 828;
			7062: out = -65;
			7063: out = -1336;
			7064: out = 370;
			7065: out = -4019;
			7066: out = -7792;
			7067: out = -7991;
			7068: out = -1671;
			7069: out = 4479;
			7070: out = 6299;
			7071: out = -247;
			7072: out = -1733;
			7073: out = -309;
			7074: out = 3268;
			7075: out = 3006;
			7076: out = 2464;
			7077: out = 1038;
			7078: out = -728;
			7079: out = -1233;
			7080: out = -609;
			7081: out = -177;
			7082: out = 3604;
			7083: out = 4140;
			7084: out = 3006;
			7085: out = 457;
			7086: out = 1483;
			7087: out = 1374;
			7088: out = -1653;
			7089: out = -3616;
			7090: out = -4204;
			7091: out = -953;
			7092: out = 4740;
			7093: out = 4626;
			7094: out = -2194;
			7095: out = -13459;
			7096: out = -4579;
			7097: out = 1330;
			7098: out = 3533;
			7099: out = 708;
			7100: out = -63;
			7101: out = 246;
			7102: out = 740;
			7103: out = 486;
			7104: out = -2199;
			7105: out = -3375;
			7106: out = 3081;
			7107: out = 4034;
			7108: out = 2433;
			7109: out = -3121;
			7110: out = 3369;
			7111: out = 1696;
			7112: out = -1436;
			7113: out = -5798;
			7114: out = -954;
			7115: out = 4216;
			7116: out = 6809;
			7117: out = -2075;
			7118: out = -4553;
			7119: out = -3177;
			7120: out = 441;
			7121: out = 2410;
			7122: out = 2136;
			7123: out = -805;
			7124: out = 513;
			7125: out = -1383;
			7126: out = -1150;
			7127: out = -345;
			7128: out = 5495;
			7129: out = 4388;
			7130: out = -1400;
			7131: out = -6108;
			7132: out = -4144;
			7133: out = 164;
			7134: out = -379;
			7135: out = -281;
			7136: out = -1835;
			7137: out = -1764;
			7138: out = 5471;
			7139: out = 5655;
			7140: out = 4697;
			7141: out = 5890;
			7142: out = 658;
			7143: out = -4381;
			7144: out = -7707;
			7145: out = -3969;
			7146: out = -963;
			7147: out = 1465;
			7148: out = 4456;
			7149: out = -1577;
			7150: out = 702;
			7151: out = 6618;
			7152: out = -6673;
			7153: out = -3294;
			7154: out = 2330;
			7155: out = 7636;
			7156: out = 3401;
			7157: out = -783;
			7158: out = -3856;
			7159: out = -2729;
			7160: out = -1912;
			7161: out = 323;
			7162: out = 4256;
			7163: out = 987;
			7164: out = -814;
			7165: out = -2009;
			7166: out = 787;
			7167: out = -1118;
			7168: out = -2706;
			7169: out = -5404;
			7170: out = 1951;
			7171: out = 716;
			7172: out = -3063;
			7173: out = -3252;
			7174: out = 1217;
			7175: out = 3481;
			7176: out = -91;
			7177: out = -1687;
			7178: out = -2148;
			7179: out = -936;
			7180: out = -5815;
			7181: out = -1323;
			7182: out = 2621;
			7183: out = 3961;
			7184: out = 1086;
			7185: out = -2828;
			7186: out = -4757;
			7187: out = -5049;
			7188: out = 2146;
			7189: out = 4722;
			7190: out = 239;
			7191: out = 1314;
			7192: out = 1078;
			7193: out = 802;
			7194: out = -7451;
			7195: out = -1758;
			7196: out = 2918;
			7197: out = 3929;
			7198: out = 1074;
			7199: out = -3221;
			7200: out = -4536;
			7201: out = 3213;
			7202: out = 1182;
			7203: out = -133;
			7204: out = 141;
			7205: out = -2258;
			7206: out = 27;
			7207: out = 3673;
			7208: out = 7114;
			7209: out = 3346;
			7210: out = 742;
			7211: out = 1880;
			7212: out = 1617;
			7213: out = 1658;
			7214: out = -330;
			7215: out = 1032;
			7216: out = -3099;
			7217: out = -754;
			7218: out = 4448;
			7219: out = 5770;
			7220: out = 1676;
			7221: out = -2959;
			7222: out = -2433;
			7223: out = -2234;
			7224: out = -2584;
			7225: out = -3992;
			7226: out = 1393;
			7227: out = 4402;
			7228: out = 5320;
			7229: out = 1592;
			7230: out = 1576;
			7231: out = -322;
			7232: out = -2667;
			7233: out = 4114;
			7234: out = 3351;
			7235: out = 1893;
			7236: out = 54;
			7237: out = 1775;
			7238: out = -724;
			7239: out = -4815;
			7240: out = -4713;
			7241: out = 38;
			7242: out = 2801;
			7243: out = -3335;
			7244: out = -40;
			7245: out = 392;
			7246: out = -573;
			7247: out = -814;
			7248: out = -2912;
			7249: out = -2675;
			7250: out = -211;
			7251: out = 2370;
			7252: out = 831;
			7253: out = -2454;
			7254: out = -5823;
			7255: out = -2106;
			7256: out = 1677;
			7257: out = 2657;
			7258: out = -2227;
			7259: out = -2406;
			7260: out = 348;
			7261: out = 524;
			7262: out = -3371;
			7263: out = -5049;
			7264: out = 671;
			7265: out = -1564;
			7266: out = -864;
			7267: out = 1018;
			7268: out = -668;
			7269: out = 2998;
			7270: out = 4450;
			7271: out = 6269;
			7272: out = -5167;
			7273: out = -2320;
			7274: out = 4540;
			7275: out = -134;
			7276: out = -7443;
			7277: out = -8590;
			7278: out = 5226;
			7279: out = 1018;
			7280: out = 2014;
			7281: out = 885;
			7282: out = 72;
			7283: out = -306;
			7284: out = -1910;
			7285: out = -7717;
			7286: out = 1496;
			7287: out = 5604;
			7288: out = 7572;
			7289: out = 3002;
			7290: out = 1908;
			7291: out = -2201;
			7292: out = -5449;
			7293: out = -1819;
			7294: out = 4147;
			7295: out = 6441;
			7296: out = 2073;
			7297: out = -942;
			7298: out = -2105;
			7299: out = -2115;
			7300: out = -852;
			7301: out = -3390;
			7302: out = -4655;
			7303: out = -2819;
			7304: out = 4723;
			7305: out = 6038;
			7306: out = 901;
			7307: out = -6167;
			7308: out = -5105;
			7309: out = 1494;
			7310: out = 5225;
			7311: out = 2943;
			7312: out = -3708;
			7313: out = -10106;
			7314: out = -216;
			7315: out = 1229;
			7316: out = 712;
			7317: out = 500;
			7318: out = 1628;
			7319: out = -749;
			7320: out = -5295;
			7321: out = -5564;
			7322: out = -905;
			7323: out = 3917;
			7324: out = 945;
			7325: out = 2715;
			7326: out = 1089;
			7327: out = -33;
			7328: out = -45;
			7329: out = 410;
			7330: out = -1126;
			7331: out = -5473;
			7332: out = -1437;
			7333: out = 3360;
			7334: out = 6395;
			7335: out = 212;
			7336: out = -795;
			7337: out = -156;
			7338: out = 3125;
			7339: out = -878;
			7340: out = -1867;
			7341: out = -1470;
			7342: out = 975;
			7343: out = -2550;
			7344: out = -4674;
			7345: out = -925;
			7346: out = 573;
			7347: out = 3557;
			7348: out = 4416;
			7349: out = 905;
			7350: out = -213;
			7351: out = 673;
			7352: out = 2882;
			7353: out = 3498;
			7354: out = 309;
			7355: out = -4592;
			7356: out = 2078;
			7357: out = -691;
			7358: out = -161;
			7359: out = 151;
			7360: out = 8175;
			7361: out = 2792;
			7362: out = -4976;
			7363: out = -112;
			7364: out = -329;
			7365: out = -744;
			7366: out = -700;
			7367: out = -2431;
			7368: out = 3084;
			7369: out = 6631;
			7370: out = -1508;
			7371: out = -7684;
			7372: out = -7972;
			7373: out = 1075;
			7374: out = 6207;
			7375: out = 4541;
			7376: out = -1636;
			7377: out = 1216;
			7378: out = 0;
			7379: out = -87;
			7380: out = -4786;
			7381: out = 4318;
			7382: out = 1708;
			7383: out = -1780;
			7384: out = -4248;
			7385: out = 1647;
			7386: out = 3432;
			7387: out = -793;
			7388: out = 755;
			7389: out = 178;
			7390: out = 918;
			7391: out = 235;
			7392: out = 361;
			7393: out = -1959;
			7394: out = -4018;
			7395: out = -3678;
			7396: out = -1064;
			7397: out = 687;
			7398: out = 575;
			7399: out = -1205;
			7400: out = -702;
			7401: out = 1702;
			7402: out = 749;
			7403: out = 368;
			7404: out = -141;
			7405: out = -1017;
			7406: out = -1293;
			7407: out = -2185;
			7408: out = -1783;
			7409: out = 606;
			7410: out = 5654;
			7411: out = 7665;
			7412: out = 4879;
			7413: out = -1307;
			7414: out = -2794;
			7415: out = 1226;
			7416: out = -2164;
			7417: out = -671;
			7418: out = 51;
			7419: out = 685;
			7420: out = 4225;
			7421: out = 5464;
			7422: out = 2707;
			7423: out = 1894;
			7424: out = -3287;
			7425: out = -6844;
			7426: out = -8315;
			7427: out = -4640;
			7428: out = -1100;
			7429: out = 1812;
			7430: out = -302;
			7431: out = 2251;
			7432: out = 3468;
			7433: out = 3966;
			7434: out = -2587;
			7435: out = -3697;
			7436: out = -777;
			7437: out = 5443;
			7438: out = -416;
			7439: out = -5509;
			7440: out = 41;
			7441: out = -4380;
			7442: out = -917;
			7443: out = 3133;
			7444: out = 1970;
			7445: out = 1573;
			7446: out = 1929;
			7447: out = 4619;
			7448: out = -1989;
			7449: out = -4163;
			7450: out = -4104;
			7451: out = -4828;
			7452: out = -3539;
			7453: out = 12;
			7454: out = 5408;
			7455: out = 1484;
			7456: out = -1533;
			7457: out = -2692;
			7458: out = 1956;
			7459: out = 2466;
			7460: out = -581;
			7461: out = -8613;
			7462: out = -2459;
			7463: out = 55;
			7464: out = 2216;
			7465: out = 2513;
			7466: out = 3190;
			7467: out = 2336;
			7468: out = 2889;
			7469: out = -6221;
			7470: out = -4244;
			7471: out = 1045;
			7472: out = 1915;
			7473: out = 320;
			7474: out = -1236;
			7475: out = -464;
			7476: out = 4458;
			7477: out = 3647;
			7478: out = 850;
			7479: out = 2266;
			7480: out = 2404;
			7481: out = 374;
			7482: out = -6437;
			7483: out = -1027;
			7484: out = -1210;
			7485: out = -1306;
			7486: out = -6839;
			7487: out = 1911;
			7488: out = 4576;
			7489: out = 1460;
			7490: out = -370;
			7491: out = -654;
			7492: out = 242;
			7493: out = -288;
			7494: out = -2264;
			7495: out = -2778;
			7496: out = -393;
			7497: out = -2583;
			7498: out = 1492;
			7499: out = 6272;
			7500: out = 7927;
			7501: out = 7205;
			7502: out = 3196;
			7503: out = -1151;
			7504: out = -5378;
			7505: out = -4700;
			7506: out = -1906;
			7507: out = 3583;
			7508: out = -3156;
			7509: out = -3401;
			7510: out = 1829;
			7511: out = 4953;
			7512: out = 2831;
			7513: out = -1692;
			7514: out = -2016;
			7515: out = -4215;
			7516: out = -3494;
			7517: out = -3108;
			7518: out = -205;
			7519: out = 163;
			7520: out = -180;
			7521: out = -5180;
			7522: out = 2643;
			7523: out = 4084;
			7524: out = 2353;
			7525: out = -9311;
			7526: out = -3774;
			7527: out = 2220;
			7528: out = 208;
			7529: out = 114;
			7530: out = -1854;
			7531: out = -1466;
			7532: out = 3235;
			7533: out = 2859;
			7534: out = 2238;
			7535: out = 3526;
			7536: out = 1240;
			7537: out = -749;
			7538: out = -2492;
			7539: out = -899;
			7540: out = 59;
			7541: out = -517;
			7542: out = -4899;
			7543: out = 5773;
			7544: out = 5147;
			7545: out = -88;
			7546: out = 7253;
			7547: out = -3561;
			7548: out = -8936;
			7549: out = -6537;
			7550: out = -1435;
			7551: out = 823;
			7552: out = 1438;
			7553: out = 5079;
			7554: out = 5425;
			7555: out = 2973;
			7556: out = -2118;
			7557: out = -1727;
			7558: out = -868;
			7559: out = 271;
			7560: out = 1472;
			7561: out = -409;
			7562: out = -338;
			7563: out = 1382;
			7564: out = 941;
			7565: out = -763;
			7566: out = -1450;
			7567: out = -599;
			7568: out = 3486;
			7569: out = 3133;
			7570: out = -608;
			7571: out = -5794;
			7572: out = -3002;
			7573: out = 846;
			7574: out = -4234;
			7575: out = -4407;
			7576: out = -2753;
			7577: out = 2275;
			7578: out = 602;
			7579: out = 1095;
			7580: out = 600;
			7581: out = 256;
			7582: out = -1599;
			7583: out = -1651;
			7584: out = 1013;
			7585: out = -6216;
			7586: out = 523;
			7587: out = 6921;
			7588: out = 4631;
			7589: out = 1009;
			7590: out = -894;
			7591: out = 2065;
			7592: out = -1256;
			7593: out = 153;
			7594: out = 638;
			7595: out = 2374;
			7596: out = 1611;
			7597: out = 2766;
			7598: out = 2508;
			7599: out = -1690;
			7600: out = -4355;
			7601: out = -4369;
			7602: out = -4140;
			7603: out = 1130;
			7604: out = 1691;
			7605: out = 290;
			7606: out = -2383;
			7607: out = 762;
			7608: out = 3179;
			7609: out = 3322;
			7610: out = -836;
			7611: out = -386;
			7612: out = 2238;
			7613: out = 1459;
			7614: out = -1995;
			7615: out = -3387;
			7616: out = 838;
			7617: out = 3766;
			7618: out = 1974;
			7619: out = -3269;
			7620: out = 409;
			7621: out = -479;
			7622: out = 730;
			7623: out = 1788;
			7624: out = 279;
			7625: out = -980;
			7626: out = -703;
			7627: out = 516;
			7628: out = -182;
			7629: out = -1479;
			7630: out = -1353;
			7631: out = -276;
			7632: out = 2594;
			7633: out = 4163;
			7634: out = 573;
			7635: out = -280;
			7636: out = -2568;
			7637: out = -6291;
			7638: out = -1845;
			7639: out = 781;
			7640: out = 2081;
			7641: out = -175;
			7642: out = 3474;
			7643: out = 3651;
			7644: out = -2578;
			7645: out = 2727;
			7646: out = -1013;
			7647: out = -4959;
			7648: out = -2264;
			7649: out = 1660;
			7650: out = 4615;
			7651: out = 2957;
			7652: out = 342;
			7653: out = -4251;
			7654: out = -5523;
			7655: out = -1140;
			7656: out = 2609;
			7657: out = 3593;
			7658: out = 1387;
			7659: out = -2879;
			7660: out = -3996;
			7661: out = -2793;
			7662: out = -4871;
			7663: out = -744;
			7664: out = 1256;
			7665: out = 1560;
			7666: out = 1989;
			7667: out = 1944;
			7668: out = 917;
			7669: out = 378;
			7670: out = -3423;
			7671: out = -3126;
			7672: out = 1423;
			7673: out = -1565;
			7674: out = -252;
			7675: out = 2116;
			7676: out = 7246;
			7677: out = 3566;
			7678: out = -629;
			7679: out = -4921;
			7680: out = -1721;
			7681: out = -862;
			7682: out = 894;
			7683: out = 1572;
			7684: out = 3134;
			7685: out = -956;
			7686: out = -6865;
			7687: out = 1122;
			7688: out = 3896;
			7689: out = 3634;
			7690: out = 1485;
			7691: out = -3405;
			7692: out = -3052;
			7693: out = 1251;
			7694: out = -271;
			7695: out = -1706;
			7696: out = -2750;
			7697: out = 944;
			7698: out = -80;
			7699: out = 1551;
			7700: out = 4019;
			7701: out = 561;
			7702: out = 1595;
			7703: out = 1455;
			7704: out = 546;
			7705: out = -5517;
			7706: out = -4905;
			7707: out = 818;
			7708: out = 9;
			7709: out = 1323;
			7710: out = 1473;
			7711: out = 2003;
			7712: out = 4797;
			7713: out = 2764;
			7714: out = -4005;
			7715: out = -3775;
			7716: out = -5986;
			7717: out = -3961;
			7718: out = -2647;
			7719: out = 6076;
			7720: out = 4957;
			7721: out = 477;
			7722: out = -3103;
			7723: out = 1671;
			7724: out = 2776;
			7725: out = -7265;
			7726: out = -4981;
			7727: out = -4740;
			7728: out = -1762;
			7729: out = 223;
			7730: out = 3858;
			7731: out = 3676;
			7732: out = 628;
			7733: out = -1148;
			7734: out = -379;
			7735: out = 1818;
			7736: out = -226;
			7737: out = 496;
			7738: out = -1195;
			7739: out = -3588;
			7740: out = -2845;
			7741: out = 785;
			7742: out = 3380;
			7743: out = 219;
			7744: out = -618;
			7745: out = 720;
			7746: out = 4853;
			7747: out = 926;
			7748: out = 360;
			7749: out = -54;
			7750: out = -4749;
			7751: out = -1399;
			7752: out = -791;
			7753: out = -3827;
			7754: out = 1461;
			7755: out = 3866;
			7756: out = 5138;
			7757: out = 4363;
			7758: out = -1537;
			7759: out = -5905;
			7760: out = -3675;
			7761: out = -7546;
			7762: out = -789;
			7763: out = 5258;
			7764: out = 6093;
			7765: out = 1860;
			7766: out = -52;
			7767: out = 1685;
			7768: out = -142;
			7769: out = -656;
			7770: out = -22;
			7771: out = 4532;
			7772: out = 1672;
			7773: out = -1765;
			7774: out = -4536;
			7775: out = -495;
			7776: out = 1074;
			7777: out = 773;
			7778: out = -1512;
			7779: out = -104;
			7780: out = 1861;
			7781: out = 2252;
			7782: out = 1849;
			7783: out = -1582;
			7784: out = -3108;
			7785: out = -3352;
			7786: out = 2888;
			7787: out = 142;
			7788: out = -7306;
			7789: out = 1183;
			7790: out = 3955;
			7791: out = 4980;
			7792: out = -183;
			7793: out = 1060;
			7794: out = -1015;
			7795: out = -3338;
			7796: out = -2173;
			7797: out = -2933;
			7798: out = -1586;
			7799: out = 3036;
			7800: out = 5349;
			7801: out = 4990;
			7802: out = 1404;
			7803: out = -251;
			7804: out = -5078;
			7805: out = -6484;
			7806: out = -2367;
			7807: out = 651;
			7808: out = 4062;
			7809: out = 4512;
			7810: out = 4947;
			7811: out = -3049;
			7812: out = -6659;
			7813: out = -570;
			7814: out = -834;
			7815: out = 1810;
			7816: out = 2277;
			7817: out = 1689;
			7818: out = -2039;
			7819: out = -4343;
			7820: out = -4091;
			7821: out = -157;
			7822: out = 1844;
			7823: out = 1988;
			7824: out = 2136;
			7825: out = 2057;
			7826: out = 429;
			7827: out = -5040;
			7828: out = 525;
			7829: out = -112;
			7830: out = -484;
			7831: out = -559;
			7832: out = 3644;
			7833: out = 1529;
			7834: out = -6381;
			7835: out = -712;
			7836: out = 2384;
			7837: out = 3569;
			7838: out = 1523;
			7839: out = -3674;
			7840: out = -6126;
			7841: out = -3596;
			7842: out = 2;
			7843: out = 1655;
			7844: out = 1642;
			7845: out = 2736;
			7846: out = 1706;
			7847: out = -2214;
			7848: out = -8338;
			7849: out = -420;
			7850: out = 4813;
			7851: out = 7172;
			7852: out = 216;
			7853: out = 1059;
			7854: out = 73;
			7855: out = 664;
			7856: out = -5723;
			7857: out = -2806;
			7858: out = 748;
			7859: out = 1513;
			7860: out = 1710;
			7861: out = 3368;
			7862: out = 4615;
			7863: out = 3723;
			7864: out = -1271;
			7865: out = -5331;
			7866: out = -5791;
			7867: out = 833;
			7868: out = 4433;
			7869: out = 3553;
			7870: out = -3675;
			7871: out = -2172;
			7872: out = 1299;
			7873: out = 112;
			7874: out = 403;
			7875: out = 573;
			7876: out = 2194;
			7877: out = 422;
			7878: out = -628;
			7879: out = -1629;
			7880: out = 98;
			7881: out = 47;
			7882: out = 1271;
			7883: out = 1927;
			7884: out = 1925;
			7885: out = 1162;
			7886: out = -41;
			7887: out = -1671;
			7888: out = -602;
			7889: out = -354;
			7890: out = -1086;
			7891: out = 214;
			7892: out = -774;
			7893: out = -563;
			7894: out = -376;
			7895: out = 5502;
			7896: out = 3070;
			7897: out = -3208;
			7898: out = 1625;
			7899: out = 355;
			7900: out = -699;
			7901: out = -5969;
			7902: out = 658;
			7903: out = -625;
			7904: out = -2250;
			7905: out = 6011;
			7906: out = 6091;
			7907: out = 2625;
			7908: out = -3541;
			7909: out = -6383;
			7910: out = -4937;
			7911: out = -552;
			7912: out = -86;
			7913: out = 2559;
			7914: out = 2541;
			7915: out = 302;
			7916: out = 1432;
			7917: out = -1118;
			7918: out = -3838;
			7919: out = 604;
			7920: out = -189;
			7921: out = -348;
			7922: out = -907;
			7923: out = 3141;
			7924: out = 2515;
			7925: out = -726;
			7926: out = -4770;
			7927: out = -4765;
			7928: out = -1206;
			7929: out = 3521;
			7930: out = 4131;
			7931: out = 2727;
			7932: out = -1190;
			7933: out = -7984;
			7934: out = -6235;
			7935: out = -1630;
			7936: out = 2160;
			7937: out = 1231;
			7938: out = -812;
			7939: out = -1783;
			7940: out = 936;
			7941: out = 4013;
			7942: out = 5499;
			7943: out = 2640;
			7944: out = -1404;
			7945: out = -7000;
			7946: out = -7928;
			7947: out = -1430;
			7948: out = 3059;
			7949: out = 4679;
			7950: out = 3366;
			7951: out = 641;
			7952: out = -1255;
			7953: out = -2115;
			7954: out = 569;
			7955: out = -4077;
			7956: out = -2501;
			7957: out = 3704;
			7958: out = 6076;
			7959: out = 1059;
			7960: out = -5394;
			7961: out = 1616;
			7962: out = -7831;
			7963: out = -5557;
			7964: out = 2057;
			7965: out = 8278;
			7966: out = 4475;
			7967: out = -1106;
			7968: out = -1663;
			7969: out = -273;
			7970: out = 1025;
			7971: out = -588;
			7972: out = 1242;
			7973: out = -1246;
			7974: out = -1851;
			7975: out = -755;
			7976: out = 2505;
			7977: out = 2478;
			7978: out = 304;
			7979: out = 986;
			7980: out = -408;
			7981: out = -281;
			7982: out = 2117;
			7983: out = 316;
			7984: out = -165;
			7985: out = -219;
			7986: out = 45;
			7987: out = -851;
			7988: out = -2660;
			7989: out = -5850;
			7990: out = 1567;
			7991: out = 3130;
			7992: out = 836;
			7993: out = 3061;
			7994: out = 363;
			7995: out = 703;
			7996: out = 2933;
			7997: out = 999;
			7998: out = -4644;
			7999: out = -9718;
			8000: out = 997;
			8001: out = 552;
			8002: out = 1591;
			8003: out = 2355;
			8004: out = 2549;
			8005: out = -1127;
			8006: out = -5069;
			8007: out = -7279;
			8008: out = -482;
			8009: out = 4667;
			8010: out = 2393;
			8011: out = 5140;
			8012: out = -429;
			8013: out = -5386;
			8014: out = -1811;
			8015: out = -1822;
			8016: out = -292;
			8017: out = 1482;
			8018: out = -1393;
			8019: out = -2711;
			8020: out = -1272;
			8021: out = 6009;
			8022: out = 2205;
			8023: out = -2877;
			8024: out = -7122;
			8025: out = -1473;
			8026: out = 269;
			8027: out = 1393;
			8028: out = 8398;
			8029: out = 917;
			8030: out = -4009;
			8031: out = -5053;
			8032: out = 1661;
			8033: out = 3282;
			8034: out = 2180;
			8035: out = 1708;
			8036: out = 226;
			8037: out = 13;
			8038: out = 210;
			8039: out = 714;
			8040: out = 1135;
			8041: out = 1346;
			8042: out = 412;
			8043: out = 360;
			8044: out = -592;
			8045: out = -1085;
			8046: out = 4219;
			8047: out = 4100;
			8048: out = 2525;
			8049: out = 3239;
			8050: out = -724;
			8051: out = -2608;
			8052: out = -3800;
			8053: out = 756;
			8054: out = -2794;
			8055: out = -3814;
			8056: out = 4233;
			8057: out = 693;
			8058: out = -959;
			8059: out = -2262;
			8060: out = -900;
			8061: out = 693;
			8062: out = 3066;
			8063: out = 5619;
			8064: out = 530;
			8065: out = -776;
			8066: out = 1011;
			8067: out = -9949;
			8068: out = -4207;
			8069: out = 2501;
			8070: out = 5534;
			8071: out = 3834;
			8072: out = 843;
			8073: out = -1732;
			8074: out = 3231;
			8075: out = -1660;
			8076: out = -5055;
			8077: out = -3848;
			8078: out = 2005;
			8079: out = 3126;
			8080: out = 59;
			8081: out = 4176;
			8082: out = 238;
			8083: out = -695;
			8084: out = 225;
			8085: out = 124;
			8086: out = -2055;
			8087: out = -3240;
			8088: out = 139;
			8089: out = 2740;
			8090: out = 2557;
			8091: out = -1322;
			8092: out = -1373;
			8093: out = -783;
			8094: out = 1366;
			8095: out = 3800;
			8096: out = -450;
			8097: out = -6045;
			8098: out = -7201;
			8099: out = -1697;
			8100: out = 3381;
			8101: out = 2764;
			8102: out = 4819;
			8103: out = -6966;
			8104: out = -8989;
			8105: out = 520;
			8106: out = 4799;
			8107: out = 3551;
			8108: out = -742;
			8109: out = 240;
			8110: out = -580;
			8111: out = -1959;
			8112: out = -4819;
			8113: out = -3236;
			8114: out = 1563;
			8115: out = 5906;
			8116: out = 4461;
			8117: out = -99;
			8118: out = -4490;
			8119: out = -5072;
			8120: out = -1478;
			8121: out = -228;
			8122: out = -320;
			8123: out = 2241;
			8124: out = 3273;
			8125: out = 2842;
			8126: out = -341;
			8127: out = 955;
			8128: out = 556;
			8129: out = 853;
			8130: out = 596;
			8131: out = -1080;
			8132: out = -2565;
			8133: out = -1672;
			8134: out = -3039;
			8135: out = -237;
			8136: out = 1631;
			8137: out = 777;
			8138: out = 650;
			8139: out = 269;
			8140: out = -905;
			8141: out = 2403;
			8142: out = -3790;
			8143: out = -7173;
			8144: out = 7587;
			8145: out = -457;
			8146: out = -2230;
			8147: out = -2725;
			8148: out = 1264;
			8149: out = -2526;
			8150: out = -3196;
			8151: out = 4067;
			8152: out = 4450;
			8153: out = 2415;
			8154: out = -1303;
			8155: out = -5851;
			8156: out = -2526;
			8157: out = 1588;
			8158: out = 421;
			8159: out = 904;
			8160: out = 3203;
			8161: out = 7557;
			8162: out = 375;
			8163: out = 2152;
			8164: out = 2109;
			8165: out = -2566;
			8166: out = -537;
			8167: out = 53;
			8168: out = 944;
			8169: out = 174;
			8170: out = 3662;
			8171: out = 4031;
			8172: out = -391;
			8173: out = -2021;
			8174: out = -359;
			8175: out = 3251;
			8176: out = 306;
			8177: out = -634;
			8178: out = -2394;
			8179: out = -2829;
			8180: out = -779;
			8181: out = 145;
			8182: out = 244;
			8183: out = 7033;
			8184: out = 3656;
			8185: out = -108;
			8186: out = -3131;
			8187: out = -1602;
			8188: out = 299;
			8189: out = 1743;
			8190: out = 64;
			8191: out = 133;
			8192: out = -1129;
			8193: out = -3040;
			8194: out = -967;
			8195: out = 306;
			8196: out = 794;
			8197: out = 4640;
			8198: out = -460;
			8199: out = -5111;
			8200: out = -8157;
			8201: out = -1897;
			8202: out = -1472;
			8203: out = -2139;
			8204: out = 4819;
			8205: out = 4913;
			8206: out = 3882;
			8207: out = -503;
			8208: out = -789;
			8209: out = -4447;
			8210: out = -6430;
			8211: out = -4225;
			8212: out = -909;
			8213: out = 2879;
			8214: out = 5605;
			8215: out = 1158;
			8216: out = -898;
			8217: out = -812;
			8218: out = 3699;
			8219: out = 455;
			8220: out = -2527;
			8221: out = -4811;
			8222: out = 2996;
			8223: out = 569;
			8224: out = -3259;
			8225: out = 1113;
			8226: out = 592;
			8227: out = 1476;
			8228: out = -640;
			8229: out = 3698;
			8230: out = -2592;
			8231: out = -5744;
			8232: out = 899;
			8233: out = 2804;
			8234: out = -774;
			8235: out = -9373;
			8236: out = 1750;
			8237: out = 1564;
			8238: out = 1859;
			8239: out = 2912;
			8240: out = 2097;
			8241: out = -810;
			8242: out = -3520;
			8243: out = -1018;
			8244: out = 23;
			8245: out = -827;
			8246: out = -4860;
			8247: out = -718;
			8248: out = 1916;
			8249: out = 2816;
			8250: out = 6174;
			8251: out = 3490;
			8252: out = -1687;
			8253: out = -10621;
			8254: out = -1804;
			8255: out = 3702;
			8256: out = 5267;
			8257: out = -1305;
			8258: out = 1000;
			8259: out = 2058;
			8260: out = -1083;
			8261: out = -1967;
			8262: out = 1214;
			8263: out = 6692;
			8264: out = 641;
			8265: out = 1297;
			8266: out = -972;
			8267: out = -1672;
			8268: out = -2978;
			8269: out = 1201;
			8270: out = 3619;
			8271: out = 935;
			8272: out = -4457;
			8273: out = -4855;
			8274: out = 1267;
			8275: out = 4836;
			8276: out = 2714;
			8277: out = -2711;
			8278: out = -3108;
			8279: out = 980;
			8280: out = 4795;
			8281: out = 1169;
			8282: out = 2832;
			8283: out = -2115;
			8284: out = -4531;
			8285: out = -1230;
			8286: out = 1666;
			8287: out = 1733;
			8288: out = 191;
			8289: out = -6270;
			8290: out = -4171;
			8291: out = 1596;
			8292: out = 3069;
			8293: out = 996;
			8294: out = -749;
			8295: out = 3136;
			8296: out = -3496;
			8297: out = -1443;
			8298: out = 417;
			8299: out = 4103;
			8300: out = -3890;
			8301: out = -3139;
			8302: out = 7145;
			8303: out = 653;
			8304: out = -270;
			8305: out = -1534;
			8306: out = 2234;
			8307: out = -1281;
			8308: out = -2611;
			8309: out = -3633;
			8310: out = -683;
			8311: out = -2920;
			8312: out = -4397;
			8313: out = -1188;
			8314: out = 2384;
			8315: out = 2803;
			8316: out = -1221;
			8317: out = 4340;
			8318: out = 779;
			8319: out = -3007;
			8320: out = -4538;
			8321: out = -1230;
			8322: out = 764;
			8323: out = -240;
			8324: out = 2787;
			8325: out = 276;
			8326: out = -1059;
			8327: out = 1527;
			8328: out = 516;
			8329: out = -2510;
			8330: out = -6905;
			8331: out = 1739;
			8332: out = 1098;
			8333: out = -454;
			8334: out = -1773;
			8335: out = 2275;
			8336: out = 5798;
			8337: out = 7477;
			8338: out = -328;
			8339: out = -1602;
			8340: out = -2369;
			8341: out = -1630;
			8342: out = -4216;
			8343: out = -213;
			8344: out = 5419;
			8345: out = 790;
			8346: out = -2776;
			8347: out = -3253;
			8348: out = 5427;
			8349: out = 3808;
			8350: out = 2301;
			8351: out = -2571;
			8352: out = 1381;
			8353: out = -4441;
			8354: out = -4440;
			8355: out = 2220;
			8356: out = 4656;
			8357: out = 3200;
			8358: out = 181;
			8359: out = 600;
			8360: out = 1985;
			8361: out = 2903;
			8362: out = 2682;
			8363: out = -2051;
			8364: out = -1891;
			8365: out = 443;
			8366: out = -2353;
			8367: out = -1867;
			8368: out = -971;
			8369: out = -64;
			8370: out = 2128;
			8371: out = 1067;
			8372: out = -370;
			8373: out = -584;
			8374: out = 3489;
			8375: out = 2826;
			8376: out = -4336;
			8377: out = -4670;
			8378: out = -1580;
			8379: out = 3527;
			8380: out = -2263;
			8381: out = 2240;
			8382: out = 3592;
			8383: out = 3730;
			8384: out = 152;
			8385: out = -1778;
			8386: out = -2587;
			8387: out = 3174;
			8388: out = -1037;
			8389: out = -1765;
			8390: out = 469;
			8391: out = 2077;
			8392: out = 496;
			8393: out = -331;
			8394: out = 5876;
			8395: out = 1866;
			8396: out = -1768;
			8397: out = -3659;
			8398: out = -3382;
			8399: out = -2030;
			8400: out = -1223;
			8401: out = 3360;
			8402: out = -5307;
			8403: out = -6087;
			8404: out = 1259;
			8405: out = 3071;
			8406: out = 3366;
			8407: out = -432;
			8408: out = -7719;
			8409: out = -3504;
			8410: out = -128;
			8411: out = -123;
			8412: out = 278;
			8413: out = -86;
			8414: out = -151;
			8415: out = -5;
			8416: out = -821;
			8417: out = 1073;
			8418: out = 4153;
			8419: out = 830;
			8420: out = -824;
			8421: out = -3227;
			8422: out = -6970;
			8423: out = -1568;
			8424: out = 1038;
			8425: out = 619;
			8426: out = 1511;
			8427: out = 654;
			8428: out = 101;
			8429: out = 952;
			8430: out = -63;
			8431: out = -153;
			8432: out = -580;
			8433: out = 6372;
			8434: out = -1316;
			8435: out = -6551;
			8436: out = -1127;
			8437: out = -811;
			8438: out = 2387;
			8439: out = 4534;
			8440: out = 1163;
			8441: out = 2461;
			8442: out = 1759;
			8443: out = -2329;
			8444: out = -563;
			8445: out = -1170;
			8446: out = -3723;
			8447: out = 2616;
			8448: out = -2988;
			8449: out = -2559;
			8450: out = 3715;
			8451: out = 7616;
			8452: out = 2971;
			8453: out = -4319;
			8454: out = -10092;
			8455: out = -777;
			8456: out = 4996;
			8457: out = -341;
			8458: out = -3940;
			8459: out = -3504;
			8460: out = 1916;
			8461: out = 1370;
			8462: out = 1023;
			8463: out = 263;
			8464: out = 3461;
			8465: out = 249;
			8466: out = -1109;
			8467: out = -2534;
			8468: out = 2186;
			8469: out = 329;
			8470: out = -156;
			8471: out = -143;
			8472: out = 678;
			8473: out = 276;
			8474: out = 210;
			8475: out = 3004;
			8476: out = 2787;
			8477: out = 1938;
			8478: out = -1457;
			8479: out = 3150;
			8480: out = -2021;
			8481: out = -5549;
			8482: out = 3693;
			8483: out = 3980;
			8484: out = 3069;
			8485: out = -730;
			8486: out = 1300;
			8487: out = -845;
			8488: out = -2373;
			8489: out = -802;
			8490: out = -1523;
			8491: out = -1489;
			8492: out = -1389;
			8493: out = 3078;
			8494: out = 1553;
			8495: out = -516;
			8496: out = -209;
			8497: out = -169;
			8498: out = -198;
			8499: out = -428;
			8500: out = -3449;
			8501: out = -959;
			8502: out = 1450;
			8503: out = -330;
			8504: out = 25;
			8505: out = -1227;
			8506: out = -2822;
			8507: out = 450;
			8508: out = -832;
			8509: out = -331;
			8510: out = 3972;
			8511: out = 2530;
			8512: out = -1282;
			8513: out = -5499;
			8514: out = 56;
			8515: out = 1491;
			8516: out = 1074;
			8517: out = -1444;
			8518: out = -1716;
			8519: out = 1040;
			8520: out = 4525;
			8521: out = 1266;
			8522: out = -2305;
			8523: out = -4591;
			8524: out = 652;
			8525: out = -1360;
			8526: out = 790;
			8527: out = 1874;
			8528: out = 6245;
			8529: out = -1237;
			8530: out = -6887;
			8531: out = -6374;
			8532: out = -569;
			8533: out = 2426;
			8534: out = 1098;
			8535: out = -730;
			8536: out = -1782;
			8537: out = 533;
			8538: out = 4434;
			8539: out = 1095;
			8540: out = -2507;
			8541: out = -5056;
			8542: out = 752;
			8543: out = -105;
			8544: out = 1609;
			8545: out = 5391;
			8546: out = 1166;
			8547: out = -2178;
			8548: out = -3809;
			8549: out = -2732;
			8550: out = 584;
			8551: out = 1998;
			8552: out = 1166;
			8553: out = -2076;
			8554: out = -368;
			8555: out = 2727;
			8556: out = -47;
			8557: out = -2353;
			8558: out = -2937;
			8559: out = 2936;
			8560: out = -1690;
			8561: out = 2780;
			8562: out = 6585;
			8563: out = 5093;
			8564: out = 1776;
			8565: out = -1778;
			8566: out = -3830;
			8567: out = 2258;
			8568: out = 2668;
			8569: out = 53;
			8570: out = -1776;
			8571: out = -647;
			8572: out = 1101;
			8573: out = -278;
			8574: out = 623;
			8575: out = -2300;
			8576: out = -2402;
			8577: out = 1324;
			8578: out = 4075;
			8579: out = 1244;
			8580: out = -5154;
			8581: out = -4286;
			8582: out = 345;
			8583: out = 4612;
			8584: out = -14;
			8585: out = -408;
			8586: out = -1881;
			8587: out = -285;
			8588: out = -3127;
			8589: out = 935;
			8590: out = 2752;
			8591: out = -2113;
			8592: out = -4455;
			8593: out = -2902;
			8594: out = 3947;
			8595: out = -1230;
			8596: out = 2085;
			8597: out = 2783;
			8598: out = 1560;
			8599: out = -4159;
			8600: out = -2070;
			8601: out = 4937;
			8602: out = 584;
			8603: out = -2644;
			8604: out = -5120;
			8605: out = -67;
			8606: out = 1199;
			8607: out = 2654;
			8608: out = 691;
			8609: out = 4805;
			8610: out = -288;
			8611: out = -4524;
			8612: out = -7394;
			8613: out = 867;
			8614: out = 4265;
			8615: out = 2701;
			8616: out = 1078;
			8617: out = 249;
			8618: out = 18;
			8619: out = -2257;
			8620: out = 1411;
			8621: out = 1916;
			8622: out = -462;
			8623: out = -1994;
			8624: out = -4892;
			8625: out = -3001;
			8626: out = 4600;
			8627: out = 1720;
			8628: out = -2645;
			8629: out = -6651;
			8630: out = -253;
			8631: out = 1500;
			8632: out = 3042;
			8633: out = 3725;
			8634: out = -1025;
			8635: out = -4972;
			8636: out = -5274;
			8637: out = 7610;
			8638: out = 3211;
			8639: out = -1703;
			8640: out = -1376;
			8641: out = -337;
			8642: out = 2028;
			8643: out = 2024;
			8644: out = 3871;
			8645: out = -2158;
			8646: out = -3975;
			8647: out = 1045;
			8648: out = -347;
			8649: out = -306;
			8650: out = -298;
			8651: out = 4940;
			8652: out = 2652;
			8653: out = 635;
			8654: out = -1792;
			8655: out = -748;
			8656: out = -860;
			8657: out = 232;
			8658: out = -551;
			8659: out = 3702;
			8660: out = 3436;
			8661: out = 196;
			8662: out = -2128;
			8663: out = 309;
			8664: out = 2111;
			8665: out = -3474;
			8666: out = -5039;
			8667: out = -3709;
			8668: out = 880;
			8669: out = 315;
			8670: out = -177;
			8671: out = -658;
			8672: out = 339;
			8673: out = 420;
			8674: out = -1132;
			8675: out = -2266;
			8676: out = -481;
			8677: out = 4397;
			8678: out = 5673;
			8679: out = 1248;
			8680: out = -6512;
			8681: out = -7354;
			8682: out = -106;
			8683: out = -470;
			8684: out = 414;
			8685: out = -278;
			8686: out = 33;
			8687: out = 3562;
			8688: out = 4755;
			8689: out = 2473;
			8690: out = -1348;
			8691: out = -2513;
			8692: out = -928;
			8693: out = 2981;
			8694: out = 794;
			8695: out = 2236;
			8696: out = 5278;
			8697: out = 3159;
			8698: out = 694;
			8699: out = -1313;
			8700: out = 375;
			8701: out = -1408;
			8702: out = -1354;
			8703: out = -55;
			8704: out = 67;
			8705: out = 433;
			8706: out = -949;
			8707: out = -418;
			8708: out = -8831;
			8709: out = -4547;
			8710: out = 5935;
			8711: out = 4379;
			8712: out = 2392;
			8713: out = -1388;
			8714: out = 1013;
			8715: out = -4050;
			8716: out = -1543;
			8717: out = 1935;
			8718: out = 1054;
			8719: out = -234;
			8720: out = 200;
			8721: out = 4916;
			8722: out = -3183;
			8723: out = -5403;
			8724: out = -4704;
			8725: out = -203;
			8726: out = -2116;
			8727: out = -2327;
			8728: out = 1719;
			8729: out = 106;
			8730: out = 122;
			8731: out = 710;
			8732: out = 5586;
			8733: out = 2288;
			8734: out = -3268;
			8735: out = -10097;
			8736: out = -2458;
			8737: out = 2655;
			8738: out = 4629;
			8739: out = 1809;
			8740: out = -647;
			8741: out = -1565;
			8742: out = 1827;
			8743: out = -2031;
			8744: out = -79;
			8745: out = 803;
			8746: out = -1563;
			8747: out = -3653;
			8748: out = -1767;
			8749: out = 2649;
			8750: out = 3489;
			8751: out = 206;
			8752: out = -3942;
			8753: out = -4129;
			8754: out = -970;
			8755: out = 1913;
			8756: out = 2122;
			8757: out = -1159;
			8758: out = -1471;
			8759: out = -266;
			8760: out = -642;
			8761: out = -950;
			8762: out = -528;
			8763: out = 1082;
			8764: out = 1756;
			8765: out = 1364;
			8766: out = -102;
			8767: out = -3122;
			8768: out = 974;
			8769: out = 2303;
			8770: out = 179;
			8771: out = 953;
			8772: out = 1104;
			8773: out = 2333;
			8774: out = 3133;
			8775: out = 2741;
			8776: out = 217;
			8777: out = -3533;
			8778: out = 390;
			8779: out = 102;
			8780: out = 48;
			8781: out = -1691;
			8782: out = 2911;
			8783: out = 2622;
			8784: out = 302;
			8785: out = -1532;
			8786: out = 1884;
			8787: out = 3899;
			8788: out = 1414;
			8789: out = -3252;
			8790: out = -3001;
			8791: out = 2143;
			8792: out = 3963;
			8793: out = 2183;
			8794: out = -1042;
			8795: out = 123;
			8796: out = -602;
			8797: out = 179;
			8798: out = -665;
			8799: out = -1632;
			8800: out = -3557;
			8801: out = -3126;
			8802: out = -117;
			8803: out = -1028;
			8804: out = -2673;
			8805: out = -4339;
			8806: out = 483;
			8807: out = 389;
			8808: out = 1960;
			8809: out = 5077;
			8810: out = 2654;
			8811: out = -838;
			8812: out = -3410;
			8813: out = -3453;
			8814: out = 713;
			8815: out = 2328;
			8816: out = -1851;
			8817: out = -603;
			8818: out = -522;
			8819: out = 737;
			8820: out = 3964;
			8821: out = 1807;
			8822: out = -1494;
			8823: out = -3024;
			8824: out = -3565;
			8825: out = -1022;
			8826: out = 1544;
			8827: out = 497;
			8828: out = 442;
			8829: out = -39;
			8830: out = 709;
			8831: out = -195;
			8832: out = 1317;
			8833: out = 1916;
			8834: out = 846;
			8835: out = -2237;
			8836: out = -2361;
			8837: out = 638;
			8838: out = 299;
			8839: out = -2708;
			8840: out = -5530;
			8841: out = 888;
			8842: out = 800;
			8843: out = 1905;
			8844: out = 2127;
			8845: out = 2944;
			8846: out = 1335;
			8847: out = -575;
			8848: out = -2465;
			8849: out = -1837;
			8850: out = -46;
			8851: out = 2348;
			8852: out = -2679;
			8853: out = -977;
			8854: out = 3229;
			8855: out = 5469;
			8856: out = 3537;
			8857: out = -2239;
			8858: out = -8042;
			8859: out = -2801;
			8860: out = 458;
			8861: out = 1962;
			8862: out = 2329;
			8863: out = 1639;
			8864: out = 2474;
			8865: out = 3308;
			8866: out = -695;
			8867: out = -3337;
			8868: out = -2314;
			8869: out = 4676;
			8870: out = 3633;
			8871: out = 1083;
			8872: out = -2442;
			8873: out = -299;
			8874: out = -1035;
			8875: out = -674;
			8876: out = 3974;
			8877: out = -202;
			8878: out = 253;
			8879: out = 2621;
			8880: out = 1155;
			8881: out = -3047;
			8882: out = -5692;
			8883: out = 478;
			8884: out = -788;
			8885: out = -18;
			8886: out = -918;
			8887: out = 5813;
			8888: out = -89;
			8889: out = -3211;
			8890: out = 800;
			8891: out = 322;
			8892: out = -1395;
			8893: out = -4492;
			8894: out = -4933;
			8895: out = -2721;
			8896: out = 363;
			8897: out = 356;
			8898: out = 1859;
			8899: out = 1105;
			8900: out = 824;
			8901: out = 2026;
			8902: out = 1035;
			8903: out = -1598;
			8904: out = -3580;
			8905: out = -4780;
			8906: out = -220;
			8907: out = 5147;
			8908: out = -516;
			8909: out = 1066;
			8910: out = 706;
			8911: out = 251;
			8912: out = -346;
			8913: out = 2110;
			8914: out = 3937;
			8915: out = 1054;
			8916: out = 554;
			8917: out = -759;
			8918: out = -4248;
			8919: out = 1144;
			8920: out = 771;
			8921: out = -493;
			8922: out = -2884;
			8923: out = 2767;
			8924: out = 4483;
			8925: out = 921;
			8926: out = -2458;
			8927: out = -2747;
			8928: out = -1159;
			8929: out = -2001;
			8930: out = -3303;
			8931: out = -2587;
			8932: out = 1203;
			8933: out = 3755;
			8934: out = 902;
			8935: out = -3833;
			8936: out = 879;
			8937: out = -1893;
			8938: out = -566;
			8939: out = 1071;
			8940: out = -165;
			8941: out = -1124;
			8942: out = 252;
			8943: out = 1843;
			8944: out = 5031;
			8945: out = 3876;
			8946: out = 341;
			8947: out = -7681;
			8948: out = -5193;
			8949: out = 1333;
			8950: out = 2582;
			8951: out = 3810;
			8952: out = 1605;
			8953: out = -566;
			8954: out = -5311;
			8955: out = -4287;
			8956: out = -940;
			8957: out = 2723;
			8958: out = 3884;
			8959: out = 3826;
			8960: out = 2556;
			8961: out = -1365;
			8962: out = -3020;
			8963: out = -2533;
			8964: out = -94;
			8965: out = 1231;
			8966: out = 1612;
			8967: out = 1076;
			8968: out = 4041;
			8969: out = 1521;
			8970: out = -723;
			8971: out = 491;
			8972: out = -829;
			8973: out = -1052;
			8974: out = -1504;
			8975: out = 350;
			8976: out = -211;
			8977: out = 11;
			8978: out = 338;
			8979: out = 1605;
			8980: out = -231;
			8981: out = -2926;
			8982: out = -2536;
			8983: out = -301;
			8984: out = 907;
			8985: out = -2265;
			8986: out = 427;
			8987: out = 316;
			8988: out = 289;
			8989: out = 2010;
			8990: out = 984;
			8991: out = -577;
			8992: out = -466;
			8993: out = -2068;
			8994: out = 208;
			8995: out = 2951;
			8996: out = 2472;
			8997: out = 1296;
			8998: out = 143;
			8999: out = 397;
			9000: out = -367;
			9001: out = 511;
			9002: out = 1533;
			9003: out = -296;
			9004: out = 348;
			9005: out = -805;
			9006: out = -3292;
			9007: out = -2310;
			9008: out = -874;
			9009: out = 249;
			9010: out = 2218;
			9011: out = -1073;
			9012: out = -1840;
			9013: out = 2077;
			9014: out = -63;
			9015: out = -186;
			9016: out = -1525;
			9017: out = -4687;
			9018: out = -3635;
			9019: out = -321;
			9020: out = 3461;
			9021: out = 3824;
			9022: out = 3336;
			9023: out = 352;
			9024: out = -7245;
			9025: out = -6855;
			9026: out = -2424;
			9027: out = 2999;
			9028: out = 709;
			9029: out = -1577;
			9030: out = -1897;
			9031: out = 5201;
			9032: out = 3398;
			9033: out = 1998;
			9034: out = 826;
			9035: out = -2884;
			9036: out = -4633;
			9037: out = -3411;
			9038: out = 3865;
			9039: out = 2526;
			9040: out = 2738;
			9041: out = 3928;
			9042: out = 1454;
			9043: out = -359;
			9044: out = -1341;
			9045: out = -165;
			9046: out = 155;
			9047: out = 327;
			9048: out = 445;
			9049: out = 1299;
			9050: out = 1993;
			9051: out = 1186;
			9052: out = -1883;
			9053: out = -1527;
			9054: out = 1377;
			9055: out = 4977;
			9056: out = 4189;
			9057: out = 2090;
			9058: out = -1382;
			9059: out = -5084;
			9060: out = -3903;
			9061: out = -2756;
			9062: out = -2359;
			9063: out = 27;
			9064: out = 1665;
			9065: out = 2519;
			9066: out = 1266;
			9067: out = 733;
			9068: out = -1037;
			9069: out = -2617;
			9070: out = 820;
			9071: out = -280;
			9072: out = -1619;
			9073: out = 13;
			9074: out = -612;
			9075: out = 974;
			9076: out = 2524;
			9077: out = 1548;
			9078: out = 61;
			9079: out = -1160;
			9080: out = -144;
			9081: out = -1995;
			9082: out = -122;
			9083: out = 3101;
			9084: out = -2770;
			9085: out = -1024;
			9086: out = -62;
			9087: out = -273;
			9088: out = -2851;
			9089: out = -1206;
			9090: out = 2563;
			9091: out = -413;
			9092: out = 1149;
			9093: out = 1309;
			9094: out = 894;
			9095: out = -3412;
			9096: out = -4374;
			9097: out = -2285;
			9098: out = -122;
			9099: out = 2783;
			9100: out = 3011;
			9101: out = 793;
			9102: out = 22;
			9103: out = -239;
			9104: out = -604;
			9105: out = -5629;
			9106: out = -3069;
			9107: out = 150;
			9108: out = 1583;
			9109: out = 3136;
			9110: out = 1880;
			9111: out = -151;
			9112: out = -3042;
			9113: out = -815;
			9114: out = 1709;
			9115: out = 2904;
			9116: out = -663;
			9117: out = -1226;
			9118: out = 292;
			9119: out = 193;
			9120: out = 3389;
			9121: out = 3732;
			9122: out = 916;
			9123: out = 654;
			9124: out = -467;
			9125: out = -143;
			9126: out = -705;
			9127: out = 497;
			9128: out = -180;
			9129: out = -210;
			9130: out = -4521;
			9131: out = -1253;
			9132: out = 2222;
			9133: out = 3985;
			9134: out = -1058;
			9135: out = -2011;
			9136: out = 866;
			9137: out = 4467;
			9138: out = 89;
			9139: out = -6245;
			9140: out = -8127;
			9141: out = -2304;
			9142: out = 1886;
			9143: out = 517;
			9144: out = 2068;
			9145: out = 366;
			9146: out = 554;
			9147: out = 3041;
			9148: out = -2759;
			9149: out = -6094;
			9150: out = -4799;
			9151: out = -3104;
			9152: out = 713;
			9153: out = 2439;
			9154: out = 1623;
			9155: out = 647;
			9156: out = -752;
			9157: out = -1770;
			9158: out = -1252;
			9159: out = 303;
			9160: out = 1072;
			9161: out = -1452;
			9162: out = 606;
			9163: out = -26;
			9164: out = -919;
			9165: out = 2612;
			9166: out = 1534;
			9167: out = 359;
			9168: out = 2100;
			9169: out = 809;
			9170: out = 2097;
			9171: out = 2056;
			9172: out = 986;
			9173: out = -3416;
			9174: out = -3116;
			9175: out = 3442;
			9176: out = 2821;
			9177: out = -361;
			9178: out = -4438;
			9179: out = 436;
			9180: out = 1761;
			9181: out = 2094;
			9182: out = -1178;
			9183: out = 162;
			9184: out = -171;
			9185: out = -78;
			9186: out = -2525;
			9187: out = -1626;
			9188: out = -490;
			9189: out = 1974;
			9190: out = 376;
			9191: out = 2170;
			9192: out = 2831;
			9193: out = -2209;
			9194: out = -4670;
			9195: out = -4262;
			9196: out = 638;
			9197: out = 2300;
			9198: out = 3378;
			9199: out = 2019;
			9200: out = 3028;
			9201: out = -1531;
			9202: out = -3484;
			9203: out = -3389;
			9204: out = 2660;
			9205: out = 3109;
			9206: out = 1088;
			9207: out = -3702;
			9208: out = 292;
			9209: out = 2072;
			9210: out = -169;
			9211: out = -2979;
			9212: out = -1993;
			9213: out = 1725;
			9214: out = 2020;
			9215: out = 2400;
			9216: out = -172;
			9217: out = -2384;
			9218: out = -3309;
			9219: out = 236;
			9220: out = 3294;
			9221: out = 119;
			9222: out = 1210;
			9223: out = 620;
			9224: out = 517;
			9225: out = -3503;
			9226: out = -1816;
			9227: out = 151;
			9228: out = -176;
			9229: out = -1395;
			9230: out = -1132;
			9231: out = 750;
			9232: out = 1951;
			9233: out = 1093;
			9234: out = -432;
			9235: out = -1191;
			9236: out = -269;
			9237: out = -84;
			9238: out = -761;
			9239: out = -1807;
			9240: out = 695;
			9241: out = 2690;
			9242: out = 50;
			9243: out = 144;
			9244: out = 600;
			9245: out = 2720;
			9246: out = -2453;
			9247: out = -911;
			9248: out = 305;
			9249: out = 1252;
			9250: out = 214;
			9251: out = 1870;
			9252: out = 3645;
			9253: out = 763;
			9254: out = -1570;
			9255: out = -1772;
			9256: out = 2212;
			9257: out = 1491;
			9258: out = 785;
			9259: out = -406;
			9260: out = -1339;
			9261: out = -813;
			9262: out = -146;
			9263: out = -71;
			9264: out = -418;
			9265: out = 1419;
			9266: out = 3767;
			9267: out = -266;
			9268: out = 156;
			9269: out = 754;
			9270: out = 2342;
			9271: out = -2688;
			9272: out = -4322;
			9273: out = -3071;
			9274: out = -82;
			9275: out = 456;
			9276: out = 873;
			9277: out = 4150;
			9278: out = -3375;
			9279: out = -2223;
			9280: out = 1424;
			9281: out = -233;
			9282: out = -2633;
			9283: out = -3685;
			9284: out = 1161;
			9285: out = -1724;
			9286: out = 1303;
			9287: out = 3164;
			9288: out = -99;
			9289: out = -1143;
			9290: out = -732;
			9291: out = 486;
			9292: out = 130;
			9293: out = -2264;
			9294: out = -3530;
			9295: out = 3160;
			9296: out = 1023;
			9297: out = -688;
			9298: out = -1100;
			9299: out = -575;
			9300: out = 1815;
			9301: out = 3505;
			9302: out = 1813;
			9303: out = 1003;
			9304: out = 101;
			9305: out = 119;
			9306: out = -4921;
			9307: out = -4062;
			9308: out = -981;
			9309: out = -1747;
			9310: out = 1922;
			9311: out = 1912;
			9312: out = 429;
			9313: out = -2871;
			9314: out = 651;
			9315: out = 3219;
			9316: out = -5995;
			9317: out = -1399;
			9318: out = 1392;
			9319: out = 3587;
			9320: out = -991;
			9321: out = -411;
			9322: out = 710;
			9323: out = 1665;
			9324: out = -578;
			9325: out = -887;
			9326: out = 690;
			9327: out = 1371;
			9328: out = 768;
			9329: out = -827;
			9330: out = -1634;
			9331: out = -456;
			9332: out = 1671;
			9333: out = 2748;
			9334: out = 266;
			9335: out = -572;
			9336: out = -1132;
			9337: out = -3145;
			9338: out = 472;
			9339: out = 2716;
			9340: out = 3531;
			9341: out = -613;
			9342: out = -407;
			9343: out = -310;
			9344: out = -1321;
			9345: out = -1566;
			9346: out = 770;
			9347: out = 3948;
			9348: out = -155;
			9349: out = -387;
			9350: out = -1189;
			9351: out = -1143;
			9352: out = -589;
			9353: out = 1058;
			9354: out = 1790;
			9355: out = 1131;
			9356: out = -589;
			9357: out = -2012;
			9358: out = -3762;
			9359: out = -147;
			9360: out = 643;
			9361: out = 344;
			9362: out = -1946;
			9363: out = 440;
			9364: out = 1325;
			9365: out = -93;
			9366: out = -1195;
			9367: out = 180;
			9368: out = 2094;
			9369: out = 294;
			9370: out = -492;
			9371: out = -417;
			9372: out = 493;
			9373: out = 1499;
			9374: out = 131;
			9375: out = -1838;
			9376: out = -4929;
			9377: out = 1291;
			9378: out = 4366;
			9379: out = 680;
			9380: out = -26;
			9381: out = -726;
			9382: out = 1428;
			9383: out = 3241;
			9384: out = 2895;
			9385: out = -130;
			9386: out = -3207;
			9387: out = -3278;
			9388: out = -1928;
			9389: out = -30;
			9390: out = 2844;
			9391: out = 2156;
			9392: out = 1625;
			9393: out = 1225;
			9394: out = 1016;
			9395: out = -913;
			9396: out = -2781;
			9397: out = -571;
			9398: out = -2282;
			9399: out = -1703;
			9400: out = 150;
			9401: out = 161;
			9402: out = 597;
			9403: out = 1284;
			9404: out = 2238;
			9405: out = 1032;
			9406: out = -1622;
			9407: out = -4222;
			9408: out = -1249;
			9409: out = 897;
			9410: out = 1819;
			9411: out = 110;
			9412: out = -836;
			9413: out = -1595;
			9414: out = -963;
			9415: out = 1062;
			9416: out = 1507;
			9417: out = 14;
			9418: out = -2305;
			9419: out = -1464;
			9420: out = 306;
			9421: out = 791;
			9422: out = 1378;
			9423: out = -2137;
			9424: out = -3887;
			9425: out = -983;
			9426: out = 1954;
			9427: out = 2240;
			9428: out = -1028;
			9429: out = -1754;
			9430: out = -2577;
			9431: out = -590;
			9432: out = 817;
			9433: out = 3676;
			9434: out = 2148;
			9435: out = -401;
			9436: out = -1820;
			9437: out = -468;
			9438: out = 390;
			9439: out = 57;
			9440: out = -3303;
			9441: out = -2502;
			9442: out = 735;
			9443: out = 195;
			9444: out = 585;
			9445: out = 538;
			9446: out = 1143;
			9447: out = 234;
			9448: out = -1157;
			9449: out = -1844;
			9450: out = 2368;
			9451: out = 2639;
			9452: out = 1812;
			9453: out = 246;
			9454: out = -1936;
			9455: out = -1233;
			9456: out = 933;
			9457: out = 382;
			9458: out = -150;
			9459: out = -2;
			9460: out = 3267;
			9461: out = -9;
			9462: out = -62;
			9463: out = 307;
			9464: out = 4213;
			9465: out = 1114;
			9466: out = -1148;
			9467: out = -2515;
			9468: out = 614;
			9469: out = 107;
			9470: out = -597;
			9471: out = 698;
			9472: out = 3488;
			9473: out = 3151;
			9474: out = -802;
			9475: out = -1723;
			9476: out = -332;
			9477: out = 2222;
			9478: out = 1464;
			9479: out = 144;
			9480: out = -1518;
			9481: out = -1194;
			9482: out = -725;
			9483: out = -179;
			9484: out = -421;
			9485: out = 478;
			9486: out = -120;
			9487: out = -324;
			9488: out = -960;
			9489: out = -359;
			9490: out = 382;
			9491: out = 1568;
			9492: out = 473;
			9493: out = 855;
			9494: out = -1427;
			9495: out = -4034;
			9496: out = -1022;
			9497: out = 1286;
			9498: out = 1199;
			9499: out = -508;
			9500: out = -4363;
			9501: out = -3684;
			9502: out = 1131;
			9503: out = 4593;
			9504: out = 3345;
			9505: out = -696;
			9506: out = -3771;
			9507: out = -3555;
			9508: out = -2370;
			9509: out = -2025;
			9510: out = 3647;
			9511: out = 2724;
			9512: out = -184;
			9513: out = -2007;
			9514: out = -853;
			9515: out = 1719;
			9516: out = 1769;
			9517: out = 1856;
			9518: out = -4418;
			9519: out = -6761;
			9520: out = 677;
			9521: out = 4005;
			9522: out = 2690;
			9523: out = -3440;
			9524: out = -4023;
			9525: out = -2312;
			9526: out = 2167;
			9527: out = 2205;
			9528: out = 4022;
			9529: out = 669;
			9530: out = -2450;
			9531: out = -2152;
			9532: out = 1143;
			9533: out = 3134;
			9534: out = 2696;
			9535: out = -433;
			9536: out = -1252;
			9537: out = -59;
			9538: out = -305;
			9539: out = -1531;
			9540: out = -1958;
			9541: out = 1357;
			9542: out = -570;
			9543: out = -914;
			9544: out = -1217;
			9545: out = 536;
			9546: out = 981;
			9547: out = 1494;
			9548: out = -19;
			9549: out = 3704;
			9550: out = 2503;
			9551: out = -404;
			9552: out = -3455;
			9553: out = -1024;
			9554: out = 1973;
			9555: out = 2416;
			9556: out = 610;
			9557: out = -1145;
			9558: out = -737;
			9559: out = 2919;
			9560: out = 2147;
			9561: out = 558;
			9562: out = 132;
			9563: out = -2777;
			9564: out = -2968;
			9565: out = -2029;
			9566: out = 889;
			9567: out = 319;
			9568: out = 777;
			9569: out = 2320;
			9570: out = 1880;
			9571: out = 420;
			9572: out = -807;
			9573: out = 2860;
			9574: out = -1680;
			9575: out = -4449;
			9576: out = -3204;
			9577: out = -5072;
			9578: out = -2057;
			9579: out = 1225;
			9580: out = 4135;
			9581: out = 974;
			9582: out = 45;
			9583: out = 1985;
			9584: out = -993;
			9585: out = -2650;
			9586: out = -2906;
			9587: out = 2144;
			9588: out = 618;
			9589: out = 534;
			9590: out = 1514;
			9591: out = 338;
			9592: out = 729;
			9593: out = 700;
			9594: out = 465;
			9595: out = -679;
			9596: out = -605;
			9597: out = -446;
			9598: out = 709;
			9599: out = -3181;
			9600: out = -5649;
			9601: out = -203;
			9602: out = 956;
			9603: out = 2752;
			9604: out = 2311;
			9605: out = 298;
			9606: out = -1475;
			9607: out = -1919;
			9608: out = -3094;
			9609: out = 257;
			9610: out = 751;
			9611: out = -248;
			9612: out = 462;
			9613: out = 1366;
			9614: out = 1513;
			9615: out = -949;
			9616: out = 139;
			9617: out = 407;
			9618: out = 214;
			9619: out = -2102;
			9620: out = -3753;
			9621: out = -4000;
			9622: out = -67;
			9623: out = -2321;
			9624: out = 120;
			9625: out = 3644;
			9626: out = 5968;
			9627: out = 2398;
			9628: out = -1178;
			9629: out = -252;
			9630: out = -319;
			9631: out = 822;
			9632: out = -83;
			9633: out = -132;
			9634: out = -3580;
			9635: out = -3064;
			9636: out = 1880;
			9637: out = 2236;
			9638: out = 1653;
			9639: out = 75;
			9640: out = -1081;
			9641: out = -319;
			9642: out = 526;
			9643: out = 170;
			9644: out = -1344;
			9645: out = -719;
			9646: out = 1441;
			9647: out = -559;
			9648: out = 2809;
			9649: out = 4157;
			9650: out = 3654;
			9651: out = -128;
			9652: out = -417;
			9653: out = 1010;
			9654: out = -1191;
			9655: out = -524;
			9656: out = -1858;
			9657: out = -3347;
			9658: out = -1912;
			9659: out = 806;
			9660: out = 2393;
			9661: out = 2307;
			9662: out = 1149;
			9663: out = 739;
			9664: out = -2;
			9665: out = 378;
			9666: out = -3255;
			9667: out = -5890;
			9668: out = -3962;
			9669: out = 1941;
			9670: out = 5058;
			9671: out = 3207;
			9672: out = -854;
			9673: out = -1852;
			9674: out = -214;
			9675: out = -579;
			9676: out = 473;
			9677: out = 412;
			9678: out = 1031;
			9679: out = 146;
			9680: out = 294;
			9681: out = 412;
			9682: out = 2403;
			9683: out = 546;
			9684: out = 178;
			9685: out = 284;
			9686: out = 1785;
			9687: out = -1133;
			9688: out = -3693;
			9689: out = 210;
			9690: out = -1592;
			9691: out = 729;
			9692: out = 3929;
			9693: out = 388;
			9694: out = -800;
			9695: out = -1636;
			9696: out = -1820;
			9697: out = -1217;
			9698: out = 151;
			9699: out = 1089;
			9700: out = -3595;
			9701: out = -3398;
			9702: out = -673;
			9703: out = 4061;
			9704: out = 795;
			9705: out = -839;
			9706: out = -392;
			9707: out = 1066;
			9708: out = 752;
			9709: out = -1269;
			9710: out = -2592;
			9711: out = -3720;
			9712: out = -727;
			9713: out = 3184;
			9714: out = 1357;
			9715: out = 566;
			9716: out = -444;
			9717: out = 107;
			9718: out = -1478;
			9719: out = -2023;
			9720: out = -2091;
			9721: out = 305;
			9722: out = 0;
			9723: out = 323;
			9724: out = 2032;
			9725: out = 628;
			9726: out = -397;
			9727: out = -1199;
			9728: out = 624;
			9729: out = -383;
			9730: out = 212;
			9731: out = 3423;
			9732: out = 374;
			9733: out = -26;
			9734: out = 257;
			9735: out = -243;
			9736: out = -984;
			9737: out = -195;
			9738: out = 4002;
			9739: out = -14;
			9740: out = 1065;
			9741: out = 1976;
			9742: out = 1073;
			9743: out = -3059;
			9744: out = -3331;
			9745: out = 2486;
			9746: out = 1019;
			9747: out = 859;
			9748: out = -401;
			9749: out = 2091;
			9750: out = -1014;
			9751: out = -1596;
			9752: out = -312;
			9753: out = -1113;
			9754: out = -2013;
			9755: out = -1781;
			9756: out = 1298;
			9757: out = 1450;
			9758: out = 1050;
			9759: out = 788;
			9760: out = -1620;
			9761: out = -1061;
			9762: out = 497;
			9763: out = 2625;
			9764: out = 611;
			9765: out = -1264;
			9766: out = -2224;
			9767: out = 2148;
			9768: out = 2096;
			9769: out = 630;
			9770: out = -1417;
			9771: out = -612;
			9772: out = -524;
			9773: out = -836;
			9774: out = -2467;
			9775: out = -322;
			9776: out = 1606;
			9777: out = 1252;
			9778: out = -293;
			9779: out = -580;
			9780: out = 182;
			9781: out = 48;
			9782: out = -1292;
			9783: out = -1164;
			9784: out = 1199;
			9785: out = 2350;
			9786: out = -44;
			9787: out = -3861;
			9788: out = -5244;
			9789: out = -411;
			9790: out = 3843;
			9791: out = 1834;
			9792: out = -265;
			9793: out = -453;
			9794: out = 2707;
			9795: out = -534;
			9796: out = -620;
			9797: out = -1466;
			9798: out = 335;
			9799: out = -3074;
			9800: out = -1916;
			9801: out = 1088;
			9802: out = 2844;
			9803: out = 2007;
			9804: out = -51;
			9805: out = -1141;
			9806: out = -1945;
			9807: out = -934;
			9808: out = 4;
			9809: out = 577;
			9810: out = -1936;
			9811: out = -3016;
			9812: out = 562;
			9813: out = -26;
			9814: out = 1980;
			9815: out = 2822;
			9816: out = 543;
			9817: out = -1891;
			9818: out = -2526;
			9819: out = -418;
			9820: out = -217;
			9821: out = 306;
			9822: out = 567;
			9823: out = 1424;
			9824: out = 131;
			9825: out = -1288;
			9826: out = -1425;
			9827: out = 567;
			9828: out = 3415;
			9829: out = 3536;
			9830: out = -4171;
			9831: out = -6414;
			9832: out = -5120;
			9833: out = 880;
			9834: out = -9;
			9835: out = 1336;
			9836: out = 1392;
			9837: out = 2222;
			9838: out = 580;
			9839: out = 575;
			9840: out = 210;
			9841: out = 1021;
			9842: out = -2446;
			9843: out = -5099;
			9844: out = -4429;
			9845: out = 1703;
			9846: out = 4065;
			9847: out = 815;
			9848: out = -378;
			9849: out = -1468;
			9850: out = -509;
			9851: out = 1028;
			9852: out = -730;
			9853: out = -916;
			9854: out = 2087;
			9855: out = 276;
			9856: out = 1544;
			9857: out = 1629;
			9858: out = 602;
			9859: out = 707;
			9860: out = 1156;
			9861: out = 797;
			9862: out = 2371;
			9863: out = 823;
			9864: out = -674;
			9865: out = -1798;
			9866: out = -427;
			9867: out = 176;
			9868: out = 295;
			9869: out = -3617;
			9870: out = -1988;
			9871: out = 1242;
			9872: out = 4735;
			9873: out = 1437;
			9874: out = 63;
			9875: out = 252;
			9876: out = -194;
			9877: out = -860;
			9878: out = -1890;
			9879: out = -5291;
			9880: out = 2219;
			9881: out = 2871;
			9882: out = -515;
			9883: out = 3489;
			9884: out = 2770;
			9885: out = 1079;
			9886: out = -1869;
			9887: out = -4106;
			9888: out = -3164;
			9889: out = -44;
			9890: out = 1167;
			9891: out = 661;
			9892: out = -139;
			9893: out = 555;
			9894: out = 308;
			9895: out = -1;
			9896: out = -93;
			9897: out = -438;
			9898: out = 2534;
			9899: out = 3162;
			9900: out = -226;
			9901: out = -5309;
			9902: out = -5583;
			9903: out = -852;
			9904: out = -1923;
			9905: out = 2833;
			9906: out = 3185;
			9907: out = 829;
			9908: out = -1636;
			9909: out = -2231;
			9910: out = -1703;
			9911: out = 1584;
			9912: out = 74;
			9913: out = -714;
			9914: out = -1073;
			9915: out = 3394;
			9916: out = 2449;
			9917: out = 129;
			9918: out = 349;
			9919: out = 1136;
			9920: out = 508;
			9921: out = -1857;
			9922: out = -5057;
			9923: out = -2400;
			9924: out = 2331;
			9925: out = 571;
			9926: out = 694;
			9927: out = 84;
			9928: out = 1711;
			9929: out = -2356;
			9930: out = -1465;
			9931: out = 280;
			9932: out = -73;
			9933: out = 594;
			9934: out = -118;
			9935: out = -1542;
			9936: out = 263;
			9937: out = 1190;
			9938: out = 1232;
			9939: out = 110;
			9940: out = -2;
			9941: out = -169;
			9942: out = -1142;
			9943: out = 2545;
			9944: out = 1511;
			9945: out = -318;
			9946: out = -3381;
			9947: out = 2567;
			9948: out = 3693;
			9949: out = -1006;
			9950: out = 427;
			9951: out = -176;
			9952: out = 747;
			9953: out = -619;
			9954: out = 1974;
			9955: out = 506;
			9956: out = -3017;
			9957: out = -1280;
			9958: out = -47;
			9959: out = 1230;
			9960: out = 1201;
			9961: out = 632;
			9962: out = 775;
			9963: out = 2724;
			9964: out = -3270;
			9965: out = -484;
			9966: out = 1733;
			9967: out = -960;
			9968: out = -320;
			9969: out = 44;
			9970: out = 348;
			9971: out = 2;
			9972: out = -475;
			9973: out = -1199;
			9974: out = -3965;
			9975: out = -23;
			9976: out = 1412;
			9977: out = 1557;
			9978: out = -4704;
			9979: out = -537;
			9980: out = 2980;
			9981: out = -149;
			9982: out = -1075;
			9983: out = -800;
			9984: out = 1806;
			9985: out = 306;
			9986: out = -928;
			9987: out = -1957;
			9988: out = 1986;
			9989: out = -684;
			9990: out = 193;
			9991: out = 884;
			9992: out = 2018;
			9993: out = -517;
			9994: out = -1700;
			9995: out = -571;
			9996: out = 1692;
			9997: out = 1835;
			9998: out = 412;
			9999: out = -1084;
			10000: out = -1011;
			10001: out = -856;
			10002: out = -1727;
			10003: out = 1191;
			10004: out = 1515;
			10005: out = -13;
			10006: out = 1309;
			10007: out = -1769;
			10008: out = -2556;
			10009: out = -1620;
			10010: out = 2560;
			10011: out = 1678;
			10012: out = -439;
			10013: out = -169;
			10014: out = 2445;
			10015: out = 1769;
			10016: out = -3889;
			10017: out = -2769;
			10018: out = -1293;
			10019: out = 927;
			10020: out = 799;
			10021: out = 209;
			10022: out = 365;
			10023: out = 2365;
			10024: out = 1052;
			10025: out = -662;
			10026: out = -2323;
			10027: out = -64;
			10028: out = -904;
			10029: out = -1712;
			10030: out = -2607;
			10031: out = -125;
			10032: out = 1571;
			10033: out = 2011;
			10034: out = 348;
			10035: out = -1901;
			10036: out = -1846;
			10037: out = 1505;
			10038: out = -404;
			10039: out = 1072;
			10040: out = 1817;
			10041: out = 1865;
			10042: out = -86;
			10043: out = -388;
			10044: out = 1072;
			10045: out = -764;
			10046: out = 146;
			10047: out = 956;
			10048: out = 223;
			10049: out = 210;
			10050: out = -2195;
			10051: out = -5474;
			10052: out = 1812;
			10053: out = 1497;
			10054: out = -347;
			10055: out = -2661;
			10056: out = 32;
			10057: out = 999;
			10058: out = -266;
			10059: out = 1663;
			10060: out = -803;
			10061: out = -1649;
			10062: out = 2171;
			10063: out = 941;
			10064: out = 622;
			10065: out = -303;
			10066: out = 2358;
			10067: out = 652;
			10068: out = -985;
			10069: out = -4122;
			10070: out = 1039;
			10071: out = -191;
			10072: out = -3985;
			10073: out = -647;
			10074: out = 1145;
			10075: out = 2724;
			10076: out = 2930;
			10077: out = -1130;
			10078: out = -1610;
			10079: out = 845;
			10080: out = 121;
			10081: out = 1417;
			10082: out = 2051;
			10083: out = 2918;
			10084: out = -16;
			10085: out = -1320;
			10086: out = -874;
			10087: out = -389;
			10088: out = 1311;
			10089: out = 1211;
			10090: out = 202;
			10091: out = -2956;
			10092: out = -1334;
			10093: out = 1778;
			10094: out = 1085;
			10095: out = 151;
			10096: out = -1626;
			10097: out = -3236;
			10098: out = 1102;
			10099: out = 616;
			10100: out = -1296;
			10101: out = 970;
			10102: out = 1515;
			10103: out = 78;
			10104: out = -5274;
			10105: out = -443;
			10106: out = 238;
			10107: out = 567;
			10108: out = 1748;
			10109: out = 526;
			10110: out = -372;
			10111: out = 439;
			10112: out = -2020;
			10113: out = -1408;
			10114: out = -103;
			10115: out = 2245;
			10116: out = 847;
			10117: out = 215;
			10118: out = 410;
			10119: out = 84;
			10120: out = -692;
			10121: out = -977;
			10122: out = 238;
			10123: out = 1382;
			10124: out = 1268;
			10125: out = -383;
			10126: out = -1301;
			10127: out = -2321;
			10128: out = -2338;
			10129: out = -479;
			10130: out = -1040;
			10131: out = -475;
			10132: out = 637;
			10133: out = 536;
			10134: out = 225;
			10135: out = 215;
			10136: out = 932;
			10137: out = 1532;
			10138: out = 2265;
			10139: out = 3185;
			10140: out = -2409;
			10141: out = -1177;
			10142: out = 606;
			10143: out = 903;
			10144: out = -539;
			10145: out = 871;
			10146: out = 3653;
			10147: out = 106;
			10148: out = -3022;
			10149: out = -4130;
			10150: out = 1800;
			10151: out = 1008;
			10152: out = 1211;
			10153: out = 6;
			10154: out = 1148;
			10155: out = -896;
			10156: out = -1366;
			10157: out = 238;
			10158: out = 1441;
			10159: out = 812;
			10160: out = -772;
			10161: out = 2844;
			10162: out = 1245;
			10163: out = -203;
			10164: out = 229;
			10165: out = -305;
			10166: out = -1250;
			10167: out = -2798;
			10168: out = 2646;
			10169: out = -601;
			10170: out = -2026;
			10171: out = 523;
			10172: out = 753;
			10173: out = -877;
			10174: out = -3084;
			10175: out = 3207;
			10176: out = 1553;
			10177: out = -1365;
			10178: out = -5495;
			10179: out = -1367;
			10180: out = 1907;
			10181: out = 3417;
			10182: out = -708;
			10183: out = -196;
			10184: out = 267;
			10185: out = 127;
			10186: out = -188;
			10187: out = -131;
			10188: out = 219;
			10189: out = -343;
			10190: out = -811;
			10191: out = -1028;
			10192: out = 684;
			10193: out = -3009;
			10194: out = -975;
			10195: out = 2521;
			10196: out = 3760;
			10197: out = 1751;
			10198: out = -660;
			10199: out = -1043;
			10200: out = -1092;
			10201: out = -102;
			10202: out = -83;
			10203: out = -1092;
			10204: out = -2023;
			10205: out = -1309;
			10206: out = 1175;
			10207: out = 178;
			10208: out = 1584;
			10209: out = 2079;
			10210: out = -1312;
			10211: out = -1466;
			10212: out = -2214;
			10213: out = -3069;
			10214: out = 444;
			10215: out = 1071;
			10216: out = 992;
			10217: out = 2191;
			10218: out = 2072;
			10219: out = 1093;
			10220: out = -1663;
			10221: out = 455;
			10222: out = -1815;
			10223: out = -2819;
			10224: out = 554;
			10225: out = 283;
			10226: out = 412;
			10227: out = 833;
			10228: out = -2004;
			10229: out = -1045;
			10230: out = 512;
			10231: out = 2214;
			10232: out = -434;
			10233: out = -489;
			10234: out = 1432;
			10235: out = -585;
			10236: out = -1548;
			10237: out = -1754;
			10238: out = 607;
			10239: out = 1010;
			10240: out = 1405;
			10241: out = 1069;
			10242: out = -596;
			10243: out = 362;
			10244: out = 787;
			10245: out = -3059;
			10246: out = -349;
			10247: out = -800;
			10248: out = -2007;
			10249: out = 738;
			10250: out = 1454;
			10251: out = 1505;
			10252: out = 216;
			10253: out = 72;
			10254: out = -976;
			10255: out = -1643;
			10256: out = -2291;
			10257: out = 1027;
			10258: out = 2743;
			10259: out = -1271;
			10260: out = 1423;
			10261: out = -111;
			10262: out = -1842;
			10263: out = -3707;
			10264: out = -220;
			10265: out = 2205;
			10266: out = 1026;
			10267: out = 1524;
			10268: out = 584;
			10269: out = -386;
			10270: out = -592;
			10271: out = -245;
			10272: out = 686;
			10273: out = 673;
			10274: out = 2834;
			10275: out = 1345;
			10276: out = -458;
			10277: out = -415;
			10278: out = 2146;
			10279: out = 2175;
			10280: out = -1728;
			10281: out = -2438;
			10282: out = -1524;
			10283: out = 694;
			10284: out = -1529;
			10285: out = 1374;
			10286: out = 2792;
			10287: out = 2514;
			10288: out = 752;
			10289: out = -327;
			10290: out = -574;
			10291: out = -3575;
			10292: out = -22;
			10293: out = 1068;
			10294: out = 182;
			10295: out = -2132;
			10296: out = 421;
			10297: out = 3112;
			10298: out = -1062;
			10299: out = -2114;
			10300: out = -1388;
			10301: out = 3331;
			10302: out = -3956;
			10303: out = -2258;
			10304: out = 141;
			10305: out = -364;
			10306: out = 118;
			10307: out = 578;
			10308: out = 1387;
			10309: out = 2244;
			10310: out = 1717;
			10311: out = -367;
			10312: out = -3519;
			10313: out = -3304;
			10314: out = -631;
			10315: out = 2664;
			10316: out = -72;
			10317: out = -969;
			10318: out = -2250;
			10319: out = -3988;
			10320: out = -1346;
			10321: out = 2418;
			10322: out = 4771;
			10323: out = -34;
			10324: out = -3156;
			10325: out = -4039;
			10326: out = 977;
			10327: out = -279;
			10328: out = 372;
			10329: out = 386;
			10330: out = 2389;
			10331: out = 309;
			10332: out = -466;
			10333: out = 142;
			10334: out = 2021;
			10335: out = 737;
			10336: out = -1516;
			10337: out = -5258;
			10338: out = -609;
			10339: out = 3250;
			10340: out = 1764;
			10341: out = -1391;
			10342: out = -2055;
			10343: out = 741;
			10344: out = 948;
			10345: out = 788;
			10346: out = -193;
			10347: out = 1176;
			10348: out = -574;
			10349: out = -220;
			10350: out = 105;
			10351: out = -2053;
			10352: out = -4;
			10353: out = 1539;
			10354: out = -59;
			10355: out = -157;
			10356: out = -455;
			10357: out = 707;
			10358: out = -2425;
			10359: out = 1307;
			10360: out = 1853;
			10361: out = -737;
			10362: out = -2344;
			10363: out = -280;
			10364: out = 2942;
			10365: out = 1049;
			10366: out = 1163;
			10367: out = 304;
			10368: out = -619;
			10369: out = 929;
			10370: out = 1644;
			10371: out = 2007;
			10372: out = 977;
			10373: out = 613;
			10374: out = -1414;
			10375: out = -2847;
			10376: out = -4080;
			10377: out = 694;
			10378: out = 4631;
			10379: out = 1129;
			10380: out = -1675;
			10381: out = -3174;
			10382: out = -1684;
			10383: out = 1120;
			10384: out = 1168;
			10385: out = 103;
			10386: out = 164;
			10387: out = 2196;
			10388: out = 1439;
			10389: out = -2505;
			10390: out = -3370;
			10391: out = -907;
			10392: out = 2916;
			10393: out = 2769;
			10394: out = -99;
			10395: out = -3486;
			10396: out = -3448;
			10397: out = -619;
			10398: out = 1544;
			10399: out = 1491;
			10400: out = 2311;
			10401: out = 320;
			10402: out = -208;
			10403: out = -804;
			10404: out = 936;
			10405: out = -583;
			10406: out = -1624;
			10407: out = -1688;
			10408: out = 1578;
			10409: out = 1077;
			10410: out = -2943;
			10411: out = 213;
			10412: out = 822;
			10413: out = 595;
			10414: out = -4244;
			10415: out = -1128;
			10416: out = 1494;
			10417: out = 4007;
			10418: out = -1402;
			10419: out = 639;
			10420: out = 2428;
			10421: out = -9;
			10422: out = -375;
			10423: out = -45;
			10424: out = 1732;
			10425: out = -2993;
			10426: out = -1129;
			10427: out = 697;
			10428: out = -214;
			10429: out = 1912;
			10430: out = 2117;
			10431: out = 496;
			10432: out = -3898;
			10433: out = -4190;
			10434: out = -2037;
			10435: out = -1838;
			10436: out = 2657;
			10437: out = 1968;
			10438: out = -522;
			10439: out = -2480;
			10440: out = -718;
			10441: out = 634;
			10442: out = 403;
			10443: out = -1417;
			10444: out = 614;
			10445: out = 3684;
			10446: out = 659;
			10447: out = -2667;
			10448: out = -4203;
			10449: out = 6;
			10450: out = 688;
			10451: out = 2020;
			10452: out = 1918;
			10453: out = 1410;
			10454: out = 630;
			10455: out = -108;
			10456: out = -614;
			10457: out = -1526;
			10458: out = -829;
			10459: out = 131;
			10460: out = 984;
			10461: out = -788;
			10462: out = -1015;
			10463: out = 1072;
			10464: out = 2895;
			10465: out = 1435;
			10466: out = -1997;
			10467: out = -3210;
			10468: out = -1063;
			10469: out = 2555;
			10470: out = 3855;
			10471: out = 867;
			10472: out = -2197;
			10473: out = -2210;
			10474: out = 2565;
			10475: out = 3328;
			10476: out = 1600;
			10477: out = -2048;
			10478: out = -1522;
			10479: out = -1781;
			10480: out = -1151;
			10481: out = 673;
			10482: out = 1284;
			10483: out = 62;
			10484: out = -2747;
			10485: out = 937;
			10486: out = 645;
			10487: out = 342;
			10488: out = 4377;
			10489: out = 711;
			10490: out = -2241;
			10491: out = -4023;
			10492: out = -166;
			10493: out = 1173;
			10494: out = 1518;
			10495: out = -14;
			10496: out = 2292;
			10497: out = 1245;
			10498: out = -2529;
			10499: out = 1084;
			10500: out = 472;
			10501: out = -699;
			10502: out = -2633;
			10503: out = -1639;
			10504: out = -665;
			10505: out = 123;
			10506: out = 4791;
			10507: out = 3224;
			10508: out = -595;
			10509: out = -4515;
			10510: out = -2443;
			10511: out = 412;
			10512: out = 1418;
			10513: out = 1515;
			10514: out = -1405;
			10515: out = -3275;
			10516: out = -1843;
			10517: out = 30;
			10518: out = 1060;
			10519: out = 181;
			10520: out = 1840;
			10521: out = 435;
			10522: out = -1019;
			10523: out = -4355;
			10524: out = -570;
			10525: out = -665;
			10526: out = -2007;
			10527: out = -1636;
			10528: out = 1346;
			10529: out = 2703;
			10530: out = -7;
			10531: out = -1007;
			10532: out = -1006;
			10533: out = 757;
			10534: out = 9;
			10535: out = 1736;
			10536: out = 885;
			10537: out = -3769;
			10538: out = 32;
			10539: out = 333;
			10540: out = 0;
			10541: out = -122;
			10542: out = 2100;
			10543: out = 1695;
			10544: out = -2773;
			10545: out = -292;
			10546: out = 761;
			10547: out = 1045;
			10548: out = -1357;
			10549: out = -695;
			10550: out = 1241;
			10551: out = 2961;
			10552: out = 860;
			10553: out = -2486;
			10554: out = -3944;
			10555: out = 88;
			10556: out = 3222;
			10557: out = 3205;
			10558: out = -714;
			10559: out = -2708;
			10560: out = -3296;
			10561: out = -1398;
			10562: out = 2369;
			10563: out = 1236;
			10564: out = 551;
			10565: out = 1878;
			10566: out = 349;
			10567: out = 26;
			10568: out = 157;
			10569: out = 2378;
			10570: out = 1951;
			10571: out = -4;
			10572: out = -3730;
			10573: out = 127;
			10574: out = 351;
			10575: out = 229;
			10576: out = -115;
			10577: out = 1175;
			10578: out = 1276;
			10579: out = -40;
			10580: out = -72;
			10581: out = -595;
			10582: out = -507;
			10583: out = -111;
			10584: out = 287;
			10585: out = 185;
			10586: out = -194;
			10587: out = 1412;
			10588: out = 947;
			10589: out = -201;
			10590: out = -83;
			10591: out = -347;
			10592: out = 232;
			10593: out = 195;
			10594: out = 2082;
			10595: out = -422;
			10596: out = -2158;
			10597: out = -584;
			10598: out = 1265;
			10599: out = 1353;
			10600: out = -600;
			10601: out = 394;
			10602: out = 642;
			10603: out = 617;
			10604: out = -2940;
			10605: out = 209;
			10606: out = -173;
			10607: out = -2255;
			10608: out = -40;
			10609: out = -223;
			10610: out = -84;
			10611: out = 110;
			10612: out = 1116;
			10613: out = -16;
			10614: out = -2315;
			10615: out = -524;
			10616: out = -825;
			10617: out = 84;
			10618: out = 1976;
			10619: out = 1113;
			10620: out = 192;
			10621: out = -324;
			10622: out = -1646;
			10623: out = -355;
			10624: out = 375;
			10625: out = -285;
			10626: out = -318;
			10627: out = 712;
			10628: out = 1849;
			10629: out = -1092;
			10630: out = -1242;
			10631: out = -472;
			10632: out = 1748;
			10633: out = 441;
			10634: out = 273;
			10635: out = 109;
			10636: out = 406;
			10637: out = -673;
			10638: out = -1157;
			10639: out = -577;
			10640: out = -235;
			10641: out = 171;
			10642: out = 301;
			10643: out = -110;
			10644: out = 0;
			10645: out = -940;
			10646: out = -3594;
			10647: out = -63;
			10648: out = 520;
			10649: out = 173;
			10650: out = 21;
			10651: out = -392;
			10652: out = -454;
			10653: out = 618;
			10654: out = -1494;
			10655: out = 422;
			10656: out = 2460;
			10657: out = -388;
			10658: out = 168;
			10659: out = 702;
			10660: out = 2030;
			10661: out = -1641;
			10662: out = -1737;
			10663: out = -670;
			10664: out = 345;
			10665: out = 154;
			10666: out = -156;
			10667: out = -170;
			10668: out = -1428;
			10669: out = -411;
			10670: out = 1545;
			10671: out = 2856;
			10672: out = 2495;
			10673: out = 650;
			10674: out = -1297;
			10675: out = -1166;
			10676: out = -921;
			10677: out = -110;
			10678: out = 2837;
			10679: out = -241;
			10680: out = -998;
			10681: out = 591;
			10682: out = 2598;
			10683: out = 1661;
			10684: out = -655;
			10685: out = -418;
			10686: out = -2472;
			10687: out = -1637;
			10688: out = 179;
			10689: out = 2101;
			10690: out = 1435;
			10691: out = 199;
			10692: out = -764;
			10693: out = -72;
			10694: out = -324;
			10695: out = -1263;
			10696: out = -176;
			10697: out = 317;
			10698: out = 717;
			10699: out = 160;
			10700: out = -122;
			10701: out = -274;
			10702: out = 235;
			10703: out = -269;
			10704: out = 130;
			10705: out = -31;
			10706: out = -67;
			10707: out = -1095;
			10708: out = -657;
			10709: out = 332;
			10710: out = 1443;
			10711: out = 473;
			10712: out = -253;
			10713: out = 310;
			10714: out = -549;
			10715: out = -1221;
			10716: out = -1276;
			10717: out = 2146;
			10718: out = 333;
			10719: out = -2307;
			10720: out = -3141;
			10721: out = -3112;
			10722: out = -144;
			10723: out = 2163;
			10724: out = 2467;
			10725: out = -568;
			10726: out = -2005;
			10727: out = -389;
			10728: out = 1151;
			10729: out = 1337;
			10730: out = 452;
			10731: out = -661;
			10732: out = 32;
			10733: out = 203;
			10734: out = -63;
			10735: out = -1921;
			10736: out = -822;
			10737: out = 448;
			10738: out = 418;
			10739: out = -2509;
			10740: out = -1601;
			10741: out = 3870;
			10742: out = 1054;
			10743: out = -1420;
			10744: out = -4571;
			10745: out = -4569;
			10746: out = -1800;
			10747: out = 1783;
			10748: out = 2809;
			10749: out = 228;
			10750: out = -692;
			10751: out = 481;
			10752: out = -988;
			10753: out = 2453;
			10754: out = 2354;
			10755: out = 615;
			10756: out = -2214;
			10757: out = -564;
			10758: out = 1497;
			10759: out = 242;
			10760: out = 143;
			10761: out = 433;
			10762: out = 1719;
			10763: out = 1132;
			10764: out = 684;
			10765: out = -18;
			10766: out = -224;
			10767: out = -116;
			10768: out = -163;
			10769: out = -111;
			10770: out = 513;
			10771: out = 1532;
			10772: out = 1492;
			10773: out = 197;
			10774: out = -2113;
			10775: out = -826;
			10776: out = 2942;
			10777: out = -1172;
			10778: out = -652;
			10779: out = 6;
			10780: out = 1173;
			10781: out = 299;
			10782: out = 143;
			10783: out = 232;
			10784: out = -242;
			10785: out = -1066;
			10786: out = -1475;
			10787: out = 404;
			10788: out = -2522;
			10789: out = -1849;
			10790: out = 558;
			10791: out = -344;
			10792: out = -56;
			10793: out = 413;
			10794: out = 2419;
			10795: out = 326;
			10796: out = -454;
			10797: out = -644;
			10798: out = -89;
			10799: out = -433;
			10800: out = -532;
			10801: out = 471;
			10802: out = -863;
			10803: out = -682;
			10804: out = 296;
			10805: out = 1785;
			10806: out = 1060;
			10807: out = -456;
			10808: out = -1935;
			10809: out = -903;
			10810: out = -218;
			10811: out = -209;
			10812: out = -1825;
			10813: out = -506;
			10814: out = 963;
			10815: out = 954;
			10816: out = 332;
			10817: out = -1212;
			10818: out = -1599;
			10819: out = -328;
			10820: out = 2059;
			10821: out = 2591;
			10822: out = 436;
			10823: out = 106;
			10824: out = 31;
			10825: out = 813;
			10826: out = -1290;
			10827: out = 326;
			10828: out = 490;
			10829: out = -19;
			10830: out = -16;
			10831: out = 1160;
			10832: out = 1347;
			10833: out = -1862;
			10834: out = -2143;
			10835: out = -1213;
			10836: out = -39;
			10837: out = 400;
			10838: out = -945;
			10839: out = -1685;
			10840: out = -101;
			10841: out = 2020;
			10842: out = 1449;
			10843: out = -2325;
			10844: out = -1378;
			10845: out = -57;
			10846: out = 1776;
			10847: out = -952;
			10848: out = 1203;
			10849: out = 1234;
			10850: out = 724;
			10851: out = -971;
			10852: out = -109;
			10853: out = 838;
			10854: out = 289;
			10855: out = 30;
			10856: out = 7;
			10857: out = 228;
			10858: out = 703;
			10859: out = 431;
			10860: out = -36;
			10861: out = -1161;
			10862: out = 837;
			10863: out = 1239;
			10864: out = 17;
			10865: out = -1316;
			10866: out = -427;
			10867: out = 366;
			10868: out = -4142;
			10869: out = -596;
			10870: out = 341;
			10871: out = -139;
			10872: out = -1715;
			10873: out = -921;
			10874: out = 560;
			10875: out = 1505;
			10876: out = 648;
			10877: out = 391;
			10878: out = 1255;
			10879: out = -1040;
			10880: out = -196;
			10881: out = 616;
			10882: out = 1141;
			10883: out = 108;
			10884: out = -155;
			10885: out = 240;
			10886: out = 157;
			10887: out = -348;
			10888: out = -187;
			10889: out = 2421;
			10890: out = 886;
			10891: out = 365;
			10892: out = -291;
			10893: out = 1218;
			10894: out = -1397;
			10895: out = -3183;
			10896: out = -1676;
			10897: out = -117;
			10898: out = 1950;
			10899: out = 2612;
			10900: out = 319;
			10901: out = -185;
			10902: out = -45;
			10903: out = 58;
			10904: out = 84;
			10905: out = 595;
			10906: out = 1267;
			10907: out = -2613;
			10908: out = -1015;
			10909: out = 207;
			10910: out = 705;
			10911: out = -209;
			10912: out = 144;
			10913: out = 646;
			10914: out = 712;
			10915: out = -827;
			10916: out = -1864;
			10917: out = -1974;
			10918: out = 353;
			10919: out = 8;
			10920: out = -1175;
			10921: out = 196;
			10922: out = 843;
			10923: out = 593;
			10924: out = -1282;
			10925: out = -342;
			10926: out = -20;
			10927: out = 199;
			10928: out = 392;
			10929: out = -681;
			10930: out = -1142;
			10931: out = -1029;
			10932: out = 964;
			10933: out = 319;
			10934: out = -635;
			10935: out = 319;
			10936: out = 1477;
			10937: out = 1067;
			10938: out = -1402;
			10939: out = -1013;
			10940: out = -510;
			10941: out = 78;
			10942: out = -2087;
			10943: out = -675;
			10944: out = 417;
			10945: out = 1168;
			10946: out = 351;
			10947: out = -438;
			10948: out = -1393;
			10949: out = -2308;
			10950: out = -805;
			10951: out = 1396;
			10952: out = 3161;
			10953: out = -2293;
			10954: out = -1985;
			10955: out = 476;
			10956: out = 2492;
			10957: out = 2278;
			10958: out = 1097;
			10959: out = 99;
			10960: out = -294;
			10961: out = 311;
			10962: out = 688;
			10963: out = 67;
			10964: out = -398;
			10965: out = -984;
			10966: out = -1065;
			10967: out = -1998;
			10968: out = -26;
			10969: out = 2355;
			10970: out = 3313;
			10971: out = 1889;
			10972: out = -669;
			10973: out = -2413;
			10974: out = 87;
			10975: out = 332;
			10976: out = -169;
			10977: out = -606;
			10978: out = -96;
			10979: out = 1349;
			10980: out = 2372;
			10981: out = 314;
			10982: out = 75;
			10983: out = -253;
			10984: out = -1794;
			10985: out = 70;
			10986: out = -344;
			10987: out = -1089;
			10988: out = -229;
			10989: out = 701;
			10990: out = 865;
			10991: out = 232;
			10992: out = -1304;
			10993: out = -701;
			10994: out = 1152;
			10995: out = 2591;
			10996: out = 1288;
			10997: out = -1365;
			10998: out = -4362;
			10999: out = -486;
			11000: out = 18;
			11001: out = -1295;
			11002: out = 135;
			11003: out = -352;
			11004: out = 259;
			11005: out = 1014;
			11006: out = -194;
			11007: out = -1988;
			11008: out = -3024;
			11009: out = 350;
			11010: out = -122;
			11011: out = 56;
			11012: out = 208;
			11013: out = 2672;
			11014: out = 1519;
			11015: out = -709;
			11016: out = -2731;
			11017: out = -11;
			11018: out = 1797;
			11019: out = 204;
			11020: out = -1143;
			11021: out = -2789;
			11022: out = -1722;
			11023: out = 2354;
			11024: out = 2465;
			11025: out = -186;
			11026: out = -4270;
			11027: out = 173;
			11028: out = 1433;
			11029: out = 1151;
			11030: out = -540;
			11031: out = 262;
			11032: out = 1206;
			11033: out = 1282;
			11034: out = 535;
			11035: out = -1291;
			11036: out = -2192;
			11037: out = -49;
			11038: out = -140;
			11039: out = 297;
			11040: out = 774;
			11041: out = 1107;
			11042: out = 292;
			11043: out = -1158;
			11044: out = -2166;
			11045: out = -2110;
			11046: out = -1327;
			11047: out = -679;
			11048: out = 3880;
			11049: out = 2675;
			11050: out = 338;
			11051: out = -921;
			11052: out = 198;
			11053: out = 676;
			11054: out = -216;
			11055: out = 1174;
			11056: out = 341;
			11057: out = -797;
			11058: out = -2863;
			11059: out = -118;
			11060: out = 1077;
			11061: out = 591;
			11062: out = 2326;
			11063: out = 263;
			11064: out = -1454;
			11065: out = -1335;
			11066: out = -427;
			11067: out = 81;
			11068: out = -262;
			11069: out = 436;
			11070: out = -259;
			11071: out = -497;
			11072: out = 275;
			11073: out = 118;
			11074: out = 235;
			11075: out = 269;
			11076: out = 1818;
			11077: out = 715;
			11078: out = -920;
			11079: out = -2877;
			11080: out = -1734;
			11081: out = -632;
			11082: out = 670;
			11083: out = 109;
			11084: out = 1917;
			11085: out = 2356;
			11086: out = 1721;
			11087: out = -2038;
			11088: out = -2384;
			11089: out = -398;
			11090: out = 1619;
			11091: out = 1215;
			11092: out = 310;
			11093: out = -254;
			11094: out = 1569;
			11095: out = 258;
			11096: out = -2529;
			11097: out = -2578;
			11098: out = -1387;
			11099: out = 574;
			11100: out = 471;
			11101: out = 1042;
			11102: out = -299;
			11103: out = -704;
			11104: out = 1369;
			11105: out = 1116;
			11106: out = 106;
			11107: out = -483;
			11108: out = -429;
			11109: out = 1766;
			11110: out = 3203;
			11111: out = 10;
			11112: out = -940;
			11113: out = -1768;
			11114: out = -1294;
			11115: out = -241;
			11116: out = 309;
			11117: out = -336;
			11118: out = 472;
			11119: out = -1875;
			11120: out = -1435;
			11121: out = 990;
			11122: out = 1987;
			11123: out = 1046;
			11124: out = -721;
			11125: out = -913;
			11126: out = -461;
			11127: out = -206;
			11128: out = -1117;
			11129: out = 1330;
			11130: out = 1088;
			11131: out = -43;
			11132: out = -3822;
			11133: out = -881;
			11134: out = 623;
			11135: out = 188;
			11136: out = 92;
			11137: out = 47;
			11138: out = 487;
			11139: out = 39;
			11140: out = 269;
			11141: out = -1412;
			11142: out = -3614;
			11143: out = -47;
			11144: out = 1110;
			11145: out = 1337;
			11146: out = -172;
			11147: out = 1548;
			11148: out = 940;
			11149: out = -1504;
			11150: out = -2357;
			11151: out = -2305;
			11152: out = -154;
			11153: out = 2068;
			11154: out = 2260;
			11155: out = 773;
			11156: out = -63;
			11157: out = -514;
			11158: out = 2208;
			11159: out = 3238;
			11160: out = 2010;
			11161: out = -2928;
			11162: out = -3490;
			11163: out = -270;
			11164: out = 708;
			11165: out = 607;
			11166: out = 98;
			11167: out = 2381;
			11168: out = -2205;
			11169: out = -3943;
			11170: out = -3477;
			11171: out = 833;
			11172: out = 2079;
			11173: out = 1545;
			11174: out = -704;
			11175: out = -193;
			11176: out = -311;
			11177: out = -527;
			11178: out = 870;
			11179: out = 122;
			11180: out = 379;
			11181: out = 1486;
			11182: out = 1832;
			11183: out = 981;
			11184: out = 5;
			11185: out = -314;
			11186: out = 235;
			11187: out = -274;
			11188: out = -1395;
			11189: out = -1446;
			11190: out = 1498;
			11191: out = 4101;
			11192: out = 2003;
			11193: out = -1917;
			11194: out = -5047;
			11195: out = -3464;
			11196: out = -2029;
			11197: out = 1601;
			11198: out = 2945;
			11199: out = 1574;
			11200: out = -353;
			11201: out = -1151;
			11202: out = -974;
			11203: out = 107;
			11204: out = -568;
			11205: out = -1223;
			11206: out = 1250;
			11207: out = -73;
			11208: out = -972;
			11209: out = -1310;
			11210: out = -175;
			11211: out = -343;
			11212: out = -919;
			11213: out = 1089;
			11214: out = 159;
			11215: out = 1712;
			11216: out = 3622;
			11217: out = 2281;
			11218: out = -1550;
			11219: out = -4103;
			11220: out = -319;
			11221: out = -311;
			11222: out = 88;
			11223: out = -3;
			11224: out = 1333;
			11225: out = 901;
			11226: out = -136;
			11227: out = 471;
			11228: out = -2938;
			11229: out = -2227;
			11230: out = 1039;
			11231: out = -2072;
			11232: out = -1902;
			11233: out = -204;
			11234: out = 3178;
			11235: out = 3520;
			11236: out = 2472;
			11237: out = 644;
			11238: out = -2083;
			11239: out = -1677;
			11240: out = -624;
			11241: out = 476;
			11242: out = -1247;
			11243: out = 129;
			11244: out = 2598;
			11245: out = 501;
			11246: out = -1842;
			11247: out = -2445;
			11248: out = 2240;
			11249: out = 417;
			11250: out = -271;
			11251: out = -956;
			11252: out = 743;
			11253: out = 461;
			11254: out = -208;
			11255: out = -1375;
			11256: out = -750;
			11257: out = -198;
			11258: out = 235;
			11259: out = 3094;
			11260: out = 408;
			11261: out = -2132;
			11262: out = -2450;
			11263: out = -1054;
			11264: out = -102;
			11265: out = -129;
			11266: out = 319;
			11267: out = 630;
			11268: out = 263;
			11269: out = -1877;
			11270: out = -4;
			11271: out = 739;
			11272: out = 1163;
			11273: out = 207;
			11274: out = 359;
			11275: out = -204;
			11276: out = -1312;
			11277: out = -423;
			11278: out = 1049;
			11279: out = 2038;
			11280: out = -550;
			11281: out = -338;
			11282: out = 756;
			11283: out = 3539;
			11284: out = -1528;
			11285: out = -1892;
			11286: out = -379;
			11287: out = 2051;
			11288: out = 898;
			11289: out = 434;
			11290: out = 1402;
			11291: out = -612;
			11292: out = -1810;
			11293: out = -1752;
			11294: out = 903;
			11295: out = 2503;
			11296: out = 2290;
			11297: out = -171;
			11298: out = -2845;
			11299: out = -3361;
			11300: out = -1409;
			11301: out = -523;
			11302: out = 2365;
			11303: out = 2440;
			11304: out = 376;
			11305: out = 132;
			11306: out = -283;
			11307: out = -134;
			11308: out = -323;
			11309: out = 980;
			11310: out = 993;
			11311: out = -255;
			11312: out = 918;
			11313: out = 973;
			11314: out = 659;
			11315: out = -1130;
			11316: out = -555;
			11317: out = 470;
			11318: out = 1988;
			11319: out = -2384;
			11320: out = -2014;
			11321: out = -656;
			11322: out = -123;
			11323: out = -212;
			11324: out = 315;
			11325: out = 1395;
			11326: out = 386;
			11327: out = -660;
			11328: out = -1404;
			11329: out = 86;
			11330: out = -88;
			11331: out = 1007;
			11332: out = 2337;
			11333: out = 348;
			11334: out = -77;
			11335: out = -528;
			11336: out = -615;
			11337: out = -2056;
			11338: out = -1689;
			11339: out = 102;
			11340: out = 1151;
			11341: out = 663;
			11342: out = -460;
			11343: out = -74;
			11344: out = -1668;
			11345: out = -1444;
			11346: out = -454;
			11347: out = -278;
			11348: out = 5;
			11349: out = 476;
			11350: out = 1414;
			11351: out = 193;
			11352: out = -1019;
			11353: out = -1848;
			11354: out = -631;
			11355: out = -267;
			11356: out = 206;
			11357: out = 668;
			11358: out = 342;
			11359: out = 100;
			11360: out = 4;
			11361: out = -2664;
			11362: out = -1150;
			11363: out = 998;
			11364: out = 3087;
			11365: out = 434;
			11366: out = -605;
			11367: out = -513;
			11368: out = -220;
			11369: out = -715;
			11370: out = -875;
			11371: out = -83;
			11372: out = 291;
			11373: out = -330;
			11374: out = -1470;
			11375: out = 138;
			11376: out = -189;
			11377: out = 679;
			11378: out = 2072;
			11379: out = -675;
			11380: out = -2298;
			11381: out = -2159;
			11382: out = 205;
			11383: out = 1972;
			11384: out = 1920;
			11385: out = -288;
			11386: out = 1652;
			11387: out = 1274;
			11388: out = 166;
			11389: out = -2221;
			11390: out = -1243;
			11391: out = 16;
			11392: out = 704;
			11393: out = 361;
			11394: out = 674;
			11395: out = 695;
			11396: out = -2372;
			11397: out = -1558;
			11398: out = -1281;
			11399: out = -672;
			11400: out = -18;
			11401: out = 2192;
			11402: out = 3008;
			11403: out = 282;
			11404: out = -1831;
			11405: out = -2335;
			11406: out = -2;
			11407: out = 578;
			11408: out = 1954;
			11409: out = 1730;
			11410: out = 1190;
			11411: out = -1218;
			11412: out = -1582;
			11413: out = -368;
			11414: out = 178;
			11415: out = 369;
			11416: out = 266;
			11417: out = 183;
			11418: out = 536;
			11419: out = 812;
			11420: out = 883;
			11421: out = -1305;
			11422: out = -718;
			11423: out = -80;
			11424: out = -1105;
			11425: out = -253;
			11426: out = 389;
			11427: out = 1072;
			11428: out = 181;
			11429: out = -49;
			11430: out = -448;
			11431: out = -991;
			11432: out = -293;
			11433: out = 133;
			11434: out = 158;
			11435: out = -35;
			11436: out = 746;
			11437: out = 1446;
			11438: out = 390;
			11439: out = 201;
			11440: out = -972;
			11441: out = -1356;
			11442: out = -3245;
			11443: out = 784;
			11444: out = 3338;
			11445: out = 1638;
			11446: out = 1396;
			11447: out = 406;
			11448: out = -167;
			11449: out = -3020;
			11450: out = -2357;
			11451: out = -1074;
			11452: out = 452;
			11453: out = 1433;
			11454: out = 1860;
			11455: out = 1260;
			11456: out = -835;
			11457: out = -1913;
			11458: out = -1729;
			11459: out = 207;
			11460: out = -249;
			11461: out = 742;
			11462: out = 1181;
			11463: out = -498;
			11464: out = -450;
			11465: out = -17;
			11466: out = -336;
			11467: out = 1382;
			11468: out = 16;
			11469: out = -1459;
			11470: out = -1059;
			11471: out = 1590;
			11472: out = 1732;
			11473: out = -2335;
			11474: out = -1868;
			11475: out = -1331;
			11476: out = 719;
			11477: out = -1479;
			11478: out = 3219;
			11479: out = 3276;
			11480: out = -677;
			11481: out = -3626;
			11482: out = -3186;
			11483: out = 115;
			11484: out = -207;
			11485: out = 3010;
			11486: out = 1640;
			11487: out = -1957;
			11488: out = -1469;
			11489: out = 358;
			11490: out = 1776;
			11491: out = 224;
			11492: out = -1009;
			11493: out = -2103;
			11494: out = -1840;
			11495: out = -98;
			11496: out = 736;
			11497: out = 649;
			11498: out = 441;
			11499: out = 303;
			11500: out = 5;
			11501: out = -540;
			11502: out = 212;
			11503: out = 238;
			11504: out = 403;
			11505: out = 1101;
			11506: out = 1031;
			11507: out = 950;
			11508: out = 572;
			11509: out = 1426;
			11510: out = -157;
			11511: out = -1540;
			11512: out = -393;
			11513: out = -319;
			11514: out = 195;
			11515: out = 371;
			11516: out = 2520;
			11517: out = 1189;
			11518: out = -1203;
			11519: out = -3849;
			11520: out = -2762;
			11521: out = -1129;
			11522: out = 189;
			11523: out = 1018;
			11524: out = 675;
			11525: out = -211;
			11526: out = -1306;
			11527: out = -139;
			11528: out = 472;
			11529: out = 268;
			11530: out = 498;
			11531: out = -469;
			11532: out = -731;
			11533: out = 353;
			11534: out = 1111;
			11535: out = 1668;
			11536: out = 1479;
			11537: out = 323;
			11538: out = -624;
			11539: out = -962;
			11540: out = -474;
			11541: out = 659;
			11542: out = 1191;
			11543: out = 832;
			11544: out = 1124;
			11545: out = -352;
			11546: out = -1158;
			11547: out = -932;
			11548: out = 340;
			11549: out = 592;
			11550: out = 131;
			11551: out = 215;
			11552: out = -69;
			11553: out = -23;
			11554: out = 116;
			11555: out = 141;
			11556: out = -51;
			11557: out = -248;
			11558: out = 302;
			11559: out = 120;
			11560: out = 203;
			11561: out = 159;
			11562: out = -26;
			11563: out = -1295;
			11564: out = -2017;
			11565: out = 169;
			11566: out = 954;
			11567: out = 1340;
			11568: out = 739;
			11569: out = -943;
			11570: out = -1483;
			11571: out = -597;
			11572: out = -469;
			11573: out = 901;
			11574: out = 111;
			11575: out = -1779;
			11576: out = -204;
			11577: out = 1609;
			11578: out = 2182;
			11579: out = -1048;
			11580: out = -1877;
			11581: out = -1611;
			11582: out = 555;
			11583: out = -121;
			11584: out = 1337;
			11585: out = 1738;
			11586: out = 122;
			11587: out = -176;
			11588: out = -337;
			11589: out = -700;
			11590: out = -485;
			11591: out = -934;
			11592: out = -681;
			11593: out = 87;
			11594: out = 1183;
			11595: out = 819;
			11596: out = -67;
			11597: out = 1028;
			11598: out = 2380;
			11599: out = 1571;
			11600: out = -4599;
			11601: out = -2861;
			11602: out = -834;
			11603: out = 1304;
			11604: out = 1858;
			11605: out = 1129;
			11606: out = -128;
			11607: out = -77;
			11608: out = -267;
			11609: out = -285;
			11610: out = -1047;
			11611: out = 1679;
			11612: out = 683;
			11613: out = -279;
			11614: out = -2029;
			11615: out = 1375;
			11616: out = 527;
			11617: out = -2630;
			11618: out = -865;
			11619: out = -180;
			11620: out = 1165;
			11621: out = 1463;
			11622: out = 722;
			11623: out = -484;
			11624: out = -942;
			11625: out = -733;
			11626: out = 219;
			11627: out = 611;
			11628: out = 188;
			11629: out = 300;
			11630: out = 7;
			11631: out = -199;
			11632: out = 569;
			11633: out = 433;
			11634: out = -480;
			11635: out = -2726;
			11636: out = 89;
			11637: out = 668;
			11638: out = 209;
			11639: out = 1409;
			11640: out = 251;
			11641: out = -355;
			11642: out = -65;
			11643: out = -159;
			11644: out = -312;
			11645: out = -630;
			11646: out = 356;
			11647: out = -185;
			11648: out = 277;
			11649: out = 1626;
			11650: out = 517;
			11651: out = -1179;
			11652: out = -2648;
			11653: out = -72;
			11654: out = -390;
			11655: out = 4;
			11656: out = -239;
			11657: out = 1411;
			11658: out = -607;
			11659: out = -2778;
			11660: out = -1191;
			11661: out = -520;
			11662: out = 291;
			11663: out = 362;
			11664: out = 2632;
			11665: out = 1935;
			11666: out = 62;
			11667: out = 498;
			11668: out = -2367;
			11669: out = -2131;
			11670: out = 195;
			11671: out = 888;
			11672: out = 240;
			11673: out = -633;
			11674: out = -208;
			11675: out = 989;
			11676: out = 689;
			11677: out = -1205;
			11678: out = -898;
			11679: out = -410;
			11680: out = 458;
			11681: out = 1014;
			11682: out = -186;
			11683: out = -272;
			11684: out = 756;
			11685: out = 325;
			11686: out = -773;
			11687: out = -1841;
			11688: out = -779;
			11689: out = -72;
			11690: out = 355;
			11691: out = -222;
			11692: out = 1339;
			11693: out = 740;
			11694: out = -730;
			11695: out = -4334;
			11696: out = -275;
			11697: out = 1831;
			11698: out = 1318;
			11699: out = 728;
			11700: out = -1090;
			11701: out = -1357;
			11702: out = -26;
			11703: out = 683;
			11704: out = -353;
			11705: out = -2154;
			11706: out = -17;
			11707: out = 267;
			11708: out = 340;
			11709: out = -118;
			11710: out = -637;
			11711: out = -739;
			11712: out = -164;
			11713: out = 1282;
			11714: out = 908;
			11715: out = 14;
			11716: out = -351;
			11717: out = -30;
			11718: out = 980;
			11719: out = 1606;
			11720: out = 383;
			11721: out = -182;
			11722: out = -542;
			11723: out = -20;
			11724: out = -285;
			11725: out = 331;
			11726: out = 579;
			11727: out = 84;
			11728: out = -635;
			11729: out = -859;
			11730: out = -890;
			11731: out = 808;
			11732: out = 709;
			11733: out = 229;
			11734: out = 590;
			11735: out = 1173;
			11736: out = 1030;
			11737: out = 636;
			11738: out = -2810;
			11739: out = -1403;
			11740: out = 1892;
			11741: out = 684;
			11742: out = 512;
			11743: out = -483;
			11744: out = -336;
			11745: out = -149;
			11746: out = 613;
			11747: out = 414;
			11748: out = 470;
			11749: out = -1163;
			11750: out = -1309;
			11751: out = 121;
			11752: out = 136;
			11753: out = -439;
			11754: out = -1211;
			11755: out = 1213;
			11756: out = 95;
			11757: out = 333;
			11758: out = 907;
			11759: out = 1427;
			11760: out = -250;
			11761: out = -1747;
			11762: out = -510;
			11763: out = 1128;
			11764: out = 1966;
			11765: out = 868;
			11766: out = -1107;
			11767: out = -2461;
			11768: out = -1688;
			11769: out = 1876;
			11770: out = 1105;
			11771: out = 78;
			11772: out = -540;
			11773: out = 58;
			11774: out = -169;
			11775: out = -488;
			11776: out = 724;
			11777: out = 27;
			11778: out = -92;
			11779: out = -241;
			11780: out = 309;
			11781: out = -343;
			11782: out = -1107;
			11783: out = -1234;
			11784: out = -1266;
			11785: out = -1220;
			11786: out = -1090;
			11787: out = -297;
			11788: out = 1066;
			11789: out = 2029;
			11790: out = 781;
			11791: out = 126;
			11792: out = -1548;
			11793: out = -2220;
			11794: out = -675;
			11795: out = 2465;
			11796: out = 3285;
			11797: out = -1643;
			11798: out = -249;
			11799: out = -48;
			11800: out = -49;
			11801: out = -114;
			11802: out = 130;
			11803: out = -115;
			11804: out = -1356;
			11805: out = 424;
			11806: out = 1434;
			11807: out = 1333;
			11808: out = -1031;
			11809: out = -1772;
			11810: out = -1077;
			11811: out = 1097;
			11812: out = 425;
			11813: out = 232;
			11814: out = 303;
			11815: out = 2209;
			11816: out = 403;
			11817: out = -1439;
			11818: out = -702;
			11819: out = -2443;
			11820: out = -1685;
			11821: out = -226;
			11822: out = 632;
			11823: out = 225;
			11824: out = -143;
			11825: out = 428;
			11826: out = -381;
			11827: out = -559;
			11828: out = -362;
			11829: out = 664;
			11830: out = 372;
			11831: out = 545;
			11832: out = 2094;
			11833: out = -1496;
			11834: out = -1806;
			11835: out = -497;
			11836: out = 197;
			11837: out = 422;
			11838: out = 442;
			11839: out = 1089;
			11840: out = 226;
			11841: out = 203;
			11842: out = -99;
			11843: out = -1610;
			11844: out = -628;
			11845: out = 1316;
			11846: out = 3037;
			11847: out = 1060;
			11848: out = -179;
			11849: out = -597;
			11850: out = -671;
			11851: out = -52;
			11852: out = 136;
			11853: out = 352;
			11854: out = -27;
			11855: out = 1105;
			11856: out = 1725;
			11857: out = 562;
			11858: out = -1136;
			11859: out = -1417;
			11860: out = 359;
			11861: out = -27;
			11862: out = -345;
			11863: out = -1079;
			11864: out = 327;
			11865: out = -280;
			11866: out = 774;
			11867: out = 2175;
			11868: out = 1340;
			11869: out = 144;
			11870: out = -873;
			11871: out = -619;
			11872: out = -670;
			11873: out = -998;
			11874: out = -1782;
			11875: out = -38;
			11876: out = 902;
			11877: out = 1475;
			11878: out = -436;
			11879: out = 338;
			11880: out = -850;
			11881: out = -1561;
			11882: out = -1410;
			11883: out = 2210;
			11884: out = 3630;
			11885: out = -104;
			11886: out = -1864;
			11887: out = -1963;
			11888: out = 689;
			11889: out = 486;
			11890: out = 1202;
			11891: out = 343;
			11892: out = -104;
			11893: out = -1676;
			11894: out = -913;
			11895: out = 339;
			11896: out = -117;
			11897: out = 45;
			11898: out = 119;
			11899: out = -1195;
			11900: out = 293;
			11901: out = -1077;
			11902: out = -2754;
			11903: out = -218;
			11904: out = 1281;
			11905: out = 1380;
			11906: out = -1131;
			11907: out = -856;
			11908: out = -436;
			11909: out = 428;
			11910: out = -121;
			11911: out = -253;
			11912: out = -548;
			11913: out = -112;
			11914: out = -1653;
			11915: out = -2281;
			11916: out = -2056;
			11917: out = -164;
			11918: out = 907;
			11919: out = 1684;
			11920: out = 1849;
			11921: out = 72;
			11922: out = -1363;
			11923: out = -1716;
			11924: out = 210;
			11925: out = 782;
			11926: out = 1304;
			11927: out = 1575;
			11928: out = 1121;
			11929: out = 464;
			11930: out = -442;
			11931: out = -2733;
			11932: out = -1319;
			11933: out = -24;
			11934: out = -90;
			11935: out = 1045;
			11936: out = 117;
			11937: out = -557;
			11938: out = 2937;
			11939: out = 268;
			11940: out = -1333;
			11941: out = -938;
			11942: out = 1041;
			11943: out = 2208;
			11944: out = 1621;
			11945: out = -421;
			11946: out = -990;
			11947: out = -473;
			11948: out = 280;
			11949: out = 205;
			11950: out = 79;
			11951: out = -5;
			11952: out = -1844;
			11953: out = 376;
			11954: out = 288;
			11955: out = -1867;
			11956: out = -862;
			11957: out = -253;
			11958: out = 500;
			11959: out = 226;
			11960: out = 371;
			11961: out = 279;
			11962: out = 331;
			11963: out = 184;
			11964: out = 57;
			11965: out = 51;
			11966: out = 625;
			11967: out = -126;
			11968: out = -1296;
			11969: out = -2318;
			11970: out = -42;
			11971: out = 927;
			11972: out = 1302;
			11973: out = 890;
			11974: out = 766;
			11975: out = 53;
			11976: out = -952;
			11977: out = 948;
			11978: out = -116;
			11979: out = -896;
			11980: out = 427;
			11981: out = 677;
			11982: out = 805;
			11983: out = -124;
			11984: out = 331;
			11985: out = -681;
			11986: out = -735;
			11987: out = -261;
			11988: out = 1955;
			11989: out = 1697;
			11990: out = -202;
			11991: out = -735;
			11992: out = -1143;
			11993: out = -690;
			11994: out = -236;
			11995: out = 949;
			11996: out = 1200;
			11997: out = 601;
			11998: out = -425;
			11999: out = -998;
			12000: out = -660;
			12001: out = -133;
			12002: out = 1288;
			12003: out = 997;
			12004: out = -74;
			12005: out = -1272;
			12006: out = -682;
			12007: out = -373;
			12008: out = -1373;
			12009: out = -130;
			12010: out = 616;
			12011: out = 594;
			12012: out = -1464;
			12013: out = -2821;
			12014: out = -2281;
			12015: out = 1058;
			12016: out = 1793;
			12017: out = 1784;
			12018: out = 235;
			12019: out = 1943;
			12020: out = -1495;
			12021: out = -3149;
			12022: out = -3006;
			12023: out = 1679;
			12024: out = 2101;
			12025: out = 496;
			12026: out = 94;
			12027: out = 720;
			12028: out = 881;
			12029: out = -1260;
			12030: out = 396;
			12031: out = -294;
			12032: out = -348;
			12033: out = -42;
			12034: out = 2276;
			12035: out = 2160;
			12036: out = -675;
			12037: out = -353;
			12038: out = -959;
			12039: out = -875;
			12040: out = -1433;
			12041: out = 364;
			12042: out = 950;
			12043: out = 370;
			12044: out = -2036;
			12045: out = -2232;
			12046: out = -1248;
			12047: out = -968;
			12048: out = 569;
			12049: out = 1118;
			12050: out = 797;
			12051: out = -562;
			12052: out = -1207;
			12053: out = -898;
			12054: out = -42;
			12055: out = 817;
			12056: out = 696;
			12057: out = -139;
			12058: out = -426;
			12059: out = 393;
			12060: out = 1581;
			12061: out = 1012;
			12062: out = 599;
			12063: out = -1899;
			12064: out = -4356;
			12065: out = -414;
			12066: out = 1286;
			12067: out = 2032;
			12068: out = 1836;
			12069: out = 638;
			12070: out = -155;
			12071: out = -132;
			12072: out = -592;
			12073: out = -208;
			12074: out = -43;
			12075: out = -161;
			12076: out = 174;
			12077: out = 208;
			12078: out = -115;
			12079: out = 221;
			12080: out = 108;
			12081: out = -123;
			12082: out = -1816;
			12083: out = 92;
			12084: out = -17;
			12085: out = -432;
			12086: out = -172;
			12087: out = 913;
			12088: out = 1006;
			12089: out = 175;
			12090: out = -831;
			12091: out = -190;
			12092: out = 694;
			12093: out = 1389;
			12094: out = -705;
			12095: out = -1160;
			12096: out = 1051;
			12097: out = 467;
			12098: out = -1766;
			12099: out = -3884;
			12100: out = -85;
			12101: out = 2022;
			12102: out = 2516;
			12103: out = -647;
			12104: out = -737;
			12105: out = -1847;
			12106: out = -1538;
			12107: out = 56;
			12108: out = 896;
			12109: out = 732;
			12110: out = -58;
			12111: out = 1161;
			12112: out = 528;
			12113: out = -483;
			12114: out = 2049;
			12115: out = 161;
			12116: out = -784;
			12117: out = -779;
			12118: out = 1205;
			12119: out = 1069;
			12120: out = -229;
			12121: out = 2;
			12122: out = -687;
			12123: out = 40;
			12124: out = 924;
			12125: out = 2305;
			12126: out = 1043;
			12127: out = -579;
			12128: out = -156;
			12129: out = -336;
			12130: out = -245;
			12131: out = -241;
			12132: out = 119;
			12133: out = 284;
			12134: out = -276;
			12135: out = -2403;
			12136: out = -1538;
			12137: out = 150;
			12138: out = 1524;
			12139: out = 1050;
			12140: out = -459;
			12141: out = -2401;
			12142: out = -4809;
			12143: out = -1447;
			12144: out = 1101;
			12145: out = 1461;
			12146: out = 1471;
			12147: out = 469;
			12148: out = -310;
			12149: out = -1222;
			12150: out = -70;
			12151: out = 231;
			12152: out = -650;
			12153: out = 824;
			12154: out = -715;
			12155: out = -1297;
			12156: out = 483;
			12157: out = 817;
			12158: out = 770;
			12159: out = -8;
			12160: out = -1385;
			12161: out = -513;
			12162: out = 429;
			12163: out = -986;
			12164: out = 170;
			12165: out = 251;
			12166: out = 448;
			12167: out = -82;
			12168: out = 478;
			12169: out = 786;
			12170: out = 1677;
			12171: out = -1848;
			12172: out = -1916;
			12173: out = 321;
			12174: out = -1055;
			12175: out = 831;
			12176: out = 1573;
			12177: out = 843;
			12178: out = -636;
			12179: out = -1282;
			12180: out = -406;
			12181: out = -86;
			12182: out = 2283;
			12183: out = 2706;
			12184: out = 333;
			12185: out = 345;
			12186: out = -246;
			12187: out = -562;
			12188: out = -489;
			12189: out = -225;
			12190: out = 912;
			12191: out = 2523;
			12192: out = 1550;
			12193: out = -835;
			12194: out = -3192;
			12195: out = -4;
			12196: out = 282;
			12197: out = -96;
			12198: out = -3428;
			12199: out = 2086;
			12200: out = 1016;
			12201: out = -1493;
			12202: out = 77;
			12203: out = 43;
			12204: out = 143;
			12205: out = -22;
			12206: out = 350;
			12207: out = 1607;
			12208: out = 2415;
			12209: out = 862;
			12210: out = -1515;
			12211: out = -2651;
			12212: out = -429;
			12213: out = -1289;
			12214: out = 894;
			12215: out = 2143;
			12216: out = -119;
			12217: out = -409;
			12218: out = -464;
			12219: out = -24;
			12220: out = -253;
			12221: out = 53;
			12222: out = 215;
			12223: out = 284;
			12224: out = -1034;
			12225: out = -1341;
			12226: out = 252;
			12227: out = -101;
			12228: out = 714;
			12229: out = 637;
			12230: out = 433;
			12231: out = -2438;
			12232: out = -3153;
			12233: out = -1022;
			12234: out = 430;
			12235: out = 1566;
			12236: out = 1124;
			12237: out = -38;
			12238: out = -255;
			12239: out = -156;
			12240: out = -621;
			12241: out = 389;
			12242: out = -252;
			12243: out = -172;
			12244: out = 1148;
			12245: out = 1204;
			12246: out = -432;
			12247: out = -2895;
			12248: out = -2014;
			12249: out = -779;
			12250: out = 532;
			12251: out = 209;
			12252: out = 416;
			12253: out = 373;
			12254: out = 616;
			12255: out = -1061;
			12256: out = -1038;
			12257: out = -455;
			12258: out = 726;
			12259: out = 863;
			12260: out = 921;
			12261: out = 510;
			12262: out = 1379;
			12263: out = -446;
			12264: out = -1512;
			12265: out = 405;
			12266: out = -210;
			12267: out = -447;
			12268: out = -1182;
			12269: out = 2276;
			12270: out = -556;
			12271: out = -2201;
			12272: out = 704;
			12273: out = -267;
			12274: out = 144;
			12275: out = 162;
			12276: out = 1073;
			12277: out = 173;
			12278: out = -124;
			12279: out = -84;
			12280: out = 1111;
			12281: out = 403;
			12282: out = -1193;
			12283: out = -1841;
			12284: out = -717;
			12285: out = 570;
			12286: out = 140;
			12287: out = 1274;
			12288: out = 612;
			12289: out = -82;
			12290: out = 629;
			12291: out = -439;
			12292: out = -2025;
			12293: out = -3314;
			12294: out = -819;
			12295: out = 1164;
			12296: out = 1776;
			12297: out = 1080;
			12298: out = 121;
			12299: out = 222;
			12300: out = 1309;
			12301: out = 983;
			12302: out = 216;
			12303: out = -591;
			12304: out = 213;
			12305: out = 101;
			12306: out = 72;
			12307: out = -258;
			12308: out = -454;
			12309: out = -186;
			12310: out = 367;
			12311: out = -312;
			12312: out = 681;
			12313: out = 520;
			12314: out = -584;
			12315: out = 1614;
			12316: out = 572;
			12317: out = -1293;
			12318: out = 183;
			12319: out = -2138;
			12320: out = -708;
			12321: out = 2954;
			12322: out = 1966;
			12323: out = 1316;
			12324: out = -140;
			12325: out = -1954;
			12326: out = -1333;
			12327: out = -444;
			12328: out = 168;
			12329: out = 69;
			12330: out = 391;
			12331: out = 452;
			12332: out = 288;
			12333: out = -1271;
			12334: out = -465;
			12335: out = 2337;
			12336: out = -190;
			12337: out = -422;
			12338: out = -972;
			12339: out = 529;
			12340: out = -1217;
			12341: out = -321;
			12342: out = 823;
			12343: out = 356;
			12344: out = -1617;
			12345: out = -2545;
			12346: out = -1450;
			12347: out = 1134;
			12348: out = 1328;
			12349: out = -339;
			12350: out = 5;
			12351: out = 18;
			12352: out = 426;
			12353: out = 575;
			12354: out = -276;
			12355: out = -270;
			12356: out = 472;
			12357: out = 1416;
			12358: out = 490;
			12359: out = -223;
			12360: out = 644;
			12361: out = 249;
			12362: out = -1158;
			12363: out = -3193;
			12364: out = -718;
			12365: out = -377;
			12366: out = 861;
			12367: out = 1620;
			12368: out = 1277;
			12369: out = -91;
			12370: out = -779;
			12371: out = -719;
			12372: out = 975;
			12373: out = 689;
			12374: out = -2075;
			12375: out = -1620;
			12376: out = -686;
			12377: out = 564;
			12378: out = 1181;
			12379: out = 109;
			12380: out = -158;
			12381: out = 1660;
			12382: out = -271;
			12383: out = -729;
			12384: out = -749;
			12385: out = -209;
			12386: out = 567;
			12387: out = 712;
			12388: out = -354;
			12389: out = -927;
			12390: out = -1184;
			12391: out = -300;
			12392: out = 1635;
			12393: out = 1694;
			12394: out = 1050;
			12395: out = 470;
			12396: out = -1583;
			12397: out = -1902;
			12398: out = -1166;
			12399: out = 113;
			12400: out = -2;
			12401: out = 7;
			12402: out = 730;
			12403: out = 460;
			12404: out = 709;
			12405: out = 311;
			12406: out = 113;
			12407: out = -2225;
			12408: out = -2233;
			12409: out = 685;
			12410: out = 219;
			12411: out = 2105;
			12412: out = 2588;
			12413: out = -605;
			12414: out = -1032;
			12415: out = -489;
			12416: out = 1655;
			12417: out = -2828;
			12418: out = -1172;
			12419: out = 1210;
			12420: out = 1886;
			12421: out = 311;
			12422: out = -1253;
			12423: out = -1720;
			12424: out = 911;
			12425: out = 415;
			12426: out = -464;
			12427: out = 1708;
			12428: out = 68;
			12429: out = -191;
			12430: out = -130;
			12431: out = -31;
			12432: out = -730;
			12433: out = -1091;
			12434: out = 288;
			12435: out = -705;
			12436: out = -539;
			12437: out = 171;
			12438: out = 2137;
			12439: out = 802;
			12440: out = -1201;
			12441: out = -1712;
			12442: out = -666;
			12443: out = 365;
			12444: out = 7;
			12445: out = 1375;
			12446: out = 365;
			12447: out = 227;
			12448: out = -321;
			12449: out = 2069;
			12450: out = 677;
			12451: out = -1998;
			12452: out = -3356;
			12453: out = -716;
			12454: out = 1773;
			12455: out = 1197;
			12456: out = 43;
			12457: out = -462;
			12458: out = 464;
			12459: out = -220;
			12460: out = -227;
			12461: out = -496;
			12462: out = 472;
			12463: out = 1005;
			12464: out = 1828;
			12465: out = 1008;
			12466: out = -1892;
			12467: out = -3844;
			12468: out = -3112;
			12469: out = 529;
			12470: out = 167;
			12471: out = 706;
			12472: out = 638;
			12473: out = -1391;
			12474: out = -1103;
			12475: out = -449;
			12476: out = -102;
			12477: out = 205;
			12478: out = 417;
			12479: out = 551;
			12480: out = -1167;
			12481: out = 123;
			12482: out = 673;
			12483: out = 136;
			12484: out = 340;
			12485: out = 454;
			12486: out = 594;
			12487: out = 170;
			12488: out = 209;
			12489: out = -190;
			12490: out = -1217;
			12491: out = 224;
			12492: out = 116;
			12493: out = -307;
			12494: out = -1525;
			12495: out = -268;
			12496: out = 540;
			12497: out = 956;
			12498: out = -1004;
			12499: out = 303;
			12500: out = 2157;
			12501: out = 1866;
			12502: out = 399;
			12503: out = -1071;
			12504: out = -967;
			12505: out = -1028;
			12506: out = 35;
			12507: out = 885;
			12508: out = 2030;
			12509: out = 733;
			12510: out = -44;
			12511: out = -89;
			12512: out = -1161;
			12513: out = -862;
			12514: out = -96;
			12515: out = 1512;
			12516: out = 433;
			12517: out = 24;
			12518: out = 191;
			12519: out = 1351;
			12520: out = 571;
			12521: out = -209;
			12522: out = 583;
			12523: out = -564;
			12524: out = -1274;
			12525: out = -1423;
			12526: out = -98;
			12527: out = 971;
			12528: out = 1049;
			12529: out = -1059;
			12530: out = -766;
			12531: out = -1060;
			12532: out = -1051;
			12533: out = -303;
			12534: out = 793;
			12535: out = 1679;
			12536: out = 1537;
			12537: out = 947;
			12538: out = -641;
			12539: out = -1991;
			12540: out = -1258;
			12541: out = -152;
			12542: out = 1061;
			12543: out = 1923;
			12544: out = 1748;
			12545: out = 998;
			12546: out = -364;
			12547: out = -995;
			12548: out = -2342;
			12549: out = -1931;
			12550: out = 363;
			12551: out = 1245;
			12552: out = 386;
			12553: out = -1386;
			12554: out = 681;
			12555: out = 36;
			12556: out = -240;
			12557: out = -978;
			12558: out = -207;
			12559: out = -402;
			12560: out = -386;
			12561: out = -172;
			12562: out = 831;
			12563: out = 662;
			12564: out = -1037;
			12565: out = -1328;
			12566: out = -1172;
			12567: out = -126;
			12568: out = 84;
			12569: out = 1448;
			12570: out = 968;
			12571: out = -1369;
			12572: out = -251;
			12573: out = 458;
			12574: out = 965;
			12575: out = -2431;
			12576: out = 209;
			12577: out = 1363;
			12578: out = 1013;
			12579: out = -1536;
			12580: out = -520;
			12581: out = 1405;
			12582: out = -325;
			12583: out = -352;
			12584: out = -1099;
			12585: out = -518;
			12586: out = -514;
			12587: out = 830;
			12588: out = 837;
			12589: out = 183;
			12590: out = -2317;
			12591: out = -1861;
			12592: out = 1010;
			12593: out = 1557;
			12594: out = 877;
			12595: out = -122;
			12596: out = 2248;
			12597: out = 244;
			12598: out = -384;
			12599: out = -530;
			12600: out = 239;
			12601: out = -360;
			12602: out = -767;
			12603: out = 346;
			12604: out = 170;
			12605: out = 329;
			12606: out = 149;
			12607: out = 685;
			12608: out = -818;
			12609: out = -1831;
			12610: out = -649;
			12611: out = 395;
			12612: out = 863;
			12613: out = -39;
			12614: out = 1289;
			12615: out = 74;
			12616: out = -417;
			12617: out = 114;
			12618: out = 767;
			12619: out = 320;
			12620: out = -602;
			12621: out = -835;
			12622: out = 165;
			12623: out = 546;
			12624: out = -1642;
			12625: out = 167;
			12626: out = 974;
			12627: out = 1170;
			12628: out = -1655;
			12629: out = -976;
			12630: out = 290;
			12631: out = 412;
			12632: out = 1574;
			12633: out = 925;
			12634: out = -290;
			12635: out = -462;
			12636: out = -156;
			12637: out = -80;
			12638: out = -1238;
			12639: out = 689;
			12640: out = 1122;
			12641: out = 548;
			12642: out = 314;
			12643: out = -1439;
			12644: out = -1906;
			12645: out = 32;
			12646: out = -1055;
			12647: out = -734;
			12648: out = 200;
			12649: out = 1805;
			12650: out = 1690;
			12651: out = 674;
			12652: out = -905;
			12653: out = -836;
			12654: out = -684;
			12655: out = -388;
			12656: out = 112;
			12657: out = -3;
			12658: out = 195;
			12659: out = 1166;
			12660: out = -297;
			12661: out = -310;
			12662: out = 192;
			12663: out = -263;
			12664: out = 94;
			12665: out = 632;
			12666: out = 1968;
			12667: out = -811;
			12668: out = -813;
			12669: out = 23;
			12670: out = -254;
			12671: out = -215;
			12672: out = 3;
			12673: out = 454;
			12674: out = -848;
			12675: out = -1616;
			12676: out = -1564;
			12677: out = -532;
			12678: out = 326;
			12679: out = 468;
			12680: out = 131;
			12681: out = -715;
			12682: out = -146;
			12683: out = 875;
			12684: out = 1876;
			12685: out = 581;
			12686: out = -580;
			12687: out = -1086;
			12688: out = 633;
			12689: out = -79;
			12690: out = -1138;
			12691: out = 1295;
			12692: out = 75;
			12693: out = -260;
			12694: out = -144;
			12695: out = 932;
			12696: out = 668;
			12697: out = -250;
			12698: out = -390;
			12699: out = -1678;
			12700: out = -1351;
			12701: out = 45;
			12702: out = 1760;
			12703: out = 602;
			12704: out = -1352;
			12705: out = -913;
			12706: out = -1374;
			12707: out = -735;
			12708: out = -420;
			12709: out = 1926;
			12710: out = 786;
			12711: out = -312;
			12712: out = 309;
			12713: out = 199;
			12714: out = 107;
			12715: out = -104;
			12716: out = -232;
			12717: out = 390;
			12718: out = 861;
			12719: out = 414;
			12720: out = 523;
			12721: out = 346;
			12722: out = 102;
			12723: out = -74;
			12724: out = -437;
			12725: out = -407;
			12726: out = 190;
			12727: out = 472;
			12728: out = -168;
			12729: out = -1325;
			12730: out = -186;
			12731: out = -88;
			12732: out = 180;
			12733: out = -23;
			12734: out = -36;
			12735: out = -710;
			12736: out = -1246;
			12737: out = -1876;
			12738: out = -199;
			12739: out = 1308;
			12740: out = 1203;
			12741: out = 350;
			12742: out = -390;
			12743: out = -15;
			12744: out = -758;
			12745: out = 1333;
			12746: out = 2125;
			12747: out = 1497;
			12748: out = 87;
			12749: out = -109;
			12750: out = -239;
			12751: out = -2149;
			12752: out = -2452;
			12753: out = -1285;
			12754: out = 979;
			12755: out = 1775;
			12756: out = 1071;
			12757: out = -692;
			12758: out = -2364;
			12759: out = -2057;
			12760: out = -408;
			12761: out = 1856;
			12762: out = 11;
			12763: out = 904;
			12764: out = 1703;
			12765: out = -896;
			12766: out = -1759;
			12767: out = -2050;
			12768: out = -852;
			12769: out = -304;
			12770: out = 433;
			12771: out = 575;
			12772: out = 932;
			12773: out = 187;
			12774: out = -206;
			12775: out = -493;
			12776: out = -32;
			12777: out = -445;
			12778: out = -596;
			12779: out = 936;
			12780: out = 415;
			12781: out = -81;
			12782: out = -838;
			12783: out = 785;
			12784: out = 499;
			12785: out = -220;
			12786: out = -1896;
			12787: out = -386;
			12788: out = -396;
			12789: out = -1465;
			12790: out = -508;
			12791: out = 666;
			12792: out = 1444;
			12793: out = 46;
			12794: out = 68;
			12795: out = -232;
			12796: out = -1;
			12797: out = -82;
			12798: out = 106;
			12799: out = -178;
			12800: out = -334;
			12801: out = -974;
			12802: out = -612;
			12803: out = 256;
			12804: out = 1577;
			12805: out = 929;
			12806: out = -123;
			12807: out = 33;
			12808: out = 258;
			12809: out = 961;
			12810: out = 867;
			12811: out = -196;
			12812: out = -1068;
			12813: out = -656;
			12814: out = 220;
			12815: out = 2652;
			12816: out = 1950;
			12817: out = -682;
			12818: out = -1506;
			12819: out = -1627;
			12820: out = -706;
			12821: out = -586;
			12822: out = 949;
			12823: out = 767;
			12824: out = -59;
			12825: out = -2312;
			12826: out = -1316;
			12827: out = 192;
			12828: out = 775;
			12829: out = 498;
			12830: out = 104;
			12831: out = 187;
			12832: out = -865;
			12833: out = 374;
			12834: out = 629;
			12835: out = -524;
			12836: out = -479;
			12837: out = 376;
			12838: out = 1481;
			12839: out = 163;
			12840: out = 117;
			12841: out = 26;
			12842: out = 978;
			12843: out = -182;
			12844: out = 214;
			12845: out = 469;
			12846: out = 910;
			12847: out = -797;
			12848: out = -1258;
			12849: out = -56;
			12850: out = -53;
			12851: out = -699;
			12852: out = -1317;
			12853: out = 609;
			12854: out = 329;
			12855: out = 198;
			12856: out = 79;
			12857: out = -1515;
			12858: out = -1248;
			12859: out = -87;
			12860: out = 28;
			12861: out = 781;
			12862: out = 641;
			12863: out = 108;
			12864: out = -101;
			12865: out = -180;
			12866: out = -50;
			12867: out = 239;
			12868: out = 496;
			12869: out = 251;
			12870: out = -541;
			12871: out = -167;
			12872: out = 303;
			12873: out = 966;
			12874: out = 326;
			12875: out = 1330;
			12876: out = 56;
			12877: out = -2693;
			12878: out = -627;
			12879: out = 358;
			12880: out = 1030;
			12881: out = -1049;
			12882: out = 111;
			12883: out = -489;
			12884: out = -1333;
			12885: out = -429;
			12886: out = 1294;
			12887: out = 1927;
			12888: out = 464;
			12889: out = -276;
			12890: out = -284;
			12891: out = 297;
			12892: out = 786;
			12893: out = -134;
			12894: out = -900;
			12895: out = -445;
			12896: out = 1322;
			12897: out = 1399;
			12898: out = -189;
			12899: out = 1142;
			12900: out = 324;
			12901: out = -892;
			12902: out = -3709;
			12903: out = -1263;
			12904: out = 858;
			12905: out = 2284;
			12906: out = -1072;
			12907: out = -430;
			12908: out = 367;
			12909: out = 769;
			12910: out = -1244;
			12911: out = -1508;
			12912: out = 25;
			12913: out = 1023;
			12914: out = 1645;
			12915: out = 176;
			12916: out = -2850;
			12917: out = -2094;
			12918: out = -508;
			12919: out = 935;
			12920: out = -437;
			12921: out = -451;
			12922: out = 115;
			12923: out = 2062;
			12924: out = -95;
			12925: out = -792;
			12926: out = -1032;
			12927: out = 370;
			12928: out = -497;
			12929: out = -386;
			12930: out = 641;
			12931: out = 2368;
			12932: out = 1191;
			12933: out = -1221;
			12934: out = 88;
			12935: out = -406;
			12936: out = 217;
			12937: out = 367;
			12938: out = 970;
			12939: out = -523;
			12940: out = -1766;
			12941: out = -128;
			12942: out = 257;
			12943: out = 906;
			12944: out = 1561;
			12945: out = 434;
			12946: out = -800;
			12947: out = -1710;
			12948: out = 1056;
			12949: out = -957;
			12950: out = -1073;
			12951: out = -97;
			12952: out = 1608;
			12953: out = -556;
			12954: out = -2919;
			12955: out = -552;
			12956: out = 455;
			12957: out = 1042;
			12958: out = -462;
			12959: out = 222;
			12960: out = -573;
			12961: out = -848;
			12962: out = -2210;
			12963: out = 187;
			12964: out = 949;
			12965: out = 530;
			12966: out = 822;
			12967: out = 1293;
			12968: out = 1489;
			12969: out = 421;
			12970: out = 171;
			12971: out = -743;
			12972: out = -1767;
			12973: out = 22;
			12974: out = 231;
			12975: out = 334;
			12976: out = 470;
			12977: out = 171;
			12978: out = -1127;
			12979: out = -2219;
			12980: out = 751;
			12981: out = 2042;
			12982: out = 1610;
			12983: out = -1572;
			12984: out = -1402;
			12985: out = -967;
			12986: out = 96;
			12987: out = 125;
			12988: out = 840;
			12989: out = 1060;
			12990: out = 767;
			12991: out = 52;
			12992: out = -224;
			12993: out = 14;
			12994: out = -274;
			12995: out = 303;
			12996: out = 432;
			12997: out = 101;
			12998: out = -1161;
			12999: out = -869;
			13000: out = 519;
			13001: out = 39;
			13002: out = 719;
			13003: out = 509;
			13004: out = -93;
			13005: out = -668;
			13006: out = -1051;
			13007: out = -1393;
			13008: out = 54;
			13009: out = -214;
			13010: out = 189;
			13011: out = 427;
			13012: out = 1894;
			13013: out = 216;
			13014: out = -1884;
			13015: out = -8;
			13016: out = 324;
			13017: out = 468;
			13018: out = 137;
			13019: out = 630;
			13020: out = 555;
			13021: out = -274;
			13022: out = 1699;
			13023: out = -2168;
			13024: out = -2790;
			13025: out = 292;
			13026: out = 2460;
			13027: out = 685;
			13028: out = -2637;
			13029: out = -1110;
			13030: out = -408;
			13031: out = -114;
			13032: out = -2599;
			13033: out = 1802;
			13034: out = 1826;
			13035: out = 1012;
			13036: out = -436;
			13037: out = -1048;
			13038: out = -1691;
			13039: out = -1862;
			13040: out = -52;
			13041: out = 683;
			13042: out = 368;
			13043: out = 40;
			13044: out = -259;
			13045: out = 269;
			13046: out = 447;
			13047: out = -84;
			13048: out = -1444;
			13049: out = -1486;
			13050: out = 1169;
			13051: out = 1446;
			13052: out = 856;
			13053: out = -172;
			13054: out = -439;
			13055: out = 598;
			13056: out = 1298;
			13057: out = 93;
			13058: out = -1143;
			13059: out = -1441;
			13060: out = -72;
			13061: out = -19;
			13062: out = 445;
			13063: out = 156;
			13064: out = 327;
			13065: out = -93;
			13066: out = 485;
			13067: out = 1007;
			13068: out = 46;
			13069: out = -583;
			13070: out = -653;
			13071: out = -791;
			13072: out = 793;
			13073: out = 698;
			13074: out = -205;
			13075: out = -172;
			13076: out = 1258;
			13077: out = 2261;
			13078: out = 434;
			13079: out = 593;
			13080: out = -968;
			13081: out = -2401;
			13082: out = -1738;
			13083: out = -700;
			13084: out = 416;
			13085: out = 1041;
			13086: out = 284;
			13087: out = -185;
			13088: out = 101;
			13089: out = -263;
			13090: out = 400;
			13091: out = 345;
			13092: out = 7;
			13093: out = -1452;
			13094: out = -793;
			13095: out = 829;
			13096: out = 984;
			13097: out = 47;
			13098: out = -652;
			13099: out = 1083;
			13100: out = -386;
			13101: out = -360;
			13102: out = -400;
			13103: out = 1480;
			13104: out = -844;
			13105: out = -2025;
			13106: out = -764;
			13107: out = 403;
			13108: out = 1024;
			13109: out = 631;
			13110: out = 669;
			13111: out = -149;
			13112: out = -545;
			13113: out = -723;
			13114: out = 357;
			13115: out = 347;
			13116: out = -26;
			13117: out = 1131;
			13118: out = 231;
			13119: out = -309;
			13120: out = -418;
			13121: out = 1311;
			13122: out = 619;
			13123: out = -1058;
			13124: out = 347;
			13125: out = -818;
			13126: out = -1318;
			13127: out = -2393;
			13128: out = 867;
			13129: out = -31;
			13130: out = -1339;
			13131: out = -68;
			13132: out = 1280;
			13133: out = 1530;
			13134: out = -132;
			13135: out = -452;
			13136: out = -867;
			13137: out = -517;
			13138: out = -73;
			13139: out = 60;
			13140: out = -251;
			13141: out = -640;
			13142: out = 1567;
			13143: out = 1717;
			13144: out = 903;
			13145: out = -460;
			13146: out = -48;
			13147: out = -213;
			13148: out = -1167;
			13149: out = -83;
			13150: out = -55;
			13151: out = -58;
			13152: out = -159;
			13153: out = 328;
			13154: out = 517;
			13155: out = 82;
			13156: out = -7;
			13157: out = -464;
			13158: out = -591;
			13159: out = -2265;
			13160: out = 555;
			13161: out = 345;
			13162: out = -1554;
			13163: out = -1679;
			13164: out = 302;
			13165: out = 2475;
			13166: out = 2570;
			13167: out = 1387;
			13168: out = 152;
			13169: out = -207;
			13170: out = -473;
			13171: out = -703;
			13172: out = -414;
			13173: out = 1074;
			13174: out = 1239;
			13175: out = 739;
			13176: out = -241;
			13177: out = 464;
			13178: out = 244;
			13179: out = -325;
			13180: out = -1499;
			13181: out = -1992;
			13182: out = -1258;
			13183: out = 480;
			13184: out = 320;
			13185: out = 485;
			13186: out = 24;
			13187: out = 264;
			13188: out = -528;
			13189: out = -63;
			13190: out = 235;
			13191: out = 1421;
			13192: out = -320;
			13193: out = -1025;
			13194: out = -86;
			13195: out = 1066;
			13196: out = 795;
			13197: out = 9;
			13198: out = 411;
			13199: out = 1172;
			13200: out = 1002;
			13201: out = -725;
			13202: out = -1560;
			13203: out = -1340;
			13204: out = -122;
			13205: out = 915;
			13206: out = -311;
			13207: out = -1157;
			13208: out = 94;
			13209: out = 179;
			13210: out = 686;
			13211: out = 204;
			13212: out = 258;
			13213: out = -890;
			13214: out = -899;
			13215: out = -486;
			13216: out = 123;
			13217: out = -381;
			13218: out = -887;
			13219: out = -1781;
			13220: out = 662;
			13221: out = 1350;
			13222: out = -325;
			13223: out = 264;
			13224: out = 59;
			13225: out = 444;
			13226: out = 943;
			13227: out = 490;
			13228: out = 20;
			13229: out = 132;
			13230: out = -473;
			13231: out = -792;
			13232: out = -1008;
			13233: out = 251;
			13234: out = 50;
			13235: out = 369;
			13236: out = 68;
			13237: out = 1432;
			13238: out = -744;
			13239: out = -2544;
			13240: out = -1848;
			13241: out = 44;
			13242: out = 871;
			13243: out = -127;
			13244: out = -487;
			13245: out = -389;
			13246: out = 446;
			13247: out = 69;
			13248: out = 1078;
			13249: out = 43;
			13250: out = -1776;
			13251: out = -688;
			13252: out = -316;
			13253: out = 155;
			13254: out = -81;
			13255: out = 706;
			13256: out = 777;
			13257: out = 776;
			13258: out = -428;
			13259: out = 188;
			13260: out = 397;
			13261: out = -5;
			13262: out = -1120;
			13263: out = -535;
			13264: out = 1025;
			13265: out = 724;
			13266: out = -49;
			13267: out = -778;
			13268: out = 352;
			13269: out = -680;
			13270: out = -373;
			13271: out = 29;
			13272: out = 245;
			13273: out = 180;
			13274: out = 364;
			13275: out = 1060;
			13276: out = 605;
			13277: out = -34;
			13278: out = -756;
			13279: out = 824;
			13280: out = 147;
			13281: out = 66;
			13282: out = 395;
			13283: out = 353;
			13284: out = -1310;
			13285: out = -2823;
			13286: out = 512;
			13287: out = 535;
			13288: out = 380;
			13289: out = -69;
			13290: out = 162;
			13291: out = 376;
			13292: out = 424;
			13293: out = -115;
			13294: out = -403;
			13295: out = -260;
			13296: out = 278;
			13297: out = 439;
			13298: out = 380;
			13299: out = 67;
			13300: out = -754;
			13301: out = 78;
			13302: out = 364;
			13303: out = -587;
			13304: out = -28;
			13305: out = 20;
			13306: out = 137;
			13307: out = -1453;
			13308: out = 173;
			13309: out = 690;
			13310: out = -224;
			13311: out = -773;
			13312: out = -1029;
			13313: out = -280;
			13314: out = 913;
			13315: out = 1167;
			13316: out = 477;
			13317: out = -447;
			13318: out = -18;
			13319: out = 635;
			13320: out = 886;
			13321: out = 105;
			13322: out = -733;
			13323: out = -846;
			13324: out = 125;
			13325: out = 538;
			13326: out = 567;
			13327: out = -189;
			13328: out = 7;
			13329: out = -1676;
			13330: out = -1452;
			13331: out = 128;
			13332: out = 1315;
			13333: out = 996;
			13334: out = -537;
			13335: out = -2878;
			13336: out = -1666;
			13337: out = -166;
			13338: out = 528;
			13339: out = 32;
			13340: out = -336;
			13341: out = -217;
			13342: out = 294;
			13343: out = 472;
			13344: out = 662;
			13345: out = 768;
			13346: out = 199;
			13347: out = 117;
			13348: out = 156;
			13349: out = 134;
			13350: out = 799;
			13351: out = 1077;
			13352: out = 710;
			13353: out = -1393;
			13354: out = -1883;
			13355: out = -716;
			13356: out = 2288;
			13357: out = 516;
			13358: out = -1193;
			13359: out = -2642;
			13360: out = -958;
			13361: out = -351;
			13362: out = 819;
			13363: out = 1078;
			13364: out = 2200;
			13365: out = 103;
			13366: out = -2330;
			13367: out = -253;
			13368: out = 1267;
			13369: out = 1697;
			13370: out = -72;
			13371: out = -81;
			13372: out = -24;
			13373: out = 187;
			13374: out = 10;
			13375: out = -978;
			13376: out = -698;
			13377: out = 1675;
			13378: out = 1484;
			13379: out = 297;
			13380: out = -1737;
			13381: out = -827;
			13382: out = -1584;
			13383: out = -1325;
			13384: out = -607;
			13385: out = 1157;
			13386: out = 1686;
			13387: out = 1085;
			13388: out = -895;
			13389: out = -1336;
			13390: out = -915;
			13391: out = 52;
			13392: out = 177;
			13393: out = 392;
			13394: out = 471;
			13395: out = -75;
			13396: out = 340;
			13397: out = 502;
			13398: out = 475;
			13399: out = 124;
			13400: out = 398;
			13401: out = 695;
			13402: out = 63;
			13403: out = -104;
			13404: out = -296;
			13405: out = -474;
			13406: out = 364;
			13407: out = 319;
			13408: out = -49;
			13409: out = -484;
			13410: out = -95;
			13411: out = 75;
			13412: out = -112;
			13413: out = -85;
			13414: out = -88;
			13415: out = -90;
			13416: out = 151;
			13417: out = -179;
			13418: out = -85;
			13419: out = -159;
			13420: out = 214;
			13421: out = -627;
			13422: out = -881;
			13423: out = -224;
			13424: out = 1362;
			13425: out = 1126;
			13426: out = -431;
			13427: out = -1265;
			13428: out = -278;
			13429: out = 884;
			13430: out = -49;
			13431: out = 151;
			13432: out = 46;
			13433: out = 48;
			13434: out = 44;
			13435: out = -1536;
			13436: out = -2262;
			13437: out = 808;
			13438: out = 107;
			13439: out = 286;
			13440: out = -267;
			13441: out = 202;
			13442: out = -1319;
			13443: out = -1513;
			13444: out = 367;
			13445: out = 853;
			13446: out = 988;
			13447: out = 645;
			13448: out = -7;
			13449: out = -103;
			13450: out = -138;
			13451: out = 191;
			13452: out = -420;
			13453: out = -217;
			13454: out = 49;
			13455: out = 1804;
			13456: out = 303;
			13457: out = -501;
			13458: out = -70;
			13459: out = 921;
			13460: out = -367;
			13461: out = -2387;
			13462: out = -409;
			13463: out = 162;
			13464: out = 375;
			13465: out = -530;
			13466: out = -855;
			13467: out = -785;
			13468: out = -121;
			13469: out = 1514;
			13470: out = -204;
			13471: out = -1665;
			13472: out = -1361;
			13473: out = -213;
			13474: out = 248;
			13475: out = 12;
			13476: out = 2087;
			13477: out = 961;
			13478: out = 161;
			13479: out = -431;
			13480: out = 611;
			13481: out = 510;
			13482: out = 180;
			13483: out = 1528;
			13484: out = 571;
			13485: out = -183;
			13486: out = -767;
			13487: out = 554;
			13488: out = 463;
			13489: out = -3;
			13490: out = -790;
			13491: out = 84;
			13492: out = 419;
			13493: out = -18;
			13494: out = -674;
			13495: out = -410;
			13496: out = 288;
			13497: out = 670;
			13498: out = 136;
			13499: out = -195;
			13500: out = -78;
			13501: out = -199;
			13502: out = -168;
			13503: out = -42;
			13504: out = -252;
			13505: out = 171;
			13506: out = -2;
			13507: out = -97;
			13508: out = -285;
			13509: out = 984;
			13510: out = 1351;
			13511: out = -179;
			13512: out = -1638;
			13513: out = -891;
			13514: out = 1690;
			13515: out = 40;
			13516: out = -198;
			13517: out = -527;
			13518: out = -143;
			13519: out = -237;
			13520: out = -99;
			13521: out = 104;
			13522: out = -145;
			13523: out = 247;
			13524: out = 336;
			13525: out = 134;
			13526: out = -1351;
			13527: out = -852;
			13528: out = 948;
			13529: out = 630;
			13530: out = -369;
			13531: out = -1460;
			13532: out = -195;
			13533: out = -407;
			13534: out = 67;
			13535: out = -49;
			13536: out = 2356;
			13537: out = 745;
			13538: out = -394;
			13539: out = -200;
			13540: out = 183;
			13541: out = -892;
			13542: out = -2610;
			13543: out = -142;
			13544: out = 141;
			13545: out = 866;
			13546: out = 1578;
			13547: out = 992;
			13548: out = -373;
			13549: out = -1777;
			13550: out = -934;
			13551: out = -1061;
			13552: out = -825;
			13553: out = -730;
			13554: out = 390;
			13555: out = 39;
			13556: out = -812;
			13557: out = -1209;
			13558: out = -158;
			13559: out = 795;
			13560: out = 646;
			13561: out = 377;
			13562: out = -194;
			13563: out = -434;
			13564: out = -957;
			13565: out = -240;
			13566: out = 408;
			13567: out = 468;
			13568: out = 1198;
			13569: out = 782;
			13570: out = 78;
			13571: out = -23;
			13572: out = 78;
			13573: out = 316;
			13574: out = 425;
			13575: out = -742;
			13576: out = -891;
			13577: out = 148;
			13578: out = 2592;
			13579: out = 1185;
			13580: out = -801;
			13581: out = -1770;
			13582: out = -1088;
			13583: out = 207;
			13584: out = 599;
			13585: out = 252;
			13586: out = -1830;
			13587: out = -1694;
			13588: out = 1433;
			13589: out = 491;
			13590: out = 1182;
			13591: out = 946;
			13592: out = 890;
			13593: out = -1920;
			13594: out = -2690;
			13595: out = -890;
			13596: out = 343;
			13597: out = 1142;
			13598: out = 724;
			13599: out = 639;
			13600: out = -1195;
			13601: out = -793;
			13602: out = 1521;
			13603: out = 110;
			13604: out = 309;
			13605: out = 154;
			13606: out = 1146;
			13607: out = -1533;
			13608: out = -1658;
			13609: out = 252;
			13610: out = 77;
			13611: out = 111;
			13612: out = -141;
			13613: out = 558;
			13614: out = -11;
			13615: out = -567;
			13616: out = -1283;
			13617: out = 680;
			13618: out = 331;
			13619: out = -265;
			13620: out = -652;
			13621: out = -133;
			13622: out = 660;
			13623: out = 1184;
			13624: out = -19;
			13625: out = 49;
			13626: out = 246;
			13627: out = 158;
			13628: out = 8;
			13629: out = -136;
			13630: out = -66;
			13631: out = -442;
			13632: out = -442;
			13633: out = -253;
			13634: out = 546;
			13635: out = 111;
			13636: out = 53;
			13637: out = -329;
			13638: out = -253;
			13639: out = -1489;
			13640: out = -1463;
			13641: out = 51;
			13642: out = 294;
			13643: out = -637;
			13644: out = -1800;
			13645: out = 291;
			13646: out = 467;
			13647: out = 281;
			13648: out = -686;
			13649: out = -100;
			13650: out = 306;
			13651: out = 469;
			13652: out = 89;
			13653: out = -1038;
			13654: out = -1041;
			13655: out = 1076;
			13656: out = -16;
			13657: out = 408;
			13658: out = 912;
			13659: out = 1476;
			13660: out = 663;
			13661: out = -509;
			13662: out = -1586;
			13663: out = -1612;
			13664: out = -556;
			13665: out = 802;
			13666: out = -2;
			13667: out = 756;
			13668: out = 604;
			13669: out = 536;
			13670: out = -1685;
			13671: out = -939;
			13672: out = 206;
			13673: out = 197;
			13674: out = -855;
			13675: out = -353;
			13676: out = 2265;
			13677: out = 8;
			13678: out = 422;
			13679: out = 676;
			13680: out = -141;
			13681: out = 483;
			13682: out = 897;
			13683: out = 824;
			13684: out = -736;
			13685: out = -858;
			13686: out = 32;
			13687: out = 1125;
			13688: out = 398;
			13689: out = -381;
			13690: out = -373;
			13691: out = -2072;
			13692: out = -1159;
			13693: out = -95;
			13694: out = 262;
			13695: out = -403;
			13696: out = -198;
			13697: out = 941;
			13698: out = 194;
			13699: out = 243;
			13700: out = 284;
			13701: out = 1318;
			13702: out = 220;
			13703: out = -501;
			13704: out = -1276;
			13705: out = 533;
			13706: out = -374;
			13707: out = -770;
			13708: out = 319;
			13709: out = 982;
			13710: out = 1084;
			13711: out = 559;
			13712: out = -57;
			13713: out = -135;
			13714: out = -17;
			13715: out = 136;
			13716: out = -785;
			13717: out = -782;
			13718: out = -295;
			13719: out = -25;
			13720: out = -421;
			13721: out = -488;
			13722: out = 299;
			13723: out = 995;
			13724: out = 1080;
			13725: out = 391;
			13726: out = -1378;
			13727: out = -1446;
			13728: out = -842;
			13729: out = 264;
			13730: out = -345;
			13731: out = -133;
			13732: out = -52;
			13733: out = 419;
			13734: out = -975;
			13735: out = -1010;
			13736: out = 628;
			13737: out = 1563;
			13738: out = 713;
			13739: out = -1048;
			13740: out = -2290;
			13741: out = -559;
			13742: out = 623;
			13743: out = -817;
			13744: out = 495;
			13745: out = 814;
			13746: out = 1225;
			13747: out = -161;
			13748: out = 353;
			13749: out = 440;
			13750: out = 83;
			13751: out = -247;
			13752: out = -450;
			13753: out = -232;
			13754: out = -224;
			13755: out = 1585;
			13756: out = 2063;
			13757: out = 636;
			13758: out = -80;
			13759: out = -998;
			13760: out = -1119;
			13761: out = -441;
			13762: out = -119;
			13763: out = -2;
			13764: out = -41;
			13765: out = 116;
			13766: out = 388;
			13767: out = 842;
			13768: out = 809;
			13769: out = 372;
			13770: out = -604;
			13771: out = -836;
			13772: out = -2025;
			13773: out = 65;
			13774: out = 1672;
			13775: out = 143;
			13776: out = -1467;
			13777: out = -1542;
			13778: out = 937;
			13779: out = 1113;
			13780: out = 1003;
			13781: out = -186;
			13782: out = 1300;
			13783: out = -1607;
			13784: out = -1587;
			13785: out = -216;
			13786: out = 1361;
			13787: out = 276;
			13788: out = -737;
			13789: out = 196;
			13790: out = 1040;
			13791: out = 1317;
			13792: out = 656;
			13793: out = -1083;
			13794: out = -785;
			13795: out = 69;
			13796: out = 91;
			13797: out = -226;
			13798: out = -524;
			13799: out = -267;
			13800: out = 1028;
			13801: out = 798;
			13802: out = 86;
			13803: out = -746;
			13804: out = 407;
			13805: out = 138;
			13806: out = -1132;
			13807: out = 101;
			13808: out = 110;
			13809: out = 144;
			13810: out = -220;
			13811: out = -152;
			13812: out = -207;
			13813: out = -88;
			13814: out = 644;
			13815: out = 364;
			13816: out = -294;
			13817: out = -1323;
			13818: out = -41;
			13819: out = -94;
			13820: out = -764;
			13821: out = 137;
			13822: out = 308;
			13823: out = 306;
			13824: out = -527;
			13825: out = 373;
			13826: out = 217;
			13827: out = -192;
			13828: out = -942;
			13829: out = -101;
			13830: out = 505;
			13831: out = -217;
			13832: out = 261;
			13833: out = 205;
			13834: out = 325;
			13835: out = -2257;
			13836: out = 293;
			13837: out = 1286;
			13838: out = -313;
			13839: out = -1188;
			13840: out = -1063;
			13841: out = 0;
			13842: out = -2262;
			13843: out = 213;
			13844: out = 1598;
			13845: out = 1501;
			13846: out = 211;
			13847: out = -262;
			13848: out = 128;
			13849: out = 85;
			13850: out = 679;
			13851: out = 303;
			13852: out = -458;
			13853: out = -1434;
			13854: out = -823;
			13855: out = 189;
			13856: out = 160;
			13857: out = 253;
			13858: out = 276;
			13859: out = 465;
			13860: out = 192;
			13861: out = -442;
			13862: out = -1058;
			13863: out = -871;
			13864: out = -315;
			13865: out = 177;
			13866: out = 91;
			13867: out = 73;
			13868: out = 54;
			13869: out = 284;
			13870: out = -114;
			13871: out = 603;
			13872: out = 619;
			13873: out = 357;
			13874: out = -1337;
			13875: out = -861;
			13876: out = 259;
			13877: out = 626;
			13878: out = 1139;
			13879: out = 742;
			13880: out = -120;
			13881: out = 1115;
			13882: out = 565;
			13883: out = -154;
			13884: out = -431;
			13885: out = -453;
			13886: out = -242;
			13887: out = 267;
			13888: out = -538;
			13889: out = 550;
			13890: out = 1008;
			13891: out = 0;
			13892: out = -1590;
			13893: out = -1806;
			13894: out = -305;
			13895: out = -289;
			13896: out = 709;
			13897: out = 695;
			13898: out = -64;
			13899: out = -765;
			13900: out = -692;
			13901: out = 75;
			13902: out = 330;
			13903: out = 845;
			13904: out = 668;
			13905: out = -199;
			13906: out = -162;
			13907: out = -243;
			13908: out = -389;
			13909: out = 466;
			13910: out = 393;
			13911: out = 306;
			13912: out = -604;
			13913: out = 102;
			13914: out = -1044;
			13915: out = -1901;
			13916: out = -178;
			13917: out = 1030;
			13918: out = 917;
			13919: out = -741;
			13920: out = -301;
			13921: out = 741;
			13922: out = 1501;
			13923: out = 164;
			13924: out = -847;
			13925: out = -1031;
			13926: out = -12;
			13927: out = 949;
			13928: out = 675;
			13929: out = -484;
			13930: out = -1980;
			13931: out = -911;
			13932: out = 606;
			13933: out = 1602;
			13934: out = 361;
			13935: out = 382;
			13936: out = 580;
			13937: out = 188;
			13938: out = -1913;
			13939: out = -1951;
			13940: out = 1154;
			13941: out = 441;
			13942: out = 678;
			13943: out = -254;
			13944: out = -673;
			13945: out = -2181;
			13946: out = -1445;
			13947: out = 695;
			13948: out = 236;
			13949: out = 148;
			13950: out = -26;
			13951: out = 23;
			13952: out = -41;
			13953: out = -267;
			13954: out = -590;
			13955: out = -160;
			13956: out = 599;
			13957: out = 1235;
			13958: out = 336;
			13959: out = 591;
			13960: out = 151;
			13961: out = -107;
			13962: out = -1226;
			13963: out = 98;
			13964: out = 1334;
			13965: out = 774;
			13966: out = 245;
			13967: out = -500;
			13968: out = -561;
			13969: out = -17;
			13970: out = 371;
			13971: out = 381;
			13972: out = 165;
			13973: out = -5;
			13974: out = -735;
			13975: out = -1799;
			13976: out = -56;
			13977: out = -47;
			13978: out = 97;
			13979: out = 146;
			13980: out = 867;
			13981: out = 430;
			13982: out = -464;
			13983: out = -35;
			13984: out = 109;
			13985: out = 206;
			13986: out = 207;
			13987: out = -96;
			13988: out = -26;
			13989: out = 83;
			13990: out = 19;
			13991: out = -464;
			13992: out = -494;
			13993: out = -44;
			13994: out = 968;
			13995: out = 474;
			13996: out = -854;
			13997: out = -312;
			13998: out = -451;
			13999: out = -163;
			14000: out = 491;
			14001: out = -669;
			14002: out = -618;
			14003: out = 123;
			14004: out = 86;
			14005: out = -131;
			14006: out = -439;
			14007: out = -283;
			14008: out = 249;
			14009: out = 843;
			14010: out = 895;
			14011: out = -1384;
			14012: out = -665;
			14013: out = 196;
			14014: out = 472;
			14015: out = 1128;
			14016: out = 1804;
			14017: out = 1655;
			14018: out = -1626;
			14019: out = -2118;
			14020: out = -1035;
			14021: out = 1764;
			14022: out = -171;
			14023: out = -446;
			14024: out = -418;
			14025: out = -610;
			14026: out = -672;
			14027: out = -367;
			14028: out = 316;
			14029: out = 775;
			14030: out = 989;
			14031: out = 528;
			14032: out = -1374;
			14033: out = -1056;
			14034: out = -41;
			14035: out = 917;
			14036: out = 294;
			14037: out = -460;
			14038: out = -900;
			14039: out = -101;
			14040: out = 83;
			14041: out = 410;
			14042: out = 580;
			14043: out = -1107;
			14044: out = -1955;
			14045: out = -1410;
			14046: out = 1406;
			14047: out = 1475;
			14048: out = 824;
			14049: out = -535;
			14050: out = 719;
			14051: out = 95;
			14052: out = -394;
			14053: out = 114;
			14054: out = 220;
			14055: out = -180;
			14056: out = -944;
			14057: out = 138;
			14058: out = 196;
			14059: out = 221;
			14060: out = 968;
			14061: out = 317;
			14062: out = 2;
			14063: out = -507;
			14064: out = 547;
			14065: out = -1160;
			14066: out = -2231;
			14067: out = -169;
			14068: out = 177;
			14069: out = 548;
			14070: out = 88;
			14071: out = 338;
			14072: out = -196;
			14073: out = -415;
			14074: out = -665;
			14075: out = 779;
			14076: out = 1116;
			14077: out = 435;
			14078: out = -464;
			14079: out = -825;
			14080: out = -337;
			14081: out = 50;
			14082: out = 1398;
			14083: out = 1034;
			14084: out = -16;
			14085: out = -373;
			14086: out = 221;
			14087: out = 434;
			14088: out = -1120;
			14089: out = -1108;
			14090: out = -545;
			14091: out = 945;
			14092: out = -904;
			14093: out = 669;
			14094: out = 1035;
			14095: out = 951;
			14096: out = -1924;
			14097: out = -1405;
			14098: out = 536;
			14099: out = 1521;
			14100: out = -503;
			14101: out = -1614;
			14102: out = 862;
			14103: out = -26;
			14104: out = 402;
			14105: out = 96;
			14106: out = 1333;
			14107: out = -405;
			14108: out = -651;
			14109: out = 478;
			14110: out = 234;
			14111: out = -28;
			14112: out = -117;
			14113: out = 21;
			14114: out = 225;
			14115: out = -80;
			14116: out = -350;
			14117: out = -328;
			14118: out = 285;
			14119: out = 168;
			14120: out = -199;
			14121: out = -2173;
			14122: out = -1608;
			14123: out = 1195;
			14124: out = 1113;
			14125: out = 7;
			14126: out = -1286;
			14127: out = -7;
			14128: out = 734;
			14129: out = 894;
			14130: out = -352;
			14131: out = 165;
			14132: out = 365;
			14133: out = 337;
			14134: out = -2472;
			14135: out = -466;
			14136: out = 906;
			14137: out = 1696;
			14138: out = 89;
			14139: out = -2;
			14140: out = -105;
			14141: out = -1524;
			14142: out = 118;
			14143: out = 872;
			14144: out = 471;
			14145: out = 295;
			14146: out = -585;
			14147: out = -640;
			14148: out = 667;
			14149: out = 534;
			14150: out = -170;
			14151: out = -1284;
			14152: out = -601;
			14153: out = -553;
			14154: out = -161;
			14155: out = 183;
			14156: out = 477;
			14157: out = -45;
			14158: out = -888;
			14159: out = 637;
			14160: out = 399;
			14161: out = -50;
			14162: out = -351;
			14163: out = 238;
			14164: out = 516;
			14165: out = 319;
			14166: out = -52;
			14167: out = 228;
			14168: out = 877;
			14169: out = 678;
			14170: out = 706;
			14171: out = -752;
			14172: out = -2019;
			14173: out = -1550;
			14174: out = -73;
			14175: out = 713;
			14176: out = 133;
			14177: out = -893;
			14178: out = -589;
			14179: out = 637;
			14180: out = -448;
			14181: out = 30;
			14182: out = 491;
			14183: out = 1354;
			14184: out = 142;
			14185: out = -451;
			14186: out = -797;
			14187: out = -2518;
			14188: out = -930;
			14189: out = 941;
			14190: out = 1880;
			14191: out = 937;
			14192: out = 442;
			14193: out = 380;
			14194: out = -61;
			14195: out = -898;
			14196: out = -1426;
			14197: out = -340;
			14198: out = -453;
			14199: out = 1131;
			14200: out = 1863;
			14201: out = -313;
			14202: out = -815;
			14203: out = -558;
			14204: out = 247;
			14205: out = 7;
			14206: out = -150;
			14207: out = 32;
			14208: out = 328;
			14209: out = 544;
			14210: out = 58;
			14211: out = -334;
			14212: out = -1705;
			14213: out = -482;
			14214: out = 781;
			14215: out = 233;
			14216: out = -1149;
			14217: out = -1048;
			14218: out = 1211;
			14219: out = 1187;
			14220: out = 474;
			14221: out = -893;
			14222: out = 191;
			14223: out = -303;
			14224: out = 262;
			14225: out = 566;
			14226: out = 563;
			14227: out = -121;
			14228: out = -252;
			14229: out = 346;
			14230: out = 554;
			14231: out = -538;
			14232: out = -2283;
			14233: out = 362;
			14234: out = 1417;
			14235: out = 1690;
			14236: out = 4;
			14237: out = 49;
			14238: out = -657;
			14239: out = -1109;
			14240: out = -284;
			14241: out = 587;
			14242: out = 643;
			14243: out = -32;
			14244: out = -1565;
			14245: out = -1446;
			14246: out = 256;
			14247: out = 41;
			14248: out = 174;
			14249: out = -127;
			14250: out = 227;
			14251: out = -114;
			14252: out = 111;
			14253: out = 17;
			14254: out = 213;
			14255: out = -156;
			14256: out = -26;
			14257: out = -273;
			14258: out = 1145;
			14259: out = 964;
			14260: out = 499;
			14261: out = -1811;
			14262: out = 471;
			14263: out = 1731;
			14264: out = -324;
			14265: out = -1314;
			14266: out = -1406;
			14267: out = -109;
			14268: out = -295;
			14269: out = 81;
			14270: out = 253;
			14271: out = 906;
			14272: out = 231;
			14273: out = -95;
			14274: out = -206;
			14275: out = -1245;
			14276: out = -70;
			14277: out = 131;
			14278: out = -1215;
			14279: out = -980;
			14280: out = -41;
			14281: out = 950;
			14282: out = 240;
			14283: out = -668;
			14284: out = -899;
			14285: out = 390;
			14286: out = 528;
			14287: out = 547;
			14288: out = -33;
			14289: out = -1060;
			14290: out = -459;
			14291: out = 115;
			14292: out = -201;
			14293: out = -678;
			14294: out = -572;
			14295: out = 344;
			14296: out = 983;
			14297: out = 979;
			14298: out = 39;
			14299: out = -1136;
			14300: out = -64;
			14301: out = 131;
			14302: out = -214;
			14303: out = 4;
			14304: out = -164;
			14305: out = 317;
			14306: out = 593;
			14307: out = 821;
			14308: out = -453;
			14309: out = -1359;
			14310: out = 32;
			14311: out = 609;
			14312: out = 768;
			14313: out = -57;
			14314: out = 85;
			14315: out = -72;
			14316: out = 374;
			14317: out = 975;
			14318: out = 878;
			14319: out = -5;
			14320: out = -957;
			14321: out = -1221;
			14322: out = -203;
			14323: out = 822;
			14324: out = 252;
			14325: out = 356;
			14326: out = -824;
			14327: out = -2150;
			14328: out = 1000;
			14329: out = 1454;
			14330: out = 687;
			14331: out = -1769;
			14332: out = -318;
			14333: out = 359;
			14334: out = 17;
			14335: out = -709;
			14336: out = -718;
			14337: out = -193;
			14338: out = -471;
			14339: out = 1175;
			14340: out = 1415;
			14341: out = 861;
			14342: out = -768;
			14343: out = -492;
			14344: out = 121;
			14345: out = 111;
			14346: out = -45;
			14347: out = -98;
			14348: out = 119;
			14349: out = -175;
			14350: out = 42;
			14351: out = 312;
			14352: out = 591;
			14353: out = 443;
			14354: out = 222;
			14355: out = 26;
			14356: out = -194;
			14357: out = -168;
			14358: out = -228;
			14359: out = -118;
			14360: out = -464;
			14361: out = 0;
			14362: out = 280;
			14363: out = -515;
			14364: out = -1449;
			14365: out = -932;
			14366: out = 1885;
			14367: out = 156;
			14368: out = -162;
			14369: out = -201;
			14370: out = -920;
			14371: out = -334;
			14372: out = 137;
			14373: out = 408;
			14374: out = -1131;
			14375: out = -904;
			14376: out = 273;
			14377: out = 273;
			14378: out = 575;
			14379: out = -4;
			14380: out = -874;
			14381: out = -253;
			14382: out = 70;
			14383: out = 93;
			14384: out = -16;
			14385: out = 579;
			14386: out = 465;
			14387: out = -1378;
			14388: out = 466;
			14389: out = -186;
			14390: out = -464;
			14391: out = -12;
			14392: out = 1271;
			14393: out = 903;
			14394: out = -485;
			14395: out = -915;
			14396: out = 67;
			14397: out = 834;
			14398: out = 139;
			14399: out = -1575;
			14400: out = -1756;
			14401: out = 48;
			14402: out = 1866;
			14403: out = 1693;
			14404: out = 454;
			14405: out = 266;
			14406: out = -88;
			14407: out = -638;
			14408: out = -1731;
			14409: out = -457;
			14410: out = 180;
			14411: out = 861;
			14412: out = 1188;
			14413: out = 316;
			14414: out = -649;
			14415: out = -1059;
			14416: out = -141;
			14417: out = -52;
			14418: out = -141;
			14419: out = -126;
			14420: out = 783;
			14421: out = 744;
			14422: out = -257;
			14423: out = -21;
			14424: out = -375;
			14425: out = -258;
			14426: out = -77;
			14427: out = -25;
			14428: out = -7;
			14429: out = 171;
			14430: out = -850;
			14431: out = -422;
			14432: out = -186;
			14433: out = -859;
			14434: out = 110;
			14435: out = 922;
			14436: out = 1434;
			14437: out = 655;
			14438: out = 315;
			14439: out = 92;
			14440: out = 153;
			14441: out = -296;
			14442: out = -450;
			14443: out = -331;
			14444: out = -133;
			14445: out = 587;
			14446: out = 981;
			14447: out = 209;
			14448: out = 642;
			14449: out = 4;
			14450: out = -803;
			14451: out = -1130;
			14452: out = -617;
			14453: out = 211;
			14454: out = 751;
			14455: out = 262;
			14456: out = -428;
			14457: out = -898;
			14458: out = -383;
			14459: out = -416;
			14460: out = -149;
			14461: out = 430;
			14462: out = 576;
			14463: out = 189;
			14464: out = -560;
			14465: out = -527;
			14466: out = -870;
			14467: out = -536;
			14468: out = 219;
			14469: out = 187;
			14470: out = 157;
			14471: out = 11;
			14472: out = -601;
			14473: out = -251;
			14474: out = 204;
			14475: out = 611;
			14476: out = 76;
			14477: out = -541;
			14478: out = -1072;
			14479: out = 304;
			14480: out = -416;
			14481: out = -396;
			14482: out = -14;
			14483: out = 816;
			14484: out = 51;
			14485: out = -1019;
			14486: out = -796;
			14487: out = -290;
			14488: out = 51;
			14489: out = -159;
			14490: out = -972;
			14491: out = -366;
			14492: out = 663;
			14493: out = 109;
			14494: out = 488;
			14495: out = 222;
			14496: out = 6;
			14497: out = 89;
			14498: out = 313;
			14499: out = 426;
			14500: out = 155;
			14501: out = 545;
			14502: out = 440;
			14503: out = -157;
			14504: out = -294;
			14505: out = -451;
			14506: out = -217;
			14507: out = 171;
			14508: out = 240;
			14509: out = -176;
			14510: out = -918;
			14511: out = -13;
			14512: out = -475;
			14513: out = -735;
			14514: out = 209;
			14515: out = 91;
			14516: out = 200;
			14517: out = 251;
			14518: out = 805;
			14519: out = 673;
			14520: out = -8;
			14521: out = -1409;
			14522: out = -823;
			14523: out = -197;
			14524: out = 243;
			14525: out = 8;
			14526: out = -354;
			14527: out = -195;
			14528: out = 2069;
			14529: out = 153;
			14530: out = -98;
			14531: out = -26;
			14532: out = 1310;
			14533: out = 39;
			14534: out = -560;
			14535: out = 187;
			14536: out = 932;
			14537: out = 157;
			14538: out = -1295;
			14539: out = -405;
			14540: out = 484;
			14541: out = 921;
			14542: out = -230;
			14543: out = 92;
			14544: out = 171;
			14545: out = 296;
			14546: out = -330;
			14547: out = -1554;
			14548: out = -2024;
			14549: out = -336;
			14550: out = -356;
			14551: out = 106;
			14552: out = 23;
			14553: out = 1990;
			14554: out = 165;
			14555: out = -747;
			14556: out = -289;
			14557: out = 31;
			14558: out = -180;
			14559: out = -658;
			14560: out = -341;
			14561: out = 446;
			14562: out = 729;
			14563: out = -275;
			14564: out = 616;
			14565: out = 655;
			14566: out = 680;
			14567: out = -1267;
			14568: out = 157;
			14569: out = 415;
			14570: out = -472;
			14571: out = -407;
			14572: out = 119;
			14573: out = 642;
			14574: out = 116;
			14575: out = -19;
			14576: out = -405;
			14577: out = -893;
			14578: out = 102;
			14579: out = 28;
			14580: out = -235;
			14581: out = -925;
			14582: out = 444;
			14583: out = 540;
			14584: out = -508;
			14585: out = -543;
			14586: out = 103;
			14587: out = 1098;
			14588: out = 1093;
			14589: out = 415;
			14590: out = -927;
			14591: out = -2092;
			14592: out = -68;
			14593: out = 173;
			14594: out = 192;
			14595: out = 633;
			14596: out = 1087;
			14597: out = 778;
			14598: out = -218;
			14599: out = 160;
			14600: out = -480;
			14601: out = -917;
			14602: out = -509;
			14603: out = -1451;
			14604: out = -961;
			14605: out = 444;
			14606: out = 535;
			14607: out = 302;
			14608: out = -276;
			14609: out = 17;
			14610: out = -209;
			14611: out = 72;
			14612: out = 31;
			14613: out = 230;
			14614: out = -387;
			14615: out = -389;
			14616: out = 198;
			14617: out = 1201;
			14618: out = 1072;
			14619: out = 130;
			14620: out = -708;
			14621: out = -543;
			14622: out = 187;
			14623: out = 553;
			14624: out = 792;
			14625: out = 488;
			14626: out = -60;
			14627: out = -73;
			14628: out = -542;
			14629: out = -328;
			14630: out = 614;
			14631: out = 735;
			14632: out = 483;
			14633: out = -154;
			14634: out = -1067;
			14635: out = -584;
			14636: out = 25;
			14637: out = 0;
			14638: out = -5;
			14639: out = -58;
			14640: out = 109;
			14641: out = -141;
			14642: out = 124;
			14643: out = -125;
			14644: out = -873;
			14645: out = -79;
			14646: out = 135;
			14647: out = 104;
			14648: out = 608;
			14649: out = 485;
			14650: out = 845;
			14651: out = 1482;
			14652: out = 544;
			14653: out = -454;
			14654: out = -1176;
			14655: out = 102;
			14656: out = -502;
			14657: out = -514;
			14658: out = -55;
			14659: out = 453;
			14660: out = 229;
			14661: out = -244;
			14662: out = 388;
			14663: out = -42;
			14664: out = -123;
			14665: out = -142;
			14666: out = 103;
			14667: out = -153;
			14668: out = -634;
			14669: out = -1625;
			14670: out = -859;
			14671: out = 235;
			14672: out = 1195;
			14673: out = 34;
			14674: out = -38;
			14675: out = 137;
			14676: out = -221;
			14677: out = -75;
			14678: out = -208;
			14679: out = -387;
			14680: out = -207;
			14681: out = -53;
			14682: out = 73;
			14683: out = -99;
			14684: out = 42;
			14685: out = 74;
			14686: out = 169;
			14687: out = 18;
			14688: out = 117;
			14689: out = -295;
			14690: out = -1619;
			14691: out = -1665;
			14692: out = -944;
			14693: out = 481;
			14694: out = 1366;
			14695: out = 1338;
			14696: out = 190;
			14697: out = -962;
			14698: out = -1675;
			14699: out = -626;
			14700: out = 948;
			14701: out = 136;
			14702: out = -63;
			14703: out = -51;
			14704: out = 174;
			14705: out = 687;
			14706: out = 485;
			14707: out = -242;
			14708: out = 119;
			14709: out = 29;
			14710: out = 197;
			14711: out = 600;
			14712: out = -383;
			14713: out = -471;
			14714: out = 248;
			14715: out = 8;
			14716: out = 833;
			14717: out = 1015;
			14718: out = 236;
			14719: out = -197;
			14720: out = -713;
			14721: out = -834;
			14722: out = -709;
			14723: out = -159;
			14724: out = 97;
			14725: out = 61;
			14726: out = -308;
			14727: out = -205;
			14728: out = 228;
			14729: out = -141;
			14730: out = 500;
			14731: out = 628;
			14732: out = -301;
			14733: out = 376;
			14734: out = -114;
			14735: out = -626;
			14736: out = 25;
			14737: out = 409;
			14738: out = 463;
			14739: out = -5;
			14740: out = 35;
			14741: out = -12;
			14742: out = -153;
			14743: out = -42;
			14744: out = -967;
			14745: out = -1149;
			14746: out = 64;
			14747: out = 515;
			14748: out = 865;
			14749: out = 258;
			14750: out = 113;
			14751: out = -1481;
			14752: out = -1074;
			14753: out = 1222;
			14754: out = 521;
			14755: out = 358;
			14756: out = -52;
			14757: out = 208;
			14758: out = -161;
			14759: out = -80;
			14760: out = -10;
			14761: out = 119;
			14762: out = -472;
			14763: out = -675;
			14764: out = 1019;
			14765: out = 167;
			14766: out = -384;
			14767: out = -354;
			14768: out = -702;
			14769: out = -226;
			14770: out = 142;
			14771: out = 384;
			14772: out = 66;
			14773: out = 375;
			14774: out = 968;
			14775: out = 596;
			14776: out = -134;
			14777: out = -749;
			14778: out = -358;
			14779: out = -247;
			14780: out = 97;
			14781: out = 295;
			14782: out = -372;
			14783: out = -46;
			14784: out = 470;
			14785: out = 459;
			14786: out = 262;
			14787: out = -172;
			14788: out = -472;
			14789: out = -889;
			14790: out = -396;
			14791: out = 204;
			14792: out = 16;
			14793: out = 386;
			14794: out = -95;
			14795: out = -637;
			14796: out = -49;
			14797: out = 628;
			14798: out = 777;
			14799: out = -207;
			14800: out = 39;
			14801: out = -339;
			14802: out = -967;
			14803: out = -103;
			14804: out = -672;
			14805: out = -690;
			14806: out = -161;
			14807: out = 1122;
			14808: out = 794;
			14809: out = -395;
			14810: out = -326;
			14811: out = -318;
			14812: out = -129;
			14813: out = -160;
			14814: out = 3;
			14815: out = 617;
			14816: out = 1019;
			14817: out = -361;
			14818: out = -1046;
			14819: out = -1383;
			14820: out = -987;
			14821: out = -290;
			14822: out = 321;
			14823: out = 527;
			14824: out = -138;
			14825: out = -279;
			14826: out = -335;
			14827: out = 214;
			14828: out = -457;
			14829: out = 283;
			14830: out = 664;
			14831: out = 312;
			14832: out = -1630;
			14833: out = -1796;
			14834: out = 491;
			14835: out = 1142;
			14836: out = 915;
			14837: out = -162;
			14838: out = 305;
			14839: out = 49;
			14840: out = 28;
			14841: out = -748;
			14842: out = -128;
			14843: out = -57;
			14844: out = 254;
			14845: out = -192;
			14846: out = 638;
			14847: out = 471;
			14848: out = -194;
			14849: out = -807;
			14850: out = 61;
			14851: out = 1083;
			14852: out = 203;
			14853: out = 720;
			14854: out = 406;
			14855: out = -283;
			14856: out = -744;
			14857: out = -588;
			14858: out = 26;
			14859: out = -225;
			14860: out = 546;
			14861: out = -125;
			14862: out = -1389;
			14863: out = -1580;
			14864: out = -288;
			14865: out = 1073;
			14866: out = 841;
			14867: out = 232;
			14868: out = -304;
			14869: out = -59;
			14870: out = -625;
			14871: out = -251;
			14872: out = 89;
			14873: out = 567;
			14874: out = 270;
			14875: out = 8;
			14876: out = -83;
			14877: out = 451;
			14878: out = 919;
			14879: out = 863;
			14880: out = -476;
			14881: out = -553;
			14882: out = -430;
			14883: out = 284;
			14884: out = -320;
			14885: out = 706;
			14886: out = 716;
			14887: out = -1174;
			14888: out = -746;
			14889: out = -58;
			14890: out = 744;
			14891: out = -792;
			14892: out = -602;
			14893: out = -222;
			14894: out = -89;
			14895: out = 76;
			14896: out = -42;
			14897: out = -89;
			14898: out = 317;
			14899: out = 245;
			14900: out = -135;
			14901: out = -313;
			14902: out = -1021;
			14903: out = -363;
			14904: out = 675;
			14905: out = 67;
			14906: out = -39;
			14907: out = 248;
			14908: out = 1350;
			14909: out = -372;
			14910: out = -1504;
			14911: out = -1782;
			14912: out = 272;
			14913: out = 606;
			14914: out = 264;
			14915: out = -608;
			14916: out = -1133;
			14917: out = -1006;
			14918: out = -219;
			14919: out = 904;
			14920: out = 718;
			14921: out = -20;
			14922: out = -747;
			14923: out = -157;
			14924: out = 99;
			14925: out = 190;
			14926: out = 803;
			14927: out = 503;
			14928: out = 268;
			14929: out = 161;
			14930: out = 94;
			14931: out = 64;
			14932: out = 106;
			14933: out = 358;
			14934: out = 192;
			14935: out = 158;
			14936: out = 331;
			14937: out = -683;
			14938: out = -796;
			14939: out = -529;
			14940: out = -660;
			14941: out = -14;
			14942: out = 199;
			14943: out = 152;
			14944: out = -93;
			14945: out = -50;
			14946: out = 99;
			14947: out = -55;
			14948: out = -115;
			14949: out = -44;
			14950: out = 155;
			14951: out = -481;
			14952: out = -743;
			14953: out = -617;
			14954: out = 436;
			14955: out = 222;
			14956: out = 168;
			14957: out = 215;
			14958: out = 1075;
			14959: out = 1010;
			14960: out = 403;
			14961: out = -874;
			14962: out = -682;
			14963: out = -439;
			14964: out = -46;
			14965: out = 42;
			14966: out = 778;
			14967: out = 808;
			14968: out = -1187;
			14969: out = -282;
			14970: out = 56;
			14971: out = 96;
			14972: out = -522;
			14973: out = -394;
			14974: out = -37;
			14975: out = -193;
			14976: out = 910;
			14977: out = 1130;
			14978: out = 762;
			14979: out = -522;
			14980: out = -251;
			14981: out = 190;
			14982: out = -194;
			14983: out = -251;
			14984: out = -575;
			14985: out = -470;
			14986: out = 247;
			14987: out = 539;
			14988: out = 303;
			14989: out = -426;
			14990: out = -585;
			14991: out = -440;
			14992: out = -90;
			14993: out = -196;
			14994: out = 191;
			14995: out = 427;
			14996: out = 519;
			14997: out = -741;
			14998: out = -1137;
			14999: out = -518;
			15000: out = 178;
			15001: out = 1155;
			15002: out = 782;
			15003: out = -965;
			15004: out = -1019;
			15005: out = -569;
			15006: out = 381;
			15007: out = 21;
			15008: out = 305;
			15009: out = -52;
			15010: out = -12;
			15011: out = -711;
			15012: out = 267;
			15013: out = 968;
			15014: out = 850;
			15015: out = -710;
			15016: out = -1230;
			15017: out = -426;
			15018: out = 1551;
			15019: out = 1130;
			15020: out = -434;
			15021: out = -1473;
			15022: out = -187;
			15023: out = 716;
			15024: out = -70;
			15025: out = 210;
			15026: out = 105;
			15027: out = 282;
			15028: out = -1211;
			15029: out = -471;
			15030: out = -229;
			15031: out = 234;
			15032: out = -1260;
			15033: out = -353;
			15034: out = 529;
			15035: out = 578;
			15036: out = -396;
			15037: out = -661;
			15038: out = 20;
			15039: out = 24;
			15040: out = 178;
			15041: out = -82;
			15042: out = -1034;
			15043: out = 207;
			15044: out = 568;
			15045: out = 65;
			15046: out = -221;
			15047: out = -140;
			15048: out = 205;
			15049: out = 60;
			15050: out = 26;
			15051: out = 151;
			15052: out = 567;
			15053: out = -932;
			15054: out = -549;
			15055: out = 137;
			15056: out = 332;
			15057: out = 850;
			15058: out = 958;
			15059: out = 716;
			15060: out = -2019;
			15061: out = -1552;
			15062: out = -198;
			15063: out = 732;
			15064: out = 174;
			15065: out = -201;
			15066: out = 122;
			15067: out = 245;
			15068: out = 709;
			15069: out = 506;
			15070: out = -104;
			15071: out = -373;
			15072: out = 48;
			15073: out = 535;
			15074: out = -516;
			15075: out = -505;
			15076: out = 109;
			15077: out = 1326;
			15078: out = 534;
			15079: out = -12;
			15080: out = -485;
			15081: out = -1225;
			15082: out = -749;
			15083: out = -33;
			15084: out = 352;
			15085: out = 45;
			15086: out = -33;
			15087: out = 148;
			15088: out = 129;
			15089: out = 14;
			15090: out = -195;
			15091: out = -51;
			15092: out = 42;
			15093: out = 130;
			15094: out = -196;
			15095: out = 699;
			15096: out = -587;
			15097: out = -784;
			15098: out = 188;
			15099: out = 1425;
			15100: out = 940;
			15101: out = -389;
			15102: out = -467;
			15103: out = -325;
			15104: out = -130;
			15105: out = -906;
			15106: out = 303;
			15107: out = 122;
			15108: out = 12;
			15109: out = 506;
			15110: out = 540;
			15111: out = 551;
			15112: out = 688;
			15113: out = -1;
			15114: out = -379;
			15115: out = -642;
			15116: out = -326;
			15117: out = -143;
			15118: out = 96;
			15119: out = -308;
			15120: out = 74;
			15121: out = -694;
			15122: out = -966;
			15123: out = -922;
			15124: out = 711;
			15125: out = 778;
			15126: out = -266;
			15127: out = -1639;
			15128: out = -250;
			15129: out = 1201;
			15130: out = -744;
			15131: out = -482;
			15132: out = -127;
			15133: out = 1144;
			15134: out = 470;
			15135: out = 444;
			15136: out = -192;
			15137: out = -952;
			15138: out = -630;
			15139: out = -28;
			15140: out = -8;
			15141: out = 113;
			15142: out = -560;
			15143: out = -418;
			15144: out = 958;
			15145: out = 878;
			15146: out = 122;
			15147: out = -823;
			15148: out = -115;
			15149: out = 345;
			15150: out = 210;
			15151: out = -1569;
			15152: out = -442;
			15153: out = 444;
			15154: out = 1184;
			15155: out = 337;
			15156: out = 255;
			15157: out = 50;
			15158: out = 128;
			15159: out = -682;
			15160: out = -455;
			15161: out = 276;
			15162: out = 501;
			15163: out = 228;
			15164: out = -323;
			15165: out = -748;
			15166: out = 516;
			15167: out = 1091;
			15168: out = 628;
			15169: out = -402;
			15170: out = -1144;
			15171: out = -1083;
			15172: out = -552;
			15173: out = -8;
			15174: out = 65;
			15175: out = -69;
			15176: out = -357;
			15177: out = 574;
			15178: out = 1115;
			15179: out = 131;
			15180: out = -46;
			15181: out = -1043;
			15182: out = -1263;
			15183: out = 24;
			15184: out = 1012;
			15185: out = 969;
			15186: out = -236;
			15187: out = -60;
			15188: out = 183;
			15189: out = 525;
			15190: out = -94;
			15191: out = 0;
			15192: out = 138;
			15193: out = 296;
			15194: out = -407;
			15195: out = -990;
			15196: out = -1048;
			15197: out = 328;
			15198: out = 1080;
			15199: out = 1348;
			15200: out = 478;
			15201: out = 299;
			15202: out = -877;
			15203: out = -1404;
			15204: out = -85;
			15205: out = -59;
			15206: out = -3;
			15207: out = 397;
			15208: out = -166;
			15209: out = -204;
			15210: out = -363;
			15211: out = 716;
			15212: out = -1359;
			15213: out = -1649;
			15214: out = -342;
			15215: out = 825;
			15216: out = -196;
			15217: out = -1562;
			15218: out = 232;
			15219: out = -235;
			15220: out = 257;
			15221: out = 504;
			15222: out = 299;
			15223: out = -139;
			15224: out = -360;
			15225: out = -539;
			15226: out = -59;
			15227: out = 324;
			15228: out = 567;
			15229: out = 216;
			15230: out = 17;
			15231: out = -110;
			15232: out = 114;
			15233: out = -388;
			15234: out = -654;
			15235: out = -661;
			15236: out = 303;
			15237: out = 213;
			15238: out = -117;
			15239: out = -42;
			15240: out = -54;
			15241: out = -155;
			15242: out = -499;
			15243: out = 1145;
			15244: out = 198;
			15245: out = -843;
			15246: out = -1140;
			15247: out = 167;
			15248: out = 537;
			15249: out = -294;
			15250: out = 163;
			15251: out = -324;
			15252: out = -64;
			15253: out = 110;
			15254: out = 1504;
			15255: out = 853;
			15256: out = -582;
			15257: out = -912;
			15258: out = -471;
			15259: out = 327;
			15260: out = 933;
			15261: out = 252;
			15262: out = 72;
			15263: out = 121;
			15264: out = -298;
			15265: out = -538;
			15266: out = -185;
			15267: out = 751;
			15268: out = 649;
			15269: out = -182;
			15270: out = -1001;
			15271: out = 165;
			15272: out = 520;
			15273: out = 621;
			15274: out = -41;
			15275: out = -430;
			15276: out = -332;
			15277: out = 362;
			15278: out = 583;
			15279: out = 721;
			15280: out = -13;
			15281: out = -1033;
			15282: out = -323;
			15283: out = 250;
			15284: out = 482;
			15285: out = 123;
			15286: out = 113;
			15287: out = -7;
			15288: out = -393;
			15289: out = 760;
			15290: out = 626;
			15291: out = 221;
			15292: out = 516;
			15293: out = -373;
			15294: out = -1337;
			15295: out = -1870;
			15296: out = -438;
			15297: out = 960;
			15298: out = 1264;
			15299: out = -802;
			15300: out = -1092;
			15301: out = -844;
			15302: out = 269;
			15303: out = -1536;
			15304: out = -871;
			15305: out = 334;
			15306: out = 1207;
			15307: out = 531;
			15308: out = -224;
			15309: out = -204;
			15310: out = -265;
			15311: out = 637;
			15312: out = 947;
			15313: out = 69;
			15314: out = -577;
			15315: out = -535;
			15316: out = 179;
			15317: out = -159;
			15318: out = 163;
			15319: out = 341;
			15320: out = 97;
			15321: out = 35;
			15322: out = -203;
			15323: out = -327;
			15324: out = -997;
			15325: out = -205;
			15326: out = 456;
			15327: out = 87;
			15328: out = -143;
			15329: out = -382;
			15330: out = -168;
			15331: out = 785;
			15332: out = 668;
			15333: out = 72;
			15334: out = -280;
			15335: out = -230;
			15336: out = -37;
			15337: out = -98;
			15338: out = 194;
			15339: out = -62;
			15340: out = -32;
			15341: out = 99;
			15342: out = 214;
			15343: out = -190;
			15344: out = -490;
			15345: out = -156;
			15346: out = 801;
			15347: out = 917;
			15348: out = -695;
			15349: out = -340;
			15350: out = -244;
			15351: out = -20;
			15352: out = -367;
			15353: out = -140;
			15354: out = 11;
			15355: out = 135;
			15356: out = -8;
			15357: out = -187;
			15358: out = -275;
			15359: out = 117;
			15360: out = 49;
			15361: out = -111;
			15362: out = -18;
			15363: out = -315;
			15364: out = -176;
			15365: out = 68;
			15366: out = 1095;
			15367: out = 124;
			15368: out = -337;
			15369: out = 229;
			15370: out = 396;
			15371: out = 308;
			15372: out = -312;
			15373: out = -1110;
			15374: out = -991;
			15375: out = -297;
			15376: out = 566;
			15377: out = -17;
			15378: out = -109;
			15379: out = -15;
			15380: out = 76;
			15381: out = -200;
			15382: out = -295;
			15383: out = -15;
			15384: out = -120;
			15385: out = -107;
			15386: out = -137;
			15387: out = -122;
			15388: out = 307;
			15389: out = 770;
			15390: out = 983;
			15391: out = -490;
			15392: out = -1035;
			15393: out = -790;
			15394: out = -95;
			15395: out = 143;
			15396: out = 68;
			15397: out = -39;
			15398: out = 69;
			15399: out = -16;
			15400: out = -24;
			15401: out = 977;
			15402: out = -24;
			15403: out = -426;
			15404: out = -244;
			15405: out = 941;
			15406: out = 638;
			15407: out = -121;
			15408: out = -284;
			15409: out = -227;
			15410: out = 58;
			15411: out = 88;
			15412: out = 514;
			15413: out = 150;
			15414: out = -383;
			15415: out = -1023;
			15416: out = -377;
			15417: out = -13;
			15418: out = -110;
			15419: out = -36;
			15420: out = -100;
			15421: out = 0;
			15422: out = 22;
			15423: out = 190;
			15424: out = -313;
			15425: out = -980;
			15426: out = 274;
			15427: out = 410;
			15428: out = -102;
			15429: out = -1979;
			15430: out = -147;
			15431: out = 823;
			15432: out = 940;
			15433: out = -636;
			15434: out = -575;
			15435: out = -130;
			15436: out = 50;
			15437: out = 185;
			15438: out = 56;
			15439: out = -123;
			15440: out = -25;
			15441: out = -87;
			15442: out = -81;
			15443: out = -35;
			15444: out = 129;
			15445: out = 141;
			15446: out = 50;
			15447: out = -124;
			15448: out = 61;
			15449: out = 180;
			15450: out = 139;
			15451: out = -418;
			15452: out = -500;
			15453: out = -206;
			15454: out = 51;
			15455: out = 114;
			15456: out = 134;
			15457: out = 376;
			15458: out = -228;
			15459: out = -226;
			15460: out = -4;
			15461: out = -371;
			15462: out = 416;
			15463: out = 545;
			15464: out = -442;
			15465: out = 124;
			15466: out = 532;
			15467: out = 980;
			15468: out = -1409;
			15469: out = 365;
			15470: out = 665;
			15471: out = -180;
			15472: out = -2153;
			15473: out = -1174;
			15474: out = 848;
			15475: out = 710;
			15476: out = 523;
			15477: out = -372;
			15478: out = -652;
			15479: out = -635;
			15480: out = -200;
			15481: out = 164;
			15482: out = 1321;
			15483: out = 267;
			15484: out = -462;
			15485: out = -903;
			15486: out = 411;
			15487: out = 466;
			15488: out = 339;
			15489: out = 529;
			15490: out = 222;
			15491: out = -83;
			15492: out = -78;
			15493: out = -223;
			15494: out = 300;
			15495: out = 404;
			15496: out = 121;
			15497: out = -651;
			15498: out = -238;
			15499: out = 755;
			15500: out = 373;
			15501: out = -542;
			15502: out = -1085;
			15503: out = 253;
			15504: out = -66;
			15505: out = -407;
			15506: out = -970;
			15507: out = 145;
			15508: out = 20;
			15509: out = -96;
			15510: out = 216;
			15511: out = -97;
			15512: out = 140;
			15513: out = 519;
			15514: out = 205;
			15515: out = -388;
			15516: out = -698;
			15517: out = -256;
			15518: out = 723;
			15519: out = 976;
			15520: out = 263;
			15521: out = -160;
			15522: out = -809;
			15523: out = -827;
			15524: out = -509;
			15525: out = 184;
			15526: out = 397;
			15527: out = 249;
			15528: out = -487;
			15529: out = 67;
			15530: out = 672;
			15531: out = 384;
			15532: out = 930;
			15533: out = 39;
			15534: out = -1071;
			15535: out = -308;
			15536: out = 242;
			15537: out = 846;
			15538: out = 490;
			15539: out = 533;
			15540: out = -589;
			15541: out = -1346;
			15542: out = -432;
			15543: out = 414;
			15544: out = 316;
			15545: out = -1067;
			15546: out = -920;
			15547: out = -597;
			15548: out = 90;
			15549: out = 449;
			15550: out = 474;
			15551: out = 115;
			15552: out = -315;
			15553: out = -145;
			15554: out = -68;
			15555: out = -10;
			15556: out = 64;
			15557: out = 115;
			15558: out = -113;
			15559: out = -492;
			15560: out = 13;
			15561: out = 471;
			15562: out = 590;
			15563: out = -21;
			15564: out = -531;
			15565: out = -593;
			15566: out = -40;
			15567: out = 14;
			15568: out = 152;
			15569: out = 120;
			15570: out = 80;
			15571: out = 140;
			15572: out = -108;
			15573: out = -804;
			15574: out = 34;
			15575: out = 7;
			15576: out = -246;
			15577: out = -940;
			15578: out = -192;
			15579: out = 618;
			15580: out = 1198;
			15581: out = 97;
			15582: out = -344;
			15583: out = -504;
			15584: out = -67;
			15585: out = -92;
			15586: out = 64;
			15587: out = 91;
			15588: out = 45;
			15589: out = -175;
			15590: out = 160;
			15591: out = 765;
			15592: out = 1141;
			15593: out = 165;
			15594: out = -1279;
			15595: out = -1254;
			15596: out = 96;
			15597: out = 1086;
			15598: out = -76;
			15599: out = -321;
			15600: out = -420;
			15601: out = 222;
			15602: out = 209;
			15603: out = 284;
			15604: out = -81;
			15605: out = -62;
			15606: out = -687;
			15607: out = -432;
			15608: out = 168;
			15609: out = 90;
			15610: out = 574;
			15611: out = 774;
			15612: out = -57;
			15613: out = 190;
			15614: out = 5;
			15615: out = 158;
			15616: out = -873;
			15617: out = 751;
			15618: out = 1564;
			15619: out = 252;
			15620: out = -586;
			15621: out = -1208;
			15622: out = -725;
			15623: out = -155;
			15624: out = 671;
			15625: out = 592;
			15626: out = -120;
			15627: out = -494;
			15628: out = -368;
			15629: out = -29;
			15630: out = -109;
			15631: out = -208;
			15632: out = -484;
			15633: out = -719;
			15634: out = -259;
			15635: out = 126;
			15636: out = 259;
			15637: out = -288;
			15638: out = -472;
			15639: out = -322;
			15640: out = 408;
			15641: out = -435;
			15642: out = -227;
			15643: out = 240;
			15644: out = 314;
			15645: out = 50;
			15646: out = -146;
			15647: out = -5;
			15648: out = 81;
			15649: out = 153;
			15650: out = 121;
			15651: out = 75;
			15652: out = -60;
			15653: out = -221;
			15654: out = -333;
			15655: out = -521;
			15656: out = -323;
			15657: out = -90;
			15658: out = -335;
			15659: out = 253;
			15660: out = 835;
			15661: out = 1082;
			15662: out = -403;
			15663: out = -1437;
			15664: out = -1509;
			15665: out = 179;
			15666: out = 817;
			15667: out = 793;
			15668: out = -204;
			15669: out = 413;
			15670: out = 39;
			15671: out = 20;
			15672: out = 36;
			15673: out = 528;
			15674: out = -25;
			15675: out = -1013;
			15676: out = -977;
			15677: out = -149;
			15678: out = 767;
			15679: out = 966;
			15680: out = 248;
			15681: out = -472;
			15682: out = -675;
			15683: out = -131;
			15684: out = -140;
			15685: out = -316;
			15686: out = 15;
			15687: out = -91;
			15688: out = -30;
			15689: out = -112;
			15690: out = 154;
			15691: out = 39;
			15692: out = -104;
			15693: out = -292;
			15694: out = -54;
			15695: out = 304;
			15696: out = 492;
			15697: out = 119;
			15698: out = -297;
			15699: out = -477;
			15700: out = 14;
			15701: out = 71;
			15702: out = 109;
			15703: out = -107;
			15704: out = 1044;
			15705: out = 349;
			15706: out = -366;
			15707: out = -1198;
			15708: out = -152;
			15709: out = 59;
			15710: out = -122;
			15711: out = -69;
			15712: out = 336;
			15713: out = 339;
			15714: out = -349;
			15715: out = -188;
			15716: out = 260;
			15717: out = 642;
			15718: out = 131;
			15719: out = -981;
			15720: out = -1583;
			15721: out = -717;
			15722: out = 167;
			15723: out = 955;
			15724: out = 839;
			15725: out = 59;
			15726: out = -406;
			15727: out = -594;
			15728: out = -949;
			15729: out = 197;
			15730: out = 294;
			15731: out = 38;
			15732: out = -20;
			15733: out = 193;
			15734: out = 401;
			15735: out = 271;
			15736: out = 177;
			15737: out = -341;
			15738: out = -643;
			15739: out = 365;
			15740: out = 301;
			15741: out = 261;
			15742: out = -140;
			15743: out = 241;
			15744: out = -461;
			15745: out = -847;
			15746: out = -38;
			15747: out = 609;
			15748: out = 707;
			15749: out = -4;
			15750: out = -564;
			15751: out = -710;
			15752: out = -387;
			15753: out = -332;
			15754: out = 47;
			15755: out = 359;
			15756: out = 711;
			15757: out = 508;
			15758: out = 221;
			15759: out = -63;
			15760: out = 559;
			15761: out = -164;
			15762: out = -89;
			15763: out = 548;
			15764: out = 31;
			15765: out = 201;
			15766: out = 140;
			15767: out = -771;
			15768: out = -97;
			15769: out = 130;
			15770: out = -152;
			15771: out = 111;
			15772: out = -409;
			15773: out = -631;
			15774: out = 105;
			15775: out = -254;
			15776: out = -255;
			15777: out = -61;
			15778: out = 89;
			15779: out = 157;
			15780: out = 141;
			15781: out = 327;
			15782: out = -54;
			15783: out = -136;
			15784: out = -134;
			15785: out = 146;
			15786: out = -151;
			15787: out = -269;
			15788: out = 73;
			15789: out = 59;
			15790: out = 63;
			15791: out = 176;
			15792: out = 214;
			15793: out = 655;
			15794: out = 624;
			15795: out = 55;
			15796: out = -876;
			15797: out = -1153;
			15798: out = -735;
			15799: out = 224;
			15800: out = 194;
			15801: out = 23;
			15802: out = 63;
			15803: out = 160;
			15804: out = -230;
			15805: out = -795;
			15806: out = -876;
			15807: out = -523;
			15808: out = -129;
			15809: out = 96;
			15810: out = -223;
			15811: out = -154;
			15812: out = 70;
			15813: out = 865;
			15814: out = 7;
			15815: out = -497;
			15816: out = 35;
			15817: out = 71;
			15818: out = -235;
			15819: out = -627;
			15820: out = 535;
			15821: out = 250;
			15822: out = -6;
			15823: out = -4;
			15824: out = 80;
			15825: out = 131;
			15826: out = -140;
			15827: out = 283;
			15828: out = -1065;
			15829: out = -1081;
			15830: out = 299;
			15831: out = 776;
			15832: out = 103;
			15833: out = -1029;
			15834: out = -359;
			15835: out = -88;
			15836: out = 185;
			15837: out = -331;
			15838: out = 1085;
			15839: out = 741;
			15840: out = -89;
			15841: out = -155;
			15842: out = -1289;
			15843: out = -809;
			15844: out = 1304;
			15845: out = 735;
			15846: out = 877;
			15847: out = 421;
			15848: out = 178;
			15849: out = -788;
			15850: out = -521;
			15851: out = 383;
			15852: out = 328;
			15853: out = -332;
			15854: out = -933;
			15855: out = -20;
			15856: out = -44;
			15857: out = 121;
			15858: out = -118;
			15859: out = 373;
			15860: out = -63;
			15861: out = -274;
			15862: out = 74;
			15863: out = 400;
			15864: out = 402;
			15865: out = 42;
			15866: out = -271;
			15867: out = -221;
			15868: out = 62;
			15869: out = 280;
			15870: out = 148;
			15871: out = -44;
			15872: out = -41;
			15873: out = 21;
			15874: out = 113;
			15875: out = 61;
			15876: out = -129;
			15877: out = -114;
			15878: out = 11;
			15879: out = 128;
			15880: out = 45;
			15881: out = 372;
			15882: out = 679;
			15883: out = 339;
			15884: out = 103;
			15885: out = -877;
			15886: out = -1467;
			15887: out = -236;
			15888: out = 946;
			15889: out = 1333;
			15890: out = 500;
			15891: out = -761;
			15892: out = -1369;
			15893: out = -875;
			15894: out = 139;
			15895: out = 349;
			15896: out = -397;
			15897: out = -1517;
			15898: out = -407;
			15899: out = 650;
			15900: out = 1080;
			15901: out = 125;
			15902: out = -601;
			15903: out = -876;
			15904: out = -165;
			15905: out = -90;
			15906: out = 392;
			15907: out = 390;
			15908: out = 232;
			15909: out = -624;
			15910: out = -836;
			15911: out = -424;
			15912: out = 829;
			15913: out = 649;
			15914: out = -80;
			15915: out = -5;
			15916: out = 69;
			15917: out = -243;
			15918: out = -1421;
			15919: out = -241;
			15920: out = 312;
			15921: out = 637;
			15922: out = -583;
			15923: out = 253;
			15924: out = 438;
			15925: out = 17;
			15926: out = -83;
			15927: out = -28;
			15928: out = -63;
			15929: out = -1140;
			15930: out = -273;
			15931: out = 298;
			15932: out = 284;
			15933: out = -15;
			15934: out = -32;
			15935: out = 252;
			15936: out = -9;
			15937: out = 235;
			15938: out = -87;
			15939: out = -272;
			15940: out = -1362;
			15941: out = -100;
			15942: out = 1005;
			15943: out = 419;
			15944: out = 243;
			15945: out = 7;
			15946: out = 91;
			15947: out = 100;
			15948: out = -357;
			15949: out = -615;
			15950: out = 18;
			15951: out = -24;
			15952: out = -117;
			15953: out = -280;
			15954: out = -495;
			15955: out = 289;
			15956: out = 900;
			15957: out = 403;
			15958: out = 124;
			15959: out = -119;
			15960: out = 15;
			15961: out = 281;
			15962: out = -209;
			15963: out = -698;
			15964: out = 232;
			15965: out = -156;
			15966: out = 338;
			15967: out = 576;
			15968: out = 574;
			15969: out = -305;
			15970: out = -649;
			15971: out = -297;
			15972: out = 374;
			15973: out = 172;
			15974: out = -316;
			15975: out = 44;
			15976: out = 865;
			15977: out = 994;
			15978: out = -265;
			15979: out = -464;
			15980: out = 32;
			15981: out = 1063;
			15982: out = 158;
			15983: out = 124;
			15984: out = -258;
			15985: out = -75;
			15986: out = -1074;
			15987: out = -581;
			15988: out = 224;
			15989: out = 240;
			15990: out = 42;
			15991: out = -336;
			15992: out = -696;
			15993: out = -81;
			15994: out = 52;
			15995: out = -92;
			15996: out = -52;
			15997: out = 15;
			15998: out = 48;
			15999: out = 32;
			16000: out = -104;
			16001: out = -29;
			16002: out = 130;
			16003: out = -160;
			16004: out = 270;
			16005: out = 365;
			16006: out = -193;
			16007: out = -336;
			16008: out = -818;
			16009: out = -686;
			16010: out = -44;
			16011: out = 912;
			16012: out = 499;
			16013: out = -1217;
			16014: out = 8;
			16015: out = 249;
			16016: out = 166;
			16017: out = -477;
			16018: out = -501;
			16019: out = -500;
			16020: out = -667;
			16021: out = 565;
			16022: out = 286;
			16023: out = -141;
			16024: out = -54;
			16025: out = 483;
			16026: out = 371;
			16027: out = -402;
			16028: out = -824;
			16029: out = -107;
			16030: out = 670;
			16031: out = -604;
			16032: out = -265;
			16033: out = -260;
			16034: out = 53;
			16035: out = -537;
			16036: out = 4;
			16037: out = 322;
			16038: out = -51;
			16039: out = -60;
			16040: out = -95;
			16041: out = -63;
			16042: out = 620;
			16043: out = 318;
			16044: out = -281;
			16045: out = -840;
			16046: out = -292;
			16047: out = 332;
			16048: out = 637;
			16049: out = 113;
			16050: out = 189;
			16051: out = 93;
			16052: out = -1164;
			16053: out = -237;
			16054: out = 259;
			16055: out = 596;
			16056: out = -1425;
			16057: out = -429;
			16058: out = 462;
			16059: out = -192;
			16060: out = -31;
			16061: out = -38;
			16062: out = 218;
			16063: out = -122;
			16064: out = 190;
			16065: out = 346;
			16066: out = 308;
			16067: out = 39;
			16068: out = -20;
			16069: out = 51;
			16070: out = -871;
			16071: out = -168;
			16072: out = 755;
			16073: out = 1676;
			16074: out = 90;
			16075: out = -551;
			16076: out = -452;
			16077: out = -723;
			16078: out = -254;
			16079: out = -109;
			16080: out = -723;
			16081: out = 203;
			16082: out = 260;
			16083: out = 129;
			16084: out = -142;
			16085: out = 318;
			16086: out = 432;
			16087: out = 276;
			16088: out = -873;
			16089: out = -721;
			16090: out = 199;
			16091: out = 1199;
			16092: out = 436;
			16093: out = -240;
			16094: out = -25;
			16095: out = 13;
			16096: out = 163;
			16097: out = 62;
			16098: out = 75;
			16099: out = 37;
			16100: out = -97;
			16101: out = -534;
			16102: out = 36;
			16103: out = 380;
			16104: out = 561;
			16105: out = -105;
			16106: out = -60;
			16107: out = -66;
			16108: out = 65;
			16109: out = -2;
			16110: out = 23;
			16111: out = -158;
			16112: out = -73;
			16113: out = -861;
			16114: out = -901;
			16115: out = -177;
			16116: out = -186;
			16117: out = 130;
			16118: out = 350;
			16119: out = 450;
			16120: out = 371;
			16121: out = 43;
			16122: out = -367;
			16123: out = -487;
			16124: out = -263;
			16125: out = -97;
			16126: out = -707;
			16127: out = -384;
			16128: out = -8;
			16129: out = 541;
			16130: out = -100;
			16131: out = 5;
			16132: out = 34;
			16133: out = -85;
			16134: out = -274;
			16135: out = -178;
			16136: out = -57;
			16137: out = -407;
			16138: out = -717;
			16139: out = -561;
			16140: out = 749;
			16141: out = 188;
			16142: out = 153;
			16143: out = 353;
			16144: out = 133;
			16145: out = 62;
			16146: out = -102;
			16147: out = -66;
			16148: out = -442;
			16149: out = -165;
			16150: out = 384;
			16151: out = 69;
			16152: out = 201;
			16153: out = 301;
			16154: out = 79;
			16155: out = 152;
			16156: out = -157;
			16157: out = -203;
			16158: out = 6;
			16159: out = 788;
			16160: out = 880;
			16161: out = -19;
			16162: out = -438;
			16163: out = -198;
			16164: out = 333;
			16165: out = 281;
			16166: out = -332;
			16167: out = -653;
			16168: out = -61;
			16169: out = 50;
			16170: out = -101;
			16171: out = -543;
			16172: out = -15;
			16173: out = -18;
			16174: out = 87;
			16175: out = -101;
			16176: out = 258;
			16177: out = 259;
			16178: out = 315;
			16179: out = 409;
			16180: out = 461;
			16181: out = 279;
			16182: out = 7;
			16183: out = -9;
			16184: out = 139;
			16185: out = 185;
			16186: out = -142;
			16187: out = -225;
			16188: out = 183;
			16189: out = 1059;
			16190: out = -165;
			16191: out = -631;
			16192: out = -628;
			16193: out = 69;
			16194: out = 38;
			16195: out = -164;
			16196: out = -558;
			16197: out = 337;
			16198: out = 271;
			16199: out = -43;
			16200: out = -332;
			16201: out = 52;
			16202: out = 257;
			16203: out = -23;
			16204: out = -57;
			16205: out = -615;
			16206: out = -873;
			16207: out = -312;
			16208: out = -151;
			16209: out = -10;
			16210: out = 48;
			16211: out = 271;
			16212: out = 91;
			16213: out = -242;
			16214: out = -838;
			16215: out = -316;
			16216: out = 258;
			16217: out = 548;
			16218: out = -186;
			16219: out = -370;
			16220: out = -240;
			16221: out = -352;
			16222: out = 113;
			16223: out = -290;
			16224: out = -1051;
			16225: out = -119;
			16226: out = 615;
			16227: out = 933;
			16228: out = -655;
			16229: out = 174;
			16230: out = -779;
			16231: out = -2207;
			16232: out = 630;
			16233: out = 978;
			16234: out = 670;
			16235: out = -314;
			16236: out = 0;
			16237: out = 80;
			16238: out = 95;
			16239: out = 447;
			16240: out = 141;
			16241: out = -208;
			16242: out = -41;
			16243: out = -616;
			16244: out = -269;
			16245: out = 369;
			16246: out = 108;
			16247: out = -8;
			16248: out = -28;
			16249: out = 499;
			16250: out = 20;
			16251: out = -167;
			16252: out = -304;
			16253: out = -89;
			16254: out = -120;
			16255: out = -123;
			16256: out = -325;
			16257: out = 230;
			16258: out = 212;
			16259: out = 152;
			16260: out = 407;
			16261: out = 164;
			16262: out = -181;
			16263: out = -42;
			16264: out = -973;
			16265: out = -623;
			16266: out = -3;
			16267: out = 161;
			16268: out = -170;
			16269: out = -67;
			16270: out = 468;
			16271: out = 1041;
			16272: out = 352;
			16273: out = -572;
			16274: out = -127;
			16275: out = 563;
			16276: out = 575;
			16277: out = -823;
			16278: out = -168;
			16279: out = 114;
			16280: out = 468;
			16281: out = 225;
			16282: out = -114;
			16283: out = -304;
			16284: out = 99;
			16285: out = 61;
			16286: out = -74;
			16287: out = -359;
			16288: out = -44;
			16289: out = -94;
			16290: out = -201;
			16291: out = -712;
			16292: out = -9;
			16293: out = 61;
			16294: out = 259;
			16295: out = 846;
			16296: out = 727;
			16297: out = 129;
			16298: out = -789;
			16299: out = -876;
			16300: out = -555;
			16301: out = 22;
			16302: out = -46;
			16303: out = 283;
			16304: out = 112;
			16305: out = -49;
			16306: out = -210;
			16307: out = 380;
			16308: out = 670;
			16309: out = 74;
			16310: out = -634;
			16311: out = -747;
			16312: out = -4;
			16313: out = -165;
			16314: out = 67;
			16315: out = -7;
			16316: out = 85;
			16317: out = 158;
			16318: out = 221;
			16319: out = -179;
			16320: out = 532;
			16321: out = -471;
			16322: out = -1189;
			16323: out = -1043;
			16324: out = 92;
			16325: out = 390;
			16326: out = -234;
			16327: out = 192;
			16328: out = -27;
			16329: out = 30;
			16330: out = 279;
			16331: out = 9;
			16332: out = -35;
			16333: out = 28;
			16334: out = -476;
			16335: out = -294;
			16336: out = 1;
			16337: out = 94;
			16338: out = 550;
			16339: out = 342;
			16340: out = -206;
			16341: out = -826;
			16342: out = -391;
			16343: out = -88;
			16344: out = -974;
			16345: out = -9;
			16346: out = -62;
			16347: out = -239;
			16348: out = -69;
			16349: out = 416;
			16350: out = 515;
			16351: out = -184;
			16352: out = 93;
			16353: out = -9;
			16354: out = 20;
			16355: out = 434;
			16356: out = 189;
			16357: out = -259;
			16358: out = -425;
			16359: out = -543;
			16360: out = -78;
			16361: out = 313;
			16362: out = -41;
			16363: out = 46;
			16364: out = 218;
			16365: out = 239;
			16366: out = 174;
			16367: out = -350;
			16368: out = -603;
			16369: out = -142;
			16370: out = 328;
			16371: out = 316;
			16372: out = -157;
			16373: out = -291;
			16374: out = 80;
			16375: out = 473;
			16376: out = 88;
			16377: out = -43;
			16378: out = -79;
			16379: out = 72;
			16380: out = 258;
			16381: out = 78;
			16382: out = -203;
			16383: out = -512;
			16384: out = 84;
			16385: out = 217;
			16386: out = -71;
			16387: out = 227;
			16388: out = 407;
			16389: out = 208;
			16390: out = -624;
			16391: out = -1178;
			16392: out = -789;
			16393: out = 279;
			16394: out = 416;
			16395: out = 117;
			16396: out = -472;
			16397: out = -771;
			16398: out = -135;
			16399: out = 310;
			16400: out = 246;
			16401: out = 169;
			16402: out = 216;
			16403: out = 231;
			16404: out = -109;
			16405: out = -394;
			16406: out = -154;
			16407: out = 538;
			16408: out = 99;
			16409: out = 30;
			16410: out = -142;
			16411: out = 111;
			16412: out = -115;
			16413: out = -40;
			16414: out = 66;
			16415: out = 138;
			16416: out = 76;
			16417: out = 234;
			16418: out = 546;
			16419: out = 88;
			16420: out = -504;
			16421: out = -742;
			16422: out = 21;
			16423: out = 539;
			16424: out = 595;
			16425: out = 1;
			16426: out = -376;
			16427: out = -353;
			16428: out = 6;
			16429: out = -111;
			16430: out = 47;
			16431: out = 66;
			16432: out = 294;
			16433: out = -505;
			16434: out = -389;
			16435: out = 233;
			16436: out = -34;
			16437: out = 250;
			16438: out = 215;
			16439: out = 288;
			16440: out = -693;
			16441: out = -565;
			16442: out = -18;
			16443: out = 22;
			16444: out = -159;
			16445: out = -179;
			16446: out = 347;
			16447: out = 360;
			16448: out = 323;
			16449: out = -97;
			16450: out = -732;
			16451: out = -824;
			16452: out = -155;
			16453: out = 933;
			16454: out = 89;
			16455: out = -230;
			16456: out = -211;
			16457: out = 272;
			16458: out = 53;
			16459: out = -202;
			16460: out = -470;
			16461: out = 37;
			16462: out = 46;
			16463: out = -199;
			16464: out = -438;
			16465: out = -199;
			16466: out = 19;
			16467: out = -122;
			16468: out = 398;
			16469: out = 288;
			16470: out = 58;
			16471: out = 73;
			16472: out = -179;
			16473: out = -418;
			16474: out = -617;
			16475: out = -149;
			16476: out = -149;
			16477: out = -250;
			16478: out = 194;
			16479: out = -75;
			16480: out = 140;
			16481: out = 622;
			16482: out = 156;
			16483: out = 63;
			16484: out = 34;
			16485: out = -153;
			16486: out = 34;
			16487: out = -16;
			16488: out = -138;
			16489: out = -644;
			16490: out = -144;
			16491: out = 365;
			16492: out = 55;
			16493: out = 274;
			16494: out = 173;
			16495: out = 24;
			16496: out = -101;
			16497: out = -102;
			16498: out = -29;
			16499: out = -120;
			16500: out = 17;
			16501: out = -444;
			16502: out = -959;
			16503: out = -5;
			16504: out = 642;
			16505: out = 710;
			16506: out = -346;
			16507: out = -95;
			16508: out = -43;
			16509: out = -52;
			16510: out = 277;
			16511: out = 153;
			16512: out = -217;
			16513: out = -1252;
			16514: out = 770;
			16515: out = 1461;
			16516: out = 1010;
			16517: out = -529;
			16518: out = -536;
			16519: out = -311;
			16520: out = -701;
			16521: out = -235;
			16522: out = 196;
			16523: out = 568;
			16524: out = 58;
			16525: out = -388;
			16526: out = -707;
			16527: out = -389;
			16528: out = 207;
			16529: out = 604;
			16530: out = 446;
			16531: out = 124;
			16532: out = -254;
			16533: out = -305;
			16534: out = -306;
			16535: out = 314;
			16536: out = 425;
			16537: out = 346;
			16538: out = -111;
			16539: out = 54;
			16540: out = -86;
			16541: out = -506;
			16542: out = -518;
			16543: out = -123;
			16544: out = 303;
			16545: out = 12;
			16546: out = -194;
			16547: out = -284;
			16548: out = -98;
			16549: out = 3;
			16550: out = 5;
			16551: out = -66;
			16552: out = 106;
			16553: out = 67;
			16554: out = -37;
			16555: out = -125;
			16556: out = -314;
			16557: out = -17;
			16558: out = 310;
			16559: out = 216;
			16560: out = 139;
			16561: out = -209;
			16562: out = -719;
			16563: out = -794;
			16564: out = -523;
			16565: out = 115;
			16566: out = 129;
			16567: out = 793;
			16568: out = 41;
			16569: out = -1285;
			16570: out = -928;
			16571: out = -2;
			16572: out = 744;
			16573: out = 897;
			16574: out = -478;
			16575: out = -1038;
			16576: out = -404;
			16577: out = 1097;
			16578: out = 793;
			16579: out = -264;
			16580: out = -717;
			16581: out = -377;
			16582: out = 70;
			16583: out = 13;
			16584: out = 154;
			16585: out = 347;
			16586: out = 564;
			16587: out = -171;
			16588: out = 25;
			16589: out = -279;
			16590: out = -370;
			16591: out = 156;
			16592: out = 381;
			16593: out = -5;
			16594: out = -564;
			16595: out = -1181;
			16596: out = -546;
			16597: out = 603;
			16598: out = 416;
			16599: out = 278;
			16600: out = 15;
			16601: out = -96;
			16602: out = 24;
			16603: out = 51;
			16604: out = 49;
			16605: out = -496;
			16606: out = 458;
			16607: out = 927;
			16608: out = -277;
			16609: out = 263;
			16610: out = 210;
			16611: out = 260;
			16612: out = -138;
			16613: out = 250;
			16614: out = 334;
			16615: out = -33;
			16616: out = -230;
			16617: out = -361;
			16618: out = -282;
			16619: out = -343;
			16620: out = 59;
			16621: out = 330;
			16622: out = 353;
			16623: out = -426;
			16624: out = -992;
			16625: out = -1093;
			16626: out = -49;
			16627: out = 19;
			16628: out = 130;
			16629: out = 103;
			16630: out = 794;
			16631: out = 501;
			16632: out = -89;
			16633: out = -273;
			16634: out = 155;
			16635: out = 387;
			16636: out = -77;
			16637: out = -348;
			16638: out = -485;
			16639: out = -192;
			16640: out = -366;
			16641: out = 334;
			16642: out = 628;
			16643: out = 677;
			16644: out = -353;
			16645: out = -295;
			16646: out = 50;
			16647: out = -370;
			16648: out = -43;
			16649: out = 10;
			16650: out = -88;
			16651: out = -121;
			16652: out = -157;
			16653: out = -137;
			16654: out = -319;
			16655: out = -37;
			16656: out = -46;
			16657: out = -307;
			16658: out = 79;
			16659: out = 40;
			16660: out = -128;
			16661: out = -246;
			16662: out = -145;
			16663: out = 109;
			16664: out = 268;
			16665: out = 820;
			16666: out = 432;
			16667: out = -17;
			16668: out = -134;
			16669: out = -6;
			16670: out = -140;
			16671: out = -524;
			16672: out = -792;
			16673: out = -171;
			16674: out = 588;
			16675: out = 272;
			16676: out = 618;
			16677: out = 166;
			16678: out = -364;
			16679: out = -806;
			16680: out = -219;
			16681: out = 333;
			16682: out = -45;
			16683: out = 104;
			16684: out = -87;
			16685: out = -79;
			16686: out = 0;
			16687: out = 567;
			16688: out = 661;
			16689: out = -223;
			16690: out = -496;
			16691: out = -774;
			16692: out = -689;
			16693: out = -45;
			16694: out = 316;
			16695: out = 324;
			16696: out = 27;
			16697: out = 62;
			16698: out = 261;
			16699: out = 557;
			16700: out = 344;
			16701: out = 107;
			16702: out = -416;
			16703: out = -767;
			16704: out = -1039;
			16705: out = -488;
			16706: out = 224;
			16707: out = 671;
			16708: out = 226;
			16709: out = -155;
			16710: out = -115;
			16711: out = -11;
			16712: out = -20;
			16713: out = -194;
			16714: out = -633;
			16715: out = -194;
			16716: out = 111;
			16717: out = 89;
			16718: out = -355;
			16719: out = -304;
			16720: out = 90;
			16721: out = 835;
			16722: out = 28;
			16723: out = -684;
			16724: out = -709;
			16725: out = 59;
			16726: out = 283;
			16727: out = 36;
			16728: out = 89;
			16729: out = 9;
			16730: out = 44;
			16731: out = -59;
			16732: out = 209;
			16733: out = 266;
			16734: out = 151;
			16735: out = -267;
			16736: out = -424;
			16737: out = -309;
			16738: out = 109;
			16739: out = 333;
			16740: out = 347;
			16741: out = 188;
			16742: out = 252;
			16743: out = 3;
			16744: out = -434;
			16745: out = -1023;
			16746: out = -222;
			16747: out = -75;
			16748: out = -147;
			16749: out = -96;
			16750: out = -90;
			16751: out = 110;
			16752: out = 420;
			16753: out = 86;
			16754: out = -75;
			16755: out = -122;
			16756: out = -69;
			16757: out = 268;
			16758: out = 348;
			16759: out = -51;
			16760: out = -10;
			16761: out = -182;
			16762: out = -2;
			16763: out = 187;
			16764: out = 848;
			16765: out = 601;
			16766: out = -312;
			16767: out = -417;
			16768: out = -375;
			16769: out = -52;
			16770: out = -158;
			16771: out = 50;
			16772: out = -142;
			16773: out = -266;
			16774: out = 0;
			16775: out = 223;
			16776: out = 157;
			16777: out = 42;
			16778: out = -419;
			16779: out = -323;
			16780: out = -38;
			16781: out = 388;
			16782: out = -108;
			16783: out = -571;
			16784: out = -441;
			16785: out = -27;
			16786: out = -7;
			16787: out = -362;
			16788: out = -91;
			16789: out = -95;
			16790: out = -42;
			16791: out = -72;
			16792: out = -74;
			16793: out = 68;
			16794: out = 254;
			16795: out = -81;
			16796: out = 140;
			16797: out = 163;
			16798: out = -368;
			16799: out = 88;
			16800: out = -147;
			16801: out = -524;
			16802: out = -793;
			16803: out = -129;
			16804: out = 294;
			16805: out = -123;
			16806: out = 91;
			16807: out = 105;
			16808: out = 284;
			16809: out = -166;
			16810: out = 43;
			16811: out = -24;
			16812: out = -82;
			16813: out = 1;
			16814: out = 387;
			16815: out = 453;
			16816: out = -17;
			16817: out = -409;
			16818: out = -299;
			16819: out = 50;
			16820: out = 541;
			16821: out = 57;
			16822: out = -656;
			16823: out = -1157;
			16824: out = -343;
			16825: out = 170;
			16826: out = 23;
			16827: out = -34;
			16828: out = 244;
			16829: out = 547;
			16830: out = -160;
			16831: out = -96;
			16832: out = -108;
			16833: out = -63;
			16834: out = -221;
			16835: out = -474;
			16836: out = -516;
			16837: out = 72;
			16838: out = 433;
			16839: out = 507;
			16840: out = 178;
			16841: out = 11;
			16842: out = -122;
			16843: out = -124;
			16844: out = -295;
			16845: out = -155;
			16846: out = -15;
			16847: out = 139;
			16848: out = 239;
			16849: out = 175;
			16850: out = 57;
			16851: out = 71;
			16852: out = 4;
			16853: out = 81;
			16854: out = 71;
			16855: out = -29;
			16856: out = -295;
			16857: out = -368;
			16858: out = 143;
			16859: out = -432;
			16860: out = -607;
			16861: out = -256;
			16862: out = 696;
			16863: out = 687;
			16864: out = 182;
			16865: out = 116;
			16866: out = -820;
			16867: out = -656;
			16868: out = 29;
			16869: out = 660;
			16870: out = 226;
			16871: out = -178;
			16872: out = -40;
			16873: out = 535;
			16874: out = 301;
			16875: out = -606;
			16876: out = -196;
			16877: out = -433;
			16878: out = -303;
			16879: out = 57;
			16880: out = -28;
			16881: out = -28;
			16882: out = 55;
			16883: out = 45;
			16884: out = -50;
			16885: out = -86;
			16886: out = 146;
			16887: out = 284;
			16888: out = 490;
			16889: out = 437;
			16890: out = 73;
			16891: out = -318;
			16892: out = -422;
			16893: out = -93;
			16894: out = -12;
			16895: out = -12;
			16896: out = -112;
			16897: out = 547;
			16898: out = 76;
			16899: out = -178;
			16900: out = -130;
			16901: out = 18;
			16902: out = -277;
			16903: out = -615;
			16904: out = -44;
			16905: out = -100;
			16906: out = -117;
			16907: out = -113;
			16908: out = 61;
			16909: out = 165;
			16910: out = 288;
			16911: out = 495;
			16912: out = 230;
			16913: out = -326;
			16914: out = -988;
			16915: out = -383;
			16916: out = -132;
			16917: out = 7;
			16918: out = 390;
			16919: out = 291;
			16920: out = 117;
			16921: out = -91;
			16922: out = -61;
			16923: out = -94;
			16924: out = -104;
			16925: out = 32;
			16926: out = -97;
			16927: out = -115;
			16928: out = -50;
			16929: out = -79;
			16930: out = -86;
			16931: out = -126;
			16932: out = 51;
			16933: out = -114;
			16934: out = 42;
			16935: out = 414;
			16936: out = -104;
			16937: out = -216;
			16938: out = -225;
			16939: out = 278;
			16940: out = -44;
			16941: out = 123;
			16942: out = 545;
			16943: out = 238;
			16944: out = 36;
			16945: out = -75;
			16946: out = 231;
			16947: out = 54;
			16948: out = -120;
			16949: out = -331;
			16950: out = 57;
			16951: out = -24;
			16952: out = -139;
			16953: out = -316;
			16954: out = -138;
			16955: out = -25;
			16956: out = 61;
			16957: out = -458;
			16958: out = -184;
			16959: out = 48;
			16960: out = -94;
			16961: out = 21;
			16962: out = -102;
			16963: out = -289;
			16964: out = 405;
			16965: out = -210;
			16966: out = -611;
			16967: out = 12;
			16968: out = 356;
			16969: out = 362;
			16970: out = -286;
			16971: out = 141;
			16972: out = -552;
			16973: out = -812;
			16974: out = -978;
			16975: out = 318;
			16976: out = 361;
			16977: out = -152;
			16978: out = -409;
			16979: out = 235;
			16980: out = 839;
			16981: out = 698;
			16982: out = -543;
			16983: out = -1241;
			16984: out = -865;
			16985: out = -184;
			16986: out = 533;
			16987: out = 498;
			16988: out = -139;
			16989: out = -115;
			16990: out = 11;
			16991: out = 112;
			16992: out = 85;
			16993: out = -16;
			16994: out = -186;
			16995: out = -235;
			16996: out = -17;
			16997: out = 15;
			16998: out = -123;
			16999: out = 158;
			17000: out = -49;
			17001: out = 22;
			17002: out = 82;
			17003: out = 286;
			17004: out = -88;
			17005: out = -528;
			17006: out = -754;
			17007: out = -166;
			17008: out = 210;
			17009: out = 69;
			17010: out = -47;
			17011: out = -7;
			17012: out = 118;
			17013: out = -33;
			17014: out = -324;
			17015: out = -201;
			17016: out = 506;
			17017: out = 45;
			17018: out = -68;
			17019: out = -296;
			17020: out = 205;
			17021: out = -580;
			17022: out = -437;
			17023: out = 372;
			17024: out = 238;
			17025: out = 204;
			17026: out = 64;
			17027: out = 55;
			17028: out = 55;
			17029: out = -50;
			17030: out = -276;
			17031: out = 36;
			17032: out = 154;
			17033: out = 238;
			17034: out = 83;
			17035: out = 62;
			17036: out = 146;
			17037: out = 407;
			17038: out = 60;
			17039: out = 190;
			17040: out = 149;
			17041: out = -79;
			17042: out = -478;
			17043: out = -713;
			17044: out = -679;
			17045: out = 164;
			17046: out = 195;
			17047: out = -111;
			17048: out = -609;
			17049: out = -94;
			17050: out = 134;
			17051: out = 91;
			17052: out = 55;
			17053: out = 53;
			17054: out = -11;
			17055: out = -280;
			17056: out = -261;
			17057: out = -163;
			17058: out = 24;
			17059: out = 521;
			17060: out = 281;
			17061: out = 37;
			17062: out = 65;
			17063: out = -34;
			17064: out = -278;
			17065: out = -602;
			17066: out = 78;
			17067: out = 139;
			17068: out = 290;
			17069: out = 7;
			17070: out = 793;
			17071: out = 171;
			17072: out = -674;
			17073: out = -102;
			17074: out = -78;
			17075: out = -54;
			17076: out = 78;
			17077: out = -107;
			17078: out = 201;
			17079: out = 254;
			17080: out = -355;
			17081: out = -1080;
			17082: out = -906;
			17083: out = 222;
			17084: out = 591;
			17085: out = 502;
			17086: out = 78;
			17087: out = -754;
			17088: out = -160;
			17089: out = 30;
			17090: out = -432;
			17091: out = -59;
			17092: out = 594;
			17093: out = 1017;
			17094: out = 393;
			17095: out = -412;
			17096: out = -818;
			17097: out = -502;
			17098: out = 398;
			17099: out = 370;
			17100: out = -68;
			17101: out = -596;
			17102: out = 309;
			17103: out = 530;
			17104: out = -263;
			17105: out = -487;
			17106: out = -387;
			17107: out = 15;
			17108: out = -491;
			17109: out = -109;
			17110: out = 227;
			17111: out = 827;
			17112: out = -332;
			17113: out = -364;
			17114: out = -104;
			17115: out = 544;
			17116: out = 183;
			17117: out = -41;
			17118: out = -32;
			17119: out = 13;
			17120: out = 48;
			17121: out = 10;
			17122: out = -53;
			17123: out = -102;
			17124: out = -92;
			17125: out = -45;
			17126: out = -110;
			17127: out = 67;
			17128: out = 284;
			17129: out = 171;
			17130: out = 35;
			17131: out = -480;
			17132: out = -868;
			17133: out = -190;
			17134: out = 163;
			17135: out = 136;
			17136: out = -248;
			17137: out = -641;
			17138: out = -454;
			17139: out = 150;
			17140: out = -269;
			17141: out = -111;
			17142: out = -105;
			17143: out = -216;
			17144: out = 134;
			17145: out = 422;
			17146: out = 491;
			17147: out = -5;
			17148: out = 32;
			17149: out = 84;
			17150: out = -63;
			17151: out = -27;
			17152: out = -15;
			17153: out = 52;
			17154: out = -106;
			17155: out = -169;
			17156: out = -224;
			17157: out = 113;
			17158: out = -110;
			17159: out = 18;
			17160: out = 86;
			17161: out = 450;
			17162: out = -426;
			17163: out = -875;
			17164: out = -291;
			17165: out = 75;
			17166: out = 419;
			17167: out = 332;
			17168: out = 439;
			17169: out = 120;
			17170: out = 182;
			17171: out = 619;
			17172: out = -447;
			17173: out = -1151;
			17174: out = -1132;
			17175: out = 728;
			17176: out = 679;
			17177: out = 285;
			17178: out = -110;
			17179: out = -81;
			17180: out = 35;
			17181: out = 88;
			17182: out = 51;
			17183: out = -164;
			17184: out = -226;
			17185: out = 98;
			17186: out = -396;
			17187: out = -105;
			17188: out = 315;
			17189: out = 193;
			17190: out = 258;
			17191: out = 118;
			17192: out = -131;
			17193: out = -138;
			17194: out = -85;
			17195: out = -184;
			17196: out = -1113;
			17197: out = -424;
			17198: out = 187;
			17199: out = 520;
			17200: out = -19;
			17201: out = -34;
			17202: out = 236;
			17203: out = 795;
			17204: out = 54;
			17205: out = -319;
			17206: out = 130;
			17207: out = -202;
			17208: out = 138;
			17209: out = 133;
			17210: out = 154;
			17211: out = -733;
			17212: out = -647;
			17213: out = 199;
			17214: out = -91;
			17215: out = -58;
			17216: out = -137;
			17217: out = -93;
			17218: out = -20;
			17219: out = 168;
			17220: out = 400;
			17221: out = 41;
			17222: out = -38;
			17223: out = -78;
			17224: out = 619;
			17225: out = -683;
			17226: out = -632;
			17227: out = 147;
			17228: out = 233;
			17229: out = -317;
			17230: out = -804;
			17231: out = -334;
			17232: out = 168;
			17233: out = 541;
			17234: out = 455;
			17235: out = 86;
			17236: out = 10;
			17237: out = 45;
			17238: out = 95;
			17239: out = -346;
			17240: out = -337;
			17241: out = -50;
			17242: out = 226;
			17243: out = 98;
			17244: out = 108;
			17245: out = 372;
			17246: out = 843;
			17247: out = 358;
			17248: out = -599;
			17249: out = -18;
			17250: out = -150;
			17251: out = -294;
			17252: out = -1024;
			17253: out = -48;
			17254: out = 91;
			17255: out = 7;
			17256: out = -123;
			17257: out = 15;
			17258: out = 82;
			17259: out = 83;
			17260: out = 31;
			17261: out = 73;
			17262: out = 22;
			17263: out = -256;
			17264: out = -323;
			17265: out = -208;
			17266: out = -122;
			17267: out = 332;
			17268: out = 226;
			17269: out = 43;
			17270: out = 352;
			17271: out = 168;
			17272: out = -223;
			17273: out = -602;
			17274: out = -653;
			17275: out = -100;
			17276: out = 455;
			17277: out = 187;
			17278: out = 142;
			17279: out = -11;
			17280: out = -125;
			17281: out = 58;
			17282: out = -27;
			17283: out = -155;
			17284: out = -302;
			17285: out = 0;
			17286: out = 23;
			17287: out = -136;
			17288: out = -425;
			17289: out = -31;
			17290: out = 503;
			17291: out = 621;
			17292: out = -9;
			17293: out = -399;
			17294: out = -193;
			17295: out = -2;
			17296: out = 137;
			17297: out = 10;
			17298: out = 100;
			17299: out = -77;
			17300: out = -8;
			17301: out = 28;
			17302: out = -200;
			17303: out = -591;
			17304: out = -521;
			17305: out = 537;
			17306: out = 193;
			17307: out = -226;
			17308: out = -789;
			17309: out = -70;
			17310: out = -401;
			17311: out = -445;
			17312: out = 83;
			17313: out = 774;
			17314: out = 983;
			17315: out = 505;
			17316: out = -861;
			17317: out = -1280;
			17318: out = -872;
			17319: out = 133;
			17320: out = 124;
			17321: out = 86;
			17322: out = 83;
			17323: out = 360;
			17324: out = 293;
			17325: out = 116;
			17326: out = -285;
			17327: out = 5;
			17328: out = -83;
			17329: out = -225;
			17330: out = 185;
			17331: out = 443;
			17332: out = 230;
			17333: out = -799;
			17334: out = -202;
			17335: out = 0;
			17336: out = 96;
			17337: out = -65;
			17338: out = 37;
			17339: out = -104;
			17340: out = -593;
			17341: out = -93;
			17342: out = -168;
			17343: out = -360;
			17344: out = 258;
			17345: out = 221;
			17346: out = 189;
			17347: out = -90;
			17348: out = 114;
			17349: out = -70;
			17350: out = -222;
			17351: out = 21;
			17352: out = 362;
			17353: out = 424;
			17354: out = -51;
			17355: out = -314;
			17356: out = -333;
			17357: out = 23;
			17358: out = 0;
			17359: out = 278;
			17360: out = -121;
			17361: out = -884;
			17362: out = -377;
			17363: out = 134;
			17364: out = 364;
			17365: out = 268;
			17366: out = -137;
			17367: out = -46;
			17368: out = 530;
			17369: out = 143;
			17370: out = -112;
			17371: out = -211;
			17372: out = 63;
			17373: out = 567;
			17374: out = 489;
			17375: out = -395;
			17376: out = 52;
			17377: out = -17;
			17378: out = -40;
			17379: out = -649;
			17380: out = 125;
			17381: out = 323;
			17382: out = -1;
			17383: out = -73;
			17384: out = -160;
			17385: out = -168;
			17386: out = -611;
			17387: out = -102;
			17388: out = 294;
			17389: out = 626;
			17390: out = -81;
			17391: out = -130;
			17392: out = -147;
			17393: out = -17;
			17394: out = -376;
			17395: out = -267;
			17396: out = 65;
			17397: out = 372;
			17398: out = -89;
			17399: out = -403;
			17400: out = 54;
			17401: out = 398;
			17402: out = 243;
			17403: out = -361;
			17404: out = -106;
			17405: out = 121;
			17406: out = 283;
			17407: out = -528;
			17408: out = -26;
			17409: out = 78;
			17410: out = 265;
			17411: out = -59;
			17412: out = 351;
			17413: out = 331;
			17414: out = -84;
			17415: out = -651;
			17416: out = -640;
			17417: out = -351;
			17418: out = 220;
			17419: out = -187;
			17420: out = -292;
			17421: out = 247;
			17422: out = 852;
			17423: out = 573;
			17424: out = -318;
			17425: out = -207;
			17426: out = -250;
			17427: out = -77;
			17428: out = -171;
			17429: out = 58;
			17430: out = 8;
			17431: out = -72;
			17432: out = 364;
			17433: out = -59;
			17434: out = -268;
			17435: out = 52;
			17436: out = -89;
			17437: out = -26;
			17438: out = -75;
			17439: out = -899;
			17440: out = -418;
			17441: out = 95;
			17442: out = 354;
			17443: out = -8;
			17444: out = -12;
			17445: out = 80;
			17446: out = 44;
			17447: out = -304;
			17448: out = -295;
			17449: out = 120;
			17450: out = 196;
			17451: out = -69;
			17452: out = -422;
			17453: out = 108;
			17454: out = 138;
			17455: out = 209;
			17456: out = -28;
			17457: out = 100;
			17458: out = -186;
			17459: out = -424;
			17460: out = -90;
			17461: out = -59;
			17462: out = 204;
			17463: out = 447;
			17464: out = 297;
			17465: out = -245;
			17466: out = -496;
			17467: out = 369;
			17468: out = 117;
			17469: out = -158;
			17470: out = -433;
			17471: out = -28;
			17472: out = -103;
			17473: out = -275;
			17474: out = 154;
			17475: out = -449;
			17476: out = -388;
			17477: out = 95;
			17478: out = 454;
			17479: out = 209;
			17480: out = -137;
			17481: out = -49;
			17482: out = 0;
			17483: out = -35;
			17484: out = -126;
			17485: out = -287;
			17486: out = 168;
			17487: out = 453;
			17488: out = 25;
			17489: out = -168;
			17490: out = -258;
			17491: out = -93;
			17492: out = -82;
			17493: out = -166;
			17494: out = -269;
			17495: out = -88;
			17496: out = -85;
			17497: out = -26;
			17498: out = 63;
			17499: out = 32;
			17500: out = 480;
			17501: out = 667;
			17502: out = 130;
			17503: out = 84;
			17504: out = -100;
			17505: out = -120;
			17506: out = 32;
			17507: out = -28;
			17508: out = -315;
			17509: out = -728;
			17510: out = -18;
			17511: out = 463;
			17512: out = 475;
			17513: out = -361;
			17514: out = -582;
			17515: out = -433;
			17516: out = -42;
			17517: out = 256;
			17518: out = 211;
			17519: out = -121;
			17520: out = 546;
			17521: out = -347;
			17522: out = -713;
			17523: out = -204;
			17524: out = -114;
			17525: out = -260;
			17526: out = -546;
			17527: out = 254;
			17528: out = 22;
			17529: out = -112;
			17530: out = -268;
			17531: out = -78;
			17532: out = -2;
			17533: out = 62;
			17534: out = 16;
			17535: out = -36;
			17536: out = -199;
			17537: out = -199;
			17538: out = -302;
			17539: out = 73;
			17540: out = 429;
			17541: out = 608;
			17542: out = 117;
			17543: out = -143;
			17544: out = 67;
			17545: out = 51;
			17546: out = -76;
			17547: out = -271;
			17548: out = 130;
			17549: out = -105;
			17550: out = -97;
			17551: out = -133;
			17552: out = 204;
			17553: out = 40;
			17554: out = -145;
			17555: out = -116;
			17556: out = 29;
			17557: out = -5;
			17558: out = -296;
			17559: out = 82;
			17560: out = -80;
			17561: out = -294;
			17562: out = -229;
			17563: out = -175;
			17564: out = 74;
			17565: out = 348;
			17566: out = -339;
			17567: out = -195;
			17568: out = 101;
			17569: out = -26;
			17570: out = 222;
			17571: out = 124;
			17572: out = 55;
			17573: out = -117;
			17574: out = 204;
			17575: out = 204;
			17576: out = -420;
			17577: out = -527;
			17578: out = -312;
			17579: out = 158;
			17580: out = 431;
			17581: out = 240;
			17582: out = -59;
			17583: out = -88;
			17584: out = 19;
			17585: out = 21;
			17586: out = -150;
			17587: out = -243;
			17588: out = -3;
			17589: out = 236;
			17590: out = -25;
			17591: out = -8;
			17592: out = -99;
			17593: out = -37;
			17594: out = 36;
			17595: out = 94;
			17596: out = 68;
			17597: out = 224;
			17598: out = -208;
			17599: out = -156;
			17600: out = 45;
			17601: out = 206;
			17602: out = -257;
			17603: out = -536;
			17604: out = -40;
			17605: out = -148;
			17606: out = -130;
			17607: out = -263;
			17608: out = 251;
			17609: out = -30;
			17610: out = -56;
			17611: out = 45;
			17612: out = 5;
			17613: out = -254;
			17614: out = -326;
			17615: out = -29;
			17616: out = 200;
			17617: out = 154;
			17618: out = 252;
			17619: out = -729;
			17620: out = -467;
			17621: out = 125;
			17622: out = 378;
			17623: out = -523;
			17624: out = -884;
			17625: out = 59;
			17626: out = 645;
			17627: out = 652;
			17628: out = 95;
			17629: out = 674;
			17630: out = 66;
			17631: out = -235;
			17632: out = -395;
			17633: out = -22;
			17634: out = 263;
			17635: out = 411;
			17636: out = 16;
			17637: out = -278;
			17638: out = -357;
			17639: out = 89;
			17640: out = -47;
			17641: out = 206;
			17642: out = 248;
			17643: out = -49;
			17644: out = -543;
			17645: out = -655;
			17646: out = -178;
			17647: out = -136;
			17648: out = 45;
			17649: out = 54;
			17650: out = 37;
			17651: out = -197;
			17652: out = -307;
			17653: out = -407;
			17654: out = -125;
			17655: out = -185;
			17656: out = -245;
			17657: out = -256;
			17658: out = 299;
			17659: out = 463;
			17660: out = 135;
			17661: out = 119;
			17662: out = -179;
			17663: out = -215;
			17664: out = -73;
			17665: out = 65;
			17666: out = 69;
			17667: out = 7;
			17668: out = -392;
			17669: out = -147;
			17670: out = 155;
			17671: out = 45;
			17672: out = 215;
			17673: out = 133;
			17674: out = 15;
			17675: out = -49;
			17676: out = -100;
			17677: out = -109;
			17678: out = -51;
			17679: out = 5;
			17680: out = 27;
			17681: out = 45;
			17682: out = 184;
			17683: out = 440;
			17684: out = 457;
			17685: out = -367;
			17686: out = 43;
			17687: out = 8;
			17688: out = 52;
			17689: out = -605;
			17690: out = -183;
			17691: out = 15;
			17692: out = 40;
			17693: out = -639;
			17694: out = -288;
			17695: out = 416;
			17696: out = 234;
			17697: out = -569;
			17698: out = -966;
			17699: out = 52;
			17700: out = -133;
			17701: out = 56;
			17702: out = 46;
			17703: out = 513;
			17704: out = 185;
			17705: out = -33;
			17706: out = -108;
			17707: out = 145;
			17708: out = 192;
			17709: out = 4;
			17710: out = 90;
			17711: out = -522;
			17712: out = -545;
			17713: out = 99;
			17714: out = 166;
			17715: out = 175;
			17716: out = 35;
			17717: out = -63;
			17718: out = -62;
			17719: out = -44;
			17720: out = 38;
			17721: out = -272;
			17722: out = 47;
			17723: out = 385;
			17724: out = 321;
			17725: out = 13;
			17726: out = -103;
			17727: out = 86;
			17728: out = 26;
			17729: out = -212;
			17730: out = -447;
			17731: out = -409;
			17732: out = -63;
			17733: out = 27;
			17734: out = -299;
			17735: out = -109;
			17736: out = -44;
			17737: out = 53;
			17738: out = 14;
			17739: out = -69;
			17740: out = 54;
			17741: out = 508;
			17742: out = -214;
			17743: out = -253;
			17744: out = -270;
			17745: out = -366;
			17746: out = -70;
			17747: out = 316;
			17748: out = 560;
			17749: out = 93;
			17750: out = -85;
			17751: out = -134;
			17752: out = -271;
			17753: out = -38;
			17754: out = 19;
			17755: out = -68;
			17756: out = 29;
			17757: out = 10;
			17758: out = 77;
			17759: out = 353;
			17760: out = -30;
			17761: out = -31;
			17762: out = 245;
			17763: out = 272;
			17764: out = 265;
			17765: out = 86;
			17766: out = 11;
			17767: out = -114;
			17768: out = -146;
			17769: out = -123;
			17770: out = 179;
			17771: out = -1;
			17772: out = -160;
			17773: out = 29;
			17774: out = -218;
			17775: out = -289;
			17776: out = -230;
			17777: out = 166;
			17778: out = 39;
			17779: out = -159;
			17780: out = -237;
			17781: out = -162;
			17782: out = 180;
			17783: out = 388;
			17784: out = -237;
			17785: out = -550;
			17786: out = -559;
			17787: out = 146;
			17788: out = -470;
			17789: out = -346;
			17790: out = -46;
			17791: out = 218;
			17792: out = -86;
			17793: out = -127;
			17794: out = 374;
			17795: out = 64;
			17796: out = -93;
			17797: out = -253;
			17798: out = -50;
			17799: out = 89;
			17800: out = 212;
			17801: out = 15;
			17802: out = -32;
			17803: out = -289;
			17804: out = -319;
			17805: out = -100;
			17806: out = 300;
			17807: out = 448;
			17808: out = 257;
			17809: out = -375;
			17810: out = -557;
			17811: out = -214;
			17812: out = 266;
			17813: out = 369;
			17814: out = 208;
			17815: out = 60;
			17816: out = -478;
			17817: out = -435;
			17818: out = -125;
			17819: out = 329;
			17820: out = -60;
			17821: out = -277;
			17822: out = -44;
			17823: out = -147;
			17824: out = -14;
			17825: out = 35;
			17826: out = 227;
			17827: out = -230;
			17828: out = -444;
			17829: out = -331;
			17830: out = 130;
			17831: out = 191;
			17832: out = -55;
			17833: out = -340;
			17834: out = -241;
			17835: out = 77;
			17836: out = 203;
			17837: out = 473;
			17838: out = 297;
			17839: out = 141;
			17840: out = -152;
			17841: out = 71;
			17842: out = -173;
			17843: out = -544;
			17844: out = -444;
			17845: out = 48;
			17846: out = 299;
			17847: out = -117;
			17848: out = -353;
			17849: out = -77;
			17850: out = 520;
			17851: out = 565;
			17852: out = 118;
			17853: out = -329;
			17854: out = -73;
			17855: out = 289;
			17856: out = 310;
			17857: out = -239;
			17858: out = 56;
			17859: out = -18;
			17860: out = 100;
			17861: out = -47;
			17862: out = 187;
			17863: out = 96;
			17864: out = -48;
			17865: out = -1417;
			17866: out = -881;
			17867: out = -124;
			17868: out = 189;
			17869: out = 122;
			17870: out = -2;
			17871: out = -142;
			17872: out = -352;
			17873: out = -316;
			17874: out = -130;
			17875: out = 34;
			17876: out = 427;
			17877: out = 288;
			17878: out = -76;
			17879: out = -796;
			17880: out = -274;
			17881: out = 292;
			17882: out = 433;
			17883: out = 134;
			17884: out = -53;
			17885: out = -55;
			17886: out = 462;
			17887: out = 80;
			17888: out = -100;
			17889: out = 92;
			17890: out = 299;
			17891: out = -1;
			17892: out = -431;
			17893: out = -57;
			17894: out = 172;
			17895: out = 322;
			17896: out = 150;
			17897: out = -430;
			17898: out = -346;
			17899: out = 98;
			17900: out = -120;
			17901: out = -54;
			17902: out = -184;
			17903: out = -232;
			17904: out = -98;
			17905: out = 9;
			17906: out = 153;
			17907: out = 553;
			17908: out = 172;
			17909: out = -394;
			17910: out = -824;
			17911: out = -617;
			17912: out = -171;
			17913: out = 143;
			17914: out = 370;
			17915: out = -179;
			17916: out = -425;
			17917: out = -329;
			17918: out = 500;
			17919: out = 311;
			17920: out = -173;
			17921: out = -203;
			17922: out = -154;
			17923: out = -113;
			17924: out = -251;
			17925: out = -89;
			17926: out = -7;
			17927: out = 201;
			17928: out = 587;
			17929: out = 111;
			17930: out = -116;
			17931: out = -30;
			17932: out = -84;
			17933: out = -8;
			17934: out = -20;
			17935: out = -423;
			17936: out = -9;
			17937: out = 79;
			17938: out = 17;
			17939: out = -260;
			17940: out = 162;
			17941: out = 460;
			17942: out = 171;
			17943: out = 81;
			17944: out = -9;
			17945: out = -9;
			17946: out = -74;
			17947: out = -318;
			17948: out = -269;
			17949: out = 198;
			17950: out = 424;
			17951: out = 63;
			17952: out = -603;
			17953: out = -242;
			17954: out = -19;
			17955: out = 270;
			17956: out = 144;
			17957: out = -309;
			17958: out = -801;
			17959: out = -863;
			17960: out = 5;
			17961: out = 155;
			17962: out = -8;
			17963: out = -204;
			17964: out = -85;
			17965: out = -19;
			17966: out = 0;
			17967: out = 600;
			17968: out = 253;
			17969: out = -48;
			17970: out = 68;
			17971: out = 0;
			17972: out = 82;
			17973: out = 47;
			17974: out = 248;
			17975: out = -299;
			17976: out = -430;
			17977: out = 149;
			17978: out = 40;
			17979: out = 36;
			17980: out = -151;
			17981: out = 50;
			17982: out = -83;
			17983: out = -23;
			17984: out = 200;
			17985: out = -14;
			17986: out = -113;
			17987: out = -63;
			17988: out = 183;
			17989: out = 106;
			17990: out = -25;
			17991: out = 39;
			17992: out = -393;
			17993: out = -217;
			17994: out = -35;
			17995: out = 59;
			17996: out = -322;
			17997: out = -172;
			17998: out = 365;
			17999: out = 356;
			18000: out = -236;
			18001: out = -927;
			18002: out = -431;
			18003: out = -272;
			18004: out = 234;
			18005: out = 399;
			18006: out = 183;
			18007: out = -388;
			18008: out = -557;
			18009: out = -46;
			18010: out = 510;
			18011: out = 521;
			18012: out = -64;
			18013: out = -43;
			18014: out = -203;
			18015: out = -211;
			18016: out = -236;
			18017: out = 96;
			18018: out = 266;
			18019: out = 308;
			18020: out = -28;
			18021: out = -6;
			18022: out = 62;
			18023: out = -118;
			18024: out = -3;
			18025: out = -12;
			18026: out = -120;
			18027: out = 31;
			18028: out = -117;
			18029: out = -304;
			18030: out = -511;
			18031: out = 41;
			18032: out = 179;
			18033: out = -102;
			18034: out = 356;
			18035: out = 123;
			18036: out = -14;
			18037: out = -133;
			18038: out = 172;
			18039: out = 30;
			18040: out = -266;
			18041: out = -371;
			18042: out = -282;
			18043: out = -202;
			18044: out = -55;
			18045: out = -355;
			18046: out = 20;
			18047: out = 609;
			18048: out = 197;
			18049: out = -187;
			18050: out = -534;
			18051: out = -140;
			18052: out = -137;
			18053: out = 130;
			18054: out = 160;
			18055: out = 12;
			18056: out = -292;
			18057: out = -223;
			18058: out = 100;
			18059: out = 378;
			18060: out = 351;
			18061: out = 151;
			18062: out = 86;
			18063: out = 29;
			18064: out = 20;
			18065: out = 82;
			18066: out = -66;
			18067: out = -50;
			18068: out = -114;
			18069: out = -177;
			18070: out = -551;
			18071: out = -406;
			18072: out = 367;
			18073: out = 114;
			18074: out = -353;
			18075: out = -754;
			18076: out = 102;
			18077: out = 92;
			18078: out = -10;
			18079: out = -386;
			18080: out = -49;
			18081: out = -61;
			18082: out = -48;
			18083: out = 81;
			18084: out = 87;
			18085: out = -4;
			18086: out = -19;
			18087: out = -213;
			18088: out = -57;
			18089: out = 113;
			18090: out = 37;
			18091: out = -40;
			18092: out = -72;
			18093: out = 62;
			18094: out = 26;
			18095: out = 41;
			18096: out = 39;
			18097: out = 81;
			18098: out = -12;
			18099: out = -26;
			18100: out = 95;
			18101: out = -90;
			18102: out = -44;
			18103: out = 64;
			18104: out = 54;
			18105: out = -6;
			18106: out = -84;
			18107: out = -18;
			18108: out = -1;
			18109: out = 134;
			18110: out = 189;
			18111: out = 208;
			18112: out = -126;
			18113: out = -299;
			18114: out = -199;
			18115: out = 149;
			18116: out = 217;
			18117: out = 132;
			18118: out = -83;
			18119: out = 43;
			18120: out = -4;
			18121: out = -162;
			18122: out = -491;
			18123: out = -460;
			18124: out = -327;
			18125: out = -228;
			18126: out = -132;
			18127: out = -55;
			18128: out = -36;
			18129: out = 354;
			18130: out = -68;
			18131: out = -371;
			18132: out = -7;
			18133: out = -32;
			18134: out = -368;
			18135: out = -962;
			18136: out = 116;
			18137: out = 13;
			18138: out = -68;
			18139: out = -370;
			18140: out = 432;
			18141: out = 603;
			18142: out = 335;
			18143: out = -585;
			18144: out = -341;
			18145: out = 67;
			18146: out = 211;
			18147: out = -4;
			18148: out = -84;
			18149: out = -11;
			18150: out = 61;
			18151: out = -19;
			18152: out = 38;
			18153: out = 206;
			18154: out = 158;
			18155: out = -191;
			18156: out = -544;
			18157: out = -646;
			18158: out = -58;
			18159: out = 308;
			18160: out = 180;
			18161: out = 0;
			18162: out = -85;
			18163: out = 13;
			18164: out = 361;
			18165: out = -110;
			18166: out = -324;
			18167: out = 106;
			18168: out = -214;
			18169: out = -84;
			18170: out = 82;
			18171: out = 80;
			18172: out = 26;
			18173: out = -93;
			18174: out = -22;
			18175: out = -52;
			18176: out = 485;
			18177: out = 650;
			18178: out = -499;
			18179: out = -740;
			18180: out = -549;
			18181: out = 142;
			18182: out = 81;
			18183: out = 17;
			18184: out = -41;
			18185: out = 377;
			18186: out = 236;
			18187: out = 208;
			18188: out = 204;
			18189: out = 307;
			18190: out = 222;
			18191: out = -67;
			18192: out = -318;
			18193: out = -613;
			18194: out = -325;
			18195: out = 270;
			18196: out = 521;
			18197: out = 228;
			18198: out = -120;
			18199: out = 98;
			18200: out = 27;
			18201: out = -106;
			18202: out = -405;
			18203: out = -208;
			18204: out = -232;
			18205: out = -206;
			18206: out = -65;
			18207: out = -21;
			18208: out = 179;
			18209: out = 284;
			18210: out = 80;
			18211: out = -293;
			18212: out = -402;
			18213: out = 46;
			18214: out = 165;
			18215: out = 154;
			18216: out = -10;
			18217: out = -325;
			18218: out = -191;
			18219: out = 35;
			18220: out = 198;
			18221: out = -325;
			18222: out = -436;
			18223: out = -129;
			18224: out = -68;
			18225: out = -9;
			18226: out = -28;
			18227: out = 116;
			18228: out = -145;
			18229: out = -232;
			18230: out = -150;
			18231: out = 62;
			18232: out = 263;
			18233: out = 217;
			18234: out = -249;
			18235: out = -2;
			18236: out = 166;
			18237: out = 320;
			18238: out = 58;
			18239: out = 76;
			18240: out = 1;
			18241: out = 107;
			18242: out = -212;
			18243: out = -138;
			18244: out = -25;
			18245: out = 341;
			18246: out = -216;
			18247: out = -418;
			18248: out = 84;
			18249: out = -55;
			18250: out = -40;
			18251: out = -75;
			18252: out = -362;
			18253: out = -58;
			18254: out = 114;
			18255: out = 72;
			18256: out = -298;
			18257: out = -185;
			18258: out = 200;
			18259: out = 1046;
			18260: out = 152;
			18261: out = -741;
			18262: out = -1109;
			18263: out = -132;
			18264: out = 280;
			18265: out = 272;
			18266: out = -83;
			18267: out = 18;
			18268: out = 42;
			18269: out = -102;
			18270: out = -689;
			18271: out = -357;
			18272: out = 175;
			18273: out = -50;
			18274: out = -221;
			18275: out = -131;
			18276: out = 503;
			18277: out = -168;
			18278: out = -155;
			18279: out = 33;
			18280: out = 565;
			18281: out = 320;
			18282: out = 100;
			18283: out = 26;
			18284: out = -223;
			18285: out = -143;
			18286: out = -83;
			18287: out = 65;
			18288: out = -204;
			18289: out = -56;
			18290: out = 200;
			18291: out = 123;
			18292: out = -321;
			18293: out = -603;
			18294: out = -193;
			18295: out = 278;
			18296: out = 328;
			18297: out = -144;
			18298: out = -402;
			18299: out = -372;
			18300: out = -116;
			18301: out = -108;
			18302: out = 68;
			18303: out = 177;
			18304: out = 364;
			18305: out = 417;
			18306: out = 217;
			18307: out = -32;
			18308: out = 72;
			18309: out = -327;
			18310: out = -211;
			18311: out = 94;
			18312: out = 391;
			18313: out = 1;
			18314: out = -475;
			18315: out = -255;
			18316: out = -464;
			18317: out = 125;
			18318: out = 677;
			18319: out = 663;
			18320: out = -30;
			18321: out = -619;
			18322: out = -421;
			18323: out = -93;
			18324: out = 142;
			18325: out = 40;
			18326: out = 351;
			18327: out = 34;
			18328: out = -157;
			18329: out = -233;
			18330: out = 205;
			18331: out = 375;
			18332: out = 330;
			18333: out = -352;
			18334: out = -241;
			18335: out = 54;
			18336: out = 410;
			18337: out = 103;
			18338: out = -39;
			18339: out = -118;
			18340: out = 61;
			18341: out = 8;
			18342: out = -48;
			18343: out = -290;
			18344: out = 251;
			18345: out = 0;
			18346: out = -482;
			18347: out = -615;
			18348: out = -243;
			18349: out = 207;
			18350: out = 379;
			18351: out = -241;
			18352: out = -412;
			18353: out = -299;
			18354: out = -47;
			18355: out = -264;
			18356: out = -275;
			18357: out = 77;
			18358: out = 31;
			18359: out = -81;
			18360: out = -238;
			18361: out = -70;
			18362: out = 166;
			18363: out = 443;
			18364: out = 471;
			18365: out = -219;
			18366: out = -645;
			18367: out = -638;
			18368: out = 99;
			18369: out = 61;
			18370: out = 134;
			18371: out = 200;
			18372: out = 435;
			18373: out = 11;
			18374: out = -344;
			18375: out = 359;
			18376: out = 84;
			18377: out = -192;
			18378: out = -675;
			18379: out = -45;
			18380: out = -171;
			18381: out = -156;
			18382: out = 0;
			18383: out = 376;
			18384: out = 240;
			18385: out = -131;
			18386: out = -254;
			18387: out = 198;
			18388: out = 528;
			18389: out = -6;
			18390: out = -21;
			18391: out = -262;
			18392: out = -321;
			18393: out = -119;
			18394: out = 172;
			18395: out = 277;
			18396: out = 25;
			18397: out = -18;
			18398: out = -119;
			18399: out = -72;
			18400: out = -292;
			18401: out = 184;
			18402: out = 314;
			18403: out = -281;
			18404: out = -551;
			18405: out = -454;
			18406: out = 10;
			18407: out = 135;
			18408: out = 94;
			18409: out = -174;
			18410: out = -313;
			18411: out = 42;
			18412: out = 240;
			18413: out = -33;
			18414: out = 115;
			18415: out = -301;
			18416: out = -118;
			18417: out = 389;
			18418: out = 679;
			18419: out = 9;
			18420: out = -830;
			18421: out = -244;
			18422: out = 264;
			18423: out = 473;
			18424: out = -75;
			18425: out = -151;
			18426: out = -273;
			18427: out = -180;
			18428: out = 2;
			18429: out = 16;
			18430: out = 10;
			18431: out = -80;
			18432: out = 185;
			18433: out = -134;
			18434: out = -554;
			18435: out = -467;
			18436: out = -187;
			18437: out = -7;
			18438: out = -103;
			18439: out = -207;
			18440: out = 89;
			18441: out = 475;
			18442: out = 152;
			18443: out = 112;
			18444: out = -3;
			18445: out = 87;
			18446: out = -209;
			18447: out = -155;
			18448: out = -31;
			18449: out = -128;
			18450: out = 221;
			18451: out = 156;
			18452: out = -253;
			18453: out = -87;
			18454: out = 195;
			18455: out = 354;
			18456: out = -248;
			18457: out = -308;
			18458: out = -237;
			18459: out = 142;
			18460: out = 105;
			18461: out = 283;
			18462: out = 86;
			18463: out = -854;
			18464: out = -633;
			18465: out = -203;
			18466: out = 104;
			18467: out = 415;
			18468: out = 22;
			18469: out = -363;
			18470: out = 102;
			18471: out = -111;
			18472: out = -36;
			18473: out = -68;
			18474: out = 118;
			18475: out = -183;
			18476: out = -293;
			18477: out = -83;
			18478: out = 236;
			18479: out = 172;
			18480: out = -100;
			18481: out = -58;
			18482: out = 209;
			18483: out = 350;
			18484: out = -120;
			18485: out = -90;
			18486: out = 9;
			18487: out = 178;
			18488: out = 37;
			18489: out = -200;
			18490: out = -282;
			18491: out = 97;
			18492: out = -44;
			18493: out = -102;
			18494: out = -212;
			18495: out = 23;
			18496: out = -49;
			18497: out = -82;
			18498: out = -26;
			18499: out = -4;
			18500: out = 62;
			18501: out = 82;
			18502: out = 503;
			18503: out = 129;
			18504: out = -130;
			18505: out = 82;
			18506: out = -167;
			18507: out = -322;
			18508: out = -272;
			18509: out = 240;
			18510: out = 333;
			18511: out = 98;
			18512: out = -354;
			18513: out = -495;
			18514: out = -103;
			18515: out = 446;
			18516: out = -125;
			18517: out = -166;
			18518: out = -227;
			18519: out = -58;
			18520: out = -26;
			18521: out = 24;
			18522: out = -41;
			18523: out = 536;
			18524: out = 107;
			18525: out = -137;
			18526: out = -237;
			18527: out = 228;
			18528: out = 169;
			18529: out = -19;
			18530: out = -144;
			18531: out = 95;
			18532: out = 121;
			18533: out = 56;
			18534: out = -459;
			18535: out = -85;
			18536: out = 463;
			18537: out = 576;
			18538: out = -138;
			18539: out = -506;
			18540: out = -10;
			18541: out = -246;
			18542: out = -426;
			18543: out = -616;
			18544: out = -224;
			18545: out = 102;
			18546: out = 430;
			18547: out = 460;
			18548: out = -4;
			18549: out = -282;
			18550: out = -374;
			18551: out = -209;
			18552: out = -372;
			18553: out = -110;
			18554: out = 440;
			18555: out = -32;
			18556: out = -341;
			18557: out = -444;
			18558: out = -106;
			18559: out = 292;
			18560: out = 316;
			18561: out = -68;
			18562: out = -416;
			18563: out = -397;
			18564: out = -70;
			18565: out = 281;
			18566: out = 50;
			18567: out = -97;
			18568: out = -22;
			18569: out = 135;
			18570: out = 142;
			18571: out = 18;
			18572: out = 54;
			18573: out = -147;
			18574: out = -310;
			18575: out = -328;
			18576: out = -16;
			18577: out = 136;
			18578: out = 131;
			18579: out = -65;
			18580: out = -62;
			18581: out = -32;
			18582: out = -95;
			18583: out = 101;
			18584: out = -256;
			18585: out = -498;
			18586: out = -325;
			18587: out = -6;
			18588: out = 110;
			18589: out = 60;
			18590: out = -44;
			18591: out = 25;
			18592: out = 113;
			18593: out = 184;
			18594: out = -237;
			18595: out = -380;
			18596: out = -233;
			18597: out = 609;
			18598: out = 285;
			18599: out = -33;
			18600: out = 99;
			18601: out = -63;
			18602: out = -129;
			18603: out = -225;
			18604: out = 24;
			18605: out = -9;
			18606: out = -287;
			18607: out = -1055;
			18608: out = -120;
			18609: out = 266;
			18610: out = 379;
			18611: out = -212;
			18612: out = -130;
			18613: out = 48;
			18614: out = 469;
			18615: out = 48;
			18616: out = 74;
			18617: out = 48;
			18618: out = 360;
			18619: out = -369;
			18620: out = -479;
			18621: out = 83;
			18622: out = 476;
			18623: out = 124;
			18624: out = -429;
			18625: out = -53;
			18626: out = -20;
			18627: out = 99;
			18628: out = 32;
			18629: out = -78;
			18630: out = -47;
			18631: out = 0;
			18632: out = -229;
			18633: out = -236;
			18634: out = -88;
			18635: out = 221;
			18636: out = 59;
			18637: out = 51;
			18638: out = -49;
			18639: out = -482;
			18640: out = -99;
			18641: out = 59;
			18642: out = 11;
			18643: out = -46;
			18644: out = 84;
			18645: out = 137;
			18646: out = -84;
			18647: out = -291;
			18648: out = -210;
			18649: out = 82;
			18650: out = 575;
			18651: out = 240;
			18652: out = -159;
			18653: out = 222;
			18654: out = 50;
			18655: out = -20;
			18656: out = -241;
			18657: out = 260;
			18658: out = 135;
			18659: out = -120;
			18660: out = -472;
			18661: out = -292;
			18662: out = -132;
			18663: out = -46;
			18664: out = 68;
			18665: out = -44;
			18666: out = -76;
			18667: out = 77;
			18668: out = 134;
			18669: out = 97;
			18670: out = -114;
			18671: out = -192;
			18672: out = -243;
			18673: out = -149;
			18674: out = 29;
			18675: out = 142;
			18676: out = 82;
			18677: out = -66;
			18678: out = 171;
			18679: out = 75;
			18680: out = -64;
			18681: out = -229;
			18682: out = -80;
			18683: out = -63;
			18684: out = -128;
			18685: out = -204;
			18686: out = -156;
			18687: out = -39;
			18688: out = 9;
			18689: out = 163;
			18690: out = 86;
			18691: out = -150;
			18692: out = -684;
			18693: out = -504;
			18694: out = -91;
			18695: out = 421;
			18696: out = 121;
			18697: out = 37;
			18698: out = -3;
			18699: out = -79;
			18700: out = -70;
			18701: out = -41;
			18702: out = -49;
			18703: out = 150;
			18704: out = 70;
			18705: out = -148;
			18706: out = -687;
			18707: out = -215;
			18708: out = 287;
			18709: out = 464;
			18710: out = 248;
			18711: out = 63;
			18712: out = 19;
			18713: out = 10;
			18714: out = 48;
			18715: out = -25;
			18716: out = -228;
			18717: out = -113;
			18718: out = -40;
			18719: out = 34;
			18720: out = 48;
			18721: out = 75;
			18722: out = -46;
			18723: out = -214;
			18724: out = -96;
			18725: out = 87;
			18726: out = 83;
			18727: out = -325;
			18728: out = -644;
			18729: out = -569;
			18730: out = 24;
			18731: out = 281;
			18732: out = 677;
			18733: out = 654;
			18734: out = -118;
			18735: out = -275;
			18736: out = -405;
			18737: out = -309;
			18738: out = -501;
			18739: out = -85;
			18740: out = 178;
			18741: out = -46;
			18742: out = -181;
			18743: out = 38;
			18744: out = 524;
			18745: out = -22;
			18746: out = -140;
			18747: out = -198;
			18748: out = -37;
			18749: out = 16;
			18750: out = 74;
			18751: out = 0;
			18752: out = -31;
			18753: out = -65;
			18754: out = -79;
			18755: out = -203;
			18756: out = -120;
			18757: out = 182;
			18758: out = 467;
			18759: out = -284;
			18760: out = -437;
			18761: out = -382;
			18762: out = -66;
			18763: out = -2;
			18764: out = 93;
			18765: out = 182;
			18766: out = 24;
			18767: out = 59;
			18768: out = 30;
			18769: out = -54;
			18770: out = -197;
			18771: out = -127;
			18772: out = 43;
			18773: out = 17;
			18774: out = 26;
			18775: out = 22;
			18776: out = 53;
			18777: out = 50;
			18778: out = -186;
			18779: out = -447;
			18780: out = 294;
			18781: out = 130;
			18782: out = -84;
			18783: out = -340;
			18784: out = -55;
			18785: out = 26;
			18786: out = -64;
			18787: out = -36;
			18788: out = -148;
			18789: out = -184;
			18790: out = -12;
			18791: out = -73;
			18792: out = 166;
			18793: out = 449;
			18794: out = 574;
			18795: out = 95;
			18796: out = -413;
			18797: out = -381;
			18798: out = -355;
			18799: out = 244;
			18800: out = 575;
			18801: out = 416;
			18802: out = -149;
			18803: out = -334;
			18804: out = -20;
			18805: out = 117;
			18806: out = -112;
			18807: out = -515;
			18808: out = 75;
			18809: out = -33;
			18810: out = 41;
			18811: out = -18;
			18812: out = 175;
			18813: out = 25;
			18814: out = -141;
			18815: out = -627;
			18816: out = -143;
			18817: out = 75;
			18818: out = 18;
			18819: out = -525;
			18820: out = -424;
			18821: out = -82;
			18822: out = 185;
			18823: out = 0;
			18824: out = 6;
			18825: out = 193;
			18826: out = -14;
			18827: out = -277;
			18828: out = -423;
			18829: out = 81;
			18830: out = 35;
			18831: out = 88;
			18832: out = 40;
			18833: out = -53;
			18834: out = -97;
			18835: out = 0;
			18836: out = 50;
			18837: out = 173;
			18838: out = 84;
			18839: out = -58;
			18840: out = 0;
			18841: out = -34;
			18842: out = -107;
			18843: out = 69;
			18844: out = -398;
			18845: out = -315;
			18846: out = 49;
			18847: out = 554;
			18848: out = 236;
			18849: out = -127;
			18850: out = 73;
			18851: out = -195;
			18852: out = -256;
			18853: out = -340;
			18854: out = -35;
			18855: out = -156;
			18856: out = -103;
			18857: out = 312;
			18858: out = -21;
			18859: out = -71;
			18860: out = 53;
			18861: out = 163;
			18862: out = 116;
			18863: out = 0;
			18864: out = -101;
			18865: out = -105;
			18866: out = -100;
			18867: out = -77;
			18868: out = 63;
			18869: out = -118;
			18870: out = -218;
			18871: out = -55;
			18872: out = -75;
			18873: out = -33;
			18874: out = -25;
			18875: out = 512;
			18876: out = -46;
			18877: out = -414;
			18878: out = -276;
			18879: out = 51;
			18880: out = 271;
			18881: out = 259;
			18882: out = 391;
			18883: out = 131;
			18884: out = -118;
			18885: out = -387;
			18886: out = -91;
			18887: out = -29;
			18888: out = -39;
			18889: out = -621;
			18890: out = -165;
			18891: out = 96;
			18892: out = 169;
			18893: out = -84;
			18894: out = -4;
			18895: out = 13;
			18896: out = -193;
			18897: out = -353;
			18898: out = -81;
			18899: out = 395;
			18900: out = 144;
			18901: out = -433;
			18902: out = -765;
			18903: out = 103;
			18904: out = 230;
			18905: out = 122;
			18906: out = -376;
			18907: out = 27;
			18908: out = 19;
			18909: out = 53;
			18910: out = 51;
			18911: out = 55;
			18912: out = -65;
			18913: out = -208;
			18914: out = -191;
			18915: out = -121;
			18916: out = 59;
			18917: out = 367;
			18918: out = 158;
			18919: out = -65;
			18920: out = -207;
			18921: out = -435;
			18922: out = -242;
			18923: out = 34;
			18924: out = 390;
			18925: out = 26;
			18926: out = -122;
			18927: out = -18;
			18928: out = 494;
			18929: out = 481;
			18930: out = 197;
			18931: out = -224;
			18932: out = -22;
			18933: out = -19;
			18934: out = -246;
			18935: out = -60;
			18936: out = -13;
			18937: out = 73;
			18938: out = -28;
			18939: out = -33;
			18940: out = -101;
			18941: out = -66;
			18942: out = -22;
			18943: out = 122;
			18944: out = 92;
			18945: out = 62;
			18946: out = -449;
			18947: out = -462;
			18948: out = -113;
			18949: out = 113;
			18950: out = 124;
			18951: out = 0;
			18952: out = -61;
			18953: out = 30;
			18954: out = 1;
			18955: out = -115;
			18956: out = -55;
			18957: out = -7;
			18958: out = -73;
			18959: out = -461;
			18960: out = 146;
			18961: out = 381;
			18962: out = 364;
			18963: out = -415;
			18964: out = -195;
			18965: out = 63;
			18966: out = -150;
			18967: out = 314;
			18968: out = 150;
			18969: out = -173;
			18970: out = -432;
			18971: out = -76;
			18972: out = 250;
			18973: out = 206;
			18974: out = -96;
			18975: out = -375;
			18976: out = -359;
			18977: out = 129;
			18978: out = 166;
			18979: out = 113;
			18980: out = 36;
			18981: out = -61;
			18982: out = -232;
			18983: out = -337;
			18984: out = -435;
			18985: out = -108;
			18986: out = 184;
			18987: out = 363;
			18988: out = -242;
			18989: out = -219;
			18990: out = 94;
			18991: out = 20;
			18992: out = -13;
			18993: out = -243;
			18994: out = -425;
			18995: out = -110;
			18996: out = 50;
			18997: out = 34;
			18998: out = -50;
			18999: out = -86;
			19000: out = -42;
			19001: out = 37;
			19002: out = 50;
			19003: out = 117;
			19004: out = 145;
			19005: out = -56;
			19006: out = 25;
			19007: out = -14;
			19008: out = -238;
			19009: out = 15;
			19010: out = 30;
			19011: out = 30;
			19012: out = -366;
			19013: out = 141;
			19014: out = 332;
			19015: out = 320;
			19016: out = -519;
			19017: out = -294;
			19018: out = 157;
			19019: out = 337;
			19020: out = 50;
			19021: out = -176;
			19022: out = -47;
			19023: out = 6;
			19024: out = 17;
			19025: out = -112;
			19026: out = -35;
			19027: out = -194;
			19028: out = -261;
			19029: out = -328;
			19030: out = 60;
			19031: out = -20;
			19032: out = -4;
			19033: out = 152;
			19034: out = 23;
			19035: out = -200;
			19036: out = -313;
			19037: out = -122;
			19038: out = -45;
			19039: out = -160;
			19040: out = -159;
			19041: out = -465;
			19042: out = -19;
			19043: out = 511;
			19044: out = 67;
			19045: out = -444;
			19046: out = -530;
			19047: out = 400;
			19048: out = 60;
			19049: out = 85;
			19050: out = 0;
			19051: out = 59;
			19052: out = -8;
			19053: out = 47;
			19054: out = -85;
			19055: out = 86;
			19056: out = -79;
			19057: out = -140;
			19058: out = 229;
			19059: out = 466;
			19060: out = 184;
			19061: out = -630;
			19062: out = -376;
			19063: out = -41;
			19064: out = 317;
			19065: out = -144;
			19066: out = 4;
			19067: out = 17;
			19068: out = 90;
			19069: out = -207;
			19070: out = 9;
			19071: out = 288;
			19072: out = 6;
			19073: out = -138;
			19074: out = -195;
			19075: out = -15;
			19076: out = -20;
			19077: out = 8;
			19078: out = -58;
			19079: out = 204;
			19080: out = 25;
			19081: out = 107;
			19082: out = 229;
			19083: out = 206;
			19084: out = -176;
			19085: out = -475;
			19086: out = -193;
			19087: out = -145;
			19088: out = -89;
			19089: out = -88;
			19090: out = -208;
			19091: out = -10;
			19092: out = 165;
			19093: out = -73;
			19094: out = -60;
			19095: out = -66;
			19096: out = 69;
			19097: out = -66;
			19098: out = -259;
			19099: out = -415;
			19100: out = -43;
			19101: out = 58;
			19102: out = 370;
			19103: out = 492;
			19104: out = 238;
			19105: out = -343;
			19106: out = -631;
			19107: out = 4;
			19108: out = -74;
			19109: out = -35;
			19110: out = -107;
			19111: out = 79;
			19112: out = 21;
			19113: out = 11;
			19114: out = -118;
			19115: out = 137;
			19116: out = 3;
			19117: out = -229;
			19118: out = -425;
			19119: out = -137;
			19120: out = 159;
			19121: out = 353;
			19122: out = -225;
			19123: out = -492;
			19124: out = -341;
			19125: out = 15;
			19126: out = 75;
			19127: out = 30;
			19128: out = 76;
			19129: out = 147;
			19130: out = 88;
			19131: out = -98;
			19132: out = -281;
			19133: out = -120;
			19134: out = 94;
			19135: out = 43;
			19136: out = 65;
			19137: out = 89;
			19138: out = 177;
			19139: out = 4;
			19140: out = -36;
			19141: out = -180;
			19142: out = -284;
			19143: out = -154;
			19144: out = 143;
			19145: out = 339;
			19146: out = -46;
			19147: out = -143;
			19148: out = -105;
			19149: out = 311;
			19150: out = -161;
			19151: out = -103;
			19152: out = 49;
			19153: out = 383;
			19154: out = -109;
			19155: out = -258;
			19156: out = 201;
			19157: out = -69;
			19158: out = -212;
			19159: out = -294;
			19160: out = 66;
			19161: out = 230;
			19162: out = 334;
			19163: out = 69;
			19164: out = 116;
			19165: out = -228;
			19166: out = -424;
			19167: out = -222;
			19168: out = -33;
			19169: out = 121;
			19170: out = 252;
			19171: out = -52;
			19172: out = -169;
			19173: out = -204;
			19174: out = -45;
			19175: out = -265;
			19176: out = -219;
			19177: out = 79;
			19178: out = -166;
			19179: out = -393;
			19180: out = -504;
			19181: out = 74;
			19182: out = -76;
			19183: out = -86;
			19184: out = -189;
			19185: out = 524;
			19186: out = 376;
			19187: out = 19;
			19188: out = -430;
			19189: out = -110;
			19190: out = 90;
			19191: out = 28;
			19192: out = -55;
			19193: out = -80;
			19194: out = -18;
			19195: out = 17;
			19196: out = -41;
			19197: out = 138;
			19198: out = 591;
			19199: out = -196;
			19200: out = -140;
			19201: out = -75;
			19202: out = 198;
			19203: out = -326;
			19204: out = -329;
			19205: out = -29;
			19206: out = 446;
			19207: out = 73;
			19208: out = -242;
			19209: out = 35;
			19210: out = 127;
			19211: out = -8;
			19212: out = -384;
			19213: out = -290;
			19214: out = -186;
			19215: out = 19;
			19216: out = 35;
			19217: out = 64;
			19218: out = 114;
			19219: out = 262;
			19220: out = 11;
			19221: out = 12;
			19222: out = -50;
			19223: out = -205;
			19224: out = 67;
			19225: out = 217;
			19226: out = 202;
			19227: out = -76;
			19228: out = -101;
			19229: out = -55;
			19230: out = -78;
			19231: out = 14;
			19232: out = -137;
			19233: out = -337;
			19234: out = -104;
			19235: out = -109;
			19236: out = -56;
			19237: out = 56;
			19238: out = -26;
			19239: out = -143;
			19240: out = -186;
			19241: out = -64;
			19242: out = 215;
			19243: out = 310;
			19244: out = -15;
			19245: out = 58;
			19246: out = -127;
			19247: out = -228;
			19248: out = -338;
			19249: out = -53;
			19250: out = 41;
			19251: out = -75;
			19252: out = -52;
			19253: out = -82;
			19254: out = -87;
			19255: out = -48;
			19256: out = -6;
			19257: out = 25;
			19258: out = 48;
			19259: out = 329;
			19260: out = 218;
			19261: out = -64;
			19262: out = -429;
			19263: out = -323;
			19264: out = -88;
			19265: out = 53;
			19266: out = -160;
			19267: out = -184;
			19268: out = -28;
			19269: out = 31;
			19270: out = -73;
			19271: out = -370;
			19272: out = -472;
			19273: out = 32;
			19274: out = 414;
			19275: out = 342;
			19276: out = 76;
			19277: out = -470;
			19278: out = -177;
			19279: out = 602;
			19280: out = 200;
			19281: out = -240;
			19282: out = -463;
			19283: out = 425;
			19284: out = 70;
			19285: out = -80;
			19286: out = -201;
			19287: out = 124;
			19288: out = 261;
			19289: out = 231;
			19290: out = -488;
			19291: out = -93;
			19292: out = 41;
			19293: out = 23;
			19294: out = -416;
			19295: out = -200;
			19296: out = 28;
			19297: out = -235;
			19298: out = -60;
			19299: out = -82;
			19300: out = -75;
			19301: out = -208;
			19302: out = -29;
			19303: out = 67;
			19304: out = 58;
			19305: out = -23;
			19306: out = -57;
			19307: out = -116;
			19308: out = -292;
			19309: out = -208;
			19310: out = 42;
			19311: out = 137;
			19312: out = 452;
			19313: out = 169;
			19314: out = -268;
			19315: out = -539;
			19316: out = -37;
			19317: out = 289;
			19318: out = -41;
			19319: out = -402;
			19320: out = -410;
			19321: out = 0;
			default: out = 0;
		endcase
	end
endmodule
