module kick_lookup(index, out);
	input logic unsigned [14:0] index;
	output logic signed [23:0] out;
	always_comb begin
		case(index)
			0: out = 24'(0);
			1: out = 24'(0);
			2: out = 24'(308);
			3: out = 24'(3656);
			4: out = 24'(5036);
			5: out = 24'(4516);
			6: out = 24'(4908);
			7: out = 24'(5000);
			8: out = 24'(6760);
			9: out = 24'(8196);
			10: out = 24'(10456);
			11: out = 24'(12784);
			12: out = 24'(12836);
			13: out = 24'(11256);
			14: out = 24'(11808);
			15: out = 24'(11948);
			16: out = 24'(12728);
			17: out = 24'(11964);
			18: out = 24'(10660);
			19: out = 24'(11664);
			20: out = 24'(12276);
			21: out = 24'(12944);
			22: out = 24'(14272);
			23: out = 24'(16196);
			24: out = 24'(18244);
			25: out = 24'(20016);
			26: out = 24'(20652);
			27: out = 24'(22304);
			28: out = 24'(24312);
			29: out = 24'(25916);
			30: out = 24'(26308);
			31: out = 24'(24372);
			32: out = 24'(25264);
			33: out = 24'(27064);
			34: out = 24'(28364);
			35: out = 24'(28716);
			36: out = 24'(27524);
			37: out = 24'(29136);
			38: out = 24'(29436);
			39: out = 24'(29052);
			40: out = 24'(27156);
			41: out = 24'(24452);
			42: out = 24'(22824);
			43: out = 24'(22032);
			44: out = 24'(21132);
			45: out = 24'(22016);
			46: out = 24'(21580);
			47: out = 24'(19280);
			48: out = 24'(20228);
			49: out = 24'(21660);
			50: out = 24'(21324);
			51: out = 24'(20960);
			52: out = 24'(21988);
			53: out = 24'(25460);
			54: out = 24'(28132);
			55: out = 24'(29592);
			56: out = 24'(29660);
			57: out = 24'(27252);
			58: out = 24'(28096);
			59: out = 24'(32536);
			60: out = 24'(39024);
			61: out = 24'(45388);
			62: out = 24'(52316);
			63: out = 24'(55020);
			64: out = 24'(57836);
			65: out = 24'(63608);
			66: out = 24'(68824);
			67: out = 24'(72980);
			68: out = 24'(77936);
			69: out = 24'(81372);
			70: out = 24'(88344);
			71: out = 24'(92592);
			72: out = 24'(96352);
			73: out = 24'(98692);
			74: out = 24'(109800);
			75: out = 24'(128964);
			76: out = 24'(129248);
			77: out = 24'(129648);
			78: out = 24'(129108);
			79: out = 24'(129072);
			80: out = 24'(128448);
			81: out = 24'(128436);
			82: out = 24'(128216);
			83: out = 24'(128380);
			84: out = 24'(128244);
			85: out = 24'(128284);
			86: out = 24'(128088);
			87: out = 24'(128028);
			88: out = 24'(127820);
			89: out = 24'(127736);
			90: out = 24'(127596);
			91: out = 24'(127544);
			92: out = 24'(127436);
			93: out = 24'(127384);
			94: out = 24'(127276);
			95: out = 24'(127196);
			96: out = 24'(127072);
			97: out = 24'(126980);
			98: out = 24'(126864);
			99: out = 24'(126788);
			100: out = 24'(126680);
			101: out = 24'(126604);
			102: out = 24'(126516);
			103: out = 24'(126432);
			104: out = 24'(126312);
			105: out = 24'(126244);
			106: out = 24'(126116);
			107: out = 24'(126032);
			108: out = 24'(125896);
			109: out = 24'(125872);
			110: out = 24'(125672);
			111: out = 24'(125792);
			112: out = 24'(124480);
			113: out = 24'(117560);
			114: out = 24'(111816);
			115: out = 24'(105944);
			116: out = 24'(99428);
			117: out = 24'(94876);
			118: out = 24'(93244);
			119: out = 24'(91456);
			120: out = 24'(88152);
			121: out = 24'(83112);
			122: out = 24'(79788);
			123: out = 24'(77256);
			124: out = 24'(72872);
			125: out = 24'(66276);
			126: out = 24'(60392);
			127: out = 24'(54088);
			128: out = 24'(46488);
			129: out = 24'(39028);
			130: out = 24'(33692);
			131: out = 24'(30464);
			132: out = 24'(25296);
			133: out = 24'(18876);
			134: out = 24'(14376);
			135: out = 24'(8496);
			136: out = 24'(2784);
			137: out = 24'(-4932);
			138: out = 24'(-12776);
			139: out = 24'(-19036);
			140: out = 24'(-26928);
			141: out = 24'(-35084);
			142: out = 24'(-40944);
			143: out = 24'(-45172);
			144: out = 24'(-50848);
			145: out = 24'(-54800);
			146: out = 24'(-58488);
			147: out = 24'(-62804);
			148: out = 24'(-65428);
			149: out = 24'(-67552);
			150: out = 24'(-71928);
			151: out = 24'(-75724);
			152: out = 24'(-81768);
			153: out = 24'(-87928);
			154: out = 24'(-91716);
			155: out = 24'(-94352);
			156: out = 24'(-97948);
			157: out = 24'(-104312);
			158: out = 24'(-106984);
			159: out = 24'(-110780);
			160: out = 24'(-115648);
			161: out = 24'(-120156);
			162: out = 24'(-125888);
			163: out = 24'(-129952);
			164: out = 24'(-130244);
			165: out = 24'(-130336);
			166: out = 24'(-130272);
			167: out = 24'(-130208);
			168: out = 24'(-130084);
			169: out = 24'(-130008);
			170: out = 24'(-129924);
			171: out = 24'(-129812);
			172: out = 24'(-129728);
			173: out = 24'(-129688);
			174: out = 24'(-129624);
			175: out = 24'(-129512);
			176: out = 24'(-129416);
			177: out = 24'(-129320);
			178: out = 24'(-129236);
			179: out = 24'(-129136);
			180: out = 24'(-129048);
			181: out = 24'(-128956);
			182: out = 24'(-128852);
			183: out = 24'(-128752);
			184: out = 24'(-128644);
			185: out = 24'(-128548);
			186: out = 24'(-128452);
			187: out = 24'(-128348);
			188: out = 24'(-128244);
			189: out = 24'(-128160);
			190: out = 24'(-128056);
			191: out = 24'(-127952);
			192: out = 24'(-127852);
			193: out = 24'(-127736);
			194: out = 24'(-127660);
			195: out = 24'(-127540);
			196: out = 24'(-127436);
			197: out = 24'(-127336);
			198: out = 24'(-127212);
			199: out = 24'(-127120);
			200: out = 24'(-127000);
			201: out = 24'(-126892);
			202: out = 24'(-126752);
			203: out = 24'(-126604);
			204: out = 24'(-126456);
			205: out = 24'(-126372);
			206: out = 24'(-126248);
			207: out = 24'(-125936);
			208: out = 24'(-125640);
			209: out = 24'(-125224);
			210: out = 24'(-124832);
			211: out = 24'(-120900);
			212: out = 24'(-114692);
			213: out = 24'(-111144);
			214: out = 24'(-109460);
			215: out = 24'(-110404);
			216: out = 24'(-107484);
			217: out = 24'(-104488);
			218: out = 24'(-102652);
			219: out = 24'(-101060);
			220: out = 24'(-101612);
			221: out = 24'(-101596);
			222: out = 24'(-99560);
			223: out = 24'(-97092);
			224: out = 24'(-93188);
			225: out = 24'(-89008);
			226: out = 24'(-87284);
			227: out = 24'(-82868);
			228: out = 24'(-78032);
			229: out = 24'(-74284);
			230: out = 24'(-69472);
			231: out = 24'(-63464);
			232: out = 24'(-56380);
			233: out = 24'(-49884);
			234: out = 24'(-46548);
			235: out = 24'(-41424);
			236: out = 24'(-36560);
			237: out = 24'(-33860);
			238: out = 24'(-28940);
			239: out = 24'(-21308);
			240: out = 24'(-12788);
			241: out = 24'(-5256);
			242: out = 24'(-72);
			243: out = 24'(5768);
			244: out = 24'(10132);
			245: out = 24'(14896);
			246: out = 24'(18116);
			247: out = 24'(21024);
			248: out = 24'(24700);
			249: out = 24'(26496);
			250: out = 24'(29612);
			251: out = 24'(34344);
			252: out = 24'(40268);
			253: out = 24'(45184);
			254: out = 24'(51644);
			255: out = 24'(58832);
			256: out = 24'(63920);
			257: out = 24'(70324);
			258: out = 24'(76332);
			259: out = 24'(78400);
			260: out = 24'(81124);
			261: out = 24'(84104);
			262: out = 24'(88824);
			263: out = 24'(91516);
			264: out = 24'(92960);
			265: out = 24'(94108);
			266: out = 24'(95716);
			267: out = 24'(97008);
			268: out = 24'(97952);
			269: out = 24'(100060);
			270: out = 24'(102732);
			271: out = 24'(105764);
			272: out = 24'(109448);
			273: out = 24'(113672);
			274: out = 24'(117404);
			275: out = 24'(120656);
			276: out = 24'(126672);
			277: out = 24'(130408);
			278: out = 24'(130088);
			279: out = 24'(130184);
			280: out = 24'(129924);
			281: out = 24'(129920);
			282: out = 24'(129764);
			283: out = 24'(129728);
			284: out = 24'(129584);
			285: out = 24'(129520);
			286: out = 24'(129368);
			287: out = 24'(129304);
			288: out = 24'(129176);
			289: out = 24'(129088);
			290: out = 24'(128972);
			291: out = 24'(128900);
			292: out = 24'(128784);
			293: out = 24'(128712);
			294: out = 24'(128600);
			295: out = 24'(128520);
			296: out = 24'(128404);
			297: out = 24'(128316);
			298: out = 24'(128216);
			299: out = 24'(128120);
			300: out = 24'(127996);
			301: out = 24'(127964);
			302: out = 24'(125596);
			303: out = 24'(121816);
			304: out = 24'(119256);
			305: out = 24'(116848);
			306: out = 24'(114116);
			307: out = 24'(110180);
			308: out = 24'(107932);
			309: out = 24'(107076);
			310: out = 24'(104756);
			311: out = 24'(103148);
			312: out = 24'(102768);
			313: out = 24'(100760);
			314: out = 24'(99512);
			315: out = 24'(98892);
			316: out = 24'(97356);
			317: out = 24'(95768);
			318: out = 24'(93032);
			319: out = 24'(92220);
			320: out = 24'(90768);
			321: out = 24'(88240);
			322: out = 24'(84856);
			323: out = 24'(81620);
			324: out = 24'(77488);
			325: out = 24'(73308);
			326: out = 24'(72004);
			327: out = 24'(72496);
			328: out = 24'(72712);
			329: out = 24'(71316);
			330: out = 24'(66956);
			331: out = 24'(66464);
			332: out = 24'(64692);
			333: out = 24'(61772);
			334: out = 24'(58444);
			335: out = 24'(51360);
			336: out = 24'(45184);
			337: out = 24'(40080);
			338: out = 24'(36960);
			339: out = 24'(34580);
			340: out = 24'(34368);
			341: out = 24'(30492);
			342: out = 24'(27556);
			343: out = 24'(26784);
			344: out = 24'(21136);
			345: out = 24'(15624);
			346: out = 24'(12444);
			347: out = 24'(7832);
			348: out = 24'(4928);
			349: out = 24'(-48);
			350: out = 24'(-5876);
			351: out = 24'(-13840);
			352: out = 24'(-19544);
			353: out = 24'(-24136);
			354: out = 24'(-28236);
			355: out = 24'(-33248);
			356: out = 24'(-39384);
			357: out = 24'(-42424);
			358: out = 24'(-46348);
			359: out = 24'(-51904);
			360: out = 24'(-57520);
			361: out = 24'(-62840);
			362: out = 24'(-65708);
			363: out = 24'(-68280);
			364: out = 24'(-72464);
			365: out = 24'(-77416);
			366: out = 24'(-78884);
			367: out = 24'(-80060);
			368: out = 24'(-82800);
			369: out = 24'(-88348);
			370: out = 24'(-91056);
			371: out = 24'(-92628);
			372: out = 24'(-96484);
			373: out = 24'(-99580);
			374: out = 24'(-103008);
			375: out = 24'(-104436);
			376: out = 24'(-105780);
			377: out = 24'(-106676);
			378: out = 24'(-110204);
			379: out = 24'(-113000);
			380: out = 24'(-117232);
			381: out = 24'(-123164);
			382: out = 24'(-127984);
			383: out = 24'(-128860);
			384: out = 24'(-128796);
			385: out = 24'(-128780);
			386: out = 24'(-128632);
			387: out = 24'(-128500);
			388: out = 24'(-128488);
			389: out = 24'(-128428);
			390: out = 24'(-128248);
			391: out = 24'(-128200);
			392: out = 24'(-128140);
			393: out = 24'(-128124);
			394: out = 24'(-128032);
			395: out = 24'(-127944);
			396: out = 24'(-127820);
			397: out = 24'(-127724);
			398: out = 24'(-127692);
			399: out = 24'(-127636);
			400: out = 24'(-127540);
			401: out = 24'(-127464);
			402: out = 24'(-127404);
			403: out = 24'(-127296);
			404: out = 24'(-127188);
			405: out = 24'(-127048);
			406: out = 24'(-126928);
			407: out = 24'(-126796);
			408: out = 24'(-126644);
			409: out = 24'(-126604);
			410: out = 24'(-126488);
			411: out = 24'(-126384);
			412: out = 24'(-126256);
			413: out = 24'(-126188);
			414: out = 24'(-125972);
			415: out = 24'(-125828);
			416: out = 24'(-125592);
			417: out = 24'(-125304);
			418: out = 24'(-125140);
			419: out = 24'(-125252);
			420: out = 24'(-124576);
			421: out = 24'(-123712);
			422: out = 24'(-121872);
			423: out = 24'(-118952);
			424: out = 24'(-115144);
			425: out = 24'(-112816);
			426: out = 24'(-112172);
			427: out = 24'(-108752);
			428: out = 24'(-108288);
			429: out = 24'(-107312);
			430: out = 24'(-106860);
			431: out = 24'(-106240);
			432: out = 24'(-104904);
			433: out = 24'(-105828);
			434: out = 24'(-105900);
			435: out = 24'(-106076);
			436: out = 24'(-106316);
			437: out = 24'(-105428);
			438: out = 24'(-102672);
			439: out = 24'(-98828);
			440: out = 24'(-93904);
			441: out = 24'(-90516);
			442: out = 24'(-89604);
			443: out = 24'(-86968);
			444: out = 24'(-82496);
			445: out = 24'(-80236);
			446: out = 24'(-78368);
			447: out = 24'(-75332);
			448: out = 24'(-71556);
			449: out = 24'(-69820);
			450: out = 24'(-67444);
			451: out = 24'(-64648);
			452: out = 24'(-64880);
			453: out = 24'(-64900);
			454: out = 24'(-62648);
			455: out = 24'(-58984);
			456: out = 24'(-55544);
			457: out = 24'(-52120);
			458: out = 24'(-51620);
			459: out = 24'(-49980);
			460: out = 24'(-45272);
			461: out = 24'(-42832);
			462: out = 24'(-39276);
			463: out = 24'(-36792);
			464: out = 24'(-34892);
			465: out = 24'(-32148);
			466: out = 24'(-29264);
			467: out = 24'(-25204);
			468: out = 24'(-20808);
			469: out = 24'(-17176);
			470: out = 24'(-14108);
			471: out = 24'(-11656);
			472: out = 24'(-6228);
			473: out = 24'(-2240);
			474: out = 24'(2344);
			475: out = 24'(5956);
			476: out = 24'(9836);
			477: out = 24'(13324);
			478: out = 24'(15924);
			479: out = 24'(20156);
			480: out = 24'(22108);
			481: out = 24'(23792);
			482: out = 24'(25124);
			483: out = 24'(28348);
			484: out = 24'(31328);
			485: out = 24'(34560);
			486: out = 24'(37744);
			487: out = 24'(40920);
			488: out = 24'(45128);
			489: out = 24'(49676);
			490: out = 24'(53412);
			491: out = 24'(56332);
			492: out = 24'(58808);
			493: out = 24'(61880);
			494: out = 24'(65400);
			495: out = 24'(68664);
			496: out = 24'(71400);
			497: out = 24'(72084);
			498: out = 24'(73000);
			499: out = 24'(75604);
			500: out = 24'(80164);
			501: out = 24'(85328);
			502: out = 24'(91728);
			503: out = 24'(95592);
			504: out = 24'(98772);
			505: out = 24'(102844);
			506: out = 24'(105472);
			507: out = 24'(105464);
			508: out = 24'(106240);
			509: out = 24'(109872);
			510: out = 24'(111948);
			511: out = 24'(114856);
			512: out = 24'(116116);
			513: out = 24'(117676);
			514: out = 24'(118964);
			515: out = 24'(120164);
			516: out = 24'(121004);
			517: out = 24'(121420);
			518: out = 24'(122700);
			519: out = 24'(125556);
			520: out = 24'(129716);
			521: out = 24'(131060);
			522: out = 24'(130908);
			523: out = 24'(130832);
			524: out = 24'(130716);
			525: out = 24'(130624);
			526: out = 24'(130516);
			527: out = 24'(130412);
			528: out = 24'(130328);
			529: out = 24'(130224);
			530: out = 24'(130116);
			531: out = 24'(130016);
			532: out = 24'(129916);
			533: out = 24'(129812);
			534: out = 24'(129724);
			535: out = 24'(129624);
			536: out = 24'(129532);
			537: out = 24'(129432);
			538: out = 24'(129336);
			539: out = 24'(129228);
			540: out = 24'(129156);
			541: out = 24'(129048);
			542: out = 24'(128952);
			543: out = 24'(128856);
			544: out = 24'(128756);
			545: out = 24'(128628);
			546: out = 24'(128564);
			547: out = 24'(128440);
			548: out = 24'(128392);
			549: out = 24'(128232);
			550: out = 24'(128256);
			551: out = 24'(127624);
			552: out = 24'(125372);
			553: out = 24'(123792);
			554: out = 24'(119952);
			555: out = 24'(117640);
			556: out = 24'(114632);
			557: out = 24'(112780);
			558: out = 24'(110492);
			559: out = 24'(108456);
			560: out = 24'(107364);
			561: out = 24'(105232);
			562: out = 24'(103628);
			563: out = 24'(103096);
			564: out = 24'(102304);
			565: out = 24'(101664);
			566: out = 24'(101420);
			567: out = 24'(99344);
			568: out = 24'(97244);
			569: out = 24'(96408);
			570: out = 24'(95220);
			571: out = 24'(92476);
			572: out = 24'(88124);
			573: out = 24'(85508);
			574: out = 24'(83380);
			575: out = 24'(81016);
			576: out = 24'(78472);
			577: out = 24'(77052);
			578: out = 24'(76532);
			579: out = 24'(75324);
			580: out = 24'(73216);
			581: out = 24'(70600);
			582: out = 24'(68888);
			583: out = 24'(67792);
			584: out = 24'(63584);
			585: out = 24'(59504);
			586: out = 24'(57188);
			587: out = 24'(54076);
			588: out = 24'(50656);
			589: out = 24'(48824);
			590: out = 24'(48016);
			591: out = 24'(47084);
			592: out = 24'(45448);
			593: out = 24'(42336);
			594: out = 24'(40216);
			595: out = 24'(39872);
			596: out = 24'(37604);
			597: out = 24'(35552);
			598: out = 24'(33356);
			599: out = 24'(29408);
			600: out = 24'(25120);
			601: out = 24'(22976);
			602: out = 24'(21516);
			603: out = 24'(19700);
			604: out = 24'(16916);
			605: out = 24'(13940);
			606: out = 24'(9972);
			607: out = 24'(6864);
			608: out = 24'(4916);
			609: out = 24'(4184);
			610: out = 24'(2264);
			611: out = 24'(-1172);
			612: out = 24'(-5316);
			613: out = 24'(-9440);
			614: out = 24'(-13352);
			615: out = 24'(-17300);
			616: out = 24'(-19448);
			617: out = 24'(-22568);
			618: out = 24'(-26340);
			619: out = 24'(-30096);
			620: out = 24'(-32820);
			621: out = 24'(-36044);
			622: out = 24'(-40584);
			623: out = 24'(-44244);
			624: out = 24'(-48772);
			625: out = 24'(-52596);
			626: out = 24'(-55924);
			627: out = 24'(-59312);
			628: out = 24'(-60904);
			629: out = 24'(-64436);
			630: out = 24'(-68072);
			631: out = 24'(-70792);
			632: out = 24'(-72884);
			633: out = 24'(-75020);
			634: out = 24'(-77156);
			635: out = 24'(-80172);
			636: out = 24'(-80996);
			637: out = 24'(-81900);
			638: out = 24'(-83888);
			639: out = 24'(-86772);
			640: out = 24'(-90612);
			641: out = 24'(-94116);
			642: out = 24'(-96788);
			643: out = 24'(-98908);
			644: out = 24'(-101312);
			645: out = 24'(-103648);
			646: out = 24'(-105016);
			647: out = 24'(-106436);
			648: out = 24'(-107780);
			649: out = 24'(-109712);
			650: out = 24'(-110988);
			651: out = 24'(-112216);
			652: out = 24'(-113476);
			653: out = 24'(-114612);
			654: out = 24'(-114864);
			655: out = 24'(-115412);
			656: out = 24'(-117296);
			657: out = 24'(-116940);
			658: out = 24'(-118296);
			659: out = 24'(-121784);
			660: out = 24'(-123496);
			661: out = 24'(-121948);
			662: out = 24'(-120400);
			663: out = 24'(-118912);
			664: out = 24'(-118956);
			665: out = 24'(-121656);
			666: out = 24'(-122980);
			667: out = 24'(-121560);
			668: out = 24'(-121924);
			669: out = 24'(-122884);
			670: out = 24'(-125696);
			671: out = 24'(-126864);
			672: out = 24'(-126792);
			673: out = 24'(-127028);
			674: out = 24'(-126956);
			675: out = 24'(-126872);
			676: out = 24'(-126620);
			677: out = 24'(-126388);
			678: out = 24'(-125960);
			679: out = 24'(-125596);
			680: out = 24'(-125552);
			681: out = 24'(-125484);
			682: out = 24'(-125492);
			683: out = 24'(-125620);
			684: out = 24'(-125452);
			685: out = 24'(-124900);
			686: out = 24'(-124576);
			687: out = 24'(-124140);
			688: out = 24'(-122428);
			689: out = 24'(-121488);
			690: out = 24'(-120324);
			691: out = 24'(-117132);
			692: out = 24'(-115484);
			693: out = 24'(-114708);
			694: out = 24'(-112808);
			695: out = 24'(-110540);
			696: out = 24'(-108904);
			697: out = 24'(-106952);
			698: out = 24'(-106384);
			699: out = 24'(-106992);
			700: out = 24'(-105604);
			701: out = 24'(-104340);
			702: out = 24'(-102924);
			703: out = 24'(-101444);
			704: out = 24'(-100416);
			705: out = 24'(-98672);
			706: out = 24'(-97972);
			707: out = 24'(-97692);
			708: out = 24'(-98724);
			709: out = 24'(-97952);
			710: out = 24'(-97100);
			711: out = 24'(-95968);
			712: out = 24'(-95592);
			713: out = 24'(-94908);
			714: out = 24'(-94412);
			715: out = 24'(-93808);
			716: out = 24'(-93108);
			717: out = 24'(-90556);
			718: out = 24'(-88708);
			719: out = 24'(-87644);
			720: out = 24'(-85512);
			721: out = 24'(-83328);
			722: out = 24'(-82200);
			723: out = 24'(-79684);
			724: out = 24'(-75772);
			725: out = 24'(-72268);
			726: out = 24'(-69444);
			727: out = 24'(-67960);
			728: out = 24'(-66800);
			729: out = 24'(-65156);
			730: out = 24'(-63396);
			731: out = 24'(-62440);
			732: out = 24'(-61688);
			733: out = 24'(-59988);
			734: out = 24'(-59020);
			735: out = 24'(-59068);
			736: out = 24'(-58584);
			737: out = 24'(-56928);
			738: out = 24'(-55168);
			739: out = 24'(-52876);
			740: out = 24'(-51516);
			741: out = 24'(-47808);
			742: out = 24'(-44984);
			743: out = 24'(-44472);
			744: out = 24'(-42028);
			745: out = 24'(-41276);
			746: out = 24'(-41780);
			747: out = 24'(-40736);
			748: out = 24'(-38104);
			749: out = 24'(-36012);
			750: out = 24'(-32776);
			751: out = 24'(-30032);
			752: out = 24'(-28556);
			753: out = 24'(-27068);
			754: out = 24'(-25200);
			755: out = 24'(-24244);
			756: out = 24'(-22552);
			757: out = 24'(-21420);
			758: out = 24'(-21840);
			759: out = 24'(-20236);
			760: out = 24'(-18636);
			761: out = 24'(-16392);
			762: out = 24'(-13608);
			763: out = 24'(-10620);
			764: out = 24'(-7972);
			765: out = 24'(-4904);
			766: out = 24'(-1476);
			767: out = 24'(1332);
			768: out = 24'(3292);
			769: out = 24'(5148);
			770: out = 24'(5768);
			771: out = 24'(7836);
			772: out = 24'(9800);
			773: out = 24'(10936);
			774: out = 24'(13276);
			775: out = 24'(16396);
			776: out = 24'(19540);
			777: out = 24'(22228);
			778: out = 24'(24964);
			779: out = 24'(27104);
			780: out = 24'(28856);
			781: out = 24'(32360);
			782: out = 24'(34544);
			783: out = 24'(36472);
			784: out = 24'(37560);
			785: out = 24'(40120);
			786: out = 24'(43196);
			787: out = 24'(44040);
			788: out = 24'(45228);
			789: out = 24'(46080);
			790: out = 24'(48032);
			791: out = 24'(50072);
			792: out = 24'(52148);
			793: out = 24'(53992);
			794: out = 24'(54648);
			795: out = 24'(55992);
			796: out = 24'(57304);
			797: out = 24'(59548);
			798: out = 24'(61352);
			799: out = 24'(62352);
			800: out = 24'(63044);
			801: out = 24'(65576);
			802: out = 24'(68572);
			803: out = 24'(71228);
			804: out = 24'(74304);
			805: out = 24'(75388);
			806: out = 24'(76092);
			807: out = 24'(78828);
			808: out = 24'(81564);
			809: out = 24'(84708);
			810: out = 24'(88168);
			811: out = 24'(89968);
			812: out = 24'(90048);
			813: out = 24'(91884);
			814: out = 24'(95128);
			815: out = 24'(96500);
			816: out = 24'(98656);
			817: out = 24'(98540);
			818: out = 24'(98780);
			819: out = 24'(100096);
			820: out = 24'(100100);
			821: out = 24'(100668);
			822: out = 24'(101524);
			823: out = 24'(103216);
			824: out = 24'(105392);
			825: out = 24'(106804);
			826: out = 24'(107884);
			827: out = 24'(109184);
			828: out = 24'(110304);
			829: out = 24'(110368);
			830: out = 24'(110972);
			831: out = 24'(112436);
			832: out = 24'(114596);
			833: out = 24'(116104);
			834: out = 24'(117660);
			835: out = 24'(119220);
			836: out = 24'(120168);
			837: out = 24'(121392);
			838: out = 24'(122852);
			839: out = 24'(124072);
			840: out = 24'(125472);
			841: out = 24'(125736);
			842: out = 24'(126076);
			843: out = 24'(126548);
			844: out = 24'(126452);
			845: out = 24'(126064);
			846: out = 24'(125712);
			847: out = 24'(124872);
			848: out = 24'(124416);
			849: out = 24'(123100);
			850: out = 24'(122384);
			851: out = 24'(121872);
			852: out = 24'(121128);
			853: out = 24'(121292);
			854: out = 24'(121200);
			855: out = 24'(119928);
			856: out = 24'(118728);
			857: out = 24'(118100);
			858: out = 24'(118492);
			859: out = 24'(117872);
			860: out = 24'(117324);
			861: out = 24'(117000);
			862: out = 24'(115876);
			863: out = 24'(114556);
			864: out = 24'(113612);
			865: out = 24'(113332);
			866: out = 24'(112108);
			867: out = 24'(110512);
			868: out = 24'(108128);
			869: out = 24'(107212);
			870: out = 24'(106348);
			871: out = 24'(105384);
			872: out = 24'(103928);
			873: out = 24'(102412);
			874: out = 24'(101884);
			875: out = 24'(100476);
			876: out = 24'(98720);
			877: out = 24'(96992);
			878: out = 24'(96272);
			879: out = 24'(96008);
			880: out = 24'(94968);
			881: out = 24'(92804);
			882: out = 24'(90352);
			883: out = 24'(89016);
			884: out = 24'(87368);
			885: out = 24'(86536);
			886: out = 24'(85232);
			887: out = 24'(84192);
			888: out = 24'(83396);
			889: out = 24'(81276);
			890: out = 24'(79768);
			891: out = 24'(77760);
			892: out = 24'(76012);
			893: out = 24'(74648);
			894: out = 24'(73296);
			895: out = 24'(72288);
			896: out = 24'(70284);
			897: out = 24'(67888);
			898: out = 24'(66204);
			899: out = 24'(64284);
			900: out = 24'(62364);
			901: out = 24'(61264);
			902: out = 24'(60420);
			903: out = 24'(58580);
			904: out = 24'(57340);
			905: out = 24'(56132);
			906: out = 24'(55064);
			907: out = 24'(53828);
			908: out = 24'(52404);
			909: out = 24'(50164);
			910: out = 24'(48784);
			911: out = 24'(48128);
			912: out = 24'(47312);
			913: out = 24'(46140);
			914: out = 24'(44972);
			915: out = 24'(43088);
			916: out = 24'(40748);
			917: out = 24'(39500);
			918: out = 24'(39660);
			919: out = 24'(39732);
			920: out = 24'(39460);
			921: out = 24'(38832);
			922: out = 24'(36564);
			923: out = 24'(34528);
			924: out = 24'(33476);
			925: out = 24'(33448);
			926: out = 24'(33584);
			927: out = 24'(32460);
			928: out = 24'(30264);
			929: out = 24'(27840);
			930: out = 24'(26660);
			931: out = 24'(26204);
			932: out = 24'(25928);
			933: out = 24'(24536);
			934: out = 24'(21856);
			935: out = 24'(20004);
			936: out = 24'(18604);
			937: out = 24'(17160);
			938: out = 24'(16284);
			939: out = 24'(14544);
			940: out = 24'(11872);
			941: out = 24'(9424);
			942: out = 24'(6976);
			943: out = 24'(5624);
			944: out = 24'(4348);
			945: out = 24'(2728);
			946: out = 24'(904);
			947: out = 24'(-1876);
			948: out = 24'(-4748);
			949: out = 24'(-7296);
			950: out = 24'(-9092);
			951: out = 24'(-11692);
			952: out = 24'(-14532);
			953: out = 24'(-16908);
			954: out = 24'(-18720);
			955: out = 24'(-20864);
			956: out = 24'(-23520);
			957: out = 24'(-26472);
			958: out = 24'(-29352);
			959: out = 24'(-31916);
			960: out = 24'(-35572);
			961: out = 24'(-39372);
			962: out = 24'(-42068);
			963: out = 24'(-44580);
			964: out = 24'(-47112);
			965: out = 24'(-49488);
			966: out = 24'(-51200);
			967: out = 24'(-53112);
			968: out = 24'(-55452);
			969: out = 24'(-57376);
			970: out = 24'(-59504);
			971: out = 24'(-61656);
			972: out = 24'(-63744);
			973: out = 24'(-65024);
			974: out = 24'(-66732);
			975: out = 24'(-68408);
			976: out = 24'(-70272);
			977: out = 24'(-71828);
			978: out = 24'(-73180);
			979: out = 24'(-74936);
			980: out = 24'(-76648);
			981: out = 24'(-78484);
			982: out = 24'(-80744);
			983: out = 24'(-82244);
			984: out = 24'(-82748);
			985: out = 24'(-82952);
			986: out = 24'(-83532);
			987: out = 24'(-85448);
			988: out = 24'(-86460);
			989: out = 24'(-86600);
			990: out = 24'(-87936);
			991: out = 24'(-88860);
			992: out = 24'(-90016);
			993: out = 24'(-91420);
			994: out = 24'(-92268);
			995: out = 24'(-92748);
			996: out = 24'(-93992);
			997: out = 24'(-94792);
			998: out = 24'(-95052);
			999: out = 24'(-96572);
			1000: out = 24'(-96832);
			1001: out = 24'(-98004);
			1002: out = 24'(-98952);
			1003: out = 24'(-99816);
			1004: out = 24'(-101692);
			1005: out = 24'(-103320);
			1006: out = 24'(-104656);
			1007: out = 24'(-105996);
			1008: out = 24'(-107012);
			1009: out = 24'(-107960);
			1010: out = 24'(-108688);
			1011: out = 24'(-108636);
			1012: out = 24'(-108976);
			1013: out = 24'(-109392);
			1014: out = 24'(-109248);
			1015: out = 24'(-109168);
			1016: out = 24'(-109588);
			1017: out = 24'(-109680);
			1018: out = 24'(-109752);
			1019: out = 24'(-110876);
			1020: out = 24'(-112028);
			1021: out = 24'(-111876);
			1022: out = 24'(-111500);
			1023: out = 24'(-111956);
			1024: out = 24'(-111924);
			1025: out = 24'(-111636);
			1026: out = 24'(-112924);
			1027: out = 24'(-113244);
			1028: out = 24'(-113244);
			1029: out = 24'(-112980);
			1030: out = 24'(-113124);
			1031: out = 24'(-113776);
			1032: out = 24'(-113936);
			1033: out = 24'(-114476);
			1034: out = 24'(-115364);
			1035: out = 24'(-115520);
			1036: out = 24'(-115212);
			1037: out = 24'(-114584);
			1038: out = 24'(-113492);
			1039: out = 24'(-113432);
			1040: out = 24'(-114012);
			1041: out = 24'(-112784);
			1042: out = 24'(-111768);
			1043: out = 24'(-111208);
			1044: out = 24'(-110748);
			1045: out = 24'(-110128);
			1046: out = 24'(-109084);
			1047: out = 24'(-108972);
			1048: out = 24'(-108476);
			1049: out = 24'(-108144);
			1050: out = 24'(-107124);
			1051: out = 24'(-105476);
			1052: out = 24'(-104340);
			1053: out = 24'(-102868);
			1054: out = 24'(-102272);
			1055: out = 24'(-101716);
			1056: out = 24'(-100880);
			1057: out = 24'(-100268);
			1058: out = 24'(-99768);
			1059: out = 24'(-98760);
			1060: out = 24'(-98148);
			1061: out = 24'(-96812);
			1062: out = 24'(-95548);
			1063: out = 24'(-94580);
			1064: out = 24'(-93712);
			1065: out = 24'(-93132);
			1066: out = 24'(-91760);
			1067: out = 24'(-90152);
			1068: out = 24'(-88284);
			1069: out = 24'(-86260);
			1070: out = 24'(-84328);
			1071: out = 24'(-83292);
			1072: out = 24'(-81976);
			1073: out = 24'(-80456);
			1074: out = 24'(-79616);
			1075: out = 24'(-79088);
			1076: out = 24'(-78560);
			1077: out = 24'(-77496);
			1078: out = 24'(-75800);
			1079: out = 24'(-74636);
			1080: out = 24'(-73804);
			1081: out = 24'(-73640);
			1082: out = 24'(-72864);
			1083: out = 24'(-72452);
			1084: out = 24'(-72180);
			1085: out = 24'(-71672);
			1086: out = 24'(-70876);
			1087: out = 24'(-69832);
			1088: out = 24'(-69028);
			1089: out = 24'(-68232);
			1090: out = 24'(-66824);
			1091: out = 24'(-65628);
			1092: out = 24'(-65016);
			1093: out = 24'(-64320);
			1094: out = 24'(-63384);
			1095: out = 24'(-62564);
			1096: out = 24'(-62044);
			1097: out = 24'(-60856);
			1098: out = 24'(-59112);
			1099: out = 24'(-57972);
			1100: out = 24'(-56980);
			1101: out = 24'(-56044);
			1102: out = 24'(-54184);
			1103: out = 24'(-52252);
			1104: out = 24'(-50428);
			1105: out = 24'(-48840);
			1106: out = 24'(-47232);
			1107: out = 24'(-45732);
			1108: out = 24'(-44576);
			1109: out = 24'(-43396);
			1110: out = 24'(-41920);
			1111: out = 24'(-40964);
			1112: out = 24'(-40108);
			1113: out = 24'(-39180);
			1114: out = 24'(-37552);
			1115: out = 24'(-36272);
			1116: out = 24'(-35272);
			1117: out = 24'(-34596);
			1118: out = 24'(-34304);
			1119: out = 24'(-33336);
			1120: out = 24'(-31876);
			1121: out = 24'(-30976);
			1122: out = 24'(-29780);
			1123: out = 24'(-28396);
			1124: out = 24'(-27528);
			1125: out = 24'(-26520);
			1126: out = 24'(-24688);
			1127: out = 24'(-24392);
			1128: out = 24'(-23560);
			1129: out = 24'(-22600);
			1130: out = 24'(-22248);
			1131: out = 24'(-21968);
			1132: out = 24'(-21516);
			1133: out = 24'(-20368);
			1134: out = 24'(-19448);
			1135: out = 24'(-18820);
			1136: out = 24'(-17924);
			1137: out = 24'(-17312);
			1138: out = 24'(-16252);
			1139: out = 24'(-15016);
			1140: out = 24'(-13544);
			1141: out = 24'(-12184);
			1142: out = 24'(-11064);
			1143: out = 24'(-10024);
			1144: out = 24'(-8604);
			1145: out = 24'(-6980);
			1146: out = 24'(-5756);
			1147: out = 24'(-4180);
			1148: out = 24'(-3024);
			1149: out = 24'(-1536);
			1150: out = 24'(196);
			1151: out = 24'(1888);
			1152: out = 24'(3192);
			1153: out = 24'(4540);
			1154: out = 24'(5776);
			1155: out = 24'(6948);
			1156: out = 24'(7756);
			1157: out = 24'(8216);
			1158: out = 24'(9472);
			1159: out = 24'(11060);
			1160: out = 24'(12760);
			1161: out = 24'(14668);
			1162: out = 24'(16984);
			1163: out = 24'(18952);
			1164: out = 24'(20808);
			1165: out = 24'(22744);
			1166: out = 24'(24968);
			1167: out = 24'(25968);
			1168: out = 24'(27336);
			1169: out = 24'(29448);
			1170: out = 24'(30916);
			1171: out = 24'(32156);
			1172: out = 24'(33872);
			1173: out = 24'(35992);
			1174: out = 24'(37276);
			1175: out = 24'(38644);
			1176: out = 24'(40504);
			1177: out = 24'(41680);
			1178: out = 24'(43032);
			1179: out = 24'(44320);
			1180: out = 24'(45376);
			1181: out = 24'(46980);
			1182: out = 24'(47800);
			1183: out = 24'(48472);
			1184: out = 24'(49784);
			1185: out = 24'(51044);
			1186: out = 24'(52488);
			1187: out = 24'(53988);
			1188: out = 24'(55512);
			1189: out = 24'(57424);
			1190: out = 24'(58744);
			1191: out = 24'(59656);
			1192: out = 24'(60516);
			1193: out = 24'(61408);
			1194: out = 24'(62500);
			1195: out = 24'(63484);
			1196: out = 24'(65100);
			1197: out = 24'(66388);
			1198: out = 24'(67412);
			1199: out = 24'(68236);
			1200: out = 24'(69872);
			1201: out = 24'(71084);
			1202: out = 24'(71872);
			1203: out = 24'(72568);
			1204: out = 24'(73520);
			1205: out = 24'(74812);
			1206: out = 24'(75984);
			1207: out = 24'(77128);
			1208: out = 24'(77784);
			1209: out = 24'(78996);
			1210: out = 24'(79904);
			1211: out = 24'(80660);
			1212: out = 24'(81428);
			1213: out = 24'(82036);
			1214: out = 24'(83004);
			1215: out = 24'(83924);
			1216: out = 24'(84948);
			1217: out = 24'(85848);
			1218: out = 24'(87088);
			1219: out = 24'(88204);
			1220: out = 24'(88700);
			1221: out = 24'(89332);
			1222: out = 24'(90288);
			1223: out = 24'(91596);
			1224: out = 24'(92844);
			1225: out = 24'(93936);
			1226: out = 24'(94292);
			1227: out = 24'(94884);
			1228: out = 24'(96200);
			1229: out = 24'(97440);
			1230: out = 24'(98620);
			1231: out = 24'(99308);
			1232: out = 24'(99792);
			1233: out = 24'(100112);
			1234: out = 24'(100784);
			1235: out = 24'(101296);
			1236: out = 24'(102196);
			1237: out = 24'(103236);
			1238: out = 24'(103948);
			1239: out = 24'(104644);
			1240: out = 24'(105180);
			1241: out = 24'(105256);
			1242: out = 24'(105640);
			1243: out = 24'(106636);
			1244: out = 24'(107032);
			1245: out = 24'(107424);
			1246: out = 24'(107804);
			1247: out = 24'(108232);
			1248: out = 24'(108620);
			1249: out = 24'(109240);
			1250: out = 24'(109972);
			1251: out = 24'(110740);
			1252: out = 24'(111488);
			1253: out = 24'(111584);
			1254: out = 24'(111324);
			1255: out = 24'(111400);
			1256: out = 24'(111488);
			1257: out = 24'(111640);
			1258: out = 24'(111568);
			1259: out = 24'(110956);
			1260: out = 24'(110388);
			1261: out = 24'(110412);
			1262: out = 24'(110304);
			1263: out = 24'(110060);
			1264: out = 24'(109316);
			1265: out = 24'(108456);
			1266: out = 24'(107896);
			1267: out = 24'(107052);
			1268: out = 24'(106068);
			1269: out = 24'(105440);
			1270: out = 24'(104724);
			1271: out = 24'(104096);
			1272: out = 24'(103648);
			1273: out = 24'(103048);
			1274: out = 24'(102160);
			1275: out = 24'(101300);
			1276: out = 24'(100976);
			1277: out = 24'(100260);
			1278: out = 24'(99088);
			1279: out = 24'(98048);
			1280: out = 24'(97408);
			1281: out = 24'(96652);
			1282: out = 24'(96236);
			1283: out = 24'(95856);
			1284: out = 24'(95232);
			1285: out = 24'(94512);
			1286: out = 24'(93600);
			1287: out = 24'(92580);
			1288: out = 24'(91332);
			1289: out = 24'(90332);
			1290: out = 24'(89380);
			1291: out = 24'(88376);
			1292: out = 24'(86940);
			1293: out = 24'(85608);
			1294: out = 24'(84728);
			1295: out = 24'(83796);
			1296: out = 24'(82800);
			1297: out = 24'(81900);
			1298: out = 24'(80876);
			1299: out = 24'(79996);
			1300: out = 24'(79228);
			1301: out = 24'(78420);
			1302: out = 24'(77428);
			1303: out = 24'(76272);
			1304: out = 24'(75288);
			1305: out = 24'(73968);
			1306: out = 24'(72640);
			1307: out = 24'(71704);
			1308: out = 24'(70864);
			1309: out = 24'(69988);
			1310: out = 24'(69412);
			1311: out = 24'(68772);
			1312: out = 24'(68032);
			1313: out = 24'(67324);
			1314: out = 24'(66664);
			1315: out = 24'(65636);
			1316: out = 24'(64408);
			1317: out = 24'(63364);
			1318: out = 24'(62504);
			1319: out = 24'(61904);
			1320: out = 24'(61216);
			1321: out = 24'(60276);
			1322: out = 24'(59080);
			1323: out = 24'(58216);
			1324: out = 24'(57412);
			1325: out = 24'(56412);
			1326: out = 24'(55312);
			1327: out = 24'(54212);
			1328: out = 24'(53428);
			1329: out = 24'(52772);
			1330: out = 24'(51976);
			1331: out = 24'(51152);
			1332: out = 24'(49956);
			1333: out = 24'(48888);
			1334: out = 24'(47656);
			1335: out = 24'(46288);
			1336: out = 24'(45068);
			1337: out = 24'(43840);
			1338: out = 24'(42476);
			1339: out = 24'(41376);
			1340: out = 24'(40348);
			1341: out = 24'(39128);
			1342: out = 24'(37980);
			1343: out = 24'(36904);
			1344: out = 24'(36056);
			1345: out = 24'(35248);
			1346: out = 24'(34500);
			1347: out = 24'(33492);
			1348: out = 24'(32484);
			1349: out = 24'(31596);
			1350: out = 24'(30768);
			1351: out = 24'(30088);
			1352: out = 24'(29216);
			1353: out = 24'(28524);
			1354: out = 24'(27448);
			1355: out = 24'(26292);
			1356: out = 24'(25568);
			1357: out = 24'(24768);
			1358: out = 24'(23796);
			1359: out = 24'(22992);
			1360: out = 24'(22076);
			1361: out = 24'(20796);
			1362: out = 24'(19860);
			1363: out = 24'(19032);
			1364: out = 24'(18452);
			1365: out = 24'(17768);
			1366: out = 24'(16556);
			1367: out = 24'(15448);
			1368: out = 24'(14428);
			1369: out = 24'(13504);
			1370: out = 24'(12716);
			1371: out = 24'(12136);
			1372: out = 24'(11540);
			1373: out = 24'(10732);
			1374: out = 24'(9572);
			1375: out = 24'(8476);
			1376: out = 24'(7452);
			1377: out = 24'(6372);
			1378: out = 24'(5320);
			1379: out = 24'(4536);
			1380: out = 24'(3960);
			1381: out = 24'(3304);
			1382: out = 24'(2524);
			1383: out = 24'(1564);
			1384: out = 24'(292);
			1385: out = 24'(-952);
			1386: out = 24'(-1948);
			1387: out = 24'(-2820);
			1388: out = 24'(-3936);
			1389: out = 24'(-5132);
			1390: out = 24'(-6088);
			1391: out = 24'(-6844);
			1392: out = 24'(-7784);
			1393: out = 24'(-8644);
			1394: out = 24'(-9800);
			1395: out = 24'(-11484);
			1396: out = 24'(-12868);
			1397: out = 24'(-14112);
			1398: out = 24'(-15568);
			1399: out = 24'(-17000);
			1400: out = 24'(-18408);
			1401: out = 24'(-19644);
			1402: out = 24'(-20652);
			1403: out = 24'(-21880);
			1404: out = 24'(-23472);
			1405: out = 24'(-25176);
			1406: out = 24'(-26216);
			1407: out = 24'(-27392);
			1408: out = 24'(-28820);
			1409: out = 24'(-30488);
			1410: out = 24'(-32296);
			1411: out = 24'(-33924);
			1412: out = 24'(-35624);
			1413: out = 24'(-37560);
			1414: out = 24'(-39124);
			1415: out = 24'(-40436);
			1416: out = 24'(-41968);
			1417: out = 24'(-43340);
			1418: out = 24'(-44788);
			1419: out = 24'(-46396);
			1420: out = 24'(-48068);
			1421: out = 24'(-49468);
			1422: out = 24'(-50576);
			1423: out = 24'(-51632);
			1424: out = 24'(-52736);
			1425: out = 24'(-54136);
			1426: out = 24'(-55544);
			1427: out = 24'(-56716);
			1428: out = 24'(-57856);
			1429: out = 24'(-59188);
			1430: out = 24'(-60496);
			1431: out = 24'(-61908);
			1432: out = 24'(-63272);
			1433: out = 24'(-64492);
			1434: out = 24'(-65420);
			1435: out = 24'(-66352);
			1436: out = 24'(-67420);
			1437: out = 24'(-68360);
			1438: out = 24'(-69428);
			1439: out = 24'(-70408);
			1440: out = 24'(-71496);
			1441: out = 24'(-72688);
			1442: out = 24'(-73748);
			1443: out = 24'(-74540);
			1444: out = 24'(-75480);
			1445: out = 24'(-76448);
			1446: out = 24'(-76996);
			1447: out = 24'(-77648);
			1448: out = 24'(-78392);
			1449: out = 24'(-79136);
			1450: out = 24'(-79968);
			1451: out = 24'(-80696);
			1452: out = 24'(-81248);
			1453: out = 24'(-82040);
			1454: out = 24'(-83036);
			1455: out = 24'(-83884);
			1456: out = 24'(-84312);
			1457: out = 24'(-84752);
			1458: out = 24'(-85444);
			1459: out = 24'(-86292);
			1460: out = 24'(-86948);
			1461: out = 24'(-87444);
			1462: out = 24'(-88160);
			1463: out = 24'(-88756);
			1464: out = 24'(-89188);
			1465: out = 24'(-89860);
			1466: out = 24'(-90392);
			1467: out = 24'(-90768);
			1468: out = 24'(-91296);
			1469: out = 24'(-91756);
			1470: out = 24'(-92232);
			1471: out = 24'(-92452);
			1472: out = 24'(-92648);
			1473: out = 24'(-92908);
			1474: out = 24'(-93168);
			1475: out = 24'(-93488);
			1476: out = 24'(-93872);
			1477: out = 24'(-94164);
			1478: out = 24'(-94156);
			1479: out = 24'(-94232);
			1480: out = 24'(-94356);
			1481: out = 24'(-94608);
			1482: out = 24'(-95004);
			1483: out = 24'(-95372);
			1484: out = 24'(-95464);
			1485: out = 24'(-95576);
			1486: out = 24'(-95652);
			1487: out = 24'(-95840);
			1488: out = 24'(-96136);
			1489: out = 24'(-96252);
			1490: out = 24'(-96412);
			1491: out = 24'(-96684);
			1492: out = 24'(-96764);
			1493: out = 24'(-96988);
			1494: out = 24'(-97200);
			1495: out = 24'(-97272);
			1496: out = 24'(-97156);
			1497: out = 24'(-96760);
			1498: out = 24'(-96948);
			1499: out = 24'(-97168);
			1500: out = 24'(-97164);
			1501: out = 24'(-97516);
			1502: out = 24'(-97924);
			1503: out = 24'(-98124);
			1504: out = 24'(-97996);
			1505: out = 24'(-97764);
			1506: out = 24'(-97704);
			1507: out = 24'(-97844);
			1508: out = 24'(-97856);
			1509: out = 24'(-97848);
			1510: out = 24'(-98084);
			1511: out = 24'(-98372);
			1512: out = 24'(-98436);
			1513: out = 24'(-98316);
			1514: out = 24'(-98132);
			1515: out = 24'(-97848);
			1516: out = 24'(-97500);
			1517: out = 24'(-97376);
			1518: out = 24'(-97340);
			1519: out = 24'(-96944);
			1520: out = 24'(-96348);
			1521: out = 24'(-95764);
			1522: out = 24'(-95304);
			1523: out = 24'(-94960);
			1524: out = 24'(-94484);
			1525: out = 24'(-93916);
			1526: out = 24'(-93404);
			1527: out = 24'(-92792);
			1528: out = 24'(-92180);
			1529: out = 24'(-91844);
			1530: out = 24'(-91432);
			1531: out = 24'(-90872);
			1532: out = 24'(-90180);
			1533: out = 24'(-89464);
			1534: out = 24'(-88756);
			1535: out = 24'(-88036);
			1536: out = 24'(-87388);
			1537: out = 24'(-86704);
			1538: out = 24'(-85844);
			1539: out = 24'(-85064);
			1540: out = 24'(-84400);
			1541: out = 24'(-83688);
			1542: out = 24'(-82908);
			1543: out = 24'(-82052);
			1544: out = 24'(-81196);
			1545: out = 24'(-80192);
			1546: out = 24'(-79280);
			1547: out = 24'(-78216);
			1548: out = 24'(-77252);
			1549: out = 24'(-76452);
			1550: out = 24'(-75700);
			1551: out = 24'(-74960);
			1552: out = 24'(-73940);
			1553: out = 24'(-72804);
			1554: out = 24'(-71764);
			1555: out = 24'(-70888);
			1556: out = 24'(-70028);
			1557: out = 24'(-69212);
			1558: out = 24'(-68344);
			1559: out = 24'(-67424);
			1560: out = 24'(-66592);
			1561: out = 24'(-65832);
			1562: out = 24'(-65116);
			1563: out = 24'(-64320);
			1564: out = 24'(-63372);
			1565: out = 24'(-62472);
			1566: out = 24'(-61652);
			1567: out = 24'(-61056);
			1568: out = 24'(-60508);
			1569: out = 24'(-59768);
			1570: out = 24'(-58988);
			1571: out = 24'(-58200);
			1572: out = 24'(-57504);
			1573: out = 24'(-56732);
			1574: out = 24'(-55864);
			1575: out = 24'(-55052);
			1576: out = 24'(-54268);
			1577: out = 24'(-53480);
			1578: out = 24'(-52940);
			1579: out = 24'(-52360);
			1580: out = 24'(-51644);
			1581: out = 24'(-51044);
			1582: out = 24'(-50384);
			1583: out = 24'(-49668);
			1584: out = 24'(-48920);
			1585: out = 24'(-48228);
			1586: out = 24'(-47596);
			1587: out = 24'(-47020);
			1588: out = 24'(-46436);
			1589: out = 24'(-45916);
			1590: out = 24'(-45384);
			1591: out = 24'(-44756);
			1592: out = 24'(-43976);
			1593: out = 24'(-43100);
			1594: out = 24'(-42432);
			1595: out = 24'(-41832);
			1596: out = 24'(-41184);
			1597: out = 24'(-40552);
			1598: out = 24'(-39876);
			1599: out = 24'(-38980);
			1600: out = 24'(-38080);
			1601: out = 24'(-37144);
			1602: out = 24'(-36212);
			1603: out = 24'(-35364);
			1604: out = 24'(-34476);
			1605: out = 24'(-33548);
			1606: out = 24'(-32640);
			1607: out = 24'(-31864);
			1608: out = 24'(-31088);
			1609: out = 24'(-30204);
			1610: out = 24'(-29276);
			1611: out = 24'(-28428);
			1612: out = 24'(-27744);
			1613: out = 24'(-27064);
			1614: out = 24'(-26280);
			1615: out = 24'(-25504);
			1616: out = 24'(-24748);
			1617: out = 24'(-24000);
			1618: out = 24'(-23252);
			1619: out = 24'(-22660);
			1620: out = 24'(-22084);
			1621: out = 24'(-21404);
			1622: out = 24'(-20700);
			1623: out = 24'(-19948);
			1624: out = 24'(-19284);
			1625: out = 24'(-18576);
			1626: out = 24'(-17816);
			1627: out = 24'(-17144);
			1628: out = 24'(-16560);
			1629: out = 24'(-15988);
			1630: out = 24'(-15316);
			1631: out = 24'(-14620);
			1632: out = 24'(-13888);
			1633: out = 24'(-13236);
			1634: out = 24'(-12548);
			1635: out = 24'(-11824);
			1636: out = 24'(-11228);
			1637: out = 24'(-10496);
			1638: out = 24'(-9628);
			1639: out = 24'(-8832);
			1640: out = 24'(-8172);
			1641: out = 24'(-7528);
			1642: out = 24'(-6836);
			1643: out = 24'(-6236);
			1644: out = 24'(-5596);
			1645: out = 24'(-4892);
			1646: out = 24'(-4252);
			1647: out = 24'(-3680);
			1648: out = 24'(-3040);
			1649: out = 24'(-2444);
			1650: out = 24'(-1832);
			1651: out = 24'(-1152);
			1652: out = 24'(-372);
			1653: out = 24'(428);
			1654: out = 24'(1120);
			1655: out = 24'(1680);
			1656: out = 24'(2300);
			1657: out = 24'(3008);
			1658: out = 24'(3780);
			1659: out = 24'(4540);
			1660: out = 24'(5072);
			1661: out = 24'(5580);
			1662: out = 24'(6260);
			1663: out = 24'(7044);
			1664: out = 24'(7840);
			1665: out = 24'(8680);
			1666: out = 24'(9516);
			1667: out = 24'(10436);
			1668: out = 24'(11352);
			1669: out = 24'(12196);
			1670: out = 24'(13076);
			1671: out = 24'(13928);
			1672: out = 24'(14816);
			1673: out = 24'(15736);
			1674: out = 24'(16720);
			1675: out = 24'(17744);
			1676: out = 24'(18724);
			1677: out = 24'(19716);
			1678: out = 24'(20704);
			1679: out = 24'(21672);
			1680: out = 24'(22660);
			1681: out = 24'(23716);
			1682: out = 24'(24812);
			1683: out = 24'(26020);
			1684: out = 24'(26996);
			1685: out = 24'(27976);
			1686: out = 24'(29052);
			1687: out = 24'(30156);
			1688: out = 24'(31208);
			1689: out = 24'(32124);
			1690: out = 24'(32992);
			1691: out = 24'(33924);
			1692: out = 24'(34900);
			1693: out = 24'(35896);
			1694: out = 24'(36844);
			1695: out = 24'(37852);
			1696: out = 24'(38816);
			1697: out = 24'(39668);
			1698: out = 24'(40684);
			1699: out = 24'(41584);
			1700: out = 24'(42404);
			1701: out = 24'(43276);
			1702: out = 24'(44260);
			1703: out = 24'(45192);
			1704: out = 24'(46112);
			1705: out = 24'(46916);
			1706: out = 24'(47704);
			1707: out = 24'(48512);
			1708: out = 24'(49288);
			1709: out = 24'(50024);
			1710: out = 24'(50820);
			1711: out = 24'(51628);
			1712: out = 24'(52376);
			1713: out = 24'(53208);
			1714: out = 24'(53980);
			1715: out = 24'(54816);
			1716: out = 24'(55596);
			1717: out = 24'(56376);
			1718: out = 24'(57180);
			1719: out = 24'(57992);
			1720: out = 24'(58780);
			1721: out = 24'(59528);
			1722: out = 24'(60156);
			1723: out = 24'(60828);
			1724: out = 24'(61648);
			1725: out = 24'(62476);
			1726: out = 24'(63252);
			1727: out = 24'(63840);
			1728: out = 24'(64412);
			1729: out = 24'(65044);
			1730: out = 24'(65672);
			1731: out = 24'(66324);
			1732: out = 24'(66936);
			1733: out = 24'(67440);
			1734: out = 24'(67996);
			1735: out = 24'(68608);
			1736: out = 24'(69168);
			1737: out = 24'(69744);
			1738: out = 24'(70340);
			1739: out = 24'(70908);
			1740: out = 24'(71408);
			1741: out = 24'(71980);
			1742: out = 24'(72428);
			1743: out = 24'(72896);
			1744: out = 24'(73468);
			1745: out = 24'(74040);
			1746: out = 24'(74528);
			1747: out = 24'(75004);
			1748: out = 24'(75548);
			1749: out = 24'(76072);
			1750: out = 24'(76500);
			1751: out = 24'(76980);
			1752: out = 24'(77460);
			1753: out = 24'(77932);
			1754: out = 24'(78444);
			1755: out = 24'(78940);
			1756: out = 24'(79512);
			1757: out = 24'(79948);
			1758: out = 24'(80508);
			1759: out = 24'(80964);
			1760: out = 24'(81480);
			1761: out = 24'(81928);
			1762: out = 24'(82328);
			1763: out = 24'(82704);
			1764: out = 24'(83064);
			1765: out = 24'(83500);
			1766: out = 24'(83904);
			1767: out = 24'(84304);
			1768: out = 24'(84764);
			1769: out = 24'(85120);
			1770: out = 24'(85472);
			1771: out = 24'(85900);
			1772: out = 24'(86276);
			1773: out = 24'(86648);
			1774: out = 24'(86920);
			1775: out = 24'(87272);
			1776: out = 24'(87604);
			1777: out = 24'(88000);
			1778: out = 24'(88316);
			1779: out = 24'(88696);
			1780: out = 24'(88968);
			1781: out = 24'(89308);
			1782: out = 24'(89640);
			1783: out = 24'(89952);
			1784: out = 24'(90276);
			1785: out = 24'(90556);
			1786: out = 24'(90860);
			1787: out = 24'(91112);
			1788: out = 24'(91472);
			1789: out = 24'(91800);
			1790: out = 24'(92040);
			1791: out = 24'(92236);
			1792: out = 24'(92476);
			1793: out = 24'(92664);
			1794: out = 24'(92808);
			1795: out = 24'(92932);
			1796: out = 24'(93084);
			1797: out = 24'(93228);
			1798: out = 24'(93284);
			1799: out = 24'(93400);
			1800: out = 24'(93336);
			1801: out = 24'(93344);
			1802: out = 24'(93304);
			1803: out = 24'(93312);
			1804: out = 24'(93112);
			1805: out = 24'(92956);
			1806: out = 24'(92660);
			1807: out = 24'(92336);
			1808: out = 24'(92164);
			1809: out = 24'(91752);
			1810: out = 24'(91360);
			1811: out = 24'(91064);
			1812: out = 24'(90712);
			1813: out = 24'(90096);
			1814: out = 24'(89708);
			1815: out = 24'(89336);
			1816: out = 24'(88820);
			1817: out = 24'(88160);
			1818: out = 24'(87644);
			1819: out = 24'(87192);
			1820: out = 24'(86624);
			1821: out = 24'(86032);
			1822: out = 24'(85476);
			1823: out = 24'(84940);
			1824: out = 24'(84224);
			1825: out = 24'(83816);
			1826: out = 24'(83084);
			1827: out = 24'(82296);
			1828: out = 24'(81688);
			1829: out = 24'(81056);
			1830: out = 24'(80416);
			1831: out = 24'(79716);
			1832: out = 24'(79008);
			1833: out = 24'(78300);
			1834: out = 24'(77560);
			1835: out = 24'(76836);
			1836: out = 24'(76140);
			1837: out = 24'(75504);
			1838: out = 24'(74700);
			1839: out = 24'(73992);
			1840: out = 24'(73292);
			1841: out = 24'(72472);
			1842: out = 24'(71880);
			1843: out = 24'(71112);
			1844: out = 24'(70428);
			1845: out = 24'(69696);
			1846: out = 24'(68996);
			1847: out = 24'(68324);
			1848: out = 24'(67636);
			1849: out = 24'(66900);
			1850: out = 24'(66156);
			1851: out = 24'(65384);
			1852: out = 24'(64660);
			1853: out = 24'(63936);
			1854: out = 24'(63296);
			1855: out = 24'(62588);
			1856: out = 24'(61788);
			1857: out = 24'(61100);
			1858: out = 24'(60488);
			1859: out = 24'(59808);
			1860: out = 24'(59116);
			1861: out = 24'(58548);
			1862: out = 24'(57904);
			1863: out = 24'(57164);
			1864: out = 24'(56472);
			1865: out = 24'(55796);
			1866: out = 24'(55180);
			1867: out = 24'(54460);
			1868: out = 24'(53896);
			1869: out = 24'(53016);
			1870: out = 24'(52192);
			1871: out = 24'(51760);
			1872: out = 24'(51188);
			1873: out = 24'(50608);
			1874: out = 24'(50052);
			1875: out = 24'(49380);
			1876: out = 24'(48776);
			1877: out = 24'(48108);
			1878: out = 24'(47516);
			1879: out = 24'(47012);
			1880: out = 24'(46300);
			1881: out = 24'(45788);
			1882: out = 24'(45228);
			1883: out = 24'(44676);
			1884: out = 24'(44152);
			1885: out = 24'(43568);
			1886: out = 24'(43056);
			1887: out = 24'(42468);
			1888: out = 24'(41980);
			1889: out = 24'(41444);
			1890: out = 24'(40916);
			1891: out = 24'(40456);
			1892: out = 24'(39916);
			1893: out = 24'(39448);
			1894: out = 24'(38892);
			1895: out = 24'(38412);
			1896: out = 24'(37964);
			1897: out = 24'(37364);
			1898: out = 24'(36908);
			1899: out = 24'(36480);
			1900: out = 24'(36056);
			1901: out = 24'(35512);
			1902: out = 24'(35064);
			1903: out = 24'(34528);
			1904: out = 24'(34112);
			1905: out = 24'(33632);
			1906: out = 24'(33168);
			1907: out = 24'(32708);
			1908: out = 24'(32276);
			1909: out = 24'(31888);
			1910: out = 24'(31500);
			1911: out = 24'(31132);
			1912: out = 24'(30664);
			1913: out = 24'(30184);
			1914: out = 24'(29756);
			1915: out = 24'(29044);
			1916: out = 24'(28144);
			1917: out = 24'(27280);
			1918: out = 24'(26480);
			1919: out = 24'(25600);
			1920: out = 24'(24792);
			1921: out = 24'(23896);
			1922: out = 24'(23264);
			1923: out = 24'(22500);
			1924: out = 24'(21648);
			1925: out = 24'(20944);
			1926: out = 24'(20168);
			1927: out = 24'(19400);
			1928: out = 24'(18656);
			1929: out = 24'(18012);
			1930: out = 24'(17332);
			1931: out = 24'(16644);
			1932: out = 24'(15952);
			1933: out = 24'(15252);
			1934: out = 24'(14596);
			1935: out = 24'(13952);
			1936: out = 24'(13384);
			1937: out = 24'(12792);
			1938: out = 24'(12224);
			1939: out = 24'(11508);
			1940: out = 24'(10844);
			1941: out = 24'(10368);
			1942: out = 24'(9636);
			1943: out = 24'(8984);
			1944: out = 24'(8440);
			1945: out = 24'(7896);
			1946: out = 24'(7248);
			1947: out = 24'(6668);
			1948: out = 24'(6124);
			1949: out = 24'(5548);
			1950: out = 24'(4904);
			1951: out = 24'(4324);
			1952: out = 24'(3796);
			1953: out = 24'(3172);
			1954: out = 24'(2852);
			1955: out = 24'(2248);
			1956: out = 24'(1648);
			1957: out = 24'(1104);
			1958: out = 24'(452);
			1959: out = 24'(-156);
			1960: out = 24'(-704);
			1961: out = 24'(-1332);
			1962: out = 24'(-1860);
			1963: out = 24'(-2340);
			1964: out = 24'(-2944);
			1965: out = 24'(-3472);
			1966: out = 24'(-4048);
			1967: out = 24'(-4560);
			1968: out = 24'(-5084);
			1969: out = 24'(-5664);
			1970: out = 24'(-6272);
			1971: out = 24'(-6692);
			1972: out = 24'(-7232);
			1973: out = 24'(-7800);
			1974: out = 24'(-8332);
			1975: out = 24'(-8920);
			1976: out = 24'(-9384);
			1977: out = 24'(-10072);
			1978: out = 24'(-10620);
			1979: out = 24'(-11212);
			1980: out = 24'(-11800);
			1981: out = 24'(-12416);
			1982: out = 24'(-12988);
			1983: out = 24'(-13604);
			1984: out = 24'(-14208);
			1985: out = 24'(-14852);
			1986: out = 24'(-15404);
			1987: out = 24'(-15956);
			1988: out = 24'(-16692);
			1989: out = 24'(-17292);
			1990: out = 24'(-18012);
			1991: out = 24'(-18680);
			1992: out = 24'(-19428);
			1993: out = 24'(-20056);
			1994: out = 24'(-20796);
			1995: out = 24'(-21604);
			1996: out = 24'(-22328);
			1997: out = 24'(-23132);
			1998: out = 24'(-23852);
			1999: out = 24'(-24720);
			2000: out = 24'(-25452);
			2001: out = 24'(-26304);
			2002: out = 24'(-27144);
			2003: out = 24'(-28004);
			2004: out = 24'(-28904);
			2005: out = 24'(-29784);
			2006: out = 24'(-30620);
			2007: out = 24'(-31536);
			2008: out = 24'(-32500);
			2009: out = 24'(-33336);
			2010: out = 24'(-34312);
			2011: out = 24'(-35236);
			2012: out = 24'(-36224);
			2013: out = 24'(-37240);
			2014: out = 24'(-38124);
			2015: out = 24'(-39080);
			2016: out = 24'(-40048);
			2017: out = 24'(-41056);
			2018: out = 24'(-42040);
			2019: out = 24'(-43036);
			2020: out = 24'(-43956);
			2021: out = 24'(-44940);
			2022: out = 24'(-45896);
			2023: out = 24'(-46808);
			2024: out = 24'(-47808);
			2025: out = 24'(-48688);
			2026: out = 24'(-49696);
			2027: out = 24'(-50628);
			2028: out = 24'(-51488);
			2029: out = 24'(-52368);
			2030: out = 24'(-53256);
			2031: out = 24'(-54168);
			2032: out = 24'(-55036);
			2033: out = 24'(-55828);
			2034: out = 24'(-56620);
			2035: out = 24'(-57496);
			2036: out = 24'(-58244);
			2037: out = 24'(-59008);
			2038: out = 24'(-59768);
			2039: out = 24'(-60564);
			2040: out = 24'(-61280);
			2041: out = 24'(-62068);
			2042: out = 24'(-62800);
			2043: out = 24'(-63400);
			2044: out = 24'(-64160);
			2045: out = 24'(-64828);
			2046: out = 24'(-65452);
			2047: out = 24'(-66100);
			2048: out = 24'(-66756);
			2049: out = 24'(-67292);
			2050: out = 24'(-67976);
			2051: out = 24'(-68544);
			2052: out = 24'(-69108);
			2053: out = 24'(-69676);
			2054: out = 24'(-70184);
			2055: out = 24'(-70872);
			2056: out = 24'(-71356);
			2057: out = 24'(-71792);
			2058: out = 24'(-72296);
			2059: out = 24'(-72664);
			2060: out = 24'(-73112);
			2061: out = 24'(-73540);
			2062: out = 24'(-73892);
			2063: out = 24'(-74368);
			2064: out = 24'(-74872);
			2065: out = 24'(-75172);
			2066: out = 24'(-75600);
			2067: out = 24'(-75908);
			2068: out = 24'(-76244);
			2069: out = 24'(-76684);
			2070: out = 24'(-76928);
			2071: out = 24'(-77312);
			2072: out = 24'(-77628);
			2073: out = 24'(-77952);
			2074: out = 24'(-78272);
			2075: out = 24'(-78600);
			2076: out = 24'(-78864);
			2077: out = 24'(-79076);
			2078: out = 24'(-79312);
			2079: out = 24'(-79564);
			2080: out = 24'(-79836);
			2081: out = 24'(-80044);
			2082: out = 24'(-80280);
			2083: out = 24'(-80524);
			2084: out = 24'(-80620);
			2085: out = 24'(-80956);
			2086: out = 24'(-81084);
			2087: out = 24'(-81344);
			2088: out = 24'(-81452);
			2089: out = 24'(-81596);
			2090: out = 24'(-81748);
			2091: out = 24'(-81908);
			2092: out = 24'(-81976);
			2093: out = 24'(-82140);
			2094: out = 24'(-82304);
			2095: out = 24'(-82340);
			2096: out = 24'(-82480);
			2097: out = 24'(-82600);
			2098: out = 24'(-82632);
			2099: out = 24'(-82764);
			2100: out = 24'(-82848);
			2101: out = 24'(-82916);
			2102: out = 24'(-82952);
			2103: out = 24'(-83000);
			2104: out = 24'(-83096);
			2105: out = 24'(-83064);
			2106: out = 24'(-83156);
			2107: out = 24'(-83236);
			2108: out = 24'(-83204);
			2109: out = 24'(-83296);
			2110: out = 24'(-83296);
			2111: out = 24'(-83276);
			2112: out = 24'(-83364);
			2113: out = 24'(-83316);
			2114: out = 24'(-83320);
			2115: out = 24'(-83412);
			2116: out = 24'(-83408);
			2117: out = 24'(-83368);
			2118: out = 24'(-83312);
			2119: out = 24'(-83272);
			2120: out = 24'(-83320);
			2121: out = 24'(-83276);
			2122: out = 24'(-83244);
			2123: out = 24'(-83200);
			2124: out = 24'(-83132);
			2125: out = 24'(-83120);
			2126: out = 24'(-83040);
			2127: out = 24'(-82960);
			2128: out = 24'(-82984);
			2129: out = 24'(-82860);
			2130: out = 24'(-82780);
			2131: out = 24'(-82672);
			2132: out = 24'(-82672);
			2133: out = 24'(-82576);
			2134: out = 24'(-82412);
			2135: out = 24'(-82268);
			2136: out = 24'(-82184);
			2137: out = 24'(-82068);
			2138: out = 24'(-81912);
			2139: out = 24'(-81804);
			2140: out = 24'(-81504);
			2141: out = 24'(-81280);
			2142: out = 24'(-81240);
			2143: out = 24'(-81048);
			2144: out = 24'(-80856);
			2145: out = 24'(-80720);
			2146: out = 24'(-80500);
			2147: out = 24'(-80344);
			2148: out = 24'(-80064);
			2149: out = 24'(-79848);
			2150: out = 24'(-79552);
			2151: out = 24'(-79248);
			2152: out = 24'(-79020);
			2153: out = 24'(-78644);
			2154: out = 24'(-78400);
			2155: out = 24'(-78080);
			2156: out = 24'(-77676);
			2157: out = 24'(-77376);
			2158: out = 24'(-76920);
			2159: out = 24'(-76540);
			2160: out = 24'(-76224);
			2161: out = 24'(-75820);
			2162: out = 24'(-75384);
			2163: out = 24'(-74860);
			2164: out = 24'(-74444);
			2165: out = 24'(-73908);
			2166: out = 24'(-73428);
			2167: out = 24'(-72936);
			2168: out = 24'(-72432);
			2169: out = 24'(-71848);
			2170: out = 24'(-71224);
			2171: out = 24'(-70740);
			2172: out = 24'(-70132);
			2173: out = 24'(-69588);
			2174: out = 24'(-68904);
			2175: out = 24'(-68320);
			2176: out = 24'(-67672);
			2177: out = 24'(-67044);
			2178: out = 24'(-66404);
			2179: out = 24'(-65784);
			2180: out = 24'(-65016);
			2181: out = 24'(-64404);
			2182: out = 24'(-63720);
			2183: out = 24'(-63052);
			2184: out = 24'(-62492);
			2185: out = 24'(-61752);
			2186: out = 24'(-61036);
			2187: out = 24'(-60400);
			2188: out = 24'(-59716);
			2189: out = 24'(-58996);
			2190: out = 24'(-58380);
			2191: out = 24'(-57680);
			2192: out = 24'(-56980);
			2193: out = 24'(-56292);
			2194: out = 24'(-55696);
			2195: out = 24'(-55056);
			2196: out = 24'(-54376);
			2197: out = 24'(-53748);
			2198: out = 24'(-53088);
			2199: out = 24'(-52388);
			2200: out = 24'(-51684);
			2201: out = 24'(-51096);
			2202: out = 24'(-50452);
			2203: out = 24'(-49800);
			2204: out = 24'(-49232);
			2205: out = 24'(-48552);
			2206: out = 24'(-47984);
			2207: out = 24'(-47404);
			2208: out = 24'(-46744);
			2209: out = 24'(-46184);
			2210: out = 24'(-45508);
			2211: out = 24'(-44988);
			2212: out = 24'(-44348);
			2213: out = 24'(-43816);
			2214: out = 24'(-43216);
			2215: out = 24'(-42612);
			2216: out = 24'(-42108);
			2217: out = 24'(-41444);
			2218: out = 24'(-40976);
			2219: out = 24'(-40412);
			2220: out = 24'(-39884);
			2221: out = 24'(-39408);
			2222: out = 24'(-38756);
			2223: out = 24'(-38280);
			2224: out = 24'(-37740);
			2225: out = 24'(-37160);
			2226: out = 24'(-36672);
			2227: out = 24'(-36184);
			2228: out = 24'(-35660);
			2229: out = 24'(-35176);
			2230: out = 24'(-34676);
			2231: out = 24'(-34168);
			2232: out = 24'(-33724);
			2233: out = 24'(-33296);
			2234: out = 24'(-32740);
			2235: out = 24'(-32256);
			2236: out = 24'(-31812);
			2237: out = 24'(-31268);
			2238: out = 24'(-30868);
			2239: out = 24'(-30404);
			2240: out = 24'(-30016);
			2241: out = 24'(-29556);
			2242: out = 24'(-29180);
			2243: out = 24'(-28748);
			2244: out = 24'(-28296);
			2245: out = 24'(-27812);
			2246: out = 24'(-27528);
			2247: out = 24'(-27152);
			2248: out = 24'(-26700);
			2249: out = 24'(-26344);
			2250: out = 24'(-25724);
			2251: out = 24'(-25044);
			2252: out = 24'(-24408);
			2253: out = 24'(-23768);
			2254: out = 24'(-23112);
			2255: out = 24'(-22484);
			2256: out = 24'(-21856);
			2257: out = 24'(-21324);
			2258: out = 24'(-20668);
			2259: out = 24'(-20056);
			2260: out = 24'(-19492);
			2261: out = 24'(-18888);
			2262: out = 24'(-18256);
			2263: out = 24'(-17772);
			2264: out = 24'(-17200);
			2265: out = 24'(-16604);
			2266: out = 24'(-16056);
			2267: out = 24'(-15580);
			2268: out = 24'(-14964);
			2269: out = 24'(-14512);
			2270: out = 24'(-14044);
			2271: out = 24'(-13472);
			2272: out = 24'(-13004);
			2273: out = 24'(-12500);
			2274: out = 24'(-12004);
			2275: out = 24'(-11540);
			2276: out = 24'(-11036);
			2277: out = 24'(-10592);
			2278: out = 24'(-10060);
			2279: out = 24'(-9580);
			2280: out = 24'(-9204);
			2281: out = 24'(-8736);
			2282: out = 24'(-8308);
			2283: out = 24'(-7828);
			2284: out = 24'(-7452);
			2285: out = 24'(-6944);
			2286: out = 24'(-6508);
			2287: out = 24'(-6136);
			2288: out = 24'(-5644);
			2289: out = 24'(-5236);
			2290: out = 24'(-4728);
			2291: out = 24'(-4376);
			2292: out = 24'(-3996);
			2293: out = 24'(-3576);
			2294: out = 24'(-3200);
			2295: out = 24'(-2668);
			2296: out = 24'(-2252);
			2297: out = 24'(-1820);
			2298: out = 24'(-1348);
			2299: out = 24'(-964);
			2300: out = 24'(-552);
			2301: out = 24'(-164);
			2302: out = 24'(260);
			2303: out = 24'(684);
			2304: out = 24'(1072);
			2305: out = 24'(1412);
			2306: out = 24'(1852);
			2307: out = 24'(2332);
			2308: out = 24'(2736);
			2309: out = 24'(3232);
			2310: out = 24'(3620);
			2311: out = 24'(4016);
			2312: out = 24'(4552);
			2313: out = 24'(4880);
			2314: out = 24'(5344);
			2315: out = 24'(5800);
			2316: out = 24'(6120);
			2317: out = 24'(6640);
			2318: out = 24'(6876);
			2319: out = 24'(7260);
			2320: out = 24'(7828);
			2321: out = 24'(8292);
			2322: out = 24'(8856);
			2323: out = 24'(9292);
			2324: out = 24'(9784);
			2325: out = 24'(10252);
			2326: out = 24'(10856);
			2327: out = 24'(11344);
			2328: out = 24'(11860);
			2329: out = 24'(12364);
			2330: out = 24'(12900);
			2331: out = 24'(13452);
			2332: out = 24'(13976);
			2333: out = 24'(14564);
			2334: out = 24'(15076);
			2335: out = 24'(15692);
			2336: out = 24'(16340);
			2337: out = 24'(16920);
			2338: out = 24'(17580);
			2339: out = 24'(18276);
			2340: out = 24'(18820);
			2341: out = 24'(19480);
			2342: out = 24'(20124);
			2343: out = 24'(20880);
			2344: out = 24'(21476);
			2345: out = 24'(22128);
			2346: out = 24'(22864);
			2347: out = 24'(23604);
			2348: out = 24'(24284);
			2349: out = 24'(25024);
			2350: out = 24'(25732);
			2351: out = 24'(26388);
			2352: out = 24'(27160);
			2353: out = 24'(27852);
			2354: out = 24'(28620);
			2355: out = 24'(29312);
			2356: out = 24'(30096);
			2357: out = 24'(30728);
			2358: out = 24'(31396);
			2359: out = 24'(32212);
			2360: out = 24'(32880);
			2361: out = 24'(33548);
			2362: out = 24'(34332);
			2363: out = 24'(35008);
			2364: out = 24'(35668);
			2365: out = 24'(36392);
			2366: out = 24'(37064);
			2367: out = 24'(37708);
			2368: out = 24'(38352);
			2369: out = 24'(39032);
			2370: out = 24'(39660);
			2371: out = 24'(40416);
			2372: out = 24'(41056);
			2373: out = 24'(41648);
			2374: out = 24'(42252);
			2375: out = 24'(42956);
			2376: out = 24'(43504);
			2377: out = 24'(44148);
			2378: out = 24'(44768);
			2379: out = 24'(45356);
			2380: out = 24'(45892);
			2381: out = 24'(46456);
			2382: out = 24'(47080);
			2383: out = 24'(47652);
			2384: out = 24'(48192);
			2385: out = 24'(48728);
			2386: out = 24'(49228);
			2387: out = 24'(49800);
			2388: out = 24'(50252);
			2389: out = 24'(50880);
			2390: out = 24'(51420);
			2391: out = 24'(51820);
			2392: out = 24'(52344);
			2393: out = 24'(52828);
			2394: out = 24'(53332);
			2395: out = 24'(53780);
			2396: out = 24'(54456);
			2397: out = 24'(54836);
			2398: out = 24'(55344);
			2399: out = 24'(55784);
			2400: out = 24'(56268);
			2401: out = 24'(56684);
			2402: out = 24'(57332);
			2403: out = 24'(57832);
			2404: out = 24'(58192);
			2405: out = 24'(58636);
			2406: out = 24'(58944);
			2407: out = 24'(59368);
			2408: out = 24'(59760);
			2409: out = 24'(60132);
			2410: out = 24'(60504);
			2411: out = 24'(60968);
			2412: out = 24'(61360);
			2413: out = 24'(61800);
			2414: out = 24'(62092);
			2415: out = 24'(62516);
			2416: out = 24'(62892);
			2417: out = 24'(63288);
			2418: out = 24'(63608);
			2419: out = 24'(64060);
			2420: out = 24'(64404);
			2421: out = 24'(64708);
			2422: out = 24'(65080);
			2423: out = 24'(65452);
			2424: out = 24'(65788);
			2425: out = 24'(66176);
			2426: out = 24'(66460);
			2427: out = 24'(66824);
			2428: out = 24'(67108);
			2429: out = 24'(67456);
			2430: out = 24'(67740);
			2431: out = 24'(68060);
			2432: out = 24'(68364);
			2433: out = 24'(68692);
			2434: out = 24'(68956);
			2435: out = 24'(69276);
			2436: out = 24'(69572);
			2437: out = 24'(69872);
			2438: out = 24'(70192);
			2439: out = 24'(70460);
			2440: out = 24'(70800);
			2441: out = 24'(71076);
			2442: out = 24'(71316);
			2443: out = 24'(71572);
			2444: out = 24'(71876);
			2445: out = 24'(72240);
			2446: out = 24'(72452);
			2447: out = 24'(72776);
			2448: out = 24'(72976);
			2449: out = 24'(73308);
			2450: out = 24'(73552);
			2451: out = 24'(73824);
			2452: out = 24'(74128);
			2453: out = 24'(74348);
			2454: out = 24'(74532);
			2455: out = 24'(74872);
			2456: out = 24'(75096);
			2457: out = 24'(75300);
			2458: out = 24'(75584);
			2459: out = 24'(75740);
			2460: out = 24'(76048);
			2461: out = 24'(76244);
			2462: out = 24'(76484);
			2463: out = 24'(76692);
			2464: out = 24'(76936);
			2465: out = 24'(77036);
			2466: out = 24'(77052);
			2467: out = 24'(77028);
			2468: out = 24'(77132);
			2469: out = 24'(77292);
			2470: out = 24'(77344);
			2471: out = 24'(77472);
			2472: out = 24'(77556);
			2473: out = 24'(77664);
			2474: out = 24'(77460);
			2475: out = 24'(77220);
			2476: out = 24'(77032);
			2477: out = 24'(76952);
			2478: out = 24'(76948);
			2479: out = 24'(76992);
			2480: out = 24'(76776);
			2481: out = 24'(76636);
			2482: out = 24'(76624);
			2483: out = 24'(76676);
			2484: out = 24'(76624);
			2485: out = 24'(76628);
			2486: out = 24'(76748);
			2487: out = 24'(76420);
			2488: out = 24'(76340);
			2489: out = 24'(76180);
			2490: out = 24'(76140);
			2491: out = 24'(76148);
			2492: out = 24'(76180);
			2493: out = 24'(76196);
			2494: out = 24'(76036);
			2495: out = 24'(75576);
			2496: out = 24'(75432);
			2497: out = 24'(75300);
			2498: out = 24'(75284);
			2499: out = 24'(75336);
			2500: out = 24'(75152);
			2501: out = 24'(74912);
			2502: out = 24'(74588);
			2503: out = 24'(74400);
			2504: out = 24'(74132);
			2505: out = 24'(74260);
			2506: out = 24'(74012);
			2507: out = 24'(73716);
			2508: out = 24'(73568);
			2509: out = 24'(73392);
			2510: out = 24'(73404);
			2511: out = 24'(73120);
			2512: out = 24'(72724);
			2513: out = 24'(72500);
			2514: out = 24'(72160);
			2515: out = 24'(72056);
			2516: out = 24'(71748);
			2517: out = 24'(71288);
			2518: out = 24'(71108);
			2519: out = 24'(70772);
			2520: out = 24'(70452);
			2521: out = 24'(70132);
			2522: out = 24'(69748);
			2523: out = 24'(69440);
			2524: out = 24'(68988);
			2525: out = 24'(68616);
			2526: out = 24'(68144);
			2527: out = 24'(67604);
			2528: out = 24'(67300);
			2529: out = 24'(66900);
			2530: out = 24'(66364);
			2531: out = 24'(66020);
			2532: out = 24'(65596);
			2533: out = 24'(65044);
			2534: out = 24'(64744);
			2535: out = 24'(64160);
			2536: out = 24'(63592);
			2537: out = 24'(63220);
			2538: out = 24'(62524);
			2539: out = 24'(62112);
			2540: out = 24'(61712);
			2541: out = 24'(61096);
			2542: out = 24'(60656);
			2543: out = 24'(60180);
			2544: out = 24'(59700);
			2545: out = 24'(59080);
			2546: out = 24'(58524);
			2547: out = 24'(58036);
			2548: out = 24'(57392);
			2549: out = 24'(57012);
			2550: out = 24'(56568);
			2551: out = 24'(56012);
			2552: out = 24'(55432);
			2553: out = 24'(54724);
			2554: out = 24'(54304);
			2555: out = 24'(53752);
			2556: out = 24'(53256);
			2557: out = 24'(52852);
			2558: out = 24'(52292);
			2559: out = 24'(51888);
			2560: out = 24'(51316);
			2561: out = 24'(50680);
			2562: out = 24'(50184);
			2563: out = 24'(49520);
			2564: out = 24'(48952);
			2565: out = 24'(48568);
			2566: out = 24'(48124);
			2567: out = 24'(47532);
			2568: out = 24'(47100);
			2569: out = 24'(46636);
			2570: out = 24'(46144);
			2571: out = 24'(45536);
			2572: out = 24'(45092);
			2573: out = 24'(44620);
			2574: out = 24'(44048);
			2575: out = 24'(43636);
			2576: out = 24'(43004);
			2577: out = 24'(42592);
			2578: out = 24'(42096);
			2579: out = 24'(41592);
			2580: out = 24'(41124);
			2581: out = 24'(40720);
			2582: out = 24'(40316);
			2583: out = 24'(39788);
			2584: out = 24'(39312);
			2585: out = 24'(38856);
			2586: out = 24'(38416);
			2587: out = 24'(37924);
			2588: out = 24'(37556);
			2589: out = 24'(37284);
			2590: out = 24'(36756);
			2591: out = 24'(36260);
			2592: out = 24'(35772);
			2593: out = 24'(35364);
			2594: out = 24'(34928);
			2595: out = 24'(34476);
			2596: out = 24'(34092);
			2597: out = 24'(33616);
			2598: out = 24'(33204);
			2599: out = 24'(32824);
			2600: out = 24'(32428);
			2601: out = 24'(32088);
			2602: out = 24'(31688);
			2603: out = 24'(31296);
			2604: out = 24'(30916);
			2605: out = 24'(30580);
			2606: out = 24'(30220);
			2607: out = 24'(29872);
			2608: out = 24'(29376);
			2609: out = 24'(29072);
			2610: out = 24'(28744);
			2611: out = 24'(28368);
			2612: out = 24'(27968);
			2613: out = 24'(27632);
			2614: out = 24'(27296);
			2615: out = 24'(26872);
			2616: out = 24'(26540);
			2617: out = 24'(26328);
			2618: out = 24'(26040);
			2619: out = 24'(25644);
			2620: out = 24'(25256);
			2621: out = 24'(24868);
			2622: out = 24'(24540);
			2623: out = 24'(24288);
			2624: out = 24'(23956);
			2625: out = 24'(23652);
			2626: out = 24'(23300);
			2627: out = 24'(22952);
			2628: out = 24'(22648);
			2629: out = 24'(22300);
			2630: out = 24'(22124);
			2631: out = 24'(21836);
			2632: out = 24'(21540);
			2633: out = 24'(21180);
			2634: out = 24'(20852);
			2635: out = 24'(20616);
			2636: out = 24'(20348);
			2637: out = 24'(20032);
			2638: out = 24'(19788);
			2639: out = 24'(19496);
			2640: out = 24'(19228);
			2641: out = 24'(18924);
			2642: out = 24'(18740);
			2643: out = 24'(18408);
			2644: out = 24'(17868);
			2645: out = 24'(17300);
			2646: out = 24'(16608);
			2647: out = 24'(15968);
			2648: out = 24'(15412);
			2649: out = 24'(14844);
			2650: out = 24'(14224);
			2651: out = 24'(13548);
			2652: out = 24'(13004);
			2653: out = 24'(12420);
			2654: out = 24'(11932);
			2655: out = 24'(11372);
			2656: out = 24'(10796);
			2657: out = 24'(10300);
			2658: out = 24'(9744);
			2659: out = 24'(9320);
			2660: out = 24'(8768);
			2661: out = 24'(8272);
			2662: out = 24'(7740);
			2663: out = 24'(7300);
			2664: out = 24'(6848);
			2665: out = 24'(6300);
			2666: out = 24'(5960);
			2667: out = 24'(5376);
			2668: out = 24'(4992);
			2669: out = 24'(4472);
			2670: out = 24'(4100);
			2671: out = 24'(3612);
			2672: out = 24'(3100);
			2673: out = 24'(2720);
			2674: out = 24'(2292);
			2675: out = 24'(1772);
			2676: out = 24'(1368);
			2677: out = 24'(916);
			2678: out = 24'(512);
			2679: out = 24'(108);
			2680: out = 24'(-332);
			2681: out = 24'(-796);
			2682: out = 24'(-1120);
			2683: out = 24'(-1544);
			2684: out = 24'(-1956);
			2685: out = 24'(-2344);
			2686: out = 24'(-2684);
			2687: out = 24'(-3132);
			2688: out = 24'(-3576);
			2689: out = 24'(-3980);
			2690: out = 24'(-4372);
			2691: out = 24'(-4768);
			2692: out = 24'(-5152);
			2693: out = 24'(-5500);
			2694: out = 24'(-5824);
			2695: out = 24'(-6268);
			2696: out = 24'(-6524);
			2697: out = 24'(-7036);
			2698: out = 24'(-7520);
			2699: out = 24'(-7792);
			2700: out = 24'(-8240);
			2701: out = 24'(-8608);
			2702: out = 24'(-9060);
			2703: out = 24'(-9448);
			2704: out = 24'(-9896);
			2705: out = 24'(-10284);
			2706: out = 24'(-10580);
			2707: out = 24'(-11040);
			2708: out = 24'(-11436);
			2709: out = 24'(-11952);
			2710: out = 24'(-12324);
			2711: out = 24'(-12680);
			2712: out = 24'(-13096);
			2713: out = 24'(-13492);
			2714: out = 24'(-13944);
			2715: out = 24'(-14312);
			2716: out = 24'(-14764);
			2717: out = 24'(-15148);
			2718: out = 24'(-15564);
			2719: out = 24'(-15940);
			2720: out = 24'(-16332);
			2721: out = 24'(-16796);
			2722: out = 24'(-17264);
			2723: out = 24'(-17644);
			2724: out = 24'(-18084);
			2725: out = 24'(-18564);
			2726: out = 24'(-19032);
			2727: out = 24'(-19420);
			2728: out = 24'(-19928);
			2729: out = 24'(-20344);
			2730: out = 24'(-20880);
			2731: out = 24'(-21332);
			2732: out = 24'(-21864);
			2733: out = 24'(-22416);
			2734: out = 24'(-22880);
			2735: out = 24'(-23352);
			2736: out = 24'(-23920);
			2737: out = 24'(-24476);
			2738: out = 24'(-25068);
			2739: out = 24'(-25536);
			2740: out = 24'(-26116);
			2741: out = 24'(-26712);
			2742: out = 24'(-27228);
			2743: out = 24'(-27772);
			2744: out = 24'(-28460);
			2745: out = 24'(-29048);
			2746: out = 24'(-29648);
			2747: out = 24'(-30356);
			2748: out = 24'(-31012);
			2749: out = 24'(-31608);
			2750: out = 24'(-32308);
			2751: out = 24'(-32876);
			2752: out = 24'(-33636);
			2753: out = 24'(-34308);
			2754: out = 24'(-34980);
			2755: out = 24'(-35752);
			2756: out = 24'(-36516);
			2757: out = 24'(-37128);
			2758: out = 24'(-37756);
			2759: out = 24'(-38492);
			2760: out = 24'(-39320);
			2761: out = 24'(-40096);
			2762: out = 24'(-40744);
			2763: out = 24'(-41548);
			2764: out = 24'(-42252);
			2765: out = 24'(-42948);
			2766: out = 24'(-43788);
			2767: out = 24'(-44640);
			2768: out = 24'(-45372);
			2769: out = 24'(-45900);
			2770: out = 24'(-46664);
			2771: out = 24'(-47364);
			2772: out = 24'(-48012);
			2773: out = 24'(-48716);
			2774: out = 24'(-49404);
			2775: out = 24'(-50080);
			2776: out = 24'(-50752);
			2777: out = 24'(-51352);
			2778: out = 24'(-52044);
			2779: out = 24'(-52724);
			2780: out = 24'(-53284);
			2781: out = 24'(-53872);
			2782: out = 24'(-54484);
			2783: out = 24'(-55088);
			2784: out = 24'(-55604);
			2785: out = 24'(-56248);
			2786: out = 24'(-56728);
			2787: out = 24'(-57336);
			2788: out = 24'(-57832);
			2789: out = 24'(-58380);
			2790: out = 24'(-58952);
			2791: out = 24'(-59380);
			2792: out = 24'(-59916);
			2793: out = 24'(-60428);
			2794: out = 24'(-60880);
			2795: out = 24'(-61272);
			2796: out = 24'(-61764);
			2797: out = 24'(-62200);
			2798: out = 24'(-62692);
			2799: out = 24'(-63060);
			2800: out = 24'(-63452);
			2801: out = 24'(-63876);
			2802: out = 24'(-64244);
			2803: out = 24'(-64652);
			2804: out = 24'(-65004);
			2805: out = 24'(-65376);
			2806: out = 24'(-65656);
			2807: out = 24'(-66044);
			2808: out = 24'(-66400);
			2809: out = 24'(-66728);
			2810: out = 24'(-67008);
			2811: out = 24'(-67324);
			2812: out = 24'(-67628);
			2813: out = 24'(-67908);
			2814: out = 24'(-68212);
			2815: out = 24'(-68480);
			2816: out = 24'(-68636);
			2817: out = 24'(-68944);
			2818: out = 24'(-69140);
			2819: out = 24'(-69480);
			2820: out = 24'(-69612);
			2821: out = 24'(-69836);
			2822: out = 24'(-70136);
			2823: out = 24'(-70296);
			2824: out = 24'(-70568);
			2825: out = 24'(-70644);
			2826: out = 24'(-70820);
			2827: out = 24'(-71052);
			2828: out = 24'(-71228);
			2829: out = 24'(-71364);
			2830: out = 24'(-71512);
			2831: out = 24'(-71592);
			2832: out = 24'(-71676);
			2833: out = 24'(-71896);
			2834: out = 24'(-72036);
			2835: out = 24'(-72140);
			2836: out = 24'(-72248);
			2837: out = 24'(-72312);
			2838: out = 24'(-72336);
			2839: out = 24'(-72528);
			2840: out = 24'(-72680);
			2841: out = 24'(-72644);
			2842: out = 24'(-72728);
			2843: out = 24'(-72808);
			2844: out = 24'(-72872);
			2845: out = 24'(-72936);
			2846: out = 24'(-73024);
			2847: out = 24'(-73068);
			2848: out = 24'(-73064);
			2849: out = 24'(-73120);
			2850: out = 24'(-73160);
			2851: out = 24'(-73000);
			2852: out = 24'(-73096);
			2853: out = 24'(-73156);
			2854: out = 24'(-73168);
			2855: out = 24'(-73280);
			2856: out = 24'(-73304);
			2857: out = 24'(-73348);
			2858: out = 24'(-73304);
			2859: out = 24'(-73260);
			2860: out = 24'(-73280);
			2861: out = 24'(-73284);
			2862: out = 24'(-73268);
			2863: out = 24'(-73348);
			2864: out = 24'(-73220);
			2865: out = 24'(-73240);
			2866: out = 24'(-73156);
			2867: out = 24'(-73164);
			2868: out = 24'(-73188);
			2869: out = 24'(-73112);
			2870: out = 24'(-73072);
			2871: out = 24'(-73104);
			2872: out = 24'(-72976);
			2873: out = 24'(-72884);
			2874: out = 24'(-72900);
			2875: out = 24'(-72820);
			2876: out = 24'(-72768);
			2877: out = 24'(-72684);
			2878: out = 24'(-72536);
			2879: out = 24'(-72472);
			2880: out = 24'(-72516);
			2881: out = 24'(-72348);
			2882: out = 24'(-72308);
			2883: out = 24'(-72180);
			2884: out = 24'(-72104);
			2885: out = 24'(-71972);
			2886: out = 24'(-71864);
			2887: out = 24'(-71760);
			2888: out = 24'(-71644);
			2889: out = 24'(-71460);
			2890: out = 24'(-71360);
			2891: out = 24'(-71224);
			2892: out = 24'(-71228);
			2893: out = 24'(-71044);
			2894: out = 24'(-70876);
			2895: out = 24'(-70804);
			2896: out = 24'(-70588);
			2897: out = 24'(-70520);
			2898: out = 24'(-70332);
			2899: out = 24'(-70236);
			2900: out = 24'(-70124);
			2901: out = 24'(-69992);
			2902: out = 24'(-69844);
			2903: out = 24'(-69700);
			2904: out = 24'(-69572);
			2905: out = 24'(-69368);
			2906: out = 24'(-69236);
			2907: out = 24'(-69032);
			2908: out = 24'(-68856);
			2909: out = 24'(-68704);
			2910: out = 24'(-68408);
			2911: out = 24'(-68320);
			2912: out = 24'(-68012);
			2913: out = 24'(-67868);
			2914: out = 24'(-67584);
			2915: out = 24'(-67412);
			2916: out = 24'(-67156);
			2917: out = 24'(-66896);
			2918: out = 24'(-66652);
			2919: out = 24'(-66348);
			2920: out = 24'(-66092);
			2921: out = 24'(-65812);
			2922: out = 24'(-65504);
			2923: out = 24'(-65188);
			2924: out = 24'(-64828);
			2925: out = 24'(-64556);
			2926: out = 24'(-64188);
			2927: out = 24'(-63868);
			2928: out = 24'(-63512);
			2929: out = 24'(-63052);
			2930: out = 24'(-62732);
			2931: out = 24'(-62248);
			2932: out = 24'(-61928);
			2933: out = 24'(-61468);
			2934: out = 24'(-61080);
			2935: out = 24'(-60600);
			2936: out = 24'(-60168);
			2937: out = 24'(-59720);
			2938: out = 24'(-59252);
			2939: out = 24'(-58840);
			2940: out = 24'(-58304);
			2941: out = 24'(-57796);
			2942: out = 24'(-57248);
			2943: out = 24'(-56792);
			2944: out = 24'(-56356);
			2945: out = 24'(-55772);
			2946: out = 24'(-55216);
			2947: out = 24'(-54728);
			2948: out = 24'(-54204);
			2949: out = 24'(-53652);
			2950: out = 24'(-53092);
			2951: out = 24'(-52592);
			2952: out = 24'(-52132);
			2953: out = 24'(-51516);
			2954: out = 24'(-50948);
			2955: out = 24'(-50352);
			2956: out = 24'(-49796);
			2957: out = 24'(-49276);
			2958: out = 24'(-48648);
			2959: out = 24'(-48084);
			2960: out = 24'(-47548);
			2961: out = 24'(-47028);
			2962: out = 24'(-46452);
			2963: out = 24'(-45872);
			2964: out = 24'(-45388);
			2965: out = 24'(-44804);
			2966: out = 24'(-44268);
			2967: out = 24'(-43788);
			2968: out = 24'(-43224);
			2969: out = 24'(-42664);
			2970: out = 24'(-42180);
			2971: out = 24'(-41616);
			2972: out = 24'(-41064);
			2973: out = 24'(-40608);
			2974: out = 24'(-40056);
			2975: out = 24'(-39552);
			2976: out = 24'(-39052);
			2977: out = 24'(-38544);
			2978: out = 24'(-38108);
			2979: out = 24'(-37596);
			2980: out = 24'(-37040);
			2981: out = 24'(-36560);
			2982: out = 24'(-36064);
			2983: out = 24'(-35556);
			2984: out = 24'(-35156);
			2985: out = 24'(-34616);
			2986: out = 24'(-34200);
			2987: out = 24'(-33720);
			2988: out = 24'(-33220);
			2989: out = 24'(-32736);
			2990: out = 24'(-32356);
			2991: out = 24'(-31868);
			2992: out = 24'(-31412);
			2993: out = 24'(-30928);
			2994: out = 24'(-30460);
			2995: out = 24'(-30048);
			2996: out = 24'(-29612);
			2997: out = 24'(-29192);
			2998: out = 24'(-28788);
			2999: out = 24'(-28264);
			3000: out = 24'(-27896);
			3001: out = 24'(-27484);
			3002: out = 24'(-27116);
			3003: out = 24'(-26728);
			3004: out = 24'(-26280);
			3005: out = 24'(-25928);
			3006: out = 24'(-25516);
			3007: out = 24'(-25112);
			3008: out = 24'(-24792);
			3009: out = 24'(-24432);
			3010: out = 24'(-24048);
			3011: out = 24'(-23676);
			3012: out = 24'(-23336);
			3013: out = 24'(-22984);
			3014: out = 24'(-22664);
			3015: out = 24'(-22304);
			3016: out = 24'(-21980);
			3017: out = 24'(-21588);
			3018: out = 24'(-21264);
			3019: out = 24'(-20936);
			3020: out = 24'(-20612);
			3021: out = 24'(-20316);
			3022: out = 24'(-19992);
			3023: out = 24'(-19544);
			3024: out = 24'(-19304);
			3025: out = 24'(-19036);
			3026: out = 24'(-18620);
			3027: out = 24'(-18404);
			3028: out = 24'(-18040);
			3029: out = 24'(-17752);
			3030: out = 24'(-17428);
			3031: out = 24'(-17024);
			3032: out = 24'(-16456);
			3033: out = 24'(-15964);
			3034: out = 24'(-15400);
			3035: out = 24'(-14900);
			3036: out = 24'(-14480);
			3037: out = 24'(-13888);
			3038: out = 24'(-13388);
			3039: out = 24'(-12984);
			3040: out = 24'(-12532);
			3041: out = 24'(-12128);
			3042: out = 24'(-11648);
			3043: out = 24'(-11236);
			3044: out = 24'(-10876);
			3045: out = 24'(-10432);
			3046: out = 24'(-10048);
			3047: out = 24'(-9588);
			3048: out = 24'(-9172);
			3049: out = 24'(-8768);
			3050: out = 24'(-8356);
			3051: out = 24'(-7976);
			3052: out = 24'(-7656);
			3053: out = 24'(-7208);
			3054: out = 24'(-6876);
			3055: out = 24'(-6552);
			3056: out = 24'(-6124);
			3057: out = 24'(-5740);
			3058: out = 24'(-5360);
			3059: out = 24'(-4984);
			3060: out = 24'(-4676);
			3061: out = 24'(-4296);
			3062: out = 24'(-3972);
			3063: out = 24'(-3636);
			3064: out = 24'(-3316);
			3065: out = 24'(-3036);
			3066: out = 24'(-2588);
			3067: out = 24'(-2308);
			3068: out = 24'(-1980);
			3069: out = 24'(-1644);
			3070: out = 24'(-1332);
			3071: out = 24'(-1068);
			3072: out = 24'(-700);
			3073: out = 24'(-388);
			3074: out = 24'(-24);
			3075: out = 24'(272);
			3076: out = 24'(560);
			3077: out = 24'(780);
			3078: out = 24'(1200);
			3079: out = 24'(1424);
			3080: out = 24'(1852);
			3081: out = 24'(2112);
			3082: out = 24'(2384);
			3083: out = 24'(2660);
			3084: out = 24'(2876);
			3085: out = 24'(3280);
			3086: out = 24'(3540);
			3087: out = 24'(3788);
			3088: out = 24'(4124);
			3089: out = 24'(4332);
			3090: out = 24'(4668);
			3091: out = 24'(4924);
			3092: out = 24'(5192);
			3093: out = 24'(5520);
			3094: out = 24'(5776);
			3095: out = 24'(6020);
			3096: out = 24'(6328);
			3097: out = 24'(6604);
			3098: out = 24'(7020);
			3099: out = 24'(7208);
			3100: out = 24'(7444);
			3101: out = 24'(7844);
			3102: out = 24'(8168);
			3103: out = 24'(8448);
			3104: out = 24'(8764);
			3105: out = 24'(9116);
			3106: out = 24'(9420);
			3107: out = 24'(9756);
			3108: out = 24'(10056);
			3109: out = 24'(10472);
			3110: out = 24'(10724);
			3111: out = 24'(11024);
			3112: out = 24'(11392);
			3113: out = 24'(11804);
			3114: out = 24'(12100);
			3115: out = 24'(12472);
			3116: out = 24'(12840);
			3117: out = 24'(13120);
			3118: out = 24'(13504);
			3119: out = 24'(13956);
			3120: out = 24'(14300);
			3121: out = 24'(14716);
			3122: out = 24'(15116);
			3123: out = 24'(15504);
			3124: out = 24'(15908);
			3125: out = 24'(16264);
			3126: out = 24'(16712);
			3127: out = 24'(17144);
			3128: out = 24'(17516);
			3129: out = 24'(17964);
			3130: out = 24'(18408);
			3131: out = 24'(18908);
			3132: out = 24'(19360);
			3133: out = 24'(19864);
			3134: out = 24'(20360);
			3135: out = 24'(20860);
			3136: out = 24'(21352);
			3137: out = 24'(21852);
			3138: out = 24'(22284);
			3139: out = 24'(22784);
			3140: out = 24'(23320);
			3141: out = 24'(23860);
			3142: out = 24'(24428);
			3143: out = 24'(24864);
			3144: out = 24'(25456);
			3145: out = 24'(25996);
			3146: out = 24'(26464);
			3147: out = 24'(27012);
			3148: out = 24'(27528);
			3149: out = 24'(28100);
			3150: out = 24'(28576);
			3151: out = 24'(29072);
			3152: out = 24'(29648);
			3153: out = 24'(30120);
			3154: out = 24'(30680);
			3155: out = 24'(31160);
			3156: out = 24'(31736);
			3157: out = 24'(32160);
			3158: out = 24'(32672);
			3159: out = 24'(33216);
			3160: out = 24'(33684);
			3161: out = 24'(34184);
			3162: out = 24'(34716);
			3163: out = 24'(35144);
			3164: out = 24'(35600);
			3165: out = 24'(36148);
			3166: out = 24'(36596);
			3167: out = 24'(37056);
			3168: out = 24'(37528);
			3169: out = 24'(37952);
			3170: out = 24'(38408);
			3171: out = 24'(38868);
			3172: out = 24'(39248);
			3173: out = 24'(39740);
			3174: out = 24'(40092);
			3175: out = 24'(40548);
			3176: out = 24'(40976);
			3177: out = 24'(41396);
			3178: out = 24'(41852);
			3179: out = 24'(42212);
			3180: out = 24'(42608);
			3181: out = 24'(42992);
			3182: out = 24'(43432);
			3183: out = 24'(43760);
			3184: out = 24'(44240);
			3185: out = 24'(44480);
			3186: out = 24'(44916);
			3187: out = 24'(45240);
			3188: out = 24'(45620);
			3189: out = 24'(45984);
			3190: out = 24'(46312);
			3191: out = 24'(46680);
			3192: out = 24'(46964);
			3193: out = 24'(47316);
			3194: out = 24'(47676);
			3195: out = 24'(48000);
			3196: out = 24'(48340);
			3197: out = 24'(48608);
			3198: out = 24'(48900);
			3199: out = 24'(49280);
			3200: out = 24'(49532);
			3201: out = 24'(49860);
			3202: out = 24'(50168);
			3203: out = 24'(50464);
			3204: out = 24'(50704);
			3205: out = 24'(51060);
			3206: out = 24'(51360);
			3207: out = 24'(51668);
			3208: out = 24'(51912);
			3209: out = 24'(52216);
			3210: out = 24'(52496);
			3211: out = 24'(52756);
			3212: out = 24'(52984);
			3213: out = 24'(53272);
			3214: out = 24'(53556);
			3215: out = 24'(53760);
			3216: out = 24'(54072);
			3217: out = 24'(54228);
			3218: out = 24'(54444);
			3219: out = 24'(54744);
			3220: out = 24'(54984);
			3221: out = 24'(55156);
			3222: out = 24'(55440);
			3223: out = 24'(55464);
			3224: out = 24'(55740);
			3225: out = 24'(55916);
			3226: out = 24'(56200);
			3227: out = 24'(56436);
			3228: out = 24'(56688);
			3229: out = 24'(56928);
			3230: out = 24'(57152);
			3231: out = 24'(57268);
			3232: out = 24'(57548);
			3233: out = 24'(57696);
			3234: out = 24'(57940);
			3235: out = 24'(58168);
			3236: out = 24'(58300);
			3237: out = 24'(58464);
			3238: out = 24'(58704);
			3239: out = 24'(58900);
			3240: out = 24'(59088);
			3241: out = 24'(59280);
			3242: out = 24'(59452);
			3243: out = 24'(59644);
			3244: out = 24'(59808);
			3245: out = 24'(60100);
			3246: out = 24'(60172);
			3247: out = 24'(60404);
			3248: out = 24'(60480);
			3249: out = 24'(60736);
			3250: out = 24'(60812);
			3251: out = 24'(61016);
			3252: out = 24'(61136);
			3253: out = 24'(61284);
			3254: out = 24'(61404);
			3255: out = 24'(61560);
			3256: out = 24'(61700);
			3257: out = 24'(61892);
			3258: out = 24'(61924);
			3259: out = 24'(61904);
			3260: out = 24'(61936);
			3261: out = 24'(61968);
			3262: out = 24'(61900);
			3263: out = 24'(61924);
			3264: out = 24'(61748);
			3265: out = 24'(61480);
			3266: out = 24'(61444);
			3267: out = 24'(61588);
			3268: out = 24'(61620);
			3269: out = 24'(61556);
			3270: out = 24'(61504);
			3271: out = 24'(61288);
			3272: out = 24'(61236);
			3273: out = 24'(61208);
			3274: out = 24'(61172);
			3275: out = 24'(61020);
			3276: out = 24'(61068);
			3277: out = 24'(60980);
			3278: out = 24'(61036);
			3279: out = 24'(61100);
			3280: out = 24'(60960);
			3281: out = 24'(60880);
			3282: out = 24'(60896);
			3283: out = 24'(60604);
			3284: out = 24'(60580);
			3285: out = 24'(60580);
			3286: out = 24'(60528);
			3287: out = 24'(60432);
			3288: out = 24'(60456);
			3289: out = 24'(60496);
			3290: out = 24'(60416);
			3291: out = 24'(60236);
			3292: out = 24'(60084);
			3293: out = 24'(60164);
			3294: out = 24'(60048);
			3295: out = 24'(60008);
			3296: out = 24'(60184);
			3297: out = 24'(60164);
			3298: out = 24'(60008);
			3299: out = 24'(59932);
			3300: out = 24'(59580);
			3301: out = 24'(59628);
			3302: out = 24'(59636);
			3303: out = 24'(59580);
			3304: out = 24'(59564);
			3305: out = 24'(59636);
			3306: out = 24'(59420);
			3307: out = 24'(59336);
			3308: out = 24'(59380);
			3309: out = 24'(59364);
			3310: out = 24'(59168);
			3311: out = 24'(59012);
			3312: out = 24'(58972);
			3313: out = 24'(58716);
			3314: out = 24'(58756);
			3315: out = 24'(58428);
			3316: out = 24'(58260);
			3317: out = 24'(58348);
			3318: out = 24'(58100);
			3319: out = 24'(57956);
			3320: out = 24'(57908);
			3321: out = 24'(57820);
			3322: out = 24'(57800);
			3323: out = 24'(57376);
			3324: out = 24'(57128);
			3325: out = 24'(56968);
			3326: out = 24'(56836);
			3327: out = 24'(56708);
			3328: out = 24'(56444);
			3329: out = 24'(56248);
			3330: out = 24'(56132);
			3331: out = 24'(55736);
			3332: out = 24'(55492);
			3333: out = 24'(55364);
			3334: out = 24'(55088);
			3335: out = 24'(54604);
			3336: out = 24'(54456);
			3337: out = 24'(54236);
			3338: out = 24'(53872);
			3339: out = 24'(53552);
			3340: out = 24'(53332);
			3341: out = 24'(53040);
			3342: out = 24'(52544);
			3343: out = 24'(52332);
			3344: out = 24'(52148);
			3345: out = 24'(51648);
			3346: out = 24'(51156);
			3347: out = 24'(50828);
			3348: out = 24'(50392);
			3349: out = 24'(50108);
			3350: out = 24'(49764);
			3351: out = 24'(49448);
			3352: out = 24'(49028);
			3353: out = 24'(48720);
			3354: out = 24'(48344);
			3355: out = 24'(48064);
			3356: out = 24'(47584);
			3357: out = 24'(47176);
			3358: out = 24'(46724);
			3359: out = 24'(46208);
			3360: out = 24'(45904);
			3361: out = 24'(45560);
			3362: out = 24'(45112);
			3363: out = 24'(44712);
			3364: out = 24'(44232);
			3365: out = 24'(43916);
			3366: out = 24'(43584);
			3367: out = 24'(43112);
			3368: out = 24'(42672);
			3369: out = 24'(42184);
			3370: out = 24'(41872);
			3371: out = 24'(41472);
			3372: out = 24'(41076);
			3373: out = 24'(40760);
			3374: out = 24'(40316);
			3375: out = 24'(39816);
			3376: out = 24'(39400);
			3377: out = 24'(38988);
			3378: out = 24'(38616);
			3379: out = 24'(38172);
			3380: out = 24'(37748);
			3381: out = 24'(37424);
			3382: out = 24'(37064);
			3383: out = 24'(36564);
			3384: out = 24'(36232);
			3385: out = 24'(35848);
			3386: out = 24'(35460);
			3387: out = 24'(35008);
			3388: out = 24'(34568);
			3389: out = 24'(34160);
			3390: out = 24'(33880);
			3391: out = 24'(33496);
			3392: out = 24'(33068);
			3393: out = 24'(32696);
			3394: out = 24'(32340);
			3395: out = 24'(31892);
			3396: out = 24'(31520);
			3397: out = 24'(31324);
			3398: out = 24'(30904);
			3399: out = 24'(30500);
			3400: out = 24'(30152);
			3401: out = 24'(29728);
			3402: out = 24'(29452);
			3403: out = 24'(29024);
			3404: out = 24'(28732);
			3405: out = 24'(28432);
			3406: out = 24'(28028);
			3407: out = 24'(27660);
			3408: out = 24'(27380);
			3409: out = 24'(27004);
			3410: out = 24'(26484);
			3411: out = 24'(26168);
			3412: out = 24'(25924);
			3413: out = 24'(25628);
			3414: out = 24'(25324);
			3415: out = 24'(25020);
			3416: out = 24'(24776);
			3417: out = 24'(24404);
			3418: out = 24'(24108);
			3419: out = 24'(23820);
			3420: out = 24'(23464);
			3421: out = 24'(23128);
			3422: out = 24'(22836);
			3423: out = 24'(22564);
			3424: out = 24'(22236);
			3425: out = 24'(22000);
			3426: out = 24'(21748);
			3427: out = 24'(21308);
			3428: out = 24'(21152);
			3429: out = 24'(20904);
			3430: out = 24'(20764);
			3431: out = 24'(20428);
			3432: out = 24'(20160);
			3433: out = 24'(19808);
			3434: out = 24'(19580);
			3435: out = 24'(19288);
			3436: out = 24'(19064);
			3437: out = 24'(18840);
			3438: out = 24'(18564);
			3439: out = 24'(18400);
			3440: out = 24'(18116);
			3441: out = 24'(17940);
			3442: out = 24'(17664);
			3443: out = 24'(17356);
			3444: out = 24'(17088);
			3445: out = 24'(16804);
			3446: out = 24'(16640);
			3447: out = 24'(16356);
			3448: out = 24'(16200);
			3449: out = 24'(16004);
			3450: out = 24'(15648);
			3451: out = 24'(15456);
			3452: out = 24'(15276);
			3453: out = 24'(15032);
			3454: out = 24'(14864);
			3455: out = 24'(14580);
			3456: out = 24'(14376);
			3457: out = 24'(14100);
			3458: out = 24'(13924);
			3459: out = 24'(13696);
			3460: out = 24'(13544);
			3461: out = 24'(13292);
			3462: out = 24'(13160);
			3463: out = 24'(12840);
			3464: out = 24'(12800);
			3465: out = 24'(12532);
			3466: out = 24'(12408);
			3467: out = 24'(12204);
			3468: out = 24'(11988);
			3469: out = 24'(11808);
			3470: out = 24'(11656);
			3471: out = 24'(11528);
			3472: out = 24'(11308);
			3473: out = 24'(10964);
			3474: out = 24'(10500);
			3475: out = 24'(10056);
			3476: out = 24'(9616);
			3477: out = 24'(9196);
			3478: out = 24'(8728);
			3479: out = 24'(8320);
			3480: out = 24'(7852);
			3481: out = 24'(7484);
			3482: out = 24'(6964);
			3483: out = 24'(6572);
			3484: out = 24'(6268);
			3485: out = 24'(5872);
			3486: out = 24'(5404);
			3487: out = 24'(4960);
			3488: out = 24'(4676);
			3489: out = 24'(4280);
			3490: out = 24'(3868);
			3491: out = 24'(3520);
			3492: out = 24'(3144);
			3493: out = 24'(2700);
			3494: out = 24'(2496);
			3495: out = 24'(2188);
			3496: out = 24'(1736);
			3497: out = 24'(1388);
			3498: out = 24'(1004);
			3499: out = 24'(640);
			3500: out = 24'(268);
			3501: out = 24'(-76);
			3502: out = 24'(-448);
			3503: out = 24'(-784);
			3504: out = 24'(-1096);
			3505: out = 24'(-1388);
			3506: out = 24'(-1652);
			3507: out = 24'(-1984);
			3508: out = 24'(-2388);
			3509: out = 24'(-2680);
			3510: out = 24'(-2988);
			3511: out = 24'(-3272);
			3512: out = 24'(-3536);
			3513: out = 24'(-3764);
			3514: out = 24'(-4120);
			3515: out = 24'(-4380);
			3516: out = 24'(-4608);
			3517: out = 24'(-4944);
			3518: out = 24'(-5232);
			3519: out = 24'(-5472);
			3520: out = 24'(-5800);
			3521: out = 24'(-6000);
			3522: out = 24'(-6368);
			3523: out = 24'(-6560);
			3524: out = 24'(-6896);
			3525: out = 24'(-7188);
			3526: out = 24'(-7452);
			3527: out = 24'(-7784);
			3528: out = 24'(-8040);
			3529: out = 24'(-8264);
			3530: out = 24'(-8628);
			3531: out = 24'(-8860);
			3532: out = 24'(-9120);
			3533: out = 24'(-9428);
			3534: out = 24'(-9664);
			3535: out = 24'(-9952);
			3536: out = 24'(-10280);
			3537: out = 24'(-10520);
			3538: out = 24'(-10788);
			3539: out = 24'(-11040);
			3540: out = 24'(-11276);
			3541: out = 24'(-11592);
			3542: out = 24'(-11924);
			3543: out = 24'(-12168);
			3544: out = 24'(-12440);
			3545: out = 24'(-12704);
			3546: out = 24'(-12980);
			3547: out = 24'(-13240);
			3548: out = 24'(-13572);
			3549: out = 24'(-13804);
			3550: out = 24'(-14072);
			3551: out = 24'(-14268);
			3552: out = 24'(-14644);
			3553: out = 24'(-14880);
			3554: out = 24'(-15228);
			3555: out = 24'(-15504);
			3556: out = 24'(-15800);
			3557: out = 24'(-16108);
			3558: out = 24'(-16380);
			3559: out = 24'(-16684);
			3560: out = 24'(-17000);
			3561: out = 24'(-17356);
			3562: out = 24'(-17636);
			3563: out = 24'(-18016);
			3564: out = 24'(-18356);
			3565: out = 24'(-18740);
			3566: out = 24'(-19000);
			3567: out = 24'(-19380);
			3568: out = 24'(-19704);
			3569: out = 24'(-20124);
			3570: out = 24'(-20544);
			3571: out = 24'(-20820);
			3572: out = 24'(-21292);
			3573: out = 24'(-21660);
			3574: out = 24'(-21996);
			3575: out = 24'(-22412);
			3576: out = 24'(-22856);
			3577: out = 24'(-23324);
			3578: out = 24'(-23732);
			3579: out = 24'(-24104);
			3580: out = 24'(-24528);
			3581: out = 24'(-24964);
			3582: out = 24'(-25448);
			3583: out = 24'(-25876);
			3584: out = 24'(-26372);
			3585: out = 24'(-26804);
			3586: out = 24'(-27384);
			3587: out = 24'(-27808);
			3588: out = 24'(-28336);
			3589: out = 24'(-28808);
			3590: out = 24'(-29292);
			3591: out = 24'(-29860);
			3592: out = 24'(-30284);
			3593: out = 24'(-30840);
			3594: out = 24'(-31384);
			3595: out = 24'(-31980);
			3596: out = 24'(-32472);
			3597: out = 24'(-32948);
			3598: out = 24'(-33560);
			3599: out = 24'(-34092);
			3600: out = 24'(-34616);
			3601: out = 24'(-35160);
			3602: out = 24'(-35696);
			3603: out = 24'(-36220);
			3604: out = 24'(-36804);
			3605: out = 24'(-37292);
			3606: out = 24'(-37868);
			3607: out = 24'(-38416);
			3608: out = 24'(-38868);
			3609: out = 24'(-39524);
			3610: out = 24'(-39936);
			3611: out = 24'(-40428);
			3612: out = 24'(-40992);
			3613: out = 24'(-41440);
			3614: out = 24'(-41908);
			3615: out = 24'(-42400);
			3616: out = 24'(-42880);
			3617: out = 24'(-43328);
			3618: out = 24'(-43744);
			3619: out = 24'(-44288);
			3620: out = 24'(-44788);
			3621: out = 24'(-45216);
			3622: out = 24'(-45656);
			3623: out = 24'(-46024);
			3624: out = 24'(-46460);
			3625: out = 24'(-46920);
			3626: out = 24'(-47288);
			3627: out = 24'(-47780);
			3628: out = 24'(-48120);
			3629: out = 24'(-48512);
			3630: out = 24'(-48884);
			3631: out = 24'(-49300);
			3632: out = 24'(-49640);
			3633: out = 24'(-50008);
			3634: out = 24'(-50284);
			3635: out = 24'(-50668);
			3636: out = 24'(-50952);
			3637: out = 24'(-51240);
			3638: out = 24'(-51616);
			3639: out = 24'(-51868);
			3640: out = 24'(-52180);
			3641: out = 24'(-52472);
			3642: out = 24'(-52756);
			3643: out = 24'(-53040);
			3644: out = 24'(-53332);
			3645: out = 24'(-53552);
			3646: out = 24'(-53740);
			3647: out = 24'(-54036);
			3648: out = 24'(-54252);
			3649: out = 24'(-54444);
			3650: out = 24'(-54712);
			3651: out = 24'(-54928);
			3652: out = 24'(-55064);
			3653: out = 24'(-55268);
			3654: out = 24'(-55496);
			3655: out = 24'(-55668);
			3656: out = 24'(-55904);
			3657: out = 24'(-56068);
			3658: out = 24'(-56200);
			3659: out = 24'(-56312);
			3660: out = 24'(-56436);
			3661: out = 24'(-56664);
			3662: out = 24'(-56796);
			3663: out = 24'(-56960);
			3664: out = 24'(-57056);
			3665: out = 24'(-57180);
			3666: out = 24'(-57336);
			3667: out = 24'(-57436);
			3668: out = 24'(-57612);
			3669: out = 24'(-57688);
			3670: out = 24'(-57784);
			3671: out = 24'(-57876);
			3672: out = 24'(-58084);
			3673: out = 24'(-58316);
			3674: out = 24'(-58300);
			3675: out = 24'(-58284);
			3676: out = 24'(-58380);
			3677: out = 24'(-58424);
			3678: out = 24'(-58404);
			3679: out = 24'(-58516);
			3680: out = 24'(-58532);
			3681: out = 24'(-58564);
			3682: out = 24'(-58696);
			3683: out = 24'(-58608);
			3684: out = 24'(-58768);
			3685: out = 24'(-58756);
			3686: out = 24'(-58828);
			3687: out = 24'(-58780);
			3688: out = 24'(-58868);
			3689: out = 24'(-58776);
			3690: out = 24'(-58804);
			3691: out = 24'(-58848);
			3692: out = 24'(-58856);
			3693: out = 24'(-58868);
			3694: out = 24'(-58920);
			3695: out = 24'(-58852);
			3696: out = 24'(-58876);
			3697: out = 24'(-58876);
			3698: out = 24'(-58844);
			3699: out = 24'(-58904);
			3700: out = 24'(-58820);
			3701: out = 24'(-58820);
			3702: out = 24'(-58804);
			3703: out = 24'(-58784);
			3704: out = 24'(-58700);
			3705: out = 24'(-58684);
			3706: out = 24'(-58600);
			3707: out = 24'(-58616);
			3708: out = 24'(-58576);
			3709: out = 24'(-58568);
			3710: out = 24'(-58464);
			3711: out = 24'(-58436);
			3712: out = 24'(-58364);
			3713: out = 24'(-58336);
			3714: out = 24'(-58340);
			3715: out = 24'(-58248);
			3716: out = 24'(-58252);
			3717: out = 24'(-58140);
			3718: out = 24'(-58080);
			3719: out = 24'(-58032);
			3720: out = 24'(-58008);
			3721: out = 24'(-57924);
			3722: out = 24'(-57852);
			3723: out = 24'(-57748);
			3724: out = 24'(-57684);
			3725: out = 24'(-57616);
			3726: out = 24'(-57448);
			3727: out = 24'(-57512);
			3728: out = 24'(-57344);
			3729: out = 24'(-57228);
			3730: out = 24'(-57104);
			3731: out = 24'(-57072);
			3732: out = 24'(-56904);
			3733: out = 24'(-56804);
			3734: out = 24'(-56820);
			3735: out = 24'(-56624);
			3736: out = 24'(-56540);
			3737: out = 24'(-56476);
			3738: out = 24'(-56340);
			3739: out = 24'(-56208);
			3740: out = 24'(-56140);
			3741: out = 24'(-56008);
			3742: out = 24'(-55944);
			3743: out = 24'(-55876);
			3744: out = 24'(-55716);
			3745: out = 24'(-55596);
			3746: out = 24'(-55460);
			3747: out = 24'(-55280);
			3748: out = 24'(-55196);
			3749: out = 24'(-55040);
			3750: out = 24'(-54916);
			3751: out = 24'(-54836);
			3752: out = 24'(-54652);
			3753: out = 24'(-54456);
			3754: out = 24'(-54372);
			3755: out = 24'(-54240);
			3756: out = 24'(-54076);
			3757: out = 24'(-53748);
			3758: out = 24'(-53584);
			3759: out = 24'(-53472);
			3760: out = 24'(-53328);
			3761: out = 24'(-53140);
			3762: out = 24'(-53032);
			3763: out = 24'(-52796);
			3764: out = 24'(-52612);
			3765: out = 24'(-52392);
			3766: out = 24'(-52128);
			3767: out = 24'(-51916);
			3768: out = 24'(-51716);
			3769: out = 24'(-51500);
			3770: out = 24'(-51232);
			3771: out = 24'(-50988);
			3772: out = 24'(-50792);
			3773: out = 24'(-50508);
			3774: out = 24'(-50276);
			3775: out = 24'(-49980);
			3776: out = 24'(-49704);
			3777: out = 24'(-49392);
			3778: out = 24'(-49056);
			3779: out = 24'(-48876);
			3780: out = 24'(-48528);
			3781: out = 24'(-48164);
			3782: out = 24'(-47908);
			3783: out = 24'(-47580);
			3784: out = 24'(-47216);
			3785: out = 24'(-46920);
			3786: out = 24'(-46500);
			3787: out = 24'(-46212);
			3788: out = 24'(-45792);
			3789: out = 24'(-45372);
			3790: out = 24'(-45048);
			3791: out = 24'(-44620);
			3792: out = 24'(-44272);
			3793: out = 24'(-43800);
			3794: out = 24'(-43488);
			3795: out = 24'(-43116);
			3796: out = 24'(-42664);
			3797: out = 24'(-42264);
			3798: out = 24'(-41824);
			3799: out = 24'(-41472);
			3800: out = 24'(-41004);
			3801: out = 24'(-40576);
			3802: out = 24'(-40196);
			3803: out = 24'(-39736);
			3804: out = 24'(-39316);
			3805: out = 24'(-38912);
			3806: out = 24'(-38464);
			3807: out = 24'(-38012);
			3808: out = 24'(-37656);
			3809: out = 24'(-37224);
			3810: out = 24'(-36756);
			3811: out = 24'(-36296);
			3812: out = 24'(-35912);
			3813: out = 24'(-35432);
			3814: out = 24'(-35060);
			3815: out = 24'(-34624);
			3816: out = 24'(-34140);
			3817: out = 24'(-33736);
			3818: out = 24'(-33324);
			3819: out = 24'(-33000);
			3820: out = 24'(-32480);
			3821: out = 24'(-32164);
			3822: out = 24'(-31736);
			3823: out = 24'(-31300);
			3824: out = 24'(-30896);
			3825: out = 24'(-30504);
			3826: out = 24'(-30096);
			3827: out = 24'(-29684);
			3828: out = 24'(-29336);
			3829: out = 24'(-28888);
			3830: out = 24'(-28596);
			3831: out = 24'(-28200);
			3832: out = 24'(-27776);
			3833: out = 24'(-27408);
			3834: out = 24'(-26984);
			3835: out = 24'(-26676);
			3836: out = 24'(-26244);
			3837: out = 24'(-25956);
			3838: out = 24'(-25548);
			3839: out = 24'(-25240);
			3840: out = 24'(-24880);
			3841: out = 24'(-24552);
			3842: out = 24'(-24160);
			3843: out = 24'(-23836);
			3844: out = 24'(-23464);
			3845: out = 24'(-23124);
			3846: out = 24'(-22820);
			3847: out = 24'(-22468);
			3848: out = 24'(-22088);
			3849: out = 24'(-21856);
			3850: out = 24'(-21476);
			3851: out = 24'(-21132);
			3852: out = 24'(-20812);
			3853: out = 24'(-20548);
			3854: out = 24'(-20272);
			3855: out = 24'(-19872);
			3856: out = 24'(-19604);
			3857: out = 24'(-19408);
			3858: out = 24'(-19160);
			3859: out = 24'(-18812);
			3860: out = 24'(-18464);
			3861: out = 24'(-18252);
			3862: out = 24'(-17916);
			3863: out = 24'(-17628);
			3864: out = 24'(-17332);
			3865: out = 24'(-17096);
			3866: out = 24'(-16788);
			3867: out = 24'(-16536);
			3868: out = 24'(-16208);
			3869: out = 24'(-15984);
			3870: out = 24'(-15768);
			3871: out = 24'(-15500);
			3872: out = 24'(-15248);
			3873: out = 24'(-14972);
			3874: out = 24'(-14756);
			3875: out = 24'(-14432);
			3876: out = 24'(-14232);
			3877: out = 24'(-14016);
			3878: out = 24'(-13804);
			3879: out = 24'(-13508);
			3880: out = 24'(-13292);
			3881: out = 24'(-13104);
			3882: out = 24'(-12852);
			3883: out = 24'(-12664);
			3884: out = 24'(-12392);
			3885: out = 24'(-12248);
			3886: out = 24'(-11996);
			3887: out = 24'(-11588);
			3888: out = 24'(-11252);
			3889: out = 24'(-10852);
			3890: out = 24'(-10488);
			3891: out = 24'(-10100);
			3892: out = 24'(-9764);
			3893: out = 24'(-9376);
			3894: out = 24'(-9080);
			3895: out = 24'(-8636);
			3896: out = 24'(-8320);
			3897: out = 24'(-7988);
			3898: out = 24'(-7612);
			3899: out = 24'(-7316);
			3900: out = 24'(-7024);
			3901: out = 24'(-6692);
			3902: out = 24'(-6300);
			3903: out = 24'(-6068);
			3904: out = 24'(-5708);
			3905: out = 24'(-5484);
			3906: out = 24'(-5136);
			3907: out = 24'(-4836);
			3908: out = 24'(-4584);
			3909: out = 24'(-4248);
			3910: out = 24'(-3972);
			3911: out = 24'(-3704);
			3912: out = 24'(-3416);
			3913: out = 24'(-3148);
			3914: out = 24'(-2892);
			3915: out = 24'(-2564);
			3916: out = 24'(-2360);
			3917: out = 24'(-2136);
			3918: out = 24'(-1900);
			3919: out = 24'(-1548);
			3920: out = 24'(-1320);
			3921: out = 24'(-1032);
			3922: out = 24'(-832);
			3923: out = 24'(-584);
			3924: out = 24'(-344);
			3925: out = 24'(-164);
			3926: out = 24'(128);
			3927: out = 24'(360);
			3928: out = 24'(544);
			3929: out = 24'(820);
			3930: out = 24'(1060);
			3931: out = 24'(1268);
			3932: out = 24'(1564);
			3933: out = 24'(1752);
			3934: out = 24'(1880);
			3935: out = 24'(2152);
			3936: out = 24'(2400);
			3937: out = 24'(2620);
			3938: out = 24'(2892);
			3939: out = 24'(3048);
			3940: out = 24'(3280);
			3941: out = 24'(3476);
			3942: out = 24'(3704);
			3943: out = 24'(4000);
			3944: out = 24'(4228);
			3945: out = 24'(4372);
			3946: out = 24'(4604);
			3947: out = 24'(4776);
			3948: out = 24'(4988);
			3949: out = 24'(5176);
			3950: out = 24'(5376);
			3951: out = 24'(5576);
			3952: out = 24'(5836);
			3953: out = 24'(6072);
			3954: out = 24'(6224);
			3955: out = 24'(6508);
			3956: out = 24'(6696);
			3957: out = 24'(6920);
			3958: out = 24'(7112);
			3959: out = 24'(7388);
			3960: out = 24'(7552);
			3961: out = 24'(7796);
			3962: out = 24'(8024);
			3963: out = 24'(8240);
			3964: out = 24'(8448);
			3965: out = 24'(8740);
			3966: out = 24'(8984);
			3967: out = 24'(9176);
			3968: out = 24'(9356);
			3969: out = 24'(9660);
			3970: out = 24'(9860);
			3971: out = 24'(10100);
			3972: out = 24'(10400);
			3973: out = 24'(10592);
			3974: out = 24'(10904);
			3975: out = 24'(11136);
			3976: out = 24'(11400);
			3977: out = 24'(11684);
			3978: out = 24'(11976);
			3979: out = 24'(12228);
			3980: out = 24'(12468);
			3981: out = 24'(12776);
			3982: out = 24'(13124);
			3983: out = 24'(13432);
			3984: out = 24'(13720);
			3985: out = 24'(14076);
			3986: out = 24'(14376);
			3987: out = 24'(14644);
			3988: out = 24'(15012);
			3989: out = 24'(15424);
			3990: out = 24'(15728);
			3991: out = 24'(16112);
			3992: out = 24'(16464);
			3993: out = 24'(16828);
			3994: out = 24'(17164);
			3995: out = 24'(17564);
			3996: out = 24'(17916);
			3997: out = 24'(18276);
			3998: out = 24'(18640);
			3999: out = 24'(19056);
			4000: out = 24'(19420);
			4001: out = 24'(19808);
			4002: out = 24'(20196);
			4003: out = 24'(20624);
			4004: out = 24'(20984);
			4005: out = 24'(21368);
			4006: out = 24'(21764);
			4007: out = 24'(22164);
			4008: out = 24'(22556);
			4009: out = 24'(22952);
			4010: out = 24'(23400);
			4011: out = 24'(23784);
			4012: out = 24'(24100);
			4013: out = 24'(24536);
			4014: out = 24'(24948);
			4015: out = 24'(25328);
			4016: out = 24'(25776);
			4017: out = 24'(26160);
			4018: out = 24'(26540);
			4019: out = 24'(26908);
			4020: out = 24'(27304);
			4021: out = 24'(27744);
			4022: out = 24'(28072);
			4023: out = 24'(28420);
			4024: out = 24'(28716);
			4025: out = 24'(29200);
			4026: out = 24'(29532);
			4027: out = 24'(29948);
			4028: out = 24'(30320);
			4029: out = 24'(30620);
			4030: out = 24'(30960);
			4031: out = 24'(31352);
			4032: out = 24'(31652);
			4033: out = 24'(31920);
			4034: out = 24'(32316);
			4035: out = 24'(32620);
			4036: out = 24'(32996);
			4037: out = 24'(33276);
			4038: out = 24'(33684);
			4039: out = 24'(33928);
			4040: out = 24'(34244);
			4041: out = 24'(34612);
			4042: out = 24'(34856);
			4043: out = 24'(35156);
			4044: out = 24'(35496);
			4045: out = 24'(35772);
			4046: out = 24'(36080);
			4047: out = 24'(36364);
			4048: out = 24'(36648);
			4049: out = 24'(36952);
			4050: out = 24'(37212);
			4051: out = 24'(37468);
			4052: out = 24'(37732);
			4053: out = 24'(37980);
			4054: out = 24'(38248);
			4055: out = 24'(38516);
			4056: out = 24'(38772);
			4057: out = 24'(39056);
			4058: out = 24'(39312);
			4059: out = 24'(39536);
			4060: out = 24'(39748);
			4061: out = 24'(40080);
			4062: out = 24'(40272);
			4063: out = 24'(40592);
			4064: out = 24'(40768);
			4065: out = 24'(40960);
			4066: out = 24'(41240);
			4067: out = 24'(41392);
			4068: out = 24'(41684);
			4069: out = 24'(41824);
			4070: out = 24'(42096);
			4071: out = 24'(42280);
			4072: out = 24'(42544);
			4073: out = 24'(42712);
			4074: out = 24'(42904);
			4075: out = 24'(43028);
			4076: out = 24'(43312);
			4077: out = 24'(43468);
			4078: out = 24'(43684);
			4079: out = 24'(43900);
			4080: out = 24'(44076);
			4081: out = 24'(44228);
			4082: out = 24'(44404);
			4083: out = 24'(44644);
			4084: out = 24'(44804);
			4085: out = 24'(44996);
			4086: out = 24'(45148);
			4087: out = 24'(45284);
			4088: out = 24'(45452);
			4089: out = 24'(45632);
			4090: out = 24'(45840);
			4091: out = 24'(46032);
			4092: out = 24'(46188);
			4093: out = 24'(46380);
			4094: out = 24'(46464);
			4095: out = 24'(46664);
			4096: out = 24'(46832);
			4097: out = 24'(46980);
			4098: out = 24'(47104);
			4099: out = 24'(47244);
			4100: out = 24'(47424);
			4101: out = 24'(47632);
			4102: out = 24'(47772);
			4103: out = 24'(47916);
			4104: out = 24'(48052);
			4105: out = 24'(48188);
			4106: out = 24'(48340);
			4107: out = 24'(48508);
			4108: out = 24'(48652);
			4109: out = 24'(48808);
			4110: out = 24'(48880);
			4111: out = 24'(49020);
			4112: out = 24'(49228);
			4113: out = 24'(49296);
			4114: out = 24'(49476);
			4115: out = 24'(49552);
			4116: out = 24'(49660);
			4117: out = 24'(49764);
			4118: out = 24'(49768);
			4119: out = 24'(49868);
			4120: out = 24'(49956);
			4121: out = 24'(49904);
			4122: out = 24'(49740);
			4123: out = 24'(49880);
			4124: out = 24'(49808);
			4125: out = 24'(49592);
			4126: out = 24'(49612);
			4127: out = 24'(49684);
			4128: out = 24'(49684);
			4129: out = 24'(49720);
			4130: out = 24'(49676);
			4131: out = 24'(49432);
			4132: out = 24'(49520);
			4133: out = 24'(49500);
			4134: out = 24'(49512);
			4135: out = 24'(49412);
			4136: out = 24'(49376);
			4137: out = 24'(49316);
			4138: out = 24'(49112);
			4139: out = 24'(48964);
			4140: out = 24'(48984);
			4141: out = 24'(48892);
			4142: out = 24'(48840);
			4143: out = 24'(48972);
			4144: out = 24'(48992);
			4145: out = 24'(48876);
			4146: out = 24'(48652);
			4147: out = 24'(48660);
			4148: out = 24'(48676);
			4149: out = 24'(48596);
			4150: out = 24'(48696);
			4151: out = 24'(48648);
			4152: out = 24'(48432);
			4153: out = 24'(48452);
			4154: out = 24'(48440);
			4155: out = 24'(48424);
			4156: out = 24'(48576);
			4157: out = 24'(48488);
			4158: out = 24'(48188);
			4159: out = 24'(48164);
			4160: out = 24'(48048);
			4161: out = 24'(48212);
			4162: out = 24'(48208);
			4163: out = 24'(48076);
			4164: out = 24'(48080);
			4165: out = 24'(48168);
			4166: out = 24'(48176);
			4167: out = 24'(48028);
			4168: out = 24'(47860);
			4169: out = 24'(47856);
			4170: out = 24'(47676);
			4171: out = 24'(47752);
			4172: out = 24'(47812);
			4173: out = 24'(47840);
			4174: out = 24'(47820);
			4175: out = 24'(47752);
			4176: out = 24'(47708);
			4177: out = 24'(47700);
			4178: out = 24'(47572);
			4179: out = 24'(47416);
			4180: out = 24'(47340);
			4181: out = 24'(47460);
			4182: out = 24'(47164);
			4183: out = 24'(46876);
			4184: out = 24'(46844);
			4185: out = 24'(46660);
			4186: out = 24'(46636);
			4187: out = 24'(46744);
			4188: out = 24'(46768);
			4189: out = 24'(46544);
			4190: out = 24'(46476);
			4191: out = 24'(46188);
			4192: out = 24'(46068);
			4193: out = 24'(46064);
			4194: out = 24'(45920);
			4195: out = 24'(45780);
			4196: out = 24'(45756);
			4197: out = 24'(45492);
			4198: out = 24'(45436);
			4199: out = 24'(45172);
			4200: out = 24'(44852);
			4201: out = 24'(44820);
			4202: out = 24'(44796);
			4203: out = 24'(44520);
			4204: out = 24'(44104);
			4205: out = 24'(44044);
			4206: out = 24'(43916);
			4207: out = 24'(43724);
			4208: out = 24'(43456);
			4209: out = 24'(43296);
			4210: out = 24'(43116);
			4211: out = 24'(42832);
			4212: out = 24'(42404);
			4213: out = 24'(42168);
			4214: out = 24'(41956);
			4215: out = 24'(41636);
			4216: out = 24'(41380);
			4217: out = 24'(41184);
			4218: out = 24'(40932);
			4219: out = 24'(40672);
			4220: out = 24'(40432);
			4221: out = 24'(40164);
			4222: out = 24'(39836);
			4223: out = 24'(39468);
			4224: out = 24'(39156);
			4225: out = 24'(38940);
			4226: out = 24'(38544);
			4227: out = 24'(38288);
			4228: out = 24'(37904);
			4229: out = 24'(37656);
			4230: out = 24'(37404);
			4231: out = 24'(37096);
			4232: out = 24'(36748);
			4233: out = 24'(36412);
			4234: out = 24'(36092);
			4235: out = 24'(35740);
			4236: out = 24'(35480);
			4237: out = 24'(35136);
			4238: out = 24'(34840);
			4239: out = 24'(34432);
			4240: out = 24'(34188);
			4241: out = 24'(33860);
			4242: out = 24'(33460);
			4243: out = 24'(33188);
			4244: out = 24'(32936);
			4245: out = 24'(32692);
			4246: out = 24'(32192);
			4247: out = 24'(31936);
			4248: out = 24'(31636);
			4249: out = 24'(31264);
			4250: out = 24'(30916);
			4251: out = 24'(30616);
			4252: out = 24'(30344);
			4253: out = 24'(30028);
			4254: out = 24'(29736);
			4255: out = 24'(29476);
			4256: out = 24'(29128);
			4257: out = 24'(28820);
			4258: out = 24'(28516);
			4259: out = 24'(28176);
			4260: out = 24'(27896);
			4261: out = 24'(27492);
			4262: out = 24'(27164);
			4263: out = 24'(26940);
			4264: out = 24'(26640);
			4265: out = 24'(26360);
			4266: out = 24'(25992);
			4267: out = 24'(25668);
			4268: out = 24'(25424);
			4269: out = 24'(25188);
			4270: out = 24'(24932);
			4271: out = 24'(24624);
			4272: out = 24'(24324);
			4273: out = 24'(23988);
			4274: out = 24'(23672);
			4275: out = 24'(23504);
			4276: out = 24'(23232);
			4277: out = 24'(22968);
			4278: out = 24'(22656);
			4279: out = 24'(22408);
			4280: out = 24'(22112);
			4281: out = 24'(21780);
			4282: out = 24'(21576);
			4283: out = 24'(21312);
			4284: out = 24'(21012);
			4285: out = 24'(20756);
			4286: out = 24'(20512);
			4287: out = 24'(20280);
			4288: out = 24'(20000);
			4289: out = 24'(19876);
			4290: out = 24'(19552);
			4291: out = 24'(19336);
			4292: out = 24'(19076);
			4293: out = 24'(18800);
			4294: out = 24'(18608);
			4295: out = 24'(18344);
			4296: out = 24'(18028);
			4297: out = 24'(17776);
			4298: out = 24'(17552);
			4299: out = 24'(17444);
			4300: out = 24'(17120);
			4301: out = 24'(16900);
			4302: out = 24'(16704);
			4303: out = 24'(16492);
			4304: out = 24'(16260);
			4305: out = 24'(16128);
			4306: out = 24'(15832);
			4307: out = 24'(15560);
			4308: out = 24'(15332);
			4309: out = 24'(15076);
			4310: out = 24'(15008);
			4311: out = 24'(14824);
			4312: out = 24'(14572);
			4313: out = 24'(14488);
			4314: out = 24'(14272);
			4315: out = 24'(14024);
			4316: out = 24'(13836);
			4317: out = 24'(13612);
			4318: out = 24'(13464);
			4319: out = 24'(13264);
			4320: out = 24'(13144);
			4321: out = 24'(12932);
			4322: out = 24'(12720);
			4323: out = 24'(12560);
			4324: out = 24'(12412);
			4325: out = 24'(12192);
			4326: out = 24'(11984);
			4327: out = 24'(11872);
			4328: out = 24'(11732);
			4329: out = 24'(11508);
			4330: out = 24'(11376);
			4331: out = 24'(11208);
			4332: out = 24'(10948);
			4333: out = 24'(10848);
			4334: out = 24'(10692);
			4335: out = 24'(10592);
			4336: out = 24'(10428);
			4337: out = 24'(10232);
			4338: out = 24'(10108);
			4339: out = 24'(9904);
			4340: out = 24'(9784);
			4341: out = 24'(9704);
			4342: out = 24'(9504);
			4343: out = 24'(9408);
			4344: out = 24'(9176);
			4345: out = 24'(9124);
			4346: out = 24'(8988);
			4347: out = 24'(8744);
			4348: out = 24'(8536);
			4349: out = 24'(8116);
			4350: out = 24'(7800);
			4351: out = 24'(7404);
			4352: out = 24'(7088);
			4353: out = 24'(6660);
			4354: out = 24'(6336);
			4355: out = 24'(5956);
			4356: out = 24'(5668);
			4357: out = 24'(5312);
			4358: out = 24'(4912);
			4359: out = 24'(4616);
			4360: out = 24'(4232);
			4361: out = 24'(3896);
			4362: out = 24'(3580);
			4363: out = 24'(3324);
			4364: out = 24'(2996);
			4365: out = 24'(2676);
			4366: out = 24'(2464);
			4367: out = 24'(2108);
			4368: out = 24'(1792);
			4369: out = 24'(1544);
			4370: out = 24'(1212);
			4371: out = 24'(984);
			4372: out = 24'(616);
			4373: out = 24'(356);
			4374: out = 24'(124);
			4375: out = 24'(-152);
			4376: out = 24'(-380);
			4377: out = 24'(-644);
			4378: out = 24'(-952);
			4379: out = 24'(-1284);
			4380: out = 24'(-1432);
			4381: out = 24'(-1692);
			4382: out = 24'(-1984);
			4383: out = 24'(-2180);
			4384: out = 24'(-2476);
			4385: out = 24'(-2728);
			4386: out = 24'(-2992);
			4387: out = 24'(-3196);
			4388: out = 24'(-3436);
			4389: out = 24'(-3652);
			4390: out = 24'(-3872);
			4391: out = 24'(-4076);
			4392: out = 24'(-4224);
			4393: out = 24'(-4480);
			4394: out = 24'(-4768);
			4395: out = 24'(-5040);
			4396: out = 24'(-5284);
			4397: out = 24'(-5508);
			4398: out = 24'(-5788);
			4399: out = 24'(-6000);
			4400: out = 24'(-6184);
			4401: out = 24'(-6364);
			4402: out = 24'(-6636);
			4403: out = 24'(-6852);
			4404: out = 24'(-7036);
			4405: out = 24'(-7236);
			4406: out = 24'(-7480);
			4407: out = 24'(-7648);
			4408: out = 24'(-7876);
			4409: out = 24'(-8100);
			4410: out = 24'(-8308);
			4411: out = 24'(-8588);
			4412: out = 24'(-8776);
			4413: out = 24'(-8936);
			4414: out = 24'(-9244);
			4415: out = 24'(-9424);
			4416: out = 24'(-9624);
			4417: out = 24'(-9812);
			4418: out = 24'(-10036);
			4419: out = 24'(-10236);
			4420: out = 24'(-10428);
			4421: out = 24'(-10604);
			4422: out = 24'(-10872);
			4423: out = 24'(-11100);
			4424: out = 24'(-11248);
			4425: out = 24'(-11488);
			4426: out = 24'(-11724);
			4427: out = 24'(-11980);
			4428: out = 24'(-12136);
			4429: out = 24'(-12336);
			4430: out = 24'(-12572);
			4431: out = 24'(-12792);
			4432: out = 24'(-13024);
			4433: out = 24'(-13276);
			4434: out = 24'(-13556);
			4435: out = 24'(-13808);
			4436: out = 24'(-14036);
			4437: out = 24'(-14384);
			4438: out = 24'(-14620);
			4439: out = 24'(-14872);
			4440: out = 24'(-15148);
			4441: out = 24'(-15408);
			4442: out = 24'(-15652);
			4443: out = 24'(-15968);
			4444: out = 24'(-16240);
			4445: out = 24'(-16572);
			4446: out = 24'(-16892);
			4447: out = 24'(-17116);
			4448: out = 24'(-17476);
			4449: out = 24'(-17784);
			4450: out = 24'(-18064);
			4451: out = 24'(-18340);
			4452: out = 24'(-18736);
			4453: out = 24'(-18972);
			4454: out = 24'(-19284);
			4455: out = 24'(-19652);
			4456: out = 24'(-19976);
			4457: out = 24'(-20296);
			4458: out = 24'(-20692);
			4459: out = 24'(-21012);
			4460: out = 24'(-21384);
			4461: out = 24'(-21808);
			4462: out = 24'(-22128);
			4463: out = 24'(-22496);
			4464: out = 24'(-22888);
			4465: out = 24'(-23260);
			4466: out = 24'(-23628);
			4467: out = 24'(-24060);
			4468: out = 24'(-24512);
			4469: out = 24'(-24852);
			4470: out = 24'(-25232);
			4471: out = 24'(-25648);
			4472: out = 24'(-26100);
			4473: out = 24'(-26524);
			4474: out = 24'(-26984);
			4475: out = 24'(-27372);
			4476: out = 24'(-27740);
			4477: out = 24'(-28192);
			4478: out = 24'(-28632);
			4479: out = 24'(-29124);
			4480: out = 24'(-29524);
			4481: out = 24'(-29980);
			4482: out = 24'(-30420);
			4483: out = 24'(-30880);
			4484: out = 24'(-31340);
			4485: out = 24'(-31768);
			4486: out = 24'(-32204);
			4487: out = 24'(-32668);
			4488: out = 24'(-33016);
			4489: out = 24'(-33448);
			4490: out = 24'(-33820);
			4491: out = 24'(-34292);
			4492: out = 24'(-34652);
			4493: out = 24'(-35096);
			4494: out = 24'(-35496);
			4495: out = 24'(-35800);
			4496: out = 24'(-36172);
			4497: out = 24'(-36556);
			4498: out = 24'(-36924);
			4499: out = 24'(-37252);
			4500: out = 24'(-37608);
			4501: out = 24'(-37904);
			4502: out = 24'(-38208);
			4503: out = 24'(-38512);
			4504: out = 24'(-38824);
			4505: out = 24'(-39120);
			4506: out = 24'(-39512);
			4507: out = 24'(-39756);
			4508: out = 24'(-40128);
			4509: out = 24'(-40432);
			4510: out = 24'(-40684);
			4511: out = 24'(-41008);
			4512: out = 24'(-41236);
			4513: out = 24'(-41588);
			4514: out = 24'(-41808);
			4515: out = 24'(-42088);
			4516: out = 24'(-42308);
			4517: out = 24'(-42596);
			4518: out = 24'(-42812);
			4519: out = 24'(-43064);
			4520: out = 24'(-43272);
			4521: out = 24'(-43556);
			4522: out = 24'(-43672);
			4523: out = 24'(-43920);
			4524: out = 24'(-44156);
			4525: out = 24'(-44360);
			4526: out = 24'(-44480);
			4527: out = 24'(-44784);
			4528: out = 24'(-44900);
			4529: out = 24'(-45008);
			4530: out = 24'(-45260);
			4531: out = 24'(-45416);
			4532: out = 24'(-45604);
			4533: out = 24'(-45708);
			4534: out = 24'(-45848);
			4535: out = 24'(-45964);
			4536: out = 24'(-46156);
			4537: out = 24'(-46308);
			4538: out = 24'(-46360);
			4539: out = 24'(-46524);
			4540: out = 24'(-46596);
			4541: out = 24'(-46728);
			4542: out = 24'(-46876);
			4543: out = 24'(-46968);
			4544: out = 24'(-47088);
			4545: out = 24'(-47124);
			4546: out = 24'(-47224);
			4547: out = 24'(-47340);
			4548: out = 24'(-47456);
			4549: out = 24'(-47480);
			4550: out = 24'(-47560);
			4551: out = 24'(-47628);
			4552: out = 24'(-47660);
			4553: out = 24'(-47676);
			4554: out = 24'(-47828);
			4555: out = 24'(-47832);
			4556: out = 24'(-47880);
			4557: out = 24'(-47876);
			4558: out = 24'(-48028);
			4559: out = 24'(-47988);
			4560: out = 24'(-48056);
			4561: out = 24'(-48056);
			4562: out = 24'(-48080);
			4563: out = 24'(-48040);
			4564: out = 24'(-48144);
			4565: out = 24'(-48144);
			4566: out = 24'(-48144);
			4567: out = 24'(-48188);
			4568: out = 24'(-48204);
			4569: out = 24'(-48220);
			4570: out = 24'(-48364);
			4571: out = 24'(-48316);
			4572: out = 24'(-48292);
			4573: out = 24'(-48256);
			4574: out = 24'(-48236);
			4575: out = 24'(-48272);
			4576: out = 24'(-48172);
			4577: out = 24'(-48196);
			4578: out = 24'(-48172);
			4579: out = 24'(-48164);
			4580: out = 24'(-48156);
			4581: out = 24'(-48084);
			4582: out = 24'(-48112);
			4583: out = 24'(-48092);
			4584: out = 24'(-48048);
			4585: out = 24'(-48052);
			4586: out = 24'(-47956);
			4587: out = 24'(-47936);
			4588: out = 24'(-47884);
			4589: out = 24'(-47892);
			4590: out = 24'(-47872);
			4591: out = 24'(-47772);
			4592: out = 24'(-47744);
			4593: out = 24'(-47676);
			4594: out = 24'(-47632);
			4595: out = 24'(-47564);
			4596: out = 24'(-47548);
			4597: out = 24'(-47396);
			4598: out = 24'(-47388);
			4599: out = 24'(-47340);
			4600: out = 24'(-47300);
			4601: out = 24'(-47248);
			4602: out = 24'(-47140);
			4603: out = 24'(-47056);
			4604: out = 24'(-47024);
			4605: out = 24'(-46928);
			4606: out = 24'(-46828);
			4607: out = 24'(-46828);
			4608: out = 24'(-46736);
			4609: out = 24'(-46608);
			4610: out = 24'(-46600);
			4611: out = 24'(-46492);
			4612: out = 24'(-46452);
			4613: out = 24'(-46348);
			4614: out = 24'(-46236);
			4615: out = 24'(-46216);
			4616: out = 24'(-46044);
			4617: out = 24'(-45972);
			4618: out = 24'(-45892);
			4619: out = 24'(-45792);
			4620: out = 24'(-45680);
			4621: out = 24'(-45624);
			4622: out = 24'(-45452);
			4623: out = 24'(-45372);
			4624: out = 24'(-45320);
			4625: out = 24'(-45212);
			4626: out = 24'(-45016);
			4627: out = 24'(-44944);
			4628: out = 24'(-44864);
			4629: out = 24'(-44720);
			4630: out = 24'(-44600);
			4631: out = 24'(-44536);
			4632: out = 24'(-44448);
			4633: out = 24'(-44300);
			4634: out = 24'(-44128);
			4635: out = 24'(-44128);
			4636: out = 24'(-43928);
			4637: out = 24'(-43772);
			4638: out = 24'(-43696);
			4639: out = 24'(-43556);
			4640: out = 24'(-43348);
			4641: out = 24'(-43272);
			4642: out = 24'(-43100);
			4643: out = 24'(-42952);
			4644: out = 24'(-42808);
			4645: out = 24'(-42648);
			4646: out = 24'(-42472);
			4647: out = 24'(-42340);
			4648: out = 24'(-42148);
			4649: out = 24'(-41956);
			4650: out = 24'(-41724);
			4651: out = 24'(-41644);
			4652: out = 24'(-41360);
			4653: out = 24'(-41208);
			4654: out = 24'(-40924);
			4655: out = 24'(-40700);
			4656: out = 24'(-40568);
			4657: out = 24'(-40316);
			4658: out = 24'(-40096);
			4659: out = 24'(-39860);
			4660: out = 24'(-39676);
			4661: out = 24'(-39352);
			4662: out = 24'(-39172);
			4663: out = 24'(-38800);
			4664: out = 24'(-38612);
			4665: out = 24'(-38344);
			4666: out = 24'(-38076);
			4667: out = 24'(-37780);
			4668: out = 24'(-37484);
			4669: out = 24'(-37200);
			4670: out = 24'(-36884);
			4671: out = 24'(-36604);
			4672: out = 24'(-36316);
			4673: out = 24'(-36008);
			4674: out = 24'(-35680);
			4675: out = 24'(-35336);
			4676: out = 24'(-35048);
			4677: out = 24'(-34704);
			4678: out = 24'(-34356);
			4679: out = 24'(-34048);
			4680: out = 24'(-33616);
			4681: out = 24'(-33380);
			4682: out = 24'(-33024);
			4683: out = 24'(-32608);
			4684: out = 24'(-32336);
			4685: out = 24'(-31944);
			4686: out = 24'(-31604);
			4687: out = 24'(-31260);
			4688: out = 24'(-30960);
			4689: out = 24'(-30584);
			4690: out = 24'(-30220);
			4691: out = 24'(-29928);
			4692: out = 24'(-29520);
			4693: out = 24'(-29192);
			4694: out = 24'(-28856);
			4695: out = 24'(-28556);
			4696: out = 24'(-28180);
			4697: out = 24'(-27884);
			4698: out = 24'(-27448);
			4699: out = 24'(-27200);
			4700: out = 24'(-26872);
			4701: out = 24'(-26512);
			4702: out = 24'(-26212);
			4703: out = 24'(-25780);
			4704: out = 24'(-25592);
			4705: out = 24'(-25208);
			4706: out = 24'(-24888);
			4707: out = 24'(-24540);
			4708: out = 24'(-24192);
			4709: out = 24'(-23892);
			4710: out = 24'(-23580);
			4711: out = 24'(-23320);
			4712: out = 24'(-22992);
			4713: out = 24'(-22656);
			4714: out = 24'(-22332);
			4715: out = 24'(-22040);
			4716: out = 24'(-21708);
			4717: out = 24'(-21428);
			4718: out = 24'(-21132);
			4719: out = 24'(-20796);
			4720: out = 24'(-20516);
			4721: out = 24'(-20244);
			4722: out = 24'(-19912);
			4723: out = 24'(-19664);
			4724: out = 24'(-19324);
			4725: out = 24'(-19064);
			4726: out = 24'(-18772);
			4727: out = 24'(-18444);
			4728: out = 24'(-18296);
			4729: out = 24'(-17932);
			4730: out = 24'(-17692);
			4731: out = 24'(-17440);
			4732: out = 24'(-17172);
			4733: out = 24'(-16908);
			4734: out = 24'(-16688);
			4735: out = 24'(-16436);
			4736: out = 24'(-16180);
			4737: out = 24'(-15928);
			4738: out = 24'(-15668);
			4739: out = 24'(-15472);
			4740: out = 24'(-15220);
			4741: out = 24'(-14968);
			4742: out = 24'(-14724);
			4743: out = 24'(-14504);
			4744: out = 24'(-14284);
			4745: out = 24'(-14068);
			4746: out = 24'(-13812);
			4747: out = 24'(-13652);
			4748: out = 24'(-13372);
			4749: out = 24'(-13160);
			4750: out = 24'(-13000);
			4751: out = 24'(-12712);
			4752: out = 24'(-12576);
			4753: out = 24'(-12312);
			4754: out = 24'(-12140);
			4755: out = 24'(-11964);
			4756: out = 24'(-11800);
			4757: out = 24'(-11552);
			4758: out = 24'(-11336);
			4759: out = 24'(-11184);
			4760: out = 24'(-10952);
			4761: out = 24'(-10728);
			4762: out = 24'(-10568);
			4763: out = 24'(-10420);
			4764: out = 24'(-10244);
			4765: out = 24'(-10012);
			4766: out = 24'(-9860);
			4767: out = 24'(-9684);
			4768: out = 24'(-9528);
			4769: out = 24'(-9356);
			4770: out = 24'(-9104);
			4771: out = 24'(-8824);
			4772: out = 24'(-8536);
			4773: out = 24'(-8176);
			4774: out = 24'(-7920);
			4775: out = 24'(-7556);
			4776: out = 24'(-7292);
			4777: out = 24'(-7016);
			4778: out = 24'(-6728);
			4779: out = 24'(-6460);
			4780: out = 24'(-6208);
			4781: out = 24'(-5896);
			4782: out = 24'(-5624);
			4783: out = 24'(-5404);
			4784: out = 24'(-5116);
			4785: out = 24'(-4900);
			4786: out = 24'(-4612);
			4787: out = 24'(-4408);
			4788: out = 24'(-4144);
			4789: out = 24'(-3892);
			4790: out = 24'(-3660);
			4791: out = 24'(-3388);
			4792: out = 24'(-3208);
			4793: out = 24'(-2960);
			4794: out = 24'(-2720);
			4795: out = 24'(-2540);
			4796: out = 24'(-2308);
			4797: out = 24'(-2064);
			4798: out = 24'(-1876);
			4799: out = 24'(-1644);
			4800: out = 24'(-1392);
			4801: out = 24'(-1224);
			4802: out = 24'(-1056);
			4803: out = 24'(-840);
			4804: out = 24'(-588);
			4805: out = 24'(-408);
			4806: out = 24'(-244);
			4807: out = 24'(-76);
			4808: out = 24'(108);
			4809: out = 24'(352);
			4810: out = 24'(500);
			4811: out = 24'(668);
			4812: out = 24'(908);
			4813: out = 24'(1080);
			4814: out = 24'(1268);
			4815: out = 24'(1396);
			4816: out = 24'(1604);
			4817: out = 24'(1752);
			4818: out = 24'(1960);
			4819: out = 24'(2116);
			4820: out = 24'(2296);
			4821: out = 24'(2500);
			4822: out = 24'(2676);
			4823: out = 24'(2828);
			4824: out = 24'(3024);
			4825: out = 24'(3184);
			4826: out = 24'(3340);
			4827: out = 24'(3560);
			4828: out = 24'(3680);
			4829: out = 24'(3844);
			4830: out = 24'(4000);
			4831: out = 24'(4188);
			4832: out = 24'(4368);
			4833: out = 24'(4532);
			4834: out = 24'(4740);
			4835: out = 24'(4852);
			4836: out = 24'(5104);
			4837: out = 24'(5164);
			4838: out = 24'(5400);
			4839: out = 24'(5560);
			4840: out = 24'(5744);
			4841: out = 24'(5940);
			4842: out = 24'(6144);
			4843: out = 24'(6284);
			4844: out = 24'(6428);
			4845: out = 24'(6592);
			4846: out = 24'(6788);
			4847: out = 24'(6896);
			4848: out = 24'(7096);
			4849: out = 24'(7292);
			4850: out = 24'(7436);
			4851: out = 24'(7700);
			4852: out = 24'(7812);
			4853: out = 24'(8056);
			4854: out = 24'(8204);
			4855: out = 24'(8420);
			4856: out = 24'(8608);
			4857: out = 24'(8792);
			4858: out = 24'(8980);
			4859: out = 24'(9172);
			4860: out = 24'(9352);
			4861: out = 24'(9588);
			4862: out = 24'(9792);
			4863: out = 24'(10056);
			4864: out = 24'(10256);
			4865: out = 24'(10512);
			4866: out = 24'(10760);
			4867: out = 24'(11024);
			4868: out = 24'(11220);
			4869: out = 24'(11492);
			4870: out = 24'(11732);
			4871: out = 24'(11976);
			4872: out = 24'(12276);
			4873: out = 24'(12516);
			4874: out = 24'(12796);
			4875: out = 24'(13104);
			4876: out = 24'(13360);
			4877: out = 24'(13616);
			4878: out = 24'(13888);
			4879: out = 24'(14224);
			4880: out = 24'(14472);
			4881: out = 24'(14704);
			4882: out = 24'(15084);
			4883: out = 24'(15368);
			4884: out = 24'(15704);
			4885: out = 24'(15976);
			4886: out = 24'(16384);
			4887: out = 24'(16604);
			4888: out = 24'(16936);
			4889: out = 24'(17272);
			4890: out = 24'(17604);
			4891: out = 24'(17852);
			4892: out = 24'(18240);
			4893: out = 24'(18524);
			4894: out = 24'(18856);
			4895: out = 24'(19180);
			4896: out = 24'(19536);
			4897: out = 24'(19852);
			4898: out = 24'(20184);
			4899: out = 24'(20472);
			4900: out = 24'(20804);
			4901: out = 24'(21140);
			4902: out = 24'(21424);
			4903: out = 24'(21768);
			4904: out = 24'(22088);
			4905: out = 24'(22332);
			4906: out = 24'(22724);
			4907: out = 24'(23052);
			4908: out = 24'(23328);
			4909: out = 24'(23676);
			4910: out = 24'(23928);
			4911: out = 24'(24244);
			4912: out = 24'(24500);
			4913: out = 24'(24824);
			4914: out = 24'(25128);
			4915: out = 24'(25384);
			4916: out = 24'(25692);
			4917: out = 24'(25880);
			4918: out = 24'(26216);
			4919: out = 24'(26484);
			4920: out = 24'(26768);
			4921: out = 24'(26964);
			4922: out = 24'(27276);
			4923: out = 24'(27532);
			4924: out = 24'(27760);
			4925: out = 24'(28056);
			4926: out = 24'(28284);
			4927: out = 24'(28584);
			4928: out = 24'(28752);
			4929: out = 24'(29008);
			4930: out = 24'(29280);
			4931: out = 24'(29472);
			4932: out = 24'(29728);
			4933: out = 24'(29928);
			4934: out = 24'(30192);
			4935: out = 24'(30452);
			4936: out = 24'(30676);
			4937: out = 24'(30872);
			4938: out = 24'(31188);
			4939: out = 24'(31336);
			4940: out = 24'(31576);
			4941: out = 24'(31764);
			4942: out = 24'(32040);
			4943: out = 24'(32240);
			4944: out = 24'(32460);
			4945: out = 24'(32632);
			4946: out = 24'(32912);
			4947: out = 24'(33040);
			4948: out = 24'(33332);
			4949: out = 24'(33444);
			4950: out = 24'(33632);
			4951: out = 24'(33832);
			4952: out = 24'(33988);
			4953: out = 24'(34200);
			4954: out = 24'(34360);
			4955: out = 24'(34520);
			4956: out = 24'(34644);
			4957: out = 24'(34868);
			4958: out = 24'(35028);
			4959: out = 24'(35184);
			4960: out = 24'(35372);
			4961: out = 24'(35456);
			4962: out = 24'(35684);
			4963: out = 24'(35776);
			4964: out = 24'(35960);
			4965: out = 24'(36180);
			4966: out = 24'(36272);
			4967: out = 24'(36392);
			4968: out = 24'(36600);
			4969: out = 24'(36772);
			4970: out = 24'(36924);
			4971: out = 24'(37084);
			4972: out = 24'(37232);
			4973: out = 24'(37408);
			4974: out = 24'(37508);
			4975: out = 24'(37636);
			4976: out = 24'(37836);
			4977: out = 24'(37936);
			4978: out = 24'(38108);
			4979: out = 24'(38172);
			4980: out = 24'(38388);
			4981: out = 24'(38540);
			4982: out = 24'(38636);
			4983: out = 24'(38768);
			4984: out = 24'(38920);
			4985: out = 24'(39060);
			4986: out = 24'(39124);
			4987: out = 24'(39264);
			4988: out = 24'(39400);
			4989: out = 24'(39528);
			4990: out = 24'(39628);
			4991: out = 24'(39736);
			4992: out = 24'(39908);
			4993: out = 24'(39984);
			4994: out = 24'(40076);
			4995: out = 24'(40220);
			4996: out = 24'(40340);
			4997: out = 24'(40416);
			4998: out = 24'(40536);
			4999: out = 24'(40628);
			5000: out = 24'(40728);
			5001: out = 24'(40864);
			5002: out = 24'(40908);
			5003: out = 24'(40976);
			5004: out = 24'(41068);
			5005: out = 24'(41140);
			5006: out = 24'(41124);
			5007: out = 24'(41060);
			5008: out = 24'(41120);
			5009: out = 24'(40924);
			5010: out = 24'(40932);
			5011: out = 24'(41088);
			5012: out = 24'(40984);
			5013: out = 24'(40916);
			5014: out = 24'(40720);
			5015: out = 24'(40768);
			5016: out = 24'(40592);
			5017: out = 24'(40636);
			5018: out = 24'(40692);
			5019: out = 24'(40604);
			5020: out = 24'(40628);
			5021: out = 24'(40524);
			5022: out = 24'(40500);
			5023: out = 24'(40424);
			5024: out = 24'(40572);
			5025: out = 24'(40496);
			5026: out = 24'(40364);
			5027: out = 24'(40456);
			5028: out = 24'(40376);
			5029: out = 24'(40444);
			5030: out = 24'(40492);
			5031: out = 24'(40360);
			5032: out = 24'(40408);
			5033: out = 24'(40336);
			5034: out = 24'(40348);
			5035: out = 24'(40296);
			5036: out = 24'(40260);
			5037: out = 24'(40216);
			5038: out = 24'(40212);
			5039: out = 24'(40100);
			5040: out = 24'(40124);
			5041: out = 24'(40100);
			5042: out = 24'(40112);
			5043: out = 24'(40144);
			5044: out = 24'(40016);
			5045: out = 24'(40084);
			5046: out = 24'(39980);
			5047: out = 24'(40036);
			5048: out = 24'(40008);
			5049: out = 24'(39880);
			5050: out = 24'(39748);
			5051: out = 24'(39764);
			5052: out = 24'(39808);
			5053: out = 24'(39896);
			5054: out = 24'(39868);
			5055: out = 24'(39936);
			5056: out = 24'(39904);
			5057: out = 24'(39764);
			5058: out = 24'(39748);
			5059: out = 24'(39708);
			5060: out = 24'(39660);
			5061: out = 24'(39580);
			5062: out = 24'(39424);
			5063: out = 24'(39316);
			5064: out = 24'(39324);
			5065: out = 24'(39280);
			5066: out = 24'(39164);
			5067: out = 24'(38992);
			5068: out = 24'(38988);
			5069: out = 24'(38980);
			5070: out = 24'(39028);
			5071: out = 24'(38984);
			5072: out = 24'(38920);
			5073: out = 24'(38804);
			5074: out = 24'(38508);
			5075: out = 24'(38620);
			5076: out = 24'(38376);
			5077: out = 24'(38360);
			5078: out = 24'(38296);
			5079: out = 24'(38112);
			5080: out = 24'(38116);
			5081: out = 24'(37948);
			5082: out = 24'(37944);
			5083: out = 24'(37804);
			5084: out = 24'(37756);
			5085: out = 24'(37648);
			5086: out = 24'(37596);
			5087: out = 24'(37332);
			5088: out = 24'(37176);
			5089: out = 24'(36988);
			5090: out = 24'(36740);
			5091: out = 24'(36672);
			5092: out = 24'(36500);
			5093: out = 24'(36236);
			5094: out = 24'(36044);
			5095: out = 24'(35960);
			5096: out = 24'(35656);
			5097: out = 24'(35560);
			5098: out = 24'(35344);
			5099: out = 24'(35128);
			5100: out = 24'(34864);
			5101: out = 24'(34636);
			5102: out = 24'(34524);
			5103: out = 24'(34332);
			5104: out = 24'(34192);
			5105: out = 24'(33912);
			5106: out = 24'(33692);
			5107: out = 24'(33448);
			5108: out = 24'(33184);
			5109: out = 24'(32948);
			5110: out = 24'(32744);
			5111: out = 24'(32496);
			5112: out = 24'(32296);
			5113: out = 24'(32000);
			5114: out = 24'(31640);
			5115: out = 24'(31408);
			5116: out = 24'(31100);
			5117: out = 24'(30888);
			5118: out = 24'(30744);
			5119: out = 24'(30348);
			5120: out = 24'(30076);
			5121: out = 24'(29860);
			5122: out = 24'(29476);
			5123: out = 24'(29260);
			5124: out = 24'(29140);
			5125: out = 24'(28820);
			5126: out = 24'(28544);
			5127: out = 24'(28320);
			5128: out = 24'(27948);
			5129: out = 24'(27752);
			5130: out = 24'(27456);
			5131: out = 24'(27180);
			5132: out = 24'(26976);
			5133: out = 24'(26776);
			5134: out = 24'(26476);
			5135: out = 24'(26216);
			5136: out = 24'(25932);
			5137: out = 24'(25716);
			5138: out = 24'(25412);
			5139: out = 24'(25116);
			5140: out = 24'(24960);
			5141: out = 24'(24632);
			5142: out = 24'(24240);
			5143: out = 24'(24084);
			5144: out = 24'(23860);
			5145: out = 24'(23640);
			5146: out = 24'(23320);
			5147: out = 24'(23124);
			5148: out = 24'(22888);
			5149: out = 24'(22552);
			5150: out = 24'(22308);
			5151: out = 24'(22200);
			5152: out = 24'(21908);
			5153: out = 24'(21600);
			5154: out = 24'(21396);
			5155: out = 24'(21136);
			5156: out = 24'(20924);
			5157: out = 24'(20688);
			5158: out = 24'(20416);
			5159: out = 24'(20200);
			5160: out = 24'(19952);
			5161: out = 24'(19752);
			5162: out = 24'(19528);
			5163: out = 24'(19408);
			5164: out = 24'(19076);
			5165: out = 24'(18840);
			5166: out = 24'(18612);
			5167: out = 24'(18476);
			5168: out = 24'(18108);
			5169: out = 24'(17880);
			5170: out = 24'(17716);
			5171: out = 24'(17488);
			5172: out = 24'(17304);
			5173: out = 24'(17144);
			5174: out = 24'(16916);
			5175: out = 24'(16732);
			5176: out = 24'(16428);
			5177: out = 24'(16320);
			5178: out = 24'(16056);
			5179: out = 24'(15876);
			5180: out = 24'(15640);
			5181: out = 24'(15488);
			5182: out = 24'(15208);
			5183: out = 24'(15060);
			5184: out = 24'(14904);
			5185: out = 24'(14712);
			5186: out = 24'(14520);
			5187: out = 24'(14320);
			5188: out = 24'(14172);
			5189: out = 24'(14004);
			5190: out = 24'(13800);
			5191: out = 24'(13564);
			5192: out = 24'(13372);
			5193: out = 24'(13336);
			5194: out = 24'(13076);
			5195: out = 24'(12852);
			5196: out = 24'(12760);
			5197: out = 24'(12556);
			5198: out = 24'(12348);
			5199: out = 24'(12252);
			5200: out = 24'(12152);
			5201: out = 24'(11904);
			5202: out = 24'(11756);
			5203: out = 24'(11584);
			5204: out = 24'(11336);
			5205: out = 24'(11212);
			5206: out = 24'(11072);
			5207: out = 24'(10968);
			5208: out = 24'(10776);
			5209: out = 24'(10716);
			5210: out = 24'(10604);
			5211: out = 24'(10408);
			5212: out = 24'(10244);
			5213: out = 24'(10096);
			5214: out = 24'(10008);
			5215: out = 24'(9876);
			5216: out = 24'(9716);
			5217: out = 24'(9532);
			5218: out = 24'(9388);
			5219: out = 24'(9300);
			5220: out = 24'(9064);
			5221: out = 24'(8960);
			5222: out = 24'(8808);
			5223: out = 24'(8720);
			5224: out = 24'(8588);
			5225: out = 24'(8432);
			5226: out = 24'(8292);
			5227: out = 24'(8204);
			5228: out = 24'(8148);
			5229: out = 24'(7928);
			5230: out = 24'(7848);
			5231: out = 24'(7672);
			5232: out = 24'(7512);
			5233: out = 24'(7468);
			5234: out = 24'(7340);
			5235: out = 24'(7264);
			5236: out = 24'(7184);
			5237: out = 24'(6916);
			5238: out = 24'(6600);
			5239: out = 24'(6304);
			5240: out = 24'(5972);
			5241: out = 24'(5700);
			5242: out = 24'(5380);
			5243: out = 24'(5040);
			5244: out = 24'(4816);
			5245: out = 24'(4460);
			5246: out = 24'(4244);
			5247: out = 24'(3940);
			5248: out = 24'(3700);
			5249: out = 24'(3448);
			5250: out = 24'(3148);
			5251: out = 24'(2880);
			5252: out = 24'(2616);
			5253: out = 24'(2384);
			5254: out = 24'(2148);
			5255: out = 24'(1900);
			5256: out = 24'(1664);
			5257: out = 24'(1488);
			5258: out = 24'(1216);
			5259: out = 24'(956);
			5260: out = 24'(808);
			5261: out = 24'(604);
			5262: out = 24'(384);
			5263: out = 24'(124);
			5264: out = 24'(-128);
			5265: out = 24'(-364);
			5266: out = 24'(-592);
			5267: out = 24'(-844);
			5268: out = 24'(-1028);
			5269: out = 24'(-1208);
			5270: out = 24'(-1460);
			5271: out = 24'(-1644);
			5272: out = 24'(-1876);
			5273: out = 24'(-2084);
			5274: out = 24'(-2264);
			5275: out = 24'(-2504);
			5276: out = 24'(-2720);
			5277: out = 24'(-2940);
			5278: out = 24'(-3148);
			5279: out = 24'(-3332);
			5280: out = 24'(-3544);
			5281: out = 24'(-3708);
			5282: out = 24'(-3912);
			5283: out = 24'(-4132);
			5284: out = 24'(-4324);
			5285: out = 24'(-4500);
			5286: out = 24'(-4700);
			5287: out = 24'(-4884);
			5288: out = 24'(-5076);
			5289: out = 24'(-5176);
			5290: out = 24'(-5256);
			5291: out = 24'(-5576);
			5292: out = 24'(-5716);
			5293: out = 24'(-5908);
			5294: out = 24'(-6116);
			5295: out = 24'(-6328);
			5296: out = 24'(-6468);
			5297: out = 24'(-6656);
			5298: out = 24'(-6796);
			5299: out = 24'(-6912);
			5300: out = 24'(-7200);
			5301: out = 24'(-7268);
			5302: out = 24'(-7480);
			5303: out = 24'(-7656);
			5304: out = 24'(-7824);
			5305: out = 24'(-7964);
			5306: out = 24'(-8204);
			5307: out = 24'(-8420);
			5308: out = 24'(-8596);
			5309: out = 24'(-8692);
			5310: out = 24'(-8908);
			5311: out = 24'(-9044);
			5312: out = 24'(-9236);
			5313: out = 24'(-9488);
			5314: out = 24'(-9668);
			5315: out = 24'(-9836);
			5316: out = 24'(-9992);
			5317: out = 24'(-10188);
			5318: out = 24'(-10472);
			5319: out = 24'(-10608);
			5320: out = 24'(-10820);
			5321: out = 24'(-11008);
			5322: out = 24'(-11184);
			5323: out = 24'(-11364);
			5324: out = 24'(-11612);
			5325: out = 24'(-11848);
			5326: out = 24'(-12076);
			5327: out = 24'(-12236);
			5328: out = 24'(-12444);
			5329: out = 24'(-12708);
			5330: out = 24'(-12912);
			5331: out = 24'(-13124);
			5332: out = 24'(-13400);
			5333: out = 24'(-13528);
			5334: out = 24'(-13832);
			5335: out = 24'(-14036);
			5336: out = 24'(-14288);
			5337: out = 24'(-14524);
			5338: out = 24'(-14784);
			5339: out = 24'(-15024);
			5340: out = 24'(-15280);
			5341: out = 24'(-15580);
			5342: out = 24'(-15852);
			5343: out = 24'(-16096);
			5344: out = 24'(-16360);
			5345: out = 24'(-16636);
			5346: out = 24'(-16900);
			5347: out = 24'(-17164);
			5348: out = 24'(-17524);
			5349: out = 24'(-17780);
			5350: out = 24'(-18076);
			5351: out = 24'(-18312);
			5352: out = 24'(-18728);
			5353: out = 24'(-19080);
			5354: out = 24'(-19324);
			5355: out = 24'(-19656);
			5356: out = 24'(-20012);
			5357: out = 24'(-20320);
			5358: out = 24'(-20664);
			5359: out = 24'(-21040);
			5360: out = 24'(-21368);
			5361: out = 24'(-21744);
			5362: out = 24'(-22040);
			5363: out = 24'(-22412);
			5364: out = 24'(-22844);
			5365: out = 24'(-23212);
			5366: out = 24'(-23500);
			5367: out = 24'(-23920);
			5368: out = 24'(-24284);
			5369: out = 24'(-24580);
			5370: out = 24'(-24940);
			5371: out = 24'(-25312);
			5372: out = 24'(-25644);
			5373: out = 24'(-26028);
			5374: out = 24'(-26332);
			5375: out = 24'(-26752);
			5376: out = 24'(-27032);
			5377: out = 24'(-27444);
			5378: out = 24'(-27796);
			5379: out = 24'(-28128);
			5380: out = 24'(-28512);
			5381: out = 24'(-28812);
			5382: out = 24'(-29168);
			5383: out = 24'(-29512);
			5384: out = 24'(-29796);
			5385: out = 24'(-30108);
			5386: out = 24'(-30416);
			5387: out = 24'(-30692);
			5388: out = 24'(-30960);
			5389: out = 24'(-31308);
			5390: out = 24'(-31496);
			5391: out = 24'(-31836);
			5392: out = 24'(-32088);
			5393: out = 24'(-32372);
			5394: out = 24'(-32644);
			5395: out = 24'(-32904);
			5396: out = 24'(-33168);
			5397: out = 24'(-33340);
			5398: out = 24'(-33588);
			5399: out = 24'(-33844);
			5400: out = 24'(-34060);
			5401: out = 24'(-34324);
			5402: out = 24'(-34576);
			5403: out = 24'(-34728);
			5404: out = 24'(-34984);
			5405: out = 24'(-35172);
			5406: out = 24'(-35384);
			5407: out = 24'(-35532);
			5408: out = 24'(-35760);
			5409: out = 24'(-35944);
			5410: out = 24'(-36108);
			5411: out = 24'(-36340);
			5412: out = 24'(-36472);
			5413: out = 24'(-36672);
			5414: out = 24'(-36784);
			5415: out = 24'(-36960);
			5416: out = 24'(-37120);
			5417: out = 24'(-37288);
			5418: out = 24'(-37408);
			5419: out = 24'(-37572);
			5420: out = 24'(-37600);
			5421: out = 24'(-37812);
			5422: out = 24'(-37904);
			5423: out = 24'(-38072);
			5424: out = 24'(-38152);
			5425: out = 24'(-38236);
			5426: out = 24'(-38380);
			5427: out = 24'(-38476);
			5428: out = 24'(-38572);
			5429: out = 24'(-38724);
			5430: out = 24'(-38760);
			5431: out = 24'(-38828);
			5432: out = 24'(-38904);
			5433: out = 24'(-38972);
			5434: out = 24'(-39088);
			5435: out = 24'(-39116);
			5436: out = 24'(-39184);
			5437: out = 24'(-39264);
			5438: out = 24'(-39316);
			5439: out = 24'(-39328);
			5440: out = 24'(-39440);
			5441: out = 24'(-39460);
			5442: out = 24'(-39468);
			5443: out = 24'(-39580);
			5444: out = 24'(-39580);
			5445: out = 24'(-39588);
			5446: out = 24'(-39696);
			5447: out = 24'(-39680);
			5448: out = 24'(-39744);
			5449: out = 24'(-39736);
			5450: out = 24'(-39744);
			5451: out = 24'(-39840);
			5452: out = 24'(-39908);
			5453: out = 24'(-39828);
			5454: out = 24'(-39868);
			5455: out = 24'(-39860);
			5456: out = 24'(-39836);
			5457: out = 24'(-39884);
			5458: out = 24'(-39888);
			5459: out = 24'(-39868);
			5460: out = 24'(-39844);
			5461: out = 24'(-39888);
			5462: out = 24'(-39872);
			5463: out = 24'(-39820);
			5464: out = 24'(-39848);
			5465: out = 24'(-39832);
			5466: out = 24'(-39808);
			5467: out = 24'(-39896);
			5468: out = 24'(-39872);
			5469: out = 24'(-39792);
			5470: out = 24'(-39772);
			5471: out = 24'(-39740);
			5472: out = 24'(-39644);
			5473: out = 24'(-39640);
			5474: out = 24'(-39612);
			5475: out = 24'(-39592);
			5476: out = 24'(-39540);
			5477: out = 24'(-39492);
			5478: out = 24'(-39460);
			5479: out = 24'(-39424);
			5480: out = 24'(-39388);
			5481: out = 24'(-39344);
			5482: out = 24'(-39356);
			5483: out = 24'(-39256);
			5484: out = 24'(-39224);
			5485: out = 24'(-39164);
			5486: out = 24'(-39132);
			5487: out = 24'(-39056);
			5488: out = 24'(-38996);
			5489: out = 24'(-38948);
			5490: out = 24'(-38912);
			5491: out = 24'(-38804);
			5492: out = 24'(-38744);
			5493: out = 24'(-38732);
			5494: out = 24'(-38628);
			5495: out = 24'(-38584);
			5496: out = 24'(-38500);
			5497: out = 24'(-38428);
			5498: out = 24'(-38364);
			5499: out = 24'(-38268);
			5500: out = 24'(-38264);
			5501: out = 24'(-38112);
			5502: out = 24'(-38116);
			5503: out = 24'(-37976);
			5504: out = 24'(-37968);
			5505: out = 24'(-37892);
			5506: out = 24'(-37824);
			5507: out = 24'(-37704);
			5508: out = 24'(-37604);
			5509: out = 24'(-37556);
			5510: out = 24'(-37444);
			5511: out = 24'(-37404);
			5512: out = 24'(-37332);
			5513: out = 24'(-37216);
			5514: out = 24'(-37084);
			5515: out = 24'(-37068);
			5516: out = 24'(-36940);
			5517: out = 24'(-36932);
			5518: out = 24'(-36744);
			5519: out = 24'(-36652);
			5520: out = 24'(-36572);
			5521: out = 24'(-36456);
			5522: out = 24'(-36340);
			5523: out = 24'(-36216);
			5524: out = 24'(-36212);
			5525: out = 24'(-36044);
			5526: out = 24'(-35888);
			5527: out = 24'(-35832);
			5528: out = 24'(-35772);
			5529: out = 24'(-35520);
			5530: out = 24'(-35484);
			5531: out = 24'(-35268);
			5532: out = 24'(-35196);
			5533: out = 24'(-35084);
			5534: out = 24'(-34916);
			5535: out = 24'(-34832);
			5536: out = 24'(-34624);
			5537: out = 24'(-34488);
			5538: out = 24'(-34396);
			5539: out = 24'(-34228);
			5540: out = 24'(-34084);
			5541: out = 24'(-33880);
			5542: out = 24'(-33724);
			5543: out = 24'(-33552);
			5544: out = 24'(-33352);
			5545: out = 24'(-33212);
			5546: out = 24'(-33064);
			5547: out = 24'(-32860);
			5548: out = 24'(-32632);
			5549: out = 24'(-32480);
			5550: out = 24'(-32236);
			5551: out = 24'(-32052);
			5552: out = 24'(-31824);
			5553: out = 24'(-31584);
			5554: out = 24'(-31340);
			5555: out = 24'(-31128);
			5556: out = 24'(-30924);
			5557: out = 24'(-30636);
			5558: out = 24'(-30492);
			5559: out = 24'(-30220);
			5560: out = 24'(-29988);
			5561: out = 24'(-29712);
			5562: out = 24'(-29500);
			5563: out = 24'(-29260);
			5564: out = 24'(-28976);
			5565: out = 24'(-28696);
			5566: out = 24'(-28476);
			5567: out = 24'(-28140);
			5568: out = 24'(-27868);
			5569: out = 24'(-27608);
			5570: out = 24'(-27328);
			5571: out = 24'(-27036);
			5572: out = 24'(-26760);
			5573: out = 24'(-26460);
			5574: out = 24'(-26140);
			5575: out = 24'(-25932);
			5576: out = 24'(-25592);
			5577: out = 24'(-25328);
			5578: out = 24'(-25064);
			5579: out = 24'(-24756);
			5580: out = 24'(-24484);
			5581: out = 24'(-24172);
			5582: out = 24'(-23892);
			5583: out = 24'(-23608);
			5584: out = 24'(-23368);
			5585: out = 24'(-23080);
			5586: out = 24'(-22804);
			5587: out = 24'(-22488);
			5588: out = 24'(-22232);
			5589: out = 24'(-22004);
			5590: out = 24'(-21700);
			5591: out = 24'(-21452);
			5592: out = 24'(-21176);
			5593: out = 24'(-20924);
			5594: out = 24'(-20632);
			5595: out = 24'(-20360);
			5596: out = 24'(-20156);
			5597: out = 24'(-19796);
			5598: out = 24'(-19592);
			5599: out = 24'(-19328);
			5600: out = 24'(-19064);
			5601: out = 24'(-18840);
			5602: out = 24'(-18536);
			5603: out = 24'(-18264);
			5604: out = 24'(-18020);
			5605: out = 24'(-17788);
			5606: out = 24'(-17500);
			5607: out = 24'(-17288);
			5608: out = 24'(-17076);
			5609: out = 24'(-16828);
			5610: out = 24'(-16548);
			5611: out = 24'(-16308);
			5612: out = 24'(-16108);
			5613: out = 24'(-15880);
			5614: out = 24'(-15604);
			5615: out = 24'(-15404);
			5616: out = 24'(-15160);
			5617: out = 24'(-14984);
			5618: out = 24'(-14700);
			5619: out = 24'(-14504);
			5620: out = 24'(-14308);
			5621: out = 24'(-14016);
			5622: out = 24'(-13844);
			5623: out = 24'(-13668);
			5624: out = 24'(-13424);
			5625: out = 24'(-13228);
			5626: out = 24'(-13024);
			5627: out = 24'(-12812);
			5628: out = 24'(-12592);
			5629: out = 24'(-12396);
			5630: out = 24'(-12244);
			5631: out = 24'(-12040);
			5632: out = 24'(-11812);
			5633: out = 24'(-11620);
			5634: out = 24'(-11456);
			5635: out = 24'(-11252);
			5636: out = 24'(-11124);
			5637: out = 24'(-10912);
			5638: out = 24'(-10728);
			5639: out = 24'(-10524);
			5640: out = 24'(-10384);
			5641: out = 24'(-10216);
			5642: out = 24'(-10040);
			5643: out = 24'(-9868);
			5644: out = 24'(-9744);
			5645: out = 24'(-9536);
			5646: out = 24'(-9376);
			5647: out = 24'(-9236);
			5648: out = 24'(-9064);
			5649: out = 24'(-8912);
			5650: out = 24'(-8772);
			5651: out = 24'(-8620);
			5652: out = 24'(-8504);
			5653: out = 24'(-8324);
			5654: out = 24'(-8232);
			5655: out = 24'(-8028);
			5656: out = 24'(-7880);
			5657: out = 24'(-7744);
			5658: out = 24'(-7600);
			5659: out = 24'(-7460);
			5660: out = 24'(-7252);
			5661: out = 24'(-6980);
			5662: out = 24'(-6728);
			5663: out = 24'(-6452);
			5664: out = 24'(-6264);
			5665: out = 24'(-5980);
			5666: out = 24'(-5768);
			5667: out = 24'(-5544);
			5668: out = 24'(-5256);
			5669: out = 24'(-5076);
			5670: out = 24'(-4812);
			5671: out = 24'(-4608);
			5672: out = 24'(-4380);
			5673: out = 24'(-4152);
			5674: out = 24'(-3956);
			5675: out = 24'(-3708);
			5676: out = 24'(-3600);
			5677: out = 24'(-3316);
			5678: out = 24'(-3120);
			5679: out = 24'(-2968);
			5680: out = 24'(-2720);
			5681: out = 24'(-2572);
			5682: out = 24'(-2380);
			5683: out = 24'(-2204);
			5684: out = 24'(-1996);
			5685: out = 24'(-1792);
			5686: out = 24'(-1644);
			5687: out = 24'(-1520);
			5688: out = 24'(-1316);
			5689: out = 24'(-1116);
			5690: out = 24'(-968);
			5691: out = 24'(-780);
			5692: out = 24'(-608);
			5693: out = 24'(-432);
			5694: out = 24'(-320);
			5695: out = 24'(-176);
			5696: out = 24'(12);
			5697: out = 24'(156);
			5698: out = 24'(400);
			5699: out = 24'(448);
			5700: out = 24'(652);
			5701: out = 24'(820);
			5702: out = 24'(924);
			5703: out = 24'(1112);
			5704: out = 24'(1268);
			5705: out = 24'(1416);
			5706: out = 24'(1528);
			5707: out = 24'(1728);
			5708: out = 24'(1848);
			5709: out = 24'(2040);
			5710: out = 24'(2132);
			5711: out = 24'(2240);
			5712: out = 24'(2384);
			5713: out = 24'(2536);
			5714: out = 24'(2728);
			5715: out = 24'(2776);
			5716: out = 24'(3040);
			5717: out = 24'(3096);
			5718: out = 24'(3252);
			5719: out = 24'(3348);
			5720: out = 24'(3520);
			5721: out = 24'(3612);
			5722: out = 24'(3780);
			5723: out = 24'(3932);
			5724: out = 24'(4024);
			5725: out = 24'(4224);
			5726: out = 24'(4360);
			5727: out = 24'(4440);
			5728: out = 24'(4572);
			5729: out = 24'(4796);
			5730: out = 24'(4864);
			5731: out = 24'(4980);
			5732: out = 24'(5196);
			5733: out = 24'(5268);
			5734: out = 24'(5432);
			5735: out = 24'(5544);
			5736: out = 24'(5708);
			5737: out = 24'(5936);
			5738: out = 24'(6052);
			5739: out = 24'(6220);
			5740: out = 24'(6360);
			5741: out = 24'(6448);
			5742: out = 24'(6648);
			5743: out = 24'(6772);
			5744: out = 24'(6892);
			5745: out = 24'(7020);
			5746: out = 24'(7244);
			5747: out = 24'(7412);
			5748: out = 24'(7540);
			5749: out = 24'(7768);
			5750: out = 24'(7924);
			5751: out = 24'(8104);
			5752: out = 24'(8272);
			5753: out = 24'(8480);
			5754: out = 24'(8608);
			5755: out = 24'(8864);
			5756: out = 24'(9064);
			5757: out = 24'(9176);
			5758: out = 24'(9424);
			5759: out = 24'(9648);
			5760: out = 24'(9868);
			5761: out = 24'(10040);
			5762: out = 24'(10244);
			5763: out = 24'(10452);
			5764: out = 24'(10660);
			5765: out = 24'(10916);
			5766: out = 24'(11128);
			5767: out = 24'(11392);
			5768: out = 24'(11612);
			5769: out = 24'(11836);
			5770: out = 24'(12112);
			5771: out = 24'(12296);
			5772: out = 24'(12556);
			5773: out = 24'(12832);
			5774: out = 24'(13040);
			5775: out = 24'(13284);
			5776: out = 24'(13560);
			5777: out = 24'(13852);
			5778: out = 24'(14112);
			5779: out = 24'(14376);
			5780: out = 24'(14604);
			5781: out = 24'(14872);
			5782: out = 24'(15140);
			5783: out = 24'(15440);
			5784: out = 24'(15636);
			5785: out = 24'(15920);
			5786: out = 24'(16160);
			5787: out = 24'(16452);
			5788: out = 24'(16744);
			5789: out = 24'(16980);
			5790: out = 24'(17292);
			5791: out = 24'(17500);
			5792: out = 24'(17764);
			5793: out = 24'(18020);
			5794: out = 24'(18280);
			5795: out = 24'(18532);
			5796: out = 24'(18772);
			5797: out = 24'(18988);
			5798: out = 24'(19236);
			5799: out = 24'(19540);
			5800: out = 24'(19776);
			5801: out = 24'(19984);
			5802: out = 24'(20268);
			5803: out = 24'(20436);
			5804: out = 24'(20692);
			5805: out = 24'(20852);
			5806: out = 24'(21164);
			5807: out = 24'(21388);
			5808: out = 24'(21588);
			5809: out = 24'(21752);
			5810: out = 24'(22080);
			5811: out = 24'(22240);
			5812: out = 24'(22468);
			5813: out = 24'(22700);
			5814: out = 24'(22912);
			5815: out = 24'(23068);
			5816: out = 24'(23312);
			5817: out = 24'(23480);
			5818: out = 24'(23772);
			5819: out = 24'(23892);
			5820: out = 24'(24068);
			5821: out = 24'(24244);
			5822: out = 24'(24544);
			5823: out = 24'(24744);
			5824: out = 24'(24872);
			5825: out = 24'(25104);
			5826: out = 24'(25260);
			5827: out = 24'(25408);
			5828: out = 24'(25624);
			5829: out = 24'(25756);
			5830: out = 24'(25932);
			5831: out = 24'(26108);
			5832: out = 24'(26284);
			5833: out = 24'(26496);
			5834: out = 24'(26608);
			5835: out = 24'(26824);
			5836: out = 24'(26984);
			5837: out = 24'(27080);
			5838: out = 24'(27304);
			5839: out = 24'(27400);
			5840: out = 24'(27564);
			5841: out = 24'(27796);
			5842: out = 24'(27800);
			5843: out = 24'(28044);
			5844: out = 24'(28192);
			5845: out = 24'(28320);
			5846: out = 24'(28468);
			5847: out = 24'(28640);
			5848: out = 24'(28780);
			5849: out = 24'(28856);
			5850: out = 24'(29036);
			5851: out = 24'(29200);
			5852: out = 24'(29356);
			5853: out = 24'(29420);
			5854: out = 24'(29608);
			5855: out = 24'(29688);
			5856: out = 24'(29872);
			5857: out = 24'(29964);
			5858: out = 24'(30088);
			5859: out = 24'(30236);
			5860: out = 24'(30300);
			5861: out = 24'(30436);
			5862: out = 24'(30592);
			5863: out = 24'(30748);
			5864: out = 24'(30824);
			5865: out = 24'(30964);
			5866: out = 24'(31064);
			5867: out = 24'(31160);
			5868: out = 24'(31292);
			5869: out = 24'(31424);
			5870: out = 24'(31516);
			5871: out = 24'(31632);
			5872: out = 24'(31736);
			5873: out = 24'(31892);
			5874: out = 24'(31912);
			5875: out = 24'(32088);
			5876: out = 24'(32248);
			5877: out = 24'(32304);
			5878: out = 24'(32380);
			5879: out = 24'(32492);
			5880: out = 24'(32596);
			5881: out = 24'(32720);
			5882: out = 24'(32780);
			5883: out = 24'(32836);
			5884: out = 24'(32984);
			5885: out = 24'(33100);
			5886: out = 24'(33216);
			5887: out = 24'(33304);
			5888: out = 24'(33384);
			5889: out = 24'(33500);
			5890: out = 24'(33528);
			5891: out = 24'(33544);
			5892: out = 24'(33708);
			5893: out = 24'(33768);
			5894: out = 24'(33712);
			5895: out = 24'(33800);
			5896: out = 24'(33868);
			5897: out = 24'(33752);
			5898: out = 24'(33708);
			5899: out = 24'(33728);
			5900: out = 24'(33620);
			5901: out = 24'(33624);
			5902: out = 24'(33708);
			5903: out = 24'(33608);
			5904: out = 24'(33776);
			5905: out = 24'(33656);
			5906: out = 24'(33668);
			5907: out = 24'(33612);
			5908: out = 24'(33472);
			5909: out = 24'(33548);
			5910: out = 24'(33592);
			5911: out = 24'(33524);
			5912: out = 24'(33488);
			5913: out = 24'(33516);
			5914: out = 24'(33440);
			5915: out = 24'(33508);
			5916: out = 24'(33216);
			5917: out = 24'(33292);
			5918: out = 24'(33396);
			5919: out = 24'(33388);
			5920: out = 24'(33328);
			5921: out = 24'(33292);
			5922: out = 24'(33324);
			5923: out = 24'(33304);
			5924: out = 24'(33168);
			5925: out = 24'(33148);
			5926: out = 24'(33100);
			5927: out = 24'(33048);
			5928: out = 24'(33076);
			5929: out = 24'(33200);
			5930: out = 24'(33088);
			5931: out = 24'(33096);
			5932: out = 24'(33124);
			5933: out = 24'(33040);
			5934: out = 24'(33064);
			5935: out = 24'(33168);
			5936: out = 24'(32872);
			5937: out = 24'(32968);
			5938: out = 24'(32792);
			5939: out = 24'(32868);
			5940: out = 24'(32952);
			5941: out = 24'(32840);
			5942: out = 24'(32904);
			5943: out = 24'(33056);
			5944: out = 24'(32992);
			5945: out = 24'(32776);
			5946: out = 24'(32740);
			5947: out = 24'(32784);
			5948: out = 24'(32636);
			5949: out = 24'(32500);
			5950: out = 24'(32588);
			5951: out = 24'(32452);
			5952: out = 24'(32408);
			5953: out = 24'(32456);
			5954: out = 24'(32424);
			5955: out = 24'(32452);
			5956: out = 24'(32452);
			5957: out = 24'(32392);
			5958: out = 24'(32304);
			5959: out = 24'(32296);
			5960: out = 24'(32320);
			5961: out = 24'(32300);
			5962: out = 24'(32040);
			5963: out = 24'(32088);
			5964: out = 24'(31992);
			5965: out = 24'(32004);
			5966: out = 24'(31908);
			5967: out = 24'(31804);
			5968: out = 24'(31656);
			5969: out = 24'(31576);
			5970: out = 24'(31576);
			5971: out = 24'(31452);
			5972: out = 24'(31396);
			5973: out = 24'(31336);
			5974: out = 24'(31372);
			5975: out = 24'(31084);
			5976: out = 24'(30948);
			5977: out = 24'(30852);
			5978: out = 24'(30724);
			5979: out = 24'(30684);
			5980: out = 24'(30548);
			5981: out = 24'(30436);
			5982: out = 24'(30320);
			5983: out = 24'(30048);
			5984: out = 24'(30016);
			5985: out = 24'(29852);
			5986: out = 24'(29584);
			5987: out = 24'(29496);
			5988: out = 24'(29328);
			5989: out = 24'(29112);
			5990: out = 24'(29004);
			5991: out = 24'(28804);
			5992: out = 24'(28584);
			5993: out = 24'(28464);
			5994: out = 24'(28276);
			5995: out = 24'(28264);
			5996: out = 24'(27840);
			5997: out = 24'(27712);
			5998: out = 24'(27480);
			5999: out = 24'(27332);
			6000: out = 24'(27304);
			6001: out = 24'(27044);
			6002: out = 24'(26808);
			6003: out = 24'(26584);
			6004: out = 24'(26408);
			6005: out = 24'(26120);
			6006: out = 24'(25880);
			6007: out = 24'(25800);
			6008: out = 24'(25504);
			6009: out = 24'(25376);
			6010: out = 24'(25136);
			6011: out = 24'(24940);
			6012: out = 24'(24728);
			6013: out = 24'(24500);
			6014: out = 24'(24296);
			6015: out = 24'(23988);
			6016: out = 24'(23816);
			6017: out = 24'(23580);
			6018: out = 24'(23360);
			6019: out = 24'(23140);
			6020: out = 24'(22992);
			6021: out = 24'(22692);
			6022: out = 24'(22464);
			6023: out = 24'(22276);
			6024: out = 24'(22080);
			6025: out = 24'(21860);
			6026: out = 24'(21564);
			6027: out = 24'(21444);
			6028: out = 24'(21148);
			6029: out = 24'(20956);
			6030: out = 24'(20784);
			6031: out = 24'(20528);
			6032: out = 24'(20288);
			6033: out = 24'(20188);
			6034: out = 24'(19868);
			6035: out = 24'(19708);
			6036: out = 24'(19468);
			6037: out = 24'(19280);
			6038: out = 24'(19044);
			6039: out = 24'(18816);
			6040: out = 24'(18624);
			6041: out = 24'(18420);
			6042: out = 24'(18184);
			6043: out = 24'(18092);
			6044: out = 24'(17768);
			6045: out = 24'(17600);
			6046: out = 24'(17404);
			6047: out = 24'(17220);
			6048: out = 24'(17056);
			6049: out = 24'(16824);
			6050: out = 24'(16600);
			6051: out = 24'(16476);
			6052: out = 24'(16284);
			6053: out = 24'(16116);
			6054: out = 24'(15908);
			6055: out = 24'(15672);
			6056: out = 24'(15584);
			6057: out = 24'(15276);
			6058: out = 24'(15152);
			6059: out = 24'(14968);
			6060: out = 24'(14852);
			6061: out = 24'(14532);
			6062: out = 24'(14404);
			6063: out = 24'(14300);
			6064: out = 24'(14128);
			6065: out = 24'(13892);
			6066: out = 24'(13768);
			6067: out = 24'(13616);
			6068: out = 24'(13316);
			6069: out = 24'(13220);
			6070: out = 24'(13140);
			6071: out = 24'(12912);
			6072: out = 24'(12728);
			6073: out = 24'(12568);
			6074: out = 24'(12392);
			6075: out = 24'(12312);
			6076: out = 24'(12136);
			6077: out = 24'(11968);
			6078: out = 24'(11808);
			6079: out = 24'(11712);
			6080: out = 24'(11556);
			6081: out = 24'(11456);
			6082: out = 24'(11308);
			6083: out = 24'(11056);
			6084: out = 24'(10964);
			6085: out = 24'(10724);
			6086: out = 24'(10668);
			6087: out = 24'(10520);
			6088: out = 24'(10404);
			6089: out = 24'(10252);
			6090: out = 24'(10132);
			6091: out = 24'(9944);
			6092: out = 24'(9812);
			6093: out = 24'(9684);
			6094: out = 24'(9496);
			6095: out = 24'(9384);
			6096: out = 24'(9320);
			6097: out = 24'(9156);
			6098: out = 24'(9044);
			6099: out = 24'(8972);
			6100: out = 24'(8768);
			6101: out = 24'(8620);
			6102: out = 24'(8440);
			6103: out = 24'(8348);
			6104: out = 24'(8308);
			6105: out = 24'(8176);
			6106: out = 24'(8072);
			6107: out = 24'(8040);
			6108: out = 24'(7852);
			6109: out = 24'(7792);
			6110: out = 24'(7652);
			6111: out = 24'(7616);
			6112: out = 24'(7472);
			6113: out = 24'(7268);
			6114: out = 24'(7204);
			6115: out = 24'(7092);
			6116: out = 24'(7044);
			6117: out = 24'(6984);
			6118: out = 24'(6808);
			6119: out = 24'(6804);
			6120: out = 24'(6640);
			6121: out = 24'(6536);
			6122: out = 24'(6448);
			6123: out = 24'(6380);
			6124: out = 24'(6204);
			6125: out = 24'(6132);
			6126: out = 24'(5988);
			6127: out = 24'(5748);
			6128: out = 24'(5504);
			6129: out = 24'(5200);
			6130: out = 24'(4952);
			6131: out = 24'(4716);
			6132: out = 24'(4432);
			6133: out = 24'(4216);
			6134: out = 24'(4028);
			6135: out = 24'(3752);
			6136: out = 24'(3488);
			6137: out = 24'(3252);
			6138: out = 24'(3072);
			6139: out = 24'(2852);
			6140: out = 24'(2680);
			6141: out = 24'(2504);
			6142: out = 24'(2276);
			6143: out = 24'(2012);
			6144: out = 24'(1876);
			6145: out = 24'(1616);
			6146: out = 24'(1380);
			6147: out = 24'(1260);
			6148: out = 24'(972);
			6149: out = 24'(828);
			6150: out = 24'(576);
			6151: out = 24'(404);
			6152: out = 24'(204);
			6153: out = 24'(108);
			6154: out = 24'(-164);
			6155: out = 24'(-300);
			6156: out = 24'(-492);
			6157: out = 24'(-716);
			6158: out = 24'(-872);
			6159: out = 24'(-1148);
			6160: out = 24'(-1304);
			6161: out = 24'(-1432);
			6162: out = 24'(-1604);
			6163: out = 24'(-1784);
			6164: out = 24'(-1912);
			6165: out = 24'(-2152);
			6166: out = 24'(-2292);
			6167: out = 24'(-2516);
			6168: out = 24'(-2588);
			6169: out = 24'(-2800);
			6170: out = 24'(-2948);
			6171: out = 24'(-3152);
			6172: out = 24'(-3268);
			6173: out = 24'(-3416);
			6174: out = 24'(-3592);
			6175: out = 24'(-3668);
			6176: out = 24'(-3956);
			6177: out = 24'(-4012);
			6178: out = 24'(-4144);
			6179: out = 24'(-4432);
			6180: out = 24'(-4428);
			6181: out = 24'(-4652);
			6182: out = 24'(-4788);
			6183: out = 24'(-4972);
			6184: out = 24'(-5144);
			6185: out = 24'(-5212);
			6186: out = 24'(-5340);
			6187: out = 24'(-5472);
			6188: out = 24'(-5616);
			6189: out = 24'(-5776);
			6190: out = 24'(-5988);
			6191: out = 24'(-6044);
			6192: out = 24'(-6264);
			6193: out = 24'(-6464);
			6194: out = 24'(-6536);
			6195: out = 24'(-6704);
			6196: out = 24'(-6852);
			6197: out = 24'(-6944);
			6198: out = 24'(-7076);
			6199: out = 24'(-7296);
			6200: out = 24'(-7376);
			6201: out = 24'(-7560);
			6202: out = 24'(-7744);
			6203: out = 24'(-7868);
			6204: out = 24'(-7968);
			6205: out = 24'(-8200);
			6206: out = 24'(-8312);
			6207: out = 24'(-8500);
			6208: out = 24'(-8684);
			6209: out = 24'(-8796);
			6210: out = 24'(-9028);
			6211: out = 24'(-9156);
			6212: out = 24'(-9328);
			6213: out = 24'(-9508);
			6214: out = 24'(-9648);
			6215: out = 24'(-9848);
			6216: out = 24'(-10004);
			6217: out = 24'(-10216);
			6218: out = 24'(-10348);
			6219: out = 24'(-10584);
			6220: out = 24'(-10712);
			6221: out = 24'(-10896);
			6222: out = 24'(-11152);
			6223: out = 24'(-11364);
			6224: out = 24'(-11508);
			6225: out = 24'(-11684);
			6226: out = 24'(-11876);
			6227: out = 24'(-12060);
			6228: out = 24'(-12344);
			6229: out = 24'(-12504);
			6230: out = 24'(-12724);
			6231: out = 24'(-12952);
			6232: out = 24'(-13144);
			6233: out = 24'(-13344);
			6234: out = 24'(-13680);
			6235: out = 24'(-13864);
			6236: out = 24'(-14060);
			6237: out = 24'(-14384);
			6238: out = 24'(-14604);
			6239: out = 24'(-14792);
			6240: out = 24'(-15088);
			6241: out = 24'(-15348);
			6242: out = 24'(-15596);
			6243: out = 24'(-15840);
			6244: out = 24'(-16184);
			6245: out = 24'(-16432);
			6246: out = 24'(-16748);
			6247: out = 24'(-16988);
			6248: out = 24'(-17256);
			6249: out = 24'(-17516);
			6250: out = 24'(-17828);
			6251: out = 24'(-18084);
			6252: out = 24'(-18408);
			6253: out = 24'(-18720);
			6254: out = 24'(-19004);
			6255: out = 24'(-19252);
			6256: out = 24'(-19584);
			6257: out = 24'(-19876);
			6258: out = 24'(-20156);
			6259: out = 24'(-20472);
			6260: out = 24'(-20748);
			6261: out = 24'(-21044);
			6262: out = 24'(-21388);
			6263: out = 24'(-21640);
			6264: out = 24'(-21892);
			6265: out = 24'(-22236);
			6266: out = 24'(-22492);
			6267: out = 24'(-22756);
			6268: out = 24'(-23108);
			6269: out = 24'(-23368);
			6270: out = 24'(-23640);
			6271: out = 24'(-23864);
			6272: out = 24'(-24176);
			6273: out = 24'(-24420);
			6274: out = 24'(-24692);
			6275: out = 24'(-24956);
			6276: out = 24'(-25248);
			6277: out = 24'(-25452);
			6278: out = 24'(-25772);
			6279: out = 24'(-26008);
			6280: out = 24'(-26216);
			6281: out = 24'(-26492);
			6282: out = 24'(-26672);
			6283: out = 24'(-26944);
			6284: out = 24'(-27108);
			6285: out = 24'(-27316);
			6286: out = 24'(-27524);
			6287: out = 24'(-27764);
			6288: out = 24'(-27940);
			6289: out = 24'(-28128);
			6290: out = 24'(-28312);
			6291: out = 24'(-28512);
			6292: out = 24'(-28640);
			6293: out = 24'(-28864);
			6294: out = 24'(-29068);
			6295: out = 24'(-29128);
			6296: out = 24'(-29356);
			6297: out = 24'(-29532);
			6298: out = 24'(-29644);
			6299: out = 24'(-29852);
			6300: out = 24'(-29944);
			6301: out = 24'(-30124);
			6302: out = 24'(-30232);
			6303: out = 24'(-30404);
			6304: out = 24'(-30520);
			6305: out = 24'(-30636);
			6306: out = 24'(-30756);
			6307: out = 24'(-30912);
			6308: out = 24'(-30980);
			6309: out = 24'(-31112);
			6310: out = 24'(-31292);
			6311: out = 24'(-31352);
			6312: out = 24'(-31456);
			6313: out = 24'(-31496);
			6314: out = 24'(-31592);
			6315: out = 24'(-31704);
			6316: out = 24'(-31772);
			6317: out = 24'(-31884);
			6318: out = 24'(-31968);
			6319: out = 24'(-32004);
			6320: out = 24'(-32108);
			6321: out = 24'(-32168);
			6322: out = 24'(-32252);
			6323: out = 24'(-32304);
			6324: out = 24'(-32364);
			6325: out = 24'(-32368);
			6326: out = 24'(-32476);
			6327: out = 24'(-32512);
			6328: out = 24'(-32560);
			6329: out = 24'(-32604);
			6330: out = 24'(-32600);
			6331: out = 24'(-32712);
			6332: out = 24'(-32712);
			6333: out = 24'(-32744);
			6334: out = 24'(-32744);
			6335: out = 24'(-32824);
			6336: out = 24'(-32796);
			6337: out = 24'(-32836);
			6338: out = 24'(-32824);
			6339: out = 24'(-32904);
			6340: out = 24'(-32880);
			6341: out = 24'(-32900);
			6342: out = 24'(-32956);
			6343: out = 24'(-32964);
			6344: out = 24'(-32908);
			6345: out = 24'(-32976);
			6346: out = 24'(-32908);
			6347: out = 24'(-32968);
			6348: out = 24'(-32892);
			6349: out = 24'(-33012);
			6350: out = 24'(-32924);
			6351: out = 24'(-32900);
			6352: out = 24'(-32904);
			6353: out = 24'(-32912);
			6354: out = 24'(-32892);
			6355: out = 24'(-32932);
			6356: out = 24'(-32824);
			6357: out = 24'(-32844);
			6358: out = 24'(-32856);
			6359: out = 24'(-32792);
			6360: out = 24'(-32828);
			6361: out = 24'(-32756);
			6362: out = 24'(-32732);
			6363: out = 24'(-32720);
			6364: out = 24'(-32736);
			6365: out = 24'(-32732);
			6366: out = 24'(-32672);
			6367: out = 24'(-32596);
			6368: out = 24'(-32532);
			6369: out = 24'(-32548);
			6370: out = 24'(-32404);
			6371: out = 24'(-32412);
			6372: out = 24'(-32384);
			6373: out = 24'(-32296);
			6374: out = 24'(-32256);
			6375: out = 24'(-32264);
			6376: out = 24'(-32196);
			6377: out = 24'(-32152);
			6378: out = 24'(-32108);
			6379: out = 24'(-32036);
			6380: out = 24'(-32020);
			6381: out = 24'(-31880);
			6382: out = 24'(-31924);
			6383: out = 24'(-31876);
			6384: out = 24'(-31788);
			6385: out = 24'(-31772);
			6386: out = 24'(-31688);
			6387: out = 24'(-31628);
			6388: out = 24'(-31548);
			6389: out = 24'(-31540);
			6390: out = 24'(-31468);
			6391: out = 24'(-31420);
			6392: out = 24'(-31292);
			6393: out = 24'(-31288);
			6394: out = 24'(-31244);
			6395: out = 24'(-31180);
			6396: out = 24'(-31032);
			6397: out = 24'(-31012);
			6398: out = 24'(-30964);
			6399: out = 24'(-30816);
			6400: out = 24'(-30808);
			6401: out = 24'(-30732);
			6402: out = 24'(-30648);
			6403: out = 24'(-30584);
			6404: out = 24'(-30496);
			6405: out = 24'(-30372);
			6406: out = 24'(-30360);
			6407: out = 24'(-30272);
			6408: out = 24'(-30192);
			6409: out = 24'(-30092);
			6410: out = 24'(-29996);
			6411: out = 24'(-29884);
			6412: out = 24'(-29828);
			6413: out = 24'(-29732);
			6414: out = 24'(-29684);
			6415: out = 24'(-29552);
			6416: out = 24'(-29404);
			6417: out = 24'(-29368);
			6418: out = 24'(-29272);
			6419: out = 24'(-29160);
			6420: out = 24'(-29024);
			6421: out = 24'(-28948);
			6422: out = 24'(-28852);
			6423: out = 24'(-28744);
			6424: out = 24'(-28600);
			6425: out = 24'(-28508);
			6426: out = 24'(-28364);
			6427: out = 24'(-28224);
			6428: out = 24'(-28156);
			6429: out = 24'(-28000);
			6430: out = 24'(-27868);
			6431: out = 24'(-27788);
			6432: out = 24'(-27580);
			6433: out = 24'(-27476);
			6434: out = 24'(-27324);
			6435: out = 24'(-27164);
			6436: out = 24'(-27040);
			6437: out = 24'(-26868);
			6438: out = 24'(-26700);
			6439: out = 24'(-26576);
			6440: out = 24'(-26312);
			6441: out = 24'(-26232);
			6442: out = 24'(-26048);
			6443: out = 24'(-25808);
			6444: out = 24'(-25664);
			6445: out = 24'(-25476);
			6446: out = 24'(-25240);
			6447: out = 24'(-25104);
			6448: out = 24'(-24816);
			6449: out = 24'(-24616);
			6450: out = 24'(-24392);
			6451: out = 24'(-24244);
			6452: out = 24'(-24048);
			6453: out = 24'(-23800);
			6454: out = 24'(-23596);
			6455: out = 24'(-23396);
			6456: out = 24'(-23208);
			6457: out = 24'(-22944);
			6458: out = 24'(-22732);
			6459: out = 24'(-22476);
			6460: out = 24'(-22312);
			6461: out = 24'(-22032);
			6462: out = 24'(-21800);
			6463: out = 24'(-21568);
			6464: out = 24'(-21368);
			6465: out = 24'(-21140);
			6466: out = 24'(-20944);
			6467: out = 24'(-20656);
			6468: out = 24'(-20396);
			6469: out = 24'(-20204);
			6470: out = 24'(-20000);
			6471: out = 24'(-19760);
			6472: out = 24'(-19472);
			6473: out = 24'(-19288);
			6474: out = 24'(-19020);
			6475: out = 24'(-18828);
			6476: out = 24'(-18560);
			6477: out = 24'(-18352);
			6478: out = 24'(-18116);
			6479: out = 24'(-17916);
			6480: out = 24'(-17664);
			6481: out = 24'(-17452);
			6482: out = 24'(-17252);
			6483: out = 24'(-17008);
			6484: out = 24'(-16776);
			6485: out = 24'(-16528);
			6486: out = 24'(-16324);
			6487: out = 24'(-16060);
			6488: out = 24'(-15932);
			6489: out = 24'(-15648);
			6490: out = 24'(-15484);
			6491: out = 24'(-15200);
			6492: out = 24'(-15024);
			6493: out = 24'(-14808);
			6494: out = 24'(-14616);
			6495: out = 24'(-14416);
			6496: out = 24'(-14184);
			6497: out = 24'(-13984);
			6498: out = 24'(-13824);
			6499: out = 24'(-13616);
			6500: out = 24'(-13380);
			6501: out = 24'(-13220);
			6502: out = 24'(-13000);
			6503: out = 24'(-12852);
			6504: out = 24'(-12676);
			6505: out = 24'(-12464);
			6506: out = 24'(-12316);
			6507: out = 24'(-12112);
			6508: out = 24'(-11944);
			6509: out = 24'(-11748);
			6510: out = 24'(-11552);
			6511: out = 24'(-11424);
			6512: out = 24'(-11220);
			6513: out = 24'(-11056);
			6514: out = 24'(-10880);
			6515: out = 24'(-10732);
			6516: out = 24'(-10540);
			6517: out = 24'(-10396);
			6518: out = 24'(-10200);
			6519: out = 24'(-10088);
			6520: out = 24'(-9836);
			6521: out = 24'(-9752);
			6522: out = 24'(-9572);
			6523: out = 24'(-9412);
			6524: out = 24'(-9268);
			6525: out = 24'(-9080);
			6526: out = 24'(-8940);
			6527: out = 24'(-8820);
			6528: out = 24'(-8700);
			6529: out = 24'(-8532);
			6530: out = 24'(-8432);
			6531: out = 24'(-8260);
			6532: out = 24'(-8064);
			6533: out = 24'(-7972);
			6534: out = 24'(-7796);
			6535: out = 24'(-7724);
			6536: out = 24'(-7564);
			6537: out = 24'(-7444);
			6538: out = 24'(-7312);
			6539: out = 24'(-7244);
			6540: out = 24'(-7112);
			6541: out = 24'(-6948);
			6542: out = 24'(-6844);
			6543: out = 24'(-6692);
			6544: out = 24'(-6608);
			6545: out = 24'(-6496);
			6546: out = 24'(-6400);
			6547: out = 24'(-6216);
			6548: out = 24'(-6140);
			6549: out = 24'(-6092);
			6550: out = 24'(-5892);
			6551: out = 24'(-5684);
			6552: out = 24'(-5500);
			6553: out = 24'(-5248);
			6554: out = 24'(-5056);
			6555: out = 24'(-4824);
			6556: out = 24'(-4664);
			6557: out = 24'(-4416);
			6558: out = 24'(-4284);
			6559: out = 24'(-4092);
			6560: out = 24'(-3912);
			6561: out = 24'(-3712);
			6562: out = 24'(-3536);
			6563: out = 24'(-3428);
			6564: out = 24'(-3180);
			6565: out = 24'(-3068);
			6566: out = 24'(-2844);
			6567: out = 24'(-2704);
			6568: out = 24'(-2544);
			6569: out = 24'(-2420);
			6570: out = 24'(-2248);
			6571: out = 24'(-2112);
			6572: out = 24'(-1932);
			6573: out = 24'(-1784);
			6574: out = 24'(-1624);
			6575: out = 24'(-1528);
			6576: out = 24'(-1384);
			6577: out = 24'(-1212);
			6578: out = 24'(-1084);
			6579: out = 24'(-960);
			6580: out = 24'(-812);
			6581: out = 24'(-696);
			6582: out = 24'(-504);
			6583: out = 24'(-428);
			6584: out = 24'(-224);
			6585: out = 24'(-172);
			6586: out = 24'(-4);
			6587: out = 24'(76);
			6588: out = 24'(240);
			6589: out = 24'(384);
			6590: out = 24'(504);
			6591: out = 24'(588);
			6592: out = 24'(732);
			6593: out = 24'(872);
			6594: out = 24'(984);
			6595: out = 24'(1108);
			6596: out = 24'(1248);
			6597: out = 24'(1368);
			6598: out = 24'(1456);
			6599: out = 24'(1580);
			6600: out = 24'(1692);
			6601: out = 24'(1824);
			6602: out = 24'(1956);
			6603: out = 24'(2004);
			6604: out = 24'(2180);
			6605: out = 24'(2248);
			6606: out = 24'(2376);
			6607: out = 24'(2540);
			6608: out = 24'(2588);
			6609: out = 24'(2688);
			6610: out = 24'(2836);
			6611: out = 24'(2944);
			6612: out = 24'(3036);
			6613: out = 24'(3156);
			6614: out = 24'(3236);
			6615: out = 24'(3364);
			6616: out = 24'(3424);
			6617: out = 24'(3580);
			6618: out = 24'(3688);
			6619: out = 24'(3828);
			6620: out = 24'(3900);
			6621: out = 24'(4064);
			6622: out = 24'(4148);
			6623: out = 24'(4268);
			6624: out = 24'(4392);
			6625: out = 24'(4516);
			6626: out = 24'(4572);
			6627: out = 24'(4716);
			6628: out = 24'(4876);
			6629: out = 24'(4964);
			6630: out = 24'(5160);
			6631: out = 24'(5232);
			6632: out = 24'(5376);
			6633: out = 24'(5460);
			6634: out = 24'(5668);
			6635: out = 24'(5776);
			6636: out = 24'(5920);
			6637: out = 24'(6060);
			6638: out = 24'(6156);
			6639: out = 24'(6308);
			6640: out = 24'(6432);
			6641: out = 24'(6560);
			6642: out = 24'(6656);
			6643: out = 24'(6836);
			6644: out = 24'(7012);
			6645: out = 24'(7124);
			6646: out = 24'(7296);
			6647: out = 24'(7488);
			6648: out = 24'(7632);
			6649: out = 24'(7780);
			6650: out = 24'(7968);
			6651: out = 24'(8120);
			6652: out = 24'(8252);
			6653: out = 24'(8516);
			6654: out = 24'(8652);
			6655: out = 24'(8816);
			6656: out = 24'(9012);
			6657: out = 24'(9216);
			6658: out = 24'(9444);
			6659: out = 24'(9592);
			6660: out = 24'(9760);
			6661: out = 24'(10012);
			6662: out = 24'(10188);
			6663: out = 24'(10388);
			6664: out = 24'(10632);
			6665: out = 24'(10784);
			6666: out = 24'(11040);
			6667: out = 24'(11192);
			6668: out = 24'(11420);
			6669: out = 24'(11632);
			6670: out = 24'(11840);
			6671: out = 24'(12072);
			6672: out = 24'(12300);
			6673: out = 24'(12476);
			6674: out = 24'(12720);
			6675: out = 24'(12904);
			6676: out = 24'(13184);
			6677: out = 24'(13304);
			6678: out = 24'(13568);
			6679: out = 24'(13780);
			6680: out = 24'(13996);
			6681: out = 24'(14204);
			6682: out = 24'(14408);
			6683: out = 24'(14652);
			6684: out = 24'(14804);
			6685: out = 24'(15012);
			6686: out = 24'(15244);
			6687: out = 24'(15468);
			6688: out = 24'(15656);
			6689: out = 24'(15840);
			6690: out = 24'(16040);
			6691: out = 24'(16224);
			6692: out = 24'(16508);
			6693: out = 24'(16608);
			6694: out = 24'(16812);
			6695: out = 24'(17076);
			6696: out = 24'(17168);
			6697: out = 24'(17388);
			6698: out = 24'(17600);
			6699: out = 24'(17764);
			6700: out = 24'(17956);
			6701: out = 24'(18096);
			6702: out = 24'(18296);
			6703: out = 24'(18464);
			6704: out = 24'(18676);
			6705: out = 24'(18832);
			6706: out = 24'(19040);
			6707: out = 24'(19204);
			6708: out = 24'(19380);
			6709: out = 24'(19536);
			6710: out = 24'(19700);
			6711: out = 24'(19916);
			6712: out = 24'(20000);
			6713: out = 24'(20184);
			6714: out = 24'(20328);
			6715: out = 24'(20504);
			6716: out = 24'(20696);
			6717: out = 24'(20752);
			6718: out = 24'(20996);
			6719: out = 24'(21072);
			6720: out = 24'(21248);
			6721: out = 24'(21408);
			6722: out = 24'(21480);
			6723: out = 24'(21668);
			6724: out = 24'(21768);
			6725: out = 24'(21896);
			6726: out = 24'(22064);
			6727: out = 24'(22204);
			6728: out = 24'(22260);
			6729: out = 24'(22456);
			6730: out = 24'(22532);
			6731: out = 24'(22652);
			6732: out = 24'(22856);
			6733: out = 24'(22916);
			6734: out = 24'(23044);
			6735: out = 24'(23212);
			6736: out = 24'(23364);
			6737: out = 24'(23420);
			6738: out = 24'(23560);
			6739: out = 24'(23700);
			6740: out = 24'(23768);
			6741: out = 24'(23968);
			6742: out = 24'(24008);
			6743: out = 24'(24104);
			6744: out = 24'(24268);
			6745: out = 24'(24292);
			6746: out = 24'(24472);
			6747: out = 24'(24552);
			6748: out = 24'(24676);
			6749: out = 24'(24788);
			6750: out = 24'(24864);
			6751: out = 24'(24980);
			6752: out = 24'(25080);
			6753: out = 24'(25220);
			6754: out = 24'(25272);
			6755: out = 24'(25328);
			6756: out = 24'(25516);
			6757: out = 24'(25540);
			6758: out = 24'(25680);
			6759: out = 24'(25772);
			6760: out = 24'(25872);
			6761: out = 24'(25940);
			6762: out = 24'(26036);
			6763: out = 24'(26140);
			6764: out = 24'(26228);
			6765: out = 24'(26344);
			6766: out = 24'(26360);
			6767: out = 24'(26452);
			6768: out = 24'(26628);
			6769: out = 24'(26628);
			6770: out = 24'(26760);
			6771: out = 24'(26848);
			6772: out = 24'(26956);
			6773: out = 24'(27000);
			6774: out = 24'(27092);
			6775: out = 24'(27204);
			6776: out = 24'(27240);
			6777: out = 24'(27436);
			6778: out = 24'(27340);
			6779: out = 24'(27512);
			6780: out = 24'(27584);
			6781: out = 24'(27588);
			6782: out = 24'(27704);
			6783: out = 24'(27776);
			6784: out = 24'(27836);
			6785: out = 24'(27836);
			6786: out = 24'(27828);
			6787: out = 24'(27840);
			6788: out = 24'(27880);
			6789: out = 24'(27928);
			6790: out = 24'(27816);
			6791: out = 24'(27812);
			6792: out = 24'(27760);
			6793: out = 24'(27728);
			6794: out = 24'(27700);
			6795: out = 24'(27700);
			6796: out = 24'(27716);
			6797: out = 24'(27632);
			6798: out = 24'(27668);
			6799: out = 24'(27540);
			6800: out = 24'(27556);
			6801: out = 24'(27512);
			6802: out = 24'(27376);
			6803: out = 24'(27484);
			6804: out = 24'(27444);
			6805: out = 24'(27440);
			6806: out = 24'(27492);
			6807: out = 24'(27536);
			6808: out = 24'(27524);
			6809: out = 24'(27596);
			6810: out = 24'(27496);
			6811: out = 24'(27564);
			6812: out = 24'(27480);
			6813: out = 24'(27528);
			6814: out = 24'(27492);
			6815: out = 24'(27364);
			6816: out = 24'(27344);
			6817: out = 24'(27428);
			6818: out = 24'(27252);
			6819: out = 24'(27260);
			6820: out = 24'(27332);
			6821: out = 24'(27300);
			6822: out = 24'(27180);
			6823: out = 24'(27188);
			6824: out = 24'(27132);
			6825: out = 24'(27096);
			6826: out = 24'(27076);
			6827: out = 24'(27228);
			6828: out = 24'(27176);
			6829: out = 24'(27208);
			6830: out = 24'(27036);
			6831: out = 24'(27112);
			6832: out = 24'(27132);
			6833: out = 24'(27088);
			6834: out = 24'(27116);
			6835: out = 24'(27180);
			6836: out = 24'(27124);
			6837: out = 24'(27048);
			6838: out = 24'(26996);
			6839: out = 24'(26832);
			6840: out = 24'(26964);
			6841: out = 24'(26852);
			6842: out = 24'(26888);
			6843: out = 24'(26852);
			6844: out = 24'(26820);
			6845: out = 24'(26824);
			6846: out = 24'(26772);
			6847: out = 24'(26804);
			6848: out = 24'(26748);
			6849: out = 24'(26804);
			6850: out = 24'(26772);
			6851: out = 24'(26684);
			6852: out = 24'(26464);
			6853: out = 24'(26376);
			6854: out = 24'(26380);
			6855: out = 24'(26336);
			6856: out = 24'(26228);
			6857: out = 24'(26296);
			6858: out = 24'(26224);
			6859: out = 24'(26144);
			6860: out = 24'(26020);
			6861: out = 24'(26044);
			6862: out = 24'(26028);
			6863: out = 24'(25780);
			6864: out = 24'(25780);
			6865: out = 24'(25760);
			6866: out = 24'(25640);
			6867: out = 24'(25556);
			6868: out = 24'(25376);
			6869: out = 24'(25296);
			6870: out = 24'(25292);
			6871: out = 24'(25072);
			6872: out = 24'(25016);
			6873: out = 24'(24884);
			6874: out = 24'(24748);
			6875: out = 24'(24692);
			6876: out = 24'(24664);
			6877: out = 24'(24356);
			6878: out = 24'(24296);
			6879: out = 24'(24208);
			6880: out = 24'(24048);
			6881: out = 24'(23924);
			6882: out = 24'(23768);
			6883: out = 24'(23608);
			6884: out = 24'(23444);
			6885: out = 24'(23392);
			6886: out = 24'(23224);
			6887: out = 24'(22996);
			6888: out = 24'(22840);
			6889: out = 24'(22604);
			6890: out = 24'(22464);
			6891: out = 24'(22408);
			6892: out = 24'(22192);
			6893: out = 24'(22108);
			6894: out = 24'(21888);
			6895: out = 24'(21700);
			6896: out = 24'(21556);
			6897: out = 24'(21304);
			6898: out = 24'(21236);
			6899: out = 24'(21012);
			6900: out = 24'(20856);
			6901: out = 24'(20648);
			6902: out = 24'(20444);
			6903: out = 24'(20356);
			6904: out = 24'(20100);
			6905: out = 24'(20040);
			6906: out = 24'(19808);
			6907: out = 24'(19620);
			6908: out = 24'(19432);
			6909: out = 24'(19224);
			6910: out = 24'(19060);
			6911: out = 24'(18936);
			6912: out = 24'(18732);
			6913: out = 24'(18452);
			6914: out = 24'(18368);
			6915: out = 24'(18092);
			6916: out = 24'(17964);
			6917: out = 24'(17788);
			6918: out = 24'(17596);
			6919: out = 24'(17444);
			6920: out = 24'(17328);
			6921: out = 24'(17056);
			6922: out = 24'(16900);
			6923: out = 24'(16732);
			6924: out = 24'(16636);
			6925: out = 24'(16352);
			6926: out = 24'(16208);
			6927: out = 24'(16040);
			6928: out = 24'(15832);
			6929: out = 24'(15716);
			6930: out = 24'(15460);
			6931: out = 24'(15392);
			6932: out = 24'(15180);
			6933: out = 24'(15056);
			6934: out = 24'(14864);
			6935: out = 24'(14660);
			6936: out = 24'(14532);
			6937: out = 24'(14332);
			6938: out = 24'(14116);
			6939: out = 24'(14080);
			6940: out = 24'(13864);
			6941: out = 24'(13640);
			6942: out = 24'(13508);
			6943: out = 24'(13448);
			6944: out = 24'(13240);
			6945: out = 24'(13148);
			6946: out = 24'(12944);
			6947: out = 24'(12728);
			6948: out = 24'(12640);
			6949: out = 24'(12444);
			6950: out = 24'(12404);
			6951: out = 24'(12220);
			6952: out = 24'(12080);
			6953: out = 24'(11912);
			6954: out = 24'(11804);
			6955: out = 24'(11612);
			6956: out = 24'(11524);
			6957: out = 24'(11308);
			6958: out = 24'(11212);
			6959: out = 24'(11096);
			6960: out = 24'(10948);
			6961: out = 24'(10812);
			6962: out = 24'(10728);
			6963: out = 24'(10504);
			6964: out = 24'(10428);
			6965: out = 24'(10272);
			6966: out = 24'(10112);
			6967: out = 24'(10048);
			6968: out = 24'(9964);
			6969: out = 24'(9836);
			6970: out = 24'(9636);
			6971: out = 24'(9548);
			6972: out = 24'(9444);
			6973: out = 24'(9260);
			6974: out = 24'(9160);
			6975: out = 24'(9100);
			6976: out = 24'(8952);
			6977: out = 24'(8856);
			6978: out = 24'(8732);
			6979: out = 24'(8584);
			6980: out = 24'(8492);
			6981: out = 24'(8388);
			6982: out = 24'(8292);
			6983: out = 24'(8132);
			6984: out = 24'(8080);
			6985: out = 24'(7940);
			6986: out = 24'(7836);
			6987: out = 24'(7716);
			6988: out = 24'(7560);
			6989: out = 24'(7504);
			6990: out = 24'(7436);
			6991: out = 24'(7268);
			6992: out = 24'(7232);
			6993: out = 24'(7092);
			6994: out = 24'(7032);
			6995: out = 24'(6852);
			6996: out = 24'(6800);
			6997: out = 24'(6764);
			6998: out = 24'(6628);
			6999: out = 24'(6476);
			7000: out = 24'(6428);
			7001: out = 24'(6328);
			7002: out = 24'(6276);
			7003: out = 24'(6136);
			7004: out = 24'(6040);
			7005: out = 24'(6024);
			7006: out = 24'(5836);
			7007: out = 24'(5736);
			7008: out = 24'(5700);
			7009: out = 24'(5596);
			7010: out = 24'(5552);
			7011: out = 24'(5480);
			7012: out = 24'(5436);
			7013: out = 24'(5352);
			7014: out = 24'(5276);
			7015: out = 24'(5128);
			7016: out = 24'(5032);
			7017: out = 24'(4948);
			7018: out = 24'(4704);
			7019: out = 24'(4512);
			7020: out = 24'(4348);
			7021: out = 24'(4124);
			7022: out = 24'(3864);
			7023: out = 24'(3696);
			7024: out = 24'(3468);
			7025: out = 24'(3252);
			7026: out = 24'(3128);
			7027: out = 24'(2864);
			7028: out = 24'(2664);
			7029: out = 24'(2476);
			7030: out = 24'(2292);
			7031: out = 24'(2148);
			7032: out = 24'(1944);
			7033: out = 24'(1768);
			7034: out = 24'(1576);
			7035: out = 24'(1468);
			7036: out = 24'(1240);
			7037: out = 24'(1080);
			7038: out = 24'(964);
			7039: out = 24'(696);
			7040: out = 24'(540);
			7041: out = 24'(428);
			7042: out = 24'(212);
			7043: out = 24'(104);
			7044: out = 24'(-40);
			7045: out = 24'(-216);
			7046: out = 24'(-368);
			7047: out = 24'(-560);
			7048: out = 24'(-692);
			7049: out = 24'(-808);
			7050: out = 24'(-968);
			7051: out = 24'(-1120);
			7052: out = 24'(-1300);
			7053: out = 24'(-1400);
			7054: out = 24'(-1556);
			7055: out = 24'(-1640);
			7056: out = 24'(-1840);
			7057: out = 24'(-1884);
			7058: out = 24'(-2152);
			7059: out = 24'(-2164);
			7060: out = 24'(-2304);
			7061: out = 24'(-2500);
			7062: out = 24'(-2640);
			7063: out = 24'(-2812);
			7064: out = 24'(-2900);
			7065: out = 24'(-3064);
			7066: out = 24'(-3156);
			7067: out = 24'(-3316);
			7068: out = 24'(-3396);
			7069: out = 24'(-3544);
			7070: out = 24'(-3672);
			7071: out = 24'(-3780);
			7072: out = 24'(-3868);
			7073: out = 24'(-4028);
			7074: out = 24'(-4200);
			7075: out = 24'(-4320);
			7076: out = 24'(-4404);
			7077: out = 24'(-4568);
			7078: out = 24'(-4632);
			7079: out = 24'(-4736);
			7080: out = 24'(-4888);
			7081: out = 24'(-5028);
			7082: out = 24'(-5104);
			7083: out = 24'(-5268);
			7084: out = 24'(-5364);
			7085: out = 24'(-5492);
			7086: out = 24'(-5664);
			7087: out = 24'(-5732);
			7088: out = 24'(-5876);
			7089: out = 24'(-5992);
			7090: out = 24'(-6084);
			7091: out = 24'(-6220);
			7092: out = 24'(-6264);
			7093: out = 24'(-6416);
			7094: out = 24'(-6592);
			7095: out = 24'(-6692);
			7096: out = 24'(-6864);
			7097: out = 24'(-7000);
			7098: out = 24'(-7160);
			7099: out = 24'(-7300);
			7100: out = 24'(-7440);
			7101: out = 24'(-7552);
			7102: out = 24'(-7672);
			7103: out = 24'(-7840);
			7104: out = 24'(-7960);
			7105: out = 24'(-8068);
			7106: out = 24'(-8256);
			7107: out = 24'(-8360);
			7108: out = 24'(-8532);
			7109: out = 24'(-8636);
			7110: out = 24'(-8864);
			7111: out = 24'(-8996);
			7112: out = 24'(-9128);
			7113: out = 24'(-9288);
			7114: out = 24'(-9500);
			7115: out = 24'(-9588);
			7116: out = 24'(-9776);
			7117: out = 24'(-9912);
			7118: out = 24'(-10084);
			7119: out = 24'(-10288);
			7120: out = 24'(-10456);
			7121: out = 24'(-10596);
			7122: out = 24'(-10784);
			7123: out = 24'(-10988);
			7124: out = 24'(-11132);
			7125: out = 24'(-11308);
			7126: out = 24'(-11556);
			7127: out = 24'(-11692);
			7128: out = 24'(-11948);
			7129: out = 24'(-12040);
			7130: out = 24'(-12348);
			7131: out = 24'(-12484);
			7132: out = 24'(-12720);
			7133: out = 24'(-12988);
			7134: out = 24'(-13152);
			7135: out = 24'(-13428);
			7136: out = 24'(-13660);
			7137: out = 24'(-13860);
			7138: out = 24'(-14076);
			7139: out = 24'(-14356);
			7140: out = 24'(-14560);
			7141: out = 24'(-14828);
			7142: out = 24'(-15076);
			7143: out = 24'(-15260);
			7144: out = 24'(-15520);
			7145: out = 24'(-15728);
			7146: out = 24'(-16064);
			7147: out = 24'(-16276);
			7148: out = 24'(-16568);
			7149: out = 24'(-16744);
			7150: out = 24'(-16988);
			7151: out = 24'(-17252);
			7152: out = 24'(-17496);
			7153: out = 24'(-17740);
			7154: out = 24'(-17928);
			7155: out = 24'(-18260);
			7156: out = 24'(-18416);
			7157: out = 24'(-18680);
			7158: out = 24'(-18900);
			7159: out = 24'(-19164);
			7160: out = 24'(-19344);
			7161: out = 24'(-19528);
			7162: out = 24'(-19824);
			7163: out = 24'(-20012);
			7164: out = 24'(-20220);
			7165: out = 24'(-20428);
			7166: out = 24'(-20676);
			7167: out = 24'(-20864);
			7168: out = 24'(-21044);
			7169: out = 24'(-21260);
			7170: out = 24'(-21508);
			7171: out = 24'(-21644);
			7172: out = 24'(-21832);
			7173: out = 24'(-22060);
			7174: out = 24'(-22176);
			7175: out = 24'(-22468);
			7176: out = 24'(-22556);
			7177: out = 24'(-22724);
			7178: out = 24'(-22964);
			7179: out = 24'(-23000);
			7180: out = 24'(-23256);
			7181: out = 24'(-23408);
			7182: out = 24'(-23576);
			7183: out = 24'(-23680);
			7184: out = 24'(-23896);
			7185: out = 24'(-23980);
			7186: out = 24'(-24176);
			7187: out = 24'(-24312);
			7188: out = 24'(-24404);
			7189: out = 24'(-24600);
			7190: out = 24'(-24684);
			7191: out = 24'(-24736);
			7192: out = 24'(-24920);
			7193: out = 24'(-25012);
			7194: out = 24'(-25148);
			7195: out = 24'(-25224);
			7196: out = 24'(-25324);
			7197: out = 24'(-25440);
			7198: out = 24'(-25520);
			7199: out = 24'(-25664);
			7200: out = 24'(-25708);
			7201: out = 24'(-25780);
			7202: out = 24'(-25880);
			7203: out = 24'(-25884);
			7204: out = 24'(-26052);
			7205: out = 24'(-26068);
			7206: out = 24'(-26152);
			7207: out = 24'(-26208);
			7208: out = 24'(-26276);
			7209: out = 24'(-26336);
			7210: out = 24'(-26392);
			7211: out = 24'(-26516);
			7212: out = 24'(-26508);
			7213: out = 24'(-26548);
			7214: out = 24'(-26612);
			7215: out = 24'(-26660);
			7216: out = 24'(-26664);
			7217: out = 24'(-26756);
			7218: out = 24'(-26728);
			7219: out = 24'(-26852);
			7220: out = 24'(-26820);
			7221: out = 24'(-26880);
			7222: out = 24'(-26952);
			7223: out = 24'(-26940);
			7224: out = 24'(-26992);
			7225: out = 24'(-26996);
			7226: out = 24'(-26992);
			7227: out = 24'(-27056);
			7228: out = 24'(-27036);
			7229: out = 24'(-27068);
			7230: out = 24'(-27124);
			7231: out = 24'(-27084);
			7232: out = 24'(-27100);
			7233: out = 24'(-27136);
			7234: out = 24'(-27148);
			7235: out = 24'(-27128);
			7236: out = 24'(-27140);
			7237: out = 24'(-27128);
			7238: out = 24'(-27112);
			7239: out = 24'(-27084);
			7240: out = 24'(-27128);
			7241: out = 24'(-27100);
			7242: out = 24'(-27048);
			7243: out = 24'(-27068);
			7244: out = 24'(-27088);
			7245: out = 24'(-27044);
			7246: out = 24'(-27044);
			7247: out = 24'(-27076);
			7248: out = 24'(-26976);
			7249: out = 24'(-26960);
			7250: out = 24'(-26984);
			7251: out = 24'(-26920);
			7252: out = 24'(-26916);
			7253: out = 24'(-26860);
			7254: out = 24'(-26896);
			7255: out = 24'(-26840);
			7256: out = 24'(-26800);
			7257: out = 24'(-26856);
			7258: out = 24'(-26776);
			7259: out = 24'(-26724);
			7260: out = 24'(-26724);
			7261: out = 24'(-26664);
			7262: out = 24'(-26652);
			7263: out = 24'(-26588);
			7264: out = 24'(-26556);
			7265: out = 24'(-26572);
			7266: out = 24'(-26512);
			7267: out = 24'(-26444);
			7268: out = 24'(-26424);
			7269: out = 24'(-26416);
			7270: out = 24'(-26392);
			7271: out = 24'(-26356);
			7272: out = 24'(-26288);
			7273: out = 24'(-26244);
			7274: out = 24'(-26184);
			7275: out = 24'(-26184);
			7276: out = 24'(-26052);
			7277: out = 24'(-26048);
			7278: out = 24'(-26000);
			7279: out = 24'(-25952);
			7280: out = 24'(-25896);
			7281: out = 24'(-25820);
			7282: out = 24'(-25816);
			7283: out = 24'(-25724);
			7284: out = 24'(-25660);
			7285: out = 24'(-25636);
			7286: out = 24'(-25608);
			7287: out = 24'(-25500);
			7288: out = 24'(-25496);
			7289: out = 24'(-25360);
			7290: out = 24'(-25328);
			7291: out = 24'(-25244);
			7292: out = 24'(-25184);
			7293: out = 24'(-25104);
			7294: out = 24'(-25116);
			7295: out = 24'(-24980);
			7296: out = 24'(-24936);
			7297: out = 24'(-24904);
			7298: out = 24'(-24832);
			7299: out = 24'(-24736);
			7300: out = 24'(-24704);
			7301: out = 24'(-24628);
			7302: out = 24'(-24500);
			7303: out = 24'(-24472);
			7304: out = 24'(-24384);
			7305: out = 24'(-24332);
			7306: out = 24'(-24244);
			7307: out = 24'(-24180);
			7308: out = 24'(-24096);
			7309: out = 24'(-24028);
			7310: out = 24'(-23968);
			7311: out = 24'(-23864);
			7312: out = 24'(-23764);
			7313: out = 24'(-23692);
			7314: out = 24'(-23576);
			7315: out = 24'(-23480);
			7316: out = 24'(-23424);
			7317: out = 24'(-23296);
			7318: out = 24'(-23200);
			7319: out = 24'(-23084);
			7320: out = 24'(-22980);
			7321: out = 24'(-22888);
			7322: out = 24'(-22784);
			7323: out = 24'(-22632);
			7324: out = 24'(-22516);
			7325: out = 24'(-22440);
			7326: out = 24'(-22252);
			7327: out = 24'(-22140);
			7328: out = 24'(-22044);
			7329: out = 24'(-21860);
			7330: out = 24'(-21768);
			7331: out = 24'(-21604);
			7332: out = 24'(-21452);
			7333: out = 24'(-21352);
			7334: out = 24'(-21180);
			7335: out = 24'(-21044);
			7336: out = 24'(-20848);
			7337: out = 24'(-20704);
			7338: out = 24'(-20544);
			7339: out = 24'(-20380);
			7340: out = 24'(-20184);
			7341: out = 24'(-20056);
			7342: out = 24'(-19848);
			7343: out = 24'(-19664);
			7344: out = 24'(-19556);
			7345: out = 24'(-19336);
			7346: out = 24'(-19152);
			7347: out = 24'(-18996);
			7348: out = 24'(-18776);
			7349: out = 24'(-18616);
			7350: out = 24'(-18424);
			7351: out = 24'(-18216);
			7352: out = 24'(-18048);
			7353: out = 24'(-17832);
			7354: out = 24'(-17624);
			7355: out = 24'(-17428);
			7356: out = 24'(-17248);
			7357: out = 24'(-17052);
			7358: out = 24'(-16900);
			7359: out = 24'(-16696);
			7360: out = 24'(-16524);
			7361: out = 24'(-16316);
			7362: out = 24'(-16172);
			7363: out = 24'(-15936);
			7364: out = 24'(-15736);
			7365: out = 24'(-15592);
			7366: out = 24'(-15364);
			7367: out = 24'(-15180);
			7368: out = 24'(-15016);
			7369: out = 24'(-14772);
			7370: out = 24'(-14612);
			7371: out = 24'(-14456);
			7372: out = 24'(-14196);
			7373: out = 24'(-14120);
			7374: out = 24'(-13948);
			7375: out = 24'(-13728);
			7376: out = 24'(-13552);
			7377: out = 24'(-13312);
			7378: out = 24'(-13180);
			7379: out = 24'(-12996);
			7380: out = 24'(-12788);
			7381: out = 24'(-12632);
			7382: out = 24'(-12472);
			7383: out = 24'(-12280);
			7384: out = 24'(-12140);
			7385: out = 24'(-11992);
			7386: out = 24'(-11788);
			7387: out = 24'(-11572);
			7388: out = 24'(-11488);
			7389: out = 24'(-11252);
			7390: out = 24'(-11116);
			7391: out = 24'(-10968);
			7392: out = 24'(-10828);
			7393: out = 24'(-10672);
			7394: out = 24'(-10484);
			7395: out = 24'(-10320);
			7396: out = 24'(-10220);
			7397: out = 24'(-10016);
			7398: out = 24'(-9920);
			7399: out = 24'(-9760);
			7400: out = 24'(-9592);
			7401: out = 24'(-9424);
			7402: out = 24'(-9292);
			7403: out = 24'(-9192);
			7404: out = 24'(-9032);
			7405: out = 24'(-8884);
			7406: out = 24'(-8732);
			7407: out = 24'(-8616);
			7408: out = 24'(-8516);
			7409: out = 24'(-8352);
			7410: out = 24'(-8204);
			7411: out = 24'(-8084);
			7412: out = 24'(-7968);
			7413: out = 24'(-7800);
			7414: out = 24'(-7696);
			7415: out = 24'(-7612);
			7416: out = 24'(-7448);
			7417: out = 24'(-7328);
			7418: out = 24'(-7216);
			7419: out = 24'(-7104);
			7420: out = 24'(-7000);
			7421: out = 24'(-6856);
			7422: out = 24'(-6776);
			7423: out = 24'(-6620);
			7424: out = 24'(-6508);
			7425: out = 24'(-6400);
			7426: out = 24'(-6304);
			7427: out = 24'(-6172);
			7428: out = 24'(-6060);
			7429: out = 24'(-6000);
			7430: out = 24'(-5860);
			7431: out = 24'(-5816);
			7432: out = 24'(-5704);
			7433: out = 24'(-5540);
			7434: out = 24'(-5480);
			7435: out = 24'(-5344);
			7436: out = 24'(-5264);
			7437: out = 24'(-5160);
			7438: out = 24'(-5076);
			7439: out = 24'(-5012);
			7440: out = 24'(-4876);
			7441: out = 24'(-4728);
			7442: out = 24'(-4584);
			7443: out = 24'(-4376);
			7444: out = 24'(-4292);
			7445: out = 24'(-4064);
			7446: out = 24'(-3916);
			7447: out = 24'(-3752);
			7448: out = 24'(-3580);
			7449: out = 24'(-3460);
			7450: out = 24'(-3328);
			7451: out = 24'(-3160);
			7452: out = 24'(-3044);
			7453: out = 24'(-2880);
			7454: out = 24'(-2728);
			7455: out = 24'(-2652);
			7456: out = 24'(-2492);
			7457: out = 24'(-2324);
			7458: out = 24'(-2184);
			7459: out = 24'(-2076);
			7460: out = 24'(-1928);
			7461: out = 24'(-1768);
			7462: out = 24'(-1716);
			7463: out = 24'(-1552);
			7464: out = 24'(-1408);
			7465: out = 24'(-1300);
			7466: out = 24'(-1160);
			7467: out = 24'(-1076);
			7468: out = 24'(-924);
			7469: out = 24'(-840);
			7470: out = 24'(-696);
			7471: out = 24'(-636);
			7472: out = 24'(-512);
			7473: out = 24'(-388);
			7474: out = 24'(-260);
			7475: out = 24'(-164);
			7476: out = 24'(-60);
			7477: out = 24'(32);
			7478: out = 24'(116);
			7479: out = 24'(264);
			7480: out = 24'(316);
			7481: out = 24'(480);
			7482: out = 24'(552);
			7483: out = 24'(604);
			7484: out = 24'(728);
			7485: out = 24'(844);
			7486: out = 24'(912);
			7487: out = 24'(1024);
			7488: out = 24'(1152);
			7489: out = 24'(1216);
			7490: out = 24'(1348);
			7491: out = 24'(1424);
			7492: out = 24'(1516);
			7493: out = 24'(1596);
			7494: out = 24'(1744);
			7495: out = 24'(1740);
			7496: out = 24'(1880);
			7497: out = 24'(1956);
			7498: out = 24'(2088);
			7499: out = 24'(2184);
			7500: out = 24'(2236);
			7501: out = 24'(2324);
			7502: out = 24'(2432);
			7503: out = 24'(2532);
			7504: out = 24'(2576);
			7505: out = 24'(2704);
			7506: out = 24'(2764);
			7507: out = 24'(2888);
			7508: out = 24'(2968);
			7509: out = 24'(3012);
			7510: out = 24'(3160);
			7511: out = 24'(3224);
			7512: out = 24'(3336);
			7513: out = 24'(3380);
			7514: out = 24'(3544);
			7515: out = 24'(3584);
			7516: out = 24'(3728);
			7517: out = 24'(3820);
			7518: out = 24'(3900);
			7519: out = 24'(3964);
			7520: out = 24'(4140);
			7521: out = 24'(4144);
			7522: out = 24'(4276);
			7523: out = 24'(4392);
			7524: out = 24'(4484);
			7525: out = 24'(4624);
			7526: out = 24'(4672);
			7527: out = 24'(4820);
			7528: out = 24'(4904);
			7529: out = 24'(5020);
			7530: out = 24'(5120);
			7531: out = 24'(5236);
			7532: out = 24'(5364);
			7533: out = 24'(5460);
			7534: out = 24'(5572);
			7535: out = 24'(5740);
			7536: out = 24'(5872);
			7537: out = 24'(5988);
			7538: out = 24'(6112);
			7539: out = 24'(6276);
			7540: out = 24'(6400);
			7541: out = 24'(6520);
			7542: out = 24'(6736);
			7543: out = 24'(6772);
			7544: out = 24'(6996);
			7545: out = 24'(7084);
			7546: out = 24'(7252);
			7547: out = 24'(7396);
			7548: out = 24'(7460);
			7549: out = 24'(7696);
			7550: out = 24'(7796);
			7551: out = 24'(7980);
			7552: out = 24'(8128);
			7553: out = 24'(8324);
			7554: out = 24'(8468);
			7555: out = 24'(8692);
			7556: out = 24'(8772);
			7557: out = 24'(8972);
			7558: out = 24'(9172);
			7559: out = 24'(9328);
			7560: out = 24'(9480);
			7561: out = 24'(9688);
			7562: out = 24'(9856);
			7563: out = 24'(10020);
			7564: out = 24'(10192);
			7565: out = 24'(10420);
			7566: out = 24'(10528);
			7567: out = 24'(10760);
			7568: out = 24'(10888);
			7569: out = 24'(11116);
			7570: out = 24'(11236);
			7571: out = 24'(11448);
			7572: out = 24'(11592);
			7573: out = 24'(11780);
			7574: out = 24'(11952);
			7575: out = 24'(12096);
			7576: out = 24'(12264);
			7577: out = 24'(12476);
			7578: out = 24'(12640);
			7579: out = 24'(12764);
			7580: out = 24'(12980);
			7581: out = 24'(13116);
			7582: out = 24'(13268);
			7583: out = 24'(13452);
			7584: out = 24'(13588);
			7585: out = 24'(13752);
			7586: out = 24'(13904);
			7587: out = 24'(14068);
			7588: out = 24'(14220);
			7589: out = 24'(14392);
			7590: out = 24'(14476);
			7591: out = 24'(14688);
			7592: out = 24'(14824);
			7593: out = 24'(14984);
			7594: out = 24'(15112);
			7595: out = 24'(15256);
			7596: out = 24'(15352);
			7597: out = 24'(15540);
			7598: out = 24'(15684);
			7599: out = 24'(15832);
			7600: out = 24'(15952);
			7601: out = 24'(16112);
			7602: out = 24'(16212);
			7603: out = 24'(16316);
			7604: out = 24'(16460);
			7605: out = 24'(16616);
			7606: out = 24'(16732);
			7607: out = 24'(16824);
			7608: out = 24'(16988);
			7609: out = 24'(17120);
			7610: out = 24'(17204);
			7611: out = 24'(17340);
			7612: out = 24'(17456);
			7613: out = 24'(17580);
			7614: out = 24'(17660);
			7615: out = 24'(17824);
			7616: out = 24'(17888);
			7617: out = 24'(18036);
			7618: out = 24'(18152);
			7619: out = 24'(18212);
			7620: out = 24'(18308);
			7621: out = 24'(18468);
			7622: out = 24'(18548);
			7623: out = 24'(18656);
			7624: out = 24'(18748);
			7625: out = 24'(18900);
			7626: out = 24'(18996);
			7627: out = 24'(19080);
			7628: out = 24'(19144);
			7629: out = 24'(19256);
			7630: out = 24'(19376);
			7631: out = 24'(19472);
			7632: out = 24'(19492);
			7633: out = 24'(19648);
			7634: out = 24'(19704);
			7635: out = 24'(19816);
			7636: out = 24'(19904);
			7637: out = 24'(19976);
			7638: out = 24'(20100);
			7639: out = 24'(20160);
			7640: out = 24'(20264);
			7641: out = 24'(20332);
			7642: out = 24'(20428);
			7643: out = 24'(20508);
			7644: out = 24'(20596);
			7645: out = 24'(20680);
			7646: out = 24'(20788);
			7647: out = 24'(20816);
			7648: out = 24'(20892);
			7649: out = 24'(21008);
			7650: out = 24'(21080);
			7651: out = 24'(21140);
			7652: out = 24'(21256);
			7653: out = 24'(21320);
			7654: out = 24'(21404);
			7655: out = 24'(21460);
			7656: out = 24'(21588);
			7657: out = 24'(21624);
			7658: out = 24'(21688);
			7659: out = 24'(21760);
			7660: out = 24'(21824);
			7661: out = 24'(21896);
			7662: out = 24'(22004);
			7663: out = 24'(22088);
			7664: out = 24'(22092);
			7665: out = 24'(22204);
			7666: out = 24'(22268);
			7667: out = 24'(22304);
			7668: out = 24'(22412);
			7669: out = 24'(22488);
			7670: out = 24'(22460);
			7671: out = 24'(22512);
			7672: out = 24'(22676);
			7673: out = 24'(22660);
			7674: out = 24'(22688);
			7675: out = 24'(22768);
			7676: out = 24'(22696);
			7677: out = 24'(22796);
			7678: out = 24'(22704);
			7679: out = 24'(22808);
			7680: out = 24'(22776);
			7681: out = 24'(22832);
			7682: out = 24'(22768);
			7683: out = 24'(22800);
			7684: out = 24'(22776);
			7685: out = 24'(22744);
			7686: out = 24'(22736);
			7687: out = 24'(22712);
			7688: out = 24'(22832);
			7689: out = 24'(22716);
			7690: out = 24'(22724);
			7691: out = 24'(22708);
			7692: out = 24'(22724);
			7693: out = 24'(22592);
			7694: out = 24'(22604);
			7695: out = 24'(22632);
			7696: out = 24'(22592);
			7697: out = 24'(22512);
			7698: out = 24'(22536);
			7699: out = 24'(22500);
			7700: out = 24'(22532);
			7701: out = 24'(22368);
			7702: out = 24'(22416);
			7703: out = 24'(22536);
			7704: out = 24'(22440);
			7705: out = 24'(22464);
			7706: out = 24'(22432);
			7707: out = 24'(22588);
			7708: out = 24'(22488);
			7709: out = 24'(22440);
			7710: out = 24'(22488);
			7711: out = 24'(22468);
			7712: out = 24'(22376);
			7713: out = 24'(22400);
			7714: out = 24'(22300);
			7715: out = 24'(22228);
			7716: out = 24'(22376);
			7717: out = 24'(22300);
			7718: out = 24'(22380);
			7719: out = 24'(22200);
			7720: out = 24'(22368);
			7721: out = 24'(22304);
			7722: out = 24'(22284);
			7723: out = 24'(22352);
			7724: out = 24'(22408);
			7725: out = 24'(22404);
			7726: out = 24'(22320);
			7727: out = 24'(22364);
			7728: out = 24'(22320);
			7729: out = 24'(22304);
			7730: out = 24'(22280);
			7731: out = 24'(22168);
			7732: out = 24'(22148);
			7733: out = 24'(22208);
			7734: out = 24'(22060);
			7735: out = 24'(22072);
			7736: out = 24'(22024);
			7737: out = 24'(22120);
			7738: out = 24'(22040);
			7739: out = 24'(22072);
			7740: out = 24'(22016);
			7741: out = 24'(21968);
			7742: out = 24'(21908);
			7743: out = 24'(21872);
			7744: out = 24'(21904);
			7745: out = 24'(21876);
			7746: out = 24'(21784);
			7747: out = 24'(21744);
			7748: out = 24'(21692);
			7749: out = 24'(21664);
			7750: out = 24'(21528);
			7751: out = 24'(21524);
			7752: out = 24'(21444);
			7753: out = 24'(21380);
			7754: out = 24'(21364);
			7755: out = 24'(21308);
			7756: out = 24'(21176);
			7757: out = 24'(21112);
			7758: out = 24'(21032);
			7759: out = 24'(20956);
			7760: out = 24'(20960);
			7761: out = 24'(20844);
			7762: out = 24'(20692);
			7763: out = 24'(20688);
			7764: out = 24'(20456);
			7765: out = 24'(20420);
			7766: out = 24'(20356);
			7767: out = 24'(20192);
			7768: out = 24'(20168);
			7769: out = 24'(20060);
			7770: out = 24'(19868);
			7771: out = 24'(19732);
			7772: out = 24'(19720);
			7773: out = 24'(19520);
			7774: out = 24'(19368);
			7775: out = 24'(19332);
			7776: out = 24'(19156);
			7777: out = 24'(19020);
			7778: out = 24'(19008);
			7779: out = 24'(18784);
			7780: out = 24'(18736);
			7781: out = 24'(18516);
			7782: out = 24'(18400);
			7783: out = 24'(18292);
			7784: out = 24'(18108);
			7785: out = 24'(18020);
			7786: out = 24'(17896);
			7787: out = 24'(17788);
			7788: out = 24'(17636);
			7789: out = 24'(17428);
			7790: out = 24'(17376);
			7791: out = 24'(17196);
			7792: out = 24'(17008);
			7793: out = 24'(16908);
			7794: out = 24'(16768);
			7795: out = 24'(16588);
			7796: out = 24'(16388);
			7797: out = 24'(16196);
			7798: out = 24'(16052);
			7799: out = 24'(15968);
			7800: out = 24'(15780);
			7801: out = 24'(15640);
			7802: out = 24'(15560);
			7803: out = 24'(15424);
			7804: out = 24'(15332);
			7805: out = 24'(15116);
			7806: out = 24'(14980);
			7807: out = 24'(14840);
			7808: out = 24'(14616);
			7809: out = 24'(14588);
			7810: out = 24'(14268);
			7811: out = 24'(14176);
			7812: out = 24'(14044);
			7813: out = 24'(13908);
			7814: out = 24'(13764);
			7815: out = 24'(13620);
			7816: out = 24'(13520);
			7817: out = 24'(13356);
			7818: out = 24'(13160);
			7819: out = 24'(13096);
			7820: out = 24'(12976);
			7821: out = 24'(12744);
			7822: out = 24'(12592);
			7823: out = 24'(12484);
			7824: out = 24'(12328);
			7825: out = 24'(12220);
			7826: out = 24'(12108);
			7827: out = 24'(11900);
			7828: out = 24'(11852);
			7829: out = 24'(11656);
			7830: out = 24'(11536);
			7831: out = 24'(11400);
			7832: out = 24'(11344);
			7833: out = 24'(11172);
			7834: out = 24'(10944);
			7835: out = 24'(10992);
			7836: out = 24'(10720);
			7837: out = 24'(10712);
			7838: out = 24'(10516);
			7839: out = 24'(10392);
			7840: out = 24'(10336);
			7841: out = 24'(10184);
			7842: out = 24'(10068);
			7843: out = 24'(9996);
			7844: out = 24'(9776);
			7845: out = 24'(9728);
			7846: out = 24'(9532);
			7847: out = 24'(9436);
			7848: out = 24'(9388);
			7849: out = 24'(9236);
			7850: out = 24'(9100);
			7851: out = 24'(9056);
			7852: out = 24'(8860);
			7853: out = 24'(8764);
			7854: out = 24'(8712);
			7855: out = 24'(8604);
			7856: out = 24'(8512);
			7857: out = 24'(8320);
			7858: out = 24'(8292);
			7859: out = 24'(8108);
			7860: out = 24'(8084);
			7861: out = 24'(8016);
			7862: out = 24'(7844);
			7863: out = 24'(7780);
			7864: out = 24'(7652);
			7865: out = 24'(7548);
			7866: out = 24'(7500);
			7867: out = 24'(7352);
			7868: out = 24'(7260);
			7869: out = 24'(7156);
			7870: out = 24'(7020);
			7871: out = 24'(7016);
			7872: out = 24'(6880);
			7873: out = 24'(6788);
			7874: out = 24'(6716);
			7875: out = 24'(6656);
			7876: out = 24'(6516);
			7877: out = 24'(6488);
			7878: out = 24'(6372);
			7879: out = 24'(6308);
			7880: out = 24'(6144);
			7881: out = 24'(6084);
			7882: out = 24'(6052);
			7883: out = 24'(5960);
			7884: out = 24'(5860);
			7885: out = 24'(5804);
			7886: out = 24'(5756);
			7887: out = 24'(5620);
			7888: out = 24'(5532);
			7889: out = 24'(5540);
			7890: out = 24'(5428);
			7891: out = 24'(5316);
			7892: out = 24'(5284);
			7893: out = 24'(5168);
			7894: out = 24'(5124);
			7895: out = 24'(5088);
			7896: out = 24'(4932);
			7897: out = 24'(4932);
			7898: out = 24'(4804);
			7899: out = 24'(4752);
			7900: out = 24'(4700);
			7901: out = 24'(4624);
			7902: out = 24'(4564);
			7903: out = 24'(4528);
			7904: out = 24'(4456);
			7905: out = 24'(4376);
			7906: out = 24'(4324);
			7907: out = 24'(4228);
			7908: out = 24'(4112);
			7909: out = 24'(3968);
			7910: out = 24'(3804);
			7911: out = 24'(3540);
			7912: out = 24'(3372);
			7913: out = 24'(3172);
			7914: out = 24'(3072);
			7915: out = 24'(2908);
			7916: out = 24'(2708);
			7917: out = 24'(2616);
			7918: out = 24'(2444);
			7919: out = 24'(2232);
			7920: out = 24'(2116);
			7921: out = 24'(1956);
			7922: out = 24'(1808);
			7923: out = 24'(1672);
			7924: out = 24'(1556);
			7925: out = 24'(1356);
			7926: out = 24'(1192);
			7927: out = 24'(1168);
			7928: out = 24'(900);
			7929: out = 24'(820);
			7930: out = 24'(652);
			7931: out = 24'(508);
			7932: out = 24'(432);
			7933: out = 24'(208);
			7934: out = 24'(148);
			7935: out = 24'(-12);
			7936: out = 24'(-144);
			7937: out = 24'(-252);
			7938: out = 24'(-404);
			7939: out = 24'(-500);
			7940: out = 24'(-604);
			7941: out = 24'(-740);
			7942: out = 24'(-916);
			7943: out = 24'(-964);
			7944: out = 24'(-1124);
			7945: out = 24'(-1224);
			7946: out = 24'(-1316);
			7947: out = 24'(-1488);
			7948: out = 24'(-1548);
			7949: out = 24'(-1692);
			7950: out = 24'(-1736);
			7951: out = 24'(-1876);
			7952: out = 24'(-1972);
			7953: out = 24'(-2132);
			7954: out = 24'(-2236);
			7955: out = 24'(-2288);
			7956: out = 24'(-2472);
			7957: out = 24'(-2512);
			7958: out = 24'(-2612);
			7959: out = 24'(-2780);
			7960: out = 24'(-2836);
			7961: out = 24'(-2956);
			7962: out = 24'(-3024);
			7963: out = 24'(-3152);
			7964: out = 24'(-3252);
			7965: out = 24'(-3420);
			7966: out = 24'(-3472);
			7967: out = 24'(-3564);
			7968: out = 24'(-3712);
			7969: out = 24'(-3780);
			7970: out = 24'(-3868);
			7971: out = 24'(-3988);
			7972: out = 24'(-4064);
			7973: out = 24'(-4172);
			7974: out = 24'(-4252);
			7975: out = 24'(-4372);
			7976: out = 24'(-4484);
			7977: out = 24'(-4568);
			7978: out = 24'(-4744);
			7979: out = 24'(-4752);
			7980: out = 24'(-4904);
			7981: out = 24'(-4980);
			7982: out = 24'(-5076);
			7983: out = 24'(-5192);
			7984: out = 24'(-5312);
			7985: out = 24'(-5408);
			7986: out = 24'(-5496);
			7987: out = 24'(-5612);
			7988: out = 24'(-5752);
			7989: out = 24'(-5744);
			7990: out = 24'(-5856);
			7991: out = 24'(-6004);
			7992: out = 24'(-6144);
			7993: out = 24'(-6244);
			7994: out = 24'(-6392);
			7995: out = 24'(-6524);
			7996: out = 24'(-6636);
			7997: out = 24'(-6744);
			7998: out = 24'(-6868);
			7999: out = 24'(-6996);
			8000: out = 24'(-7060);
			8001: out = 24'(-7236);
			8002: out = 24'(-7356);
			8003: out = 24'(-7468);
			8004: out = 24'(-7600);
			8005: out = 24'(-7756);
			8006: out = 24'(-7932);
			8007: out = 24'(-8024);
			8008: out = 24'(-8136);
			8009: out = 24'(-8308);
			8010: out = 24'(-8440);
			8011: out = 24'(-8568);
			8012: out = 24'(-8784);
			8013: out = 24'(-8864);
			8014: out = 24'(-9052);
			8015: out = 24'(-9160);
			8016: out = 24'(-9384);
			8017: out = 24'(-9492);
			8018: out = 24'(-9688);
			8019: out = 24'(-9848);
			8020: out = 24'(-10004);
			8021: out = 24'(-10160);
			8022: out = 24'(-10388);
			8023: out = 24'(-10544);
			8024: out = 24'(-10676);
			8025: out = 24'(-10892);
			8026: out = 24'(-11032);
			8027: out = 24'(-11284);
			8028: out = 24'(-11440);
			8029: out = 24'(-11652);
			8030: out = 24'(-11876);
			8031: out = 24'(-12024);
			8032: out = 24'(-12180);
			8033: out = 24'(-12436);
			8034: out = 24'(-12604);
			8035: out = 24'(-12788);
			8036: out = 24'(-13020);
			8037: out = 24'(-13232);
			8038: out = 24'(-13412);
			8039: out = 24'(-13636);
			8040: out = 24'(-13880);
			8041: out = 24'(-14020);
			8042: out = 24'(-14288);
			8043: out = 24'(-14464);
			8044: out = 24'(-14664);
			8045: out = 24'(-14848);
			8046: out = 24'(-15028);
			8047: out = 24'(-15256);
			8048: out = 24'(-15448);
			8049: out = 24'(-15640);
			8050: out = 24'(-15896);
			8051: out = 24'(-16020);
			8052: out = 24'(-16248);
			8053: out = 24'(-16380);
			8054: out = 24'(-16588);
			8055: out = 24'(-16772);
			8056: out = 24'(-16936);
			8057: out = 24'(-17136);
			8058: out = 24'(-17316);
			8059: out = 24'(-17468);
			8060: out = 24'(-17572);
			8061: out = 24'(-17808);
			8062: out = 24'(-17952);
			8063: out = 24'(-18104);
			8064: out = 24'(-18212);
			8065: out = 24'(-18432);
			8066: out = 24'(-18512);
			8067: out = 24'(-18700);
			8068: out = 24'(-18852);
			8069: out = 24'(-18944);
			8070: out = 24'(-19096);
			8071: out = 24'(-19232);
			8072: out = 24'(-19316);
			8073: out = 24'(-19516);
			8074: out = 24'(-19544);
			8075: out = 24'(-19712);
			8076: out = 24'(-19824);
			8077: out = 24'(-19968);
			8078: out = 24'(-20016);
			8079: out = 24'(-20192);
			8080: out = 24'(-20268);
			8081: out = 24'(-20408);
			8082: out = 24'(-20504);
			8083: out = 24'(-20580);
			8084: out = 24'(-20640);
			8085: out = 24'(-20760);
			8086: out = 24'(-20856);
			8087: out = 24'(-20856);
			8088: out = 24'(-21012);
			8089: out = 24'(-21088);
			8090: out = 24'(-21136);
			8091: out = 24'(-21228);
			8092: out = 24'(-21312);
			8093: out = 24'(-21368);
			8094: out = 24'(-21444);
			8095: out = 24'(-21428);
			8096: out = 24'(-21556);
			8097: out = 24'(-21556);
			8098: out = 24'(-21672);
			8099: out = 24'(-21692);
			8100: out = 24'(-21700);
			8101: out = 24'(-21788);
			8102: out = 24'(-21816);
			8103: out = 24'(-21880);
			8104: out = 24'(-21936);
			8105: out = 24'(-21968);
			8106: out = 24'(-21984);
			8107: out = 24'(-22036);
			8108: out = 24'(-22000);
			8109: out = 24'(-22124);
			8110: out = 24'(-22060);
			8111: out = 24'(-22132);
			8112: out = 24'(-22192);
			8113: out = 24'(-22168);
			8114: out = 24'(-22200);
			8115: out = 24'(-22256);
			8116: out = 24'(-22248);
			8117: out = 24'(-22252);
			8118: out = 24'(-22268);
			8119: out = 24'(-22280);
			8120: out = 24'(-22324);
			8121: out = 24'(-22324);
			8122: out = 24'(-22308);
			8123: out = 24'(-22324);
			8124: out = 24'(-22308);
			8125: out = 24'(-22348);
			8126: out = 24'(-22384);
			8127: out = 24'(-22348);
			8128: out = 24'(-22364);
			8129: out = 24'(-22324);
			8130: out = 24'(-22352);
			8131: out = 24'(-22316);
			8132: out = 24'(-22320);
			8133: out = 24'(-22384);
			8134: out = 24'(-22252);
			8135: out = 24'(-22304);
			8136: out = 24'(-22276);
			8137: out = 24'(-22296);
			8138: out = 24'(-22288);
			8139: out = 24'(-22236);
			8140: out = 24'(-22252);
			8141: out = 24'(-22192);
			8142: out = 24'(-22216);
			8143: out = 24'(-22180);
			8144: out = 24'(-22136);
			8145: out = 24'(-22140);
			8146: out = 24'(-22108);
			8147: out = 24'(-22040);
			8148: out = 24'(-22068);
			8149: out = 24'(-22076);
			8150: out = 24'(-21980);
			8151: out = 24'(-21972);
			8152: out = 24'(-22020);
			8153: out = 24'(-21896);
			8154: out = 24'(-21896);
			8155: out = 24'(-21852);
			8156: out = 24'(-21812);
			8157: out = 24'(-21828);
			8158: out = 24'(-21764);
			8159: out = 24'(-21700);
			8160: out = 24'(-21684);
			8161: out = 24'(-21656);
			8162: out = 24'(-21624);
			8163: out = 24'(-21612);
			8164: out = 24'(-21592);
			8165: out = 24'(-21464);
			8166: out = 24'(-21504);
			8167: out = 24'(-21504);
			8168: out = 24'(-21416);
			8169: out = 24'(-21396);
			8170: out = 24'(-21316);
			8171: out = 24'(-21292);
			8172: out = 24'(-21256);
			8173: out = 24'(-21192);
			8174: out = 24'(-21136);
			8175: out = 24'(-21068);
			8176: out = 24'(-21036);
			8177: out = 24'(-20948);
			8178: out = 24'(-20904);
			8179: out = 24'(-20932);
			8180: out = 24'(-20816);
			8181: out = 24'(-20736);
			8182: out = 24'(-20724);
			8183: out = 24'(-20680);
			8184: out = 24'(-20596);
			8185: out = 24'(-20552);
			8186: out = 24'(-20504);
			8187: out = 24'(-20468);
			8188: out = 24'(-20360);
			8189: out = 24'(-20380);
			8190: out = 24'(-20292);
			8191: out = 24'(-20224);
			8192: out = 24'(-20176);
			8193: out = 24'(-20120);
			8194: out = 24'(-20044);
			8195: out = 24'(-19968);
			8196: out = 24'(-19928);
			8197: out = 24'(-19868);
			8198: out = 24'(-19820);
			8199: out = 24'(-19724);
			8200: out = 24'(-19628);
			8201: out = 24'(-19600);
			8202: out = 24'(-19524);
			8203: out = 24'(-19488);
			8204: out = 24'(-19368);
			8205: out = 24'(-19324);
			8206: out = 24'(-19228);
			8207: out = 24'(-19160);
			8208: out = 24'(-19024);
			8209: out = 24'(-19060);
			8210: out = 24'(-18860);
			8211: out = 24'(-18844);
			8212: out = 24'(-18692);
			8213: out = 24'(-18668);
			8214: out = 24'(-18568);
			8215: out = 24'(-18444);
			8216: out = 24'(-18356);
			8217: out = 24'(-18244);
			8218: out = 24'(-18152);
			8219: out = 24'(-18008);
			8220: out = 24'(-17948);
			8221: out = 24'(-17800);
			8222: out = 24'(-17680);
			8223: out = 24'(-17572);
			8224: out = 24'(-17436);
			8225: out = 24'(-17380);
			8226: out = 24'(-17248);
			8227: out = 24'(-17056);
			8228: out = 24'(-17000);
			8229: out = 24'(-16776);
			8230: out = 24'(-16684);
			8231: out = 24'(-16544);
			8232: out = 24'(-16416);
			8233: out = 24'(-16216);
			8234: out = 24'(-16156);
			8235: out = 24'(-15968);
			8236: out = 24'(-15816);
			8237: out = 24'(-15700);
			8238: out = 24'(-15564);
			8239: out = 24'(-15384);
			8240: out = 24'(-15252);
			8241: out = 24'(-15048);
			8242: out = 24'(-14944);
			8243: out = 24'(-14740);
			8244: out = 24'(-14608);
			8245: out = 24'(-14488);
			8246: out = 24'(-14256);
			8247: out = 24'(-14164);
			8248: out = 24'(-14040);
			8249: out = 24'(-13816);
			8250: out = 24'(-13712);
			8251: out = 24'(-13476);
			8252: out = 24'(-13340);
			8253: out = 24'(-13200);
			8254: out = 24'(-13024);
			8255: out = 24'(-12896);
			8256: out = 24'(-12744);
			8257: out = 24'(-12584);
			8258: out = 24'(-12436);
			8259: out = 24'(-12276);
			8260: out = 24'(-12108);
			8261: out = 24'(-11964);
			8262: out = 24'(-11816);
			8263: out = 24'(-11668);
			8264: out = 24'(-11512);
			8265: out = 24'(-11380);
			8266: out = 24'(-11180);
			8267: out = 24'(-11144);
			8268: out = 24'(-10888);
			8269: out = 24'(-10784);
			8270: out = 24'(-10644);
			8271: out = 24'(-10456);
			8272: out = 24'(-10372);
			8273: out = 24'(-10168);
			8274: out = 24'(-10068);
			8275: out = 24'(-9904);
			8276: out = 24'(-9784);
			8277: out = 24'(-9632);
			8278: out = 24'(-9508);
			8279: out = 24'(-9396);
			8280: out = 24'(-9208);
			8281: out = 24'(-9096);
			8282: out = 24'(-8980);
			8283: out = 24'(-8820);
			8284: out = 24'(-8752);
			8285: out = 24'(-8568);
			8286: out = 24'(-8440);
			8287: out = 24'(-8356);
			8288: out = 24'(-8192);
			8289: out = 24'(-8088);
			8290: out = 24'(-7932);
			8291: out = 24'(-7876);
			8292: out = 24'(-7724);
			8293: out = 24'(-7608);
			8294: out = 24'(-7496);
			8295: out = 24'(-7392);
			8296: out = 24'(-7264);
			8297: out = 24'(-7160);
			8298: out = 24'(-7012);
			8299: out = 24'(-6940);
			8300: out = 24'(-6812);
			8301: out = 24'(-6688);
			8302: out = 24'(-6620);
			8303: out = 24'(-6516);
			8304: out = 24'(-6368);
			8305: out = 24'(-6352);
			8306: out = 24'(-6188);
			8307: out = 24'(-6080);
			8308: out = 24'(-5980);
			8309: out = 24'(-5884);
			8310: out = 24'(-5828);
			8311: out = 24'(-5696);
			8312: out = 24'(-5640);
			8313: out = 24'(-5444);
			8314: out = 24'(-5456);
			8315: out = 24'(-5352);
			8316: out = 24'(-5200);
			8317: out = 24'(-5168);
			8318: out = 24'(-5072);
			8319: out = 24'(-4956);
			8320: out = 24'(-4884);
			8321: out = 24'(-4792);
			8322: out = 24'(-4712);
			8323: out = 24'(-4640);
			8324: out = 24'(-4524);
			8325: out = 24'(-4472);
			8326: out = 24'(-4424);
			8327: out = 24'(-4324);
			8328: out = 24'(-4208);
			8329: out = 24'(-4172);
			8330: out = 24'(-4064);
			8331: out = 24'(-3980);
			8332: out = 24'(-3888);
			8333: out = 24'(-3792);
			8334: out = 24'(-3628);
			8335: out = 24'(-3488);
			8336: out = 24'(-3392);
			8337: out = 24'(-3212);
			8338: out = 24'(-3120);
			8339: out = 24'(-3016);
			8340: out = 24'(-2816);
			8341: out = 24'(-2752);
			8342: out = 24'(-2620);
			8343: out = 24'(-2512);
			8344: out = 24'(-2380);
			8345: out = 24'(-2260);
			8346: out = 24'(-2196);
			8347: out = 24'(-2040);
			8348: out = 24'(-1952);
			8349: out = 24'(-1820);
			8350: out = 24'(-1728);
			8351: out = 24'(-1592);
			8352: out = 24'(-1572);
			8353: out = 24'(-1440);
			8354: out = 24'(-1344);
			8355: out = 24'(-1220);
			8356: out = 24'(-1144);
			8357: out = 24'(-1008);
			8358: out = 24'(-900);
			8359: out = 24'(-864);
			8360: out = 24'(-704);
			8361: out = 24'(-624);
			8362: out = 24'(-580);
			8363: out = 24'(-476);
			8364: out = 24'(-324);
			8365: out = 24'(-288);
			8366: out = 24'(-164);
			8367: out = 24'(-120);
			8368: out = 24'(-56);
			8369: out = 24'(36);
			8370: out = 24'(200);
			8371: out = 24'(184);
			8372: out = 24'(300);
			8373: out = 24'(420);
			8374: out = 24'(456);
			8375: out = 24'(552);
			8376: out = 24'(648);
			8377: out = 24'(704);
			8378: out = 24'(776);
			8379: out = 24'(900);
			8380: out = 24'(924);
			8381: out = 24'(1048);
			8382: out = 24'(1096);
			8383: out = 24'(1212);
			8384: out = 24'(1204);
			8385: out = 24'(1364);
			8386: out = 24'(1400);
			8387: out = 24'(1456);
			8388: out = 24'(1580);
			8389: out = 24'(1616);
			8390: out = 24'(1712);
			8391: out = 24'(1772);
			8392: out = 24'(1848);
			8393: out = 24'(1936);
			8394: out = 24'(1964);
			8395: out = 24'(2088);
			8396: out = 24'(2152);
			8397: out = 24'(2200);
			8398: out = 24'(2292);
			8399: out = 24'(2328);
			8400: out = 24'(2456);
			8401: out = 24'(2520);
			8402: out = 24'(2580);
			8403: out = 24'(2612);
			8404: out = 24'(2740);
			8405: out = 24'(2808);
			8406: out = 24'(2904);
			8407: out = 24'(2924);
			8408: out = 24'(3048);
			8409: out = 24'(3084);
			8410: out = 24'(3200);
			8411: out = 24'(3284);
			8412: out = 24'(3344);
			8413: out = 24'(3464);
			8414: out = 24'(3484);
			8415: out = 24'(3624);
			8416: out = 24'(3684);
			8417: out = 24'(3760);
			8418: out = 24'(3876);
			8419: out = 24'(3932);
			8420: out = 24'(4044);
			8421: out = 24'(4140);
			8422: out = 24'(4236);
			8423: out = 24'(4292);
			8424: out = 24'(4432);
			8425: out = 24'(4484);
			8426: out = 24'(4600);
			8427: out = 24'(4692);
			8428: out = 24'(4820);
			8429: out = 24'(4932);
			8430: out = 24'(5036);
			8431: out = 24'(5160);
			8432: out = 24'(5220);
			8433: out = 24'(5376);
			8434: out = 24'(5432);
			8435: out = 24'(5592);
			8436: out = 24'(5656);
			8437: out = 24'(5844);
			8438: out = 24'(5944);
			8439: out = 24'(6092);
			8440: out = 24'(6208);
			8441: out = 24'(6304);
			8442: out = 24'(6456);
			8443: out = 24'(6560);
			8444: out = 24'(6696);
			8445: out = 24'(6772);
			8446: out = 24'(6984);
			8447: out = 24'(7076);
			8448: out = 24'(7224);
			8449: out = 24'(7388);
			8450: out = 24'(7512);
			8451: out = 24'(7652);
			8452: out = 24'(7800);
			8453: out = 24'(7960);
			8454: out = 24'(8052);
			8455: out = 24'(8212);
			8456: out = 24'(8392);
			8457: out = 24'(8496);
			8458: out = 24'(8676);
			8459: out = 24'(8788);
			8460: out = 24'(8960);
			8461: out = 24'(9060);
			8462: out = 24'(9216);
			8463: out = 24'(9384);
			8464: out = 24'(9536);
			8465: out = 24'(9624);
			8466: out = 24'(9788);
			8467: out = 24'(9916);
			8468: out = 24'(10048);
			8469: out = 24'(10216);
			8470: out = 24'(10308);
			8471: out = 24'(10472);
			8472: out = 24'(10616);
			8473: out = 24'(10732);
			8474: out = 24'(10880);
			8475: out = 24'(11048);
			8476: out = 24'(11128);
			8477: out = 24'(11260);
			8478: out = 24'(11396);
			8479: out = 24'(11528);
			8480: out = 24'(11624);
			8481: out = 24'(11800);
			8482: out = 24'(11916);
			8483: out = 24'(12032);
			8484: out = 24'(12140);
			8485: out = 24'(12284);
			8486: out = 24'(12348);
			8487: out = 24'(12508);
			8488: out = 24'(12608);
			8489: out = 24'(12664);
			8490: out = 24'(12848);
			8491: out = 24'(12908);
			8492: out = 24'(13056);
			8493: out = 24'(13184);
			8494: out = 24'(13232);
			8495: out = 24'(13380);
			8496: out = 24'(13452);
			8497: out = 24'(13572);
			8498: out = 24'(13684);
			8499: out = 24'(13764);
			8500: out = 24'(13832);
			8501: out = 24'(13956);
			8502: out = 24'(14060);
			8503: out = 24'(14116);
			8504: out = 24'(14300);
			8505: out = 24'(14332);
			8506: out = 24'(14440);
			8507: out = 24'(14560);
			8508: out = 24'(14580);
			8509: out = 24'(14728);
			8510: out = 24'(14828);
			8511: out = 24'(14868);
			8512: out = 24'(14944);
			8513: out = 24'(15048);
			8514: out = 24'(15112);
			8515: out = 24'(15264);
			8516: out = 24'(15320);
			8517: out = 24'(15396);
			8518: out = 24'(15508);
			8519: out = 24'(15520);
			8520: out = 24'(15668);
			8521: out = 24'(15728);
			8522: out = 24'(15864);
			8523: out = 24'(15920);
			8524: out = 24'(15984);
			8525: out = 24'(16072);
			8526: out = 24'(16136);
			8527: out = 24'(16168);
			8528: out = 24'(16288);
			8529: out = 24'(16304);
			8530: out = 24'(16436);
			8531: out = 24'(16488);
			8532: out = 24'(16480);
			8533: out = 24'(16636);
			8534: out = 24'(16676);
			8535: out = 24'(16740);
			8536: out = 24'(16812);
			8537: out = 24'(16900);
			8538: out = 24'(16956);
			8539: out = 24'(17020);
			8540: out = 24'(17020);
			8541: out = 24'(17160);
			8542: out = 24'(17168);
			8543: out = 24'(17268);
			8544: out = 24'(17360);
			8545: out = 24'(17424);
			8546: out = 24'(17436);
			8547: out = 24'(17528);
			8548: out = 24'(17616);
			8549: out = 24'(17620);
			8550: out = 24'(17732);
			8551: out = 24'(17756);
			8552: out = 24'(17788);
			8553: out = 24'(17916);
			8554: out = 24'(17960);
			8555: out = 24'(17988);
			8556: out = 24'(18096);
			8557: out = 24'(18112);
			8558: out = 24'(18188);
			8559: out = 24'(18208);
			8560: out = 24'(18336);
			8561: out = 24'(18344);
			8562: out = 24'(18396);
			8563: out = 24'(18416);
			8564: out = 24'(18540);
			8565: out = 24'(18524);
			8566: out = 24'(18536);
			8567: out = 24'(18620);
			8568: out = 24'(18644);
			8569: out = 24'(18624);
			8570: out = 24'(18560);
			8571: out = 24'(18628);
			8572: out = 24'(18604);
			8573: out = 24'(18532);
			8574: out = 24'(18540);
			8575: out = 24'(18632);
			8576: out = 24'(18520);
			8577: out = 24'(18528);
			8578: out = 24'(18544);
			8579: out = 24'(18516);
			8580: out = 24'(18568);
			8581: out = 24'(18500);
			8582: out = 24'(18484);
			8583: out = 24'(18468);
			8584: out = 24'(18536);
			8585: out = 24'(18544);
			8586: out = 24'(18360);
			8587: out = 24'(18428);
			8588: out = 24'(18464);
			8589: out = 24'(18468);
			8590: out = 24'(18416);
			8591: out = 24'(18472);
			8592: out = 24'(18480);
			8593: out = 24'(18448);
			8594: out = 24'(18392);
			8595: out = 24'(18492);
			8596: out = 24'(18392);
			8597: out = 24'(18384);
			8598: out = 24'(18336);
			8599: out = 24'(18376);
			8600: out = 24'(18348);
			8601: out = 24'(18336);
			8602: out = 24'(18276);
			8603: out = 24'(18352);
			8604: out = 24'(18372);
			8605: out = 24'(18296);
			8606: out = 24'(18352);
			8607: out = 24'(18372);
			8608: out = 24'(18292);
			8609: out = 24'(18340);
			8610: out = 24'(18236);
			8611: out = 24'(18252);
			8612: out = 24'(18272);
			8613: out = 24'(18292);
			8614: out = 24'(18348);
			8615: out = 24'(18300);
			8616: out = 24'(18260);
			8617: out = 24'(18248);
			8618: out = 24'(18296);
			8619: out = 24'(18312);
			8620: out = 24'(18216);
			8621: out = 24'(18212);
			8622: out = 24'(18236);
			8623: out = 24'(18184);
			8624: out = 24'(18132);
			8625: out = 24'(18124);
			8626: out = 24'(18100);
			8627: out = 24'(18088);
			8628: out = 24'(18140);
			8629: out = 24'(18116);
			8630: out = 24'(18072);
			8631: out = 24'(17972);
			8632: out = 24'(18040);
			8633: out = 24'(18012);
			8634: out = 24'(17928);
			8635: out = 24'(17988);
			8636: out = 24'(17924);
			8637: out = 24'(17996);
			8638: out = 24'(17852);
			8639: out = 24'(17784);
			8640: out = 24'(17780);
			8641: out = 24'(17788);
			8642: out = 24'(17716);
			8643: out = 24'(17692);
			8644: out = 24'(17656);
			8645: out = 24'(17616);
			8646: out = 24'(17500);
			8647: out = 24'(17476);
			8648: out = 24'(17532);
			8649: out = 24'(17388);
			8650: out = 24'(17256);
			8651: out = 24'(17268);
			8652: out = 24'(17204);
			8653: out = 24'(17080);
			8654: out = 24'(16996);
			8655: out = 24'(16936);
			8656: out = 24'(16836);
			8657: out = 24'(16732);
			8658: out = 24'(16720);
			8659: out = 24'(16664);
			8660: out = 24'(16560);
			8661: out = 24'(16480);
			8662: out = 24'(16356);
			8663: out = 24'(16264);
			8664: out = 24'(16208);
			8665: out = 24'(16108);
			8666: out = 24'(15936);
			8667: out = 24'(15836);
			8668: out = 24'(15744);
			8669: out = 24'(15684);
			8670: out = 24'(15560);
			8671: out = 24'(15444);
			8672: out = 24'(15376);
			8673: out = 24'(15232);
			8674: out = 24'(15152);
			8675: out = 24'(14984);
			8676: out = 24'(14904);
			8677: out = 24'(14772);
			8678: out = 24'(14704);
			8679: out = 24'(14560);
			8680: out = 24'(14404);
			8681: out = 24'(14296);
			8682: out = 24'(14224);
			8683: out = 24'(14080);
			8684: out = 24'(13996);
			8685: out = 24'(13792);
			8686: out = 24'(13668);
			8687: out = 24'(13576);
			8688: out = 24'(13512);
			8689: out = 24'(13356);
			8690: out = 24'(13240);
			8691: out = 24'(13112);
			8692: out = 24'(13000);
			8693: out = 24'(12908);
			8694: out = 24'(12740);
			8695: out = 24'(12592);
			8696: out = 24'(12520);
			8697: out = 24'(12360);
			8698: out = 24'(12236);
			8699: out = 24'(12188);
			8700: out = 24'(12052);
			8701: out = 24'(11976);
			8702: out = 24'(11836);
			8703: out = 24'(11696);
			8704: out = 24'(11556);
			8705: out = 24'(11368);
			8706: out = 24'(11340);
			8707: out = 24'(11200);
			8708: out = 24'(11008);
			8709: out = 24'(11016);
			8710: out = 24'(10820);
			8711: out = 24'(10764);
			8712: out = 24'(10568);
			8713: out = 24'(10520);
			8714: out = 24'(10404);
			8715: out = 24'(10232);
			8716: out = 24'(10160);
			8717: out = 24'(10056);
			8718: out = 24'(9964);
			8719: out = 24'(9804);
			8720: out = 24'(9740);
			8721: out = 24'(9600);
			8722: out = 24'(9564);
			8723: out = 24'(9384);
			8724: out = 24'(9268);
			8725: out = 24'(9168);
			8726: out = 24'(9108);
			8727: out = 24'(8924);
			8728: out = 24'(8876);
			8729: out = 24'(8732);
			8730: out = 24'(8656);
			8731: out = 24'(8544);
			8732: out = 24'(8460);
			8733: out = 24'(8368);
			8734: out = 24'(8252);
			8735: out = 24'(8196);
			8736: out = 24'(8008);
			8737: out = 24'(7968);
			8738: out = 24'(7868);
			8739: out = 24'(7788);
			8740: out = 24'(7692);
			8741: out = 24'(7612);
			8742: out = 24'(7472);
			8743: out = 24'(7400);
			8744: out = 24'(7292);
			8745: out = 24'(7248);
			8746: out = 24'(7084);
			8747: out = 24'(7016);
			8748: out = 24'(6900);
			8749: out = 24'(6852);
			8750: out = 24'(6760);
			8751: out = 24'(6708);
			8752: out = 24'(6592);
			8753: out = 24'(6520);
			8754: out = 24'(6444);
			8755: out = 24'(6344);
			8756: out = 24'(6296);
			8757: out = 24'(6220);
			8758: out = 24'(6120);
			8759: out = 24'(6024);
			8760: out = 24'(5932);
			8761: out = 24'(5860);
			8762: out = 24'(5808);
			8763: out = 24'(5660);
			8764: out = 24'(5660);
			8765: out = 24'(5500);
			8766: out = 24'(5492);
			8767: out = 24'(5400);
			8768: out = 24'(5336);
			8769: out = 24'(5240);
			8770: out = 24'(5196);
			8771: out = 24'(5060);
			8772: out = 24'(5036);
			8773: out = 24'(4940);
			8774: out = 24'(4900);
			8775: out = 24'(4824);
			8776: out = 24'(4708);
			8777: out = 24'(4676);
			8778: out = 24'(4604);
			8779: out = 24'(4600);
			8780: out = 24'(4500);
			8781: out = 24'(4424);
			8782: out = 24'(4328);
			8783: out = 24'(4308);
			8784: out = 24'(4228);
			8785: out = 24'(4188);
			8786: out = 24'(4128);
			8787: out = 24'(4060);
			8788: out = 24'(4012);
			8789: out = 24'(3988);
			8790: out = 24'(3852);
			8791: out = 24'(3852);
			8792: out = 24'(3792);
			8793: out = 24'(3668);
			8794: out = 24'(3688);
			8795: out = 24'(3640);
			8796: out = 24'(3572);
			8797: out = 24'(3516);
			8798: out = 24'(3468);
			8799: out = 24'(3424);
			8800: out = 24'(3244);
			8801: out = 24'(3084);
			8802: out = 24'(2896);
			8803: out = 24'(2772);
			8804: out = 24'(2652);
			8805: out = 24'(2496);
			8806: out = 24'(2388);
			8807: out = 24'(2220);
			8808: out = 24'(2140);
			8809: out = 24'(1960);
			8810: out = 24'(1852);
			8811: out = 24'(1684);
			8812: out = 24'(1528);
			8813: out = 24'(1428);
			8814: out = 24'(1316);
			8815: out = 24'(1196);
			8816: out = 24'(1080);
			8817: out = 24'(996);
			8818: out = 24'(796);
			8819: out = 24'(728);
			8820: out = 24'(616);
			8821: out = 24'(444);
			8822: out = 24'(392);
			8823: out = 24'(256);
			8824: out = 24'(148);
			8825: out = 24'(52);
			8826: out = 24'(-36);
			8827: out = 24'(-80);
			8828: out = 24'(-280);
			8829: out = 24'(-336);
			8830: out = 24'(-468);
			8831: out = 24'(-528);
			8832: out = 24'(-624);
			8833: out = 24'(-752);
			8834: out = 24'(-836);
			8835: out = 24'(-964);
			8836: out = 24'(-1028);
			8837: out = 24'(-1144);
			8838: out = 24'(-1216);
			8839: out = 24'(-1292);
			8840: out = 24'(-1424);
			8841: out = 24'(-1480);
			8842: out = 24'(-1616);
			8843: out = 24'(-1692);
			8844: out = 24'(-1756);
			8845: out = 24'(-1872);
			8846: out = 24'(-1980);
			8847: out = 24'(-2064);
			8848: out = 24'(-2116);
			8849: out = 24'(-2268);
			8850: out = 24'(-2288);
			8851: out = 24'(-2440);
			8852: out = 24'(-2484);
			8853: out = 24'(-2552);
			8854: out = 24'(-2720);
			8855: out = 24'(-2708);
			8856: out = 24'(-2828);
			8857: out = 24'(-2908);
			8858: out = 24'(-3036);
			8859: out = 24'(-3060);
			8860: out = 24'(-3192);
			8861: out = 24'(-3252);
			8862: out = 24'(-3324);
			8863: out = 24'(-3444);
			8864: out = 24'(-3488);
			8865: out = 24'(-3576);
			8866: out = 24'(-3664);
			8867: out = 24'(-3724);
			8868: out = 24'(-3836);
			8869: out = 24'(-3900);
			8870: out = 24'(-3992);
			8871: out = 24'(-4056);
			8872: out = 24'(-4144);
			8873: out = 24'(-4220);
			8874: out = 24'(-4308);
			8875: out = 24'(-4436);
			8876: out = 24'(-4464);
			8877: out = 24'(-4616);
			8878: out = 24'(-4632);
			8879: out = 24'(-4748);
			8880: out = 24'(-4884);
			8881: out = 24'(-4940);
			8882: out = 24'(-5072);
			8883: out = 24'(-5136);
			8884: out = 24'(-5224);
			8885: out = 24'(-5320);
			8886: out = 24'(-5400);
			8887: out = 24'(-5444);
			8888: out = 24'(-5576);
			8889: out = 24'(-5672);
			8890: out = 24'(-5812);
			8891: out = 24'(-5908);
			8892: out = 24'(-6020);
			8893: out = 24'(-6108);
			8894: out = 24'(-6260);
			8895: out = 24'(-6316);
			8896: out = 24'(-6400);
			8897: out = 24'(-6584);
			8898: out = 24'(-6612);
			8899: out = 24'(-6748);
			8900: out = 24'(-6868);
			8901: out = 24'(-7020);
			8902: out = 24'(-7096);
			8903: out = 24'(-7208);
			8904: out = 24'(-7360);
			8905: out = 24'(-7460);
			8906: out = 24'(-7576);
			8907: out = 24'(-7732);
			8908: out = 24'(-7876);
			8909: out = 24'(-8004);
			8910: out = 24'(-8120);
			8911: out = 24'(-8204);
			8912: out = 24'(-8356);
			8913: out = 24'(-8500);
			8914: out = 24'(-8624);
			8915: out = 24'(-8816);
			8916: out = 24'(-8920);
			8917: out = 24'(-9080);
			8918: out = 24'(-9224);
			8919: out = 24'(-9424);
			8920: out = 24'(-9536);
			8921: out = 24'(-9732);
			8922: out = 24'(-9884);
			8923: out = 24'(-10044);
			8924: out = 24'(-10228);
			8925: out = 24'(-10380);
			8926: out = 24'(-10520);
			8927: out = 24'(-10700);
			8928: out = 24'(-10892);
			8929: out = 24'(-11000);
			8930: out = 24'(-11180);
			8931: out = 24'(-11388);
			8932: out = 24'(-11540);
			8933: out = 24'(-11716);
			8934: out = 24'(-11856);
			8935: out = 24'(-12016);
			8936: out = 24'(-12192);
			8937: out = 24'(-12384);
			8938: out = 24'(-12504);
			8939: out = 24'(-12680);
			8940: out = 24'(-12856);
			8941: out = 24'(-12984);
			8942: out = 24'(-13128);
			8943: out = 24'(-13340);
			8944: out = 24'(-13448);
			8945: out = 24'(-13564);
			8946: out = 24'(-13784);
			8947: out = 24'(-13884);
			8948: out = 24'(-13996);
			8949: out = 24'(-14180);
			8950: out = 24'(-14336);
			8951: out = 24'(-14472);
			8952: out = 24'(-14560);
			8953: out = 24'(-14724);
			8954: out = 24'(-14900);
			8955: out = 24'(-14980);
			8956: out = 24'(-15116);
			8957: out = 24'(-15232);
			8958: out = 24'(-15340);
			8959: out = 24'(-15500);
			8960: out = 24'(-15560);
			8961: out = 24'(-15700);
			8962: out = 24'(-15852);
			8963: out = 24'(-15876);
			8964: out = 24'(-16040);
			8965: out = 24'(-16096);
			8966: out = 24'(-16236);
			8967: out = 24'(-16320);
			8968: out = 24'(-16384);
			8969: out = 24'(-16476);
			8970: out = 24'(-16596);
			8971: out = 24'(-16628);
			8972: out = 24'(-16712);
			8973: out = 24'(-16820);
			8974: out = 24'(-16912);
			8975: out = 24'(-16904);
			8976: out = 24'(-17060);
			8977: out = 24'(-17068);
			8978: out = 24'(-17192);
			8979: out = 24'(-17212);
			8980: out = 24'(-17372);
			8981: out = 24'(-17320);
			8982: out = 24'(-17452);
			8983: out = 24'(-17500);
			8984: out = 24'(-17524);
			8985: out = 24'(-17568);
			8986: out = 24'(-17600);
			8987: out = 24'(-17708);
			8988: out = 24'(-17736);
			8989: out = 24'(-17764);
			8990: out = 24'(-17812);
			8991: out = 24'(-17860);
			8992: out = 24'(-17900);
			8993: out = 24'(-17920);
			8994: out = 24'(-17960);
			8995: out = 24'(-18008);
			8996: out = 24'(-18052);
			8997: out = 24'(-18068);
			8998: out = 24'(-18092);
			8999: out = 24'(-18112);
			9000: out = 24'(-18092);
			9001: out = 24'(-18184);
			9002: out = 24'(-18168);
			9003: out = 24'(-18160);
			9004: out = 24'(-18236);
			9005: out = 24'(-18180);
			9006: out = 24'(-18228);
			9007: out = 24'(-18312);
			9008: out = 24'(-18248);
			9009: out = 24'(-18304);
			9010: out = 24'(-18248);
			9011: out = 24'(-18324);
			9012: out = 24'(-18300);
			9013: out = 24'(-18332);
			9014: out = 24'(-18280);
			9015: out = 24'(-18360);
			9016: out = 24'(-18284);
			9017: out = 24'(-18332);
			9018: out = 24'(-18324);
			9019: out = 24'(-18308);
			9020: out = 24'(-18360);
			9021: out = 24'(-18296);
			9022: out = 24'(-18284);
			9023: out = 24'(-18332);
			9024: out = 24'(-18296);
			9025: out = 24'(-18236);
			9026: out = 24'(-18332);
			9027: out = 24'(-18252);
			9028: out = 24'(-18216);
			9029: out = 24'(-18284);
			9030: out = 24'(-18256);
			9031: out = 24'(-18188);
			9032: out = 24'(-18232);
			9033: out = 24'(-18188);
			9034: out = 24'(-18184);
			9035: out = 24'(-18136);
			9036: out = 24'(-18124);
			9037: out = 24'(-18140);
			9038: out = 24'(-18104);
			9039: out = 24'(-18072);
			9040: out = 24'(-18028);
			9041: out = 24'(-18064);
			9042: out = 24'(-18028);
			9043: out = 24'(-17988);
			9044: out = 24'(-17964);
			9045: out = 24'(-17920);
			9046: out = 24'(-17964);
			9047: out = 24'(-17884);
			9048: out = 24'(-17840);
			9049: out = 24'(-17824);
			9050: out = 24'(-17820);
			9051: out = 24'(-17736);
			9052: out = 24'(-17740);
			9053: out = 24'(-17724);
			9054: out = 24'(-17688);
			9055: out = 24'(-17648);
			9056: out = 24'(-17620);
			9057: out = 24'(-17552);
			9058: out = 24'(-17532);
			9059: out = 24'(-17516);
			9060: out = 24'(-17480);
			9061: out = 24'(-17428);
			9062: out = 24'(-17428);
			9063: out = 24'(-17332);
			9064: out = 24'(-17380);
			9065: out = 24'(-17344);
			9066: out = 24'(-17240);
			9067: out = 24'(-17240);
			9068: out = 24'(-17156);
			9069: out = 24'(-17152);
			9070: out = 24'(-17076);
			9071: out = 24'(-17036);
			9072: out = 24'(-17016);
			9073: out = 24'(-16956);
			9074: out = 24'(-16892);
			9075: out = 24'(-16832);
			9076: out = 24'(-16820);
			9077: out = 24'(-16812);
			9078: out = 24'(-16736);
			9079: out = 24'(-16696);
			9080: out = 24'(-16688);
			9081: out = 24'(-16608);
			9082: out = 24'(-16580);
			9083: out = 24'(-16488);
			9084: out = 24'(-16468);
			9085: out = 24'(-16428);
			9086: out = 24'(-16384);
			9087: out = 24'(-16308);
			9088: out = 24'(-16256);
			9089: out = 24'(-16192);
			9090: out = 24'(-16160);
			9091: out = 24'(-16084);
			9092: out = 24'(-16040);
			9093: out = 24'(-15992);
			9094: out = 24'(-15928);
			9095: out = 24'(-15832);
			9096: out = 24'(-15812);
			9097: out = 24'(-15748);
			9098: out = 24'(-15660);
			9099: out = 24'(-15628);
			9100: out = 24'(-15544);
			9101: out = 24'(-15464);
			9102: out = 24'(-15400);
			9103: out = 24'(-15312);
			9104: out = 24'(-15216);
			9105: out = 24'(-15164);
			9106: out = 24'(-15084);
			9107: out = 24'(-15000);
			9108: out = 24'(-14924);
			9109: out = 24'(-14864);
			9110: out = 24'(-14764);
			9111: out = 24'(-14664);
			9112: out = 24'(-14588);
			9113: out = 24'(-14460);
			9114: out = 24'(-14380);
			9115: out = 24'(-14268);
			9116: out = 24'(-14196);
			9117: out = 24'(-14072);
			9118: out = 24'(-13972);
			9119: out = 24'(-13864);
			9120: out = 24'(-13768);
			9121: out = 24'(-13656);
			9122: out = 24'(-13560);
			9123: out = 24'(-13416);
			9124: out = 24'(-13296);
			9125: out = 24'(-13200);
			9126: out = 24'(-13072);
			9127: out = 24'(-12936);
			9128: out = 24'(-12848);
			9129: out = 24'(-12716);
			9130: out = 24'(-12576);
			9131: out = 24'(-12464);
			9132: out = 24'(-12376);
			9133: out = 24'(-12204);
			9134: out = 24'(-12108);
			9135: out = 24'(-11940);
			9136: out = 24'(-11840);
			9137: out = 24'(-11704);
			9138: out = 24'(-11588);
			9139: out = 24'(-11424);
			9140: out = 24'(-11344);
			9141: out = 24'(-11188);
			9142: out = 24'(-11068);
			9143: out = 24'(-10952);
			9144: out = 24'(-10800);
			9145: out = 24'(-10720);
			9146: out = 24'(-10568);
			9147: out = 24'(-10404);
			9148: out = 24'(-10284);
			9149: out = 24'(-10160);
			9150: out = 24'(-9972);
			9151: out = 24'(-9936);
			9152: out = 24'(-9764);
			9153: out = 24'(-9688);
			9154: out = 24'(-9532);
			9155: out = 24'(-9408);
			9156: out = 24'(-9332);
			9157: out = 24'(-9152);
			9158: out = 24'(-9076);
			9159: out = 24'(-8916);
			9160: out = 24'(-8844);
			9161: out = 24'(-8668);
			9162: out = 24'(-8588);
			9163: out = 24'(-8432);
			9164: out = 24'(-8364);
			9165: out = 24'(-8244);
			9166: out = 24'(-8116);
			9167: out = 24'(-8000);
			9168: out = 24'(-7920);
			9169: out = 24'(-7788);
			9170: out = 24'(-7644);
			9171: out = 24'(-7556);
			9172: out = 24'(-7448);
			9173: out = 24'(-7360);
			9174: out = 24'(-7224);
			9175: out = 24'(-7120);
			9176: out = 24'(-7060);
			9177: out = 24'(-6896);
			9178: out = 24'(-6832);
			9179: out = 24'(-6740);
			9180: out = 24'(-6600);
			9181: out = 24'(-6512);
			9182: out = 24'(-6432);
			9183: out = 24'(-6284);
			9184: out = 24'(-6212);
			9185: out = 24'(-6172);
			9186: out = 24'(-6036);
			9187: out = 24'(-5944);
			9188: out = 24'(-5864);
			9189: out = 24'(-5740);
			9190: out = 24'(-5668);
			9191: out = 24'(-5592);
			9192: out = 24'(-5476);
			9193: out = 24'(-5428);
			9194: out = 24'(-5304);
			9195: out = 24'(-5236);
			9196: out = 24'(-5192);
			9197: out = 24'(-5036);
			9198: out = 24'(-5020);
			9199: out = 24'(-4908);
			9200: out = 24'(-4820);
			9201: out = 24'(-4760);
			9202: out = 24'(-4628);
			9203: out = 24'(-4608);
			9204: out = 24'(-4524);
			9205: out = 24'(-4408);
			9206: out = 24'(-4344);
			9207: out = 24'(-4356);
			9208: out = 24'(-4184);
			9209: out = 24'(-4172);
			9210: out = 24'(-4012);
			9211: out = 24'(-4044);
			9212: out = 24'(-3916);
			9213: out = 24'(-3820);
			9214: out = 24'(-3824);
			9215: out = 24'(-3724);
			9216: out = 24'(-3680);
			9217: out = 24'(-3560);
			9218: out = 24'(-3540);
			9219: out = 24'(-3440);
			9220: out = 24'(-3416);
			9221: out = 24'(-3296);
			9222: out = 24'(-3288);
			9223: out = 24'(-3224);
			9224: out = 24'(-3104);
			9225: out = 24'(-2964);
			9226: out = 24'(-2900);
			9227: out = 24'(-2772);
			9228: out = 24'(-2644);
			9229: out = 24'(-2568);
			9230: out = 24'(-2452);
			9231: out = 24'(-2372);
			9232: out = 24'(-2280);
			9233: out = 24'(-2156);
			9234: out = 24'(-2072);
			9235: out = 24'(-2004);
			9236: out = 24'(-1828);
			9237: out = 24'(-1800);
			9238: out = 24'(-1692);
			9239: out = 24'(-1620);
			9240: out = 24'(-1488);
			9241: out = 24'(-1440);
			9242: out = 24'(-1384);
			9243: out = 24'(-1264);
			9244: out = 24'(-1156);
			9245: out = 24'(-1144);
			9246: out = 24'(-1044);
			9247: out = 24'(-908);
			9248: out = 24'(-872);
			9249: out = 24'(-800);
			9250: out = 24'(-772);
			9251: out = 24'(-596);
			9252: out = 24'(-592);
			9253: out = 24'(-504);
			9254: out = 24'(-404);
			9255: out = 24'(-320);
			9256: out = 24'(-280);
			9257: out = 24'(-172);
			9258: out = 24'(-152);
			9259: out = 24'(-36);
			9260: out = 24'(20);
			9261: out = 24'(84);
			9262: out = 24'(136);
			9263: out = 24'(256);
			9264: out = 24'(296);
			9265: out = 24'(356);
			9266: out = 24'(420);
			9267: out = 24'(448);
			9268: out = 24'(536);
			9269: out = 24'(644);
			9270: out = 24'(636);
			9271: out = 24'(748);
			9272: out = 24'(816);
			9273: out = 24'(800);
			9274: out = 24'(908);
			9275: out = 24'(1016);
			9276: out = 24'(1008);
			9277: out = 24'(1096);
			9278: out = 24'(1172);
			9279: out = 24'(1240);
			9280: out = 24'(1264);
			9281: out = 24'(1332);
			9282: out = 24'(1412);
			9283: out = 24'(1436);
			9284: out = 24'(1488);
			9285: out = 24'(1604);
			9286: out = 24'(1612);
			9287: out = 24'(1736);
			9288: out = 24'(1736);
			9289: out = 24'(1788);
			9290: out = 24'(1904);
			9291: out = 24'(1920);
			9292: out = 24'(2008);
			9293: out = 24'(2076);
			9294: out = 24'(2124);
			9295: out = 24'(2116);
			9296: out = 24'(2264);
			9297: out = 24'(2284);
			9298: out = 24'(2344);
			9299: out = 24'(2420);
			9300: out = 24'(2488);
			9301: out = 24'(2532);
			9302: out = 24'(2652);
			9303: out = 24'(2660);
			9304: out = 24'(2772);
			9305: out = 24'(2812);
			9306: out = 24'(2844);
			9307: out = 24'(2956);
			9308: out = 24'(3020);
			9309: out = 24'(3084);
			9310: out = 24'(3140);
			9311: out = 24'(3260);
			9312: out = 24'(3284);
			9313: out = 24'(3396);
			9314: out = 24'(3424);
			9315: out = 24'(3540);
			9316: out = 24'(3604);
			9317: out = 24'(3668);
			9318: out = 24'(3804);
			9319: out = 24'(3816);
			9320: out = 24'(3920);
			9321: out = 24'(4000);
			9322: out = 24'(4136);
			9323: out = 24'(4172);
			9324: out = 24'(4264);
			9325: out = 24'(4384);
			9326: out = 24'(4452);
			9327: out = 24'(4560);
			9328: out = 24'(4660);
			9329: out = 24'(4752);
			9330: out = 24'(4816);
			9331: out = 24'(4956);
			9332: out = 24'(5036);
			9333: out = 24'(5180);
			9334: out = 24'(5240);
			9335: out = 24'(5416);
			9336: out = 24'(5452);
			9337: out = 24'(5620);
			9338: out = 24'(5696);
			9339: out = 24'(5840);
			9340: out = 24'(5900);
			9341: out = 24'(6028);
			9342: out = 24'(6140);
			9343: out = 24'(6252);
			9344: out = 24'(6392);
			9345: out = 24'(6488);
			9346: out = 24'(6628);
			9347: out = 24'(6732);
			9348: out = 24'(6840);
			9349: out = 24'(6968);
			9350: out = 24'(7084);
			9351: out = 24'(7184);
			9352: out = 24'(7340);
			9353: out = 24'(7420);
			9354: out = 24'(7608);
			9355: out = 24'(7656);
			9356: out = 24'(7784);
			9357: out = 24'(7924);
			9358: out = 24'(8004);
			9359: out = 24'(8112);
			9360: out = 24'(8268);
			9361: out = 24'(8364);
			9362: out = 24'(8456);
			9363: out = 24'(8608);
			9364: out = 24'(8672);
			9365: out = 24'(8800);
			9366: out = 24'(8892);
			9367: out = 24'(9016);
			9368: out = 24'(9100);
			9369: out = 24'(9236);
			9370: out = 24'(9300);
			9371: out = 24'(9472);
			9372: out = 24'(9524);
			9373: out = 24'(9596);
			9374: out = 24'(9768);
			9375: out = 24'(9800);
			9376: out = 24'(9924);
			9377: out = 24'(9992);
			9378: out = 24'(10140);
			9379: out = 24'(10212);
			9380: out = 24'(10296);
			9381: out = 24'(10420);
			9382: out = 24'(10484);
			9383: out = 24'(10564);
			9384: out = 24'(10680);
			9385: out = 24'(10752);
			9386: out = 24'(10856);
			9387: out = 24'(10904);
			9388: out = 24'(11008);
			9389: out = 24'(11136);
			9390: out = 24'(11148);
			9391: out = 24'(11244);
			9392: out = 24'(11324);
			9393: out = 24'(11424);
			9394: out = 24'(11484);
			9395: out = 24'(11604);
			9396: out = 24'(11664);
			9397: out = 24'(11728);
			9398: out = 24'(11812);
			9399: out = 24'(11884);
			9400: out = 24'(11936);
			9401: out = 24'(12048);
			9402: out = 24'(12096);
			9403: out = 24'(12196);
			9404: out = 24'(12252);
			9405: out = 24'(12280);
			9406: out = 24'(12408);
			9407: out = 24'(12460);
			9408: out = 24'(12536);
			9409: out = 24'(12580);
			9410: out = 24'(12688);
			9411: out = 24'(12680);
			9412: out = 24'(12844);
			9413: out = 24'(12836);
			9414: out = 24'(12916);
			9415: out = 24'(12964);
			9416: out = 24'(13048);
			9417: out = 24'(13104);
			9418: out = 24'(13168);
			9419: out = 24'(13248);
			9420: out = 24'(13304);
			9421: out = 24'(13372);
			9422: out = 24'(13416);
			9423: out = 24'(13484);
			9424: out = 24'(13504);
			9425: out = 24'(13616);
			9426: out = 24'(13644);
			9427: out = 24'(13704);
			9428: out = 24'(13732);
			9429: out = 24'(13812);
			9430: out = 24'(13876);
			9431: out = 24'(13952);
			9432: out = 24'(13932);
			9433: out = 24'(14052);
			9434: out = 24'(14088);
			9435: out = 24'(14112);
			9436: out = 24'(14208);
			9437: out = 24'(14236);
			9438: out = 24'(14336);
			9439: out = 24'(14324);
			9440: out = 24'(14400);
			9441: out = 24'(14480);
			9442: out = 24'(14488);
			9443: out = 24'(14552);
			9444: out = 24'(14584);
			9445: out = 24'(14632);
			9446: out = 24'(14708);
			9447: out = 24'(14748);
			9448: out = 24'(14772);
			9449: out = 24'(14832);
			9450: out = 24'(14876);
			9451: out = 24'(14944);
			9452: out = 24'(14940);
			9453: out = 24'(15040);
			9454: out = 24'(15080);
			9455: out = 24'(15076);
			9456: out = 24'(15120);
			9457: out = 24'(15172);
			9458: out = 24'(15180);
			9459: out = 24'(15248);
			9460: out = 24'(15252);
			9461: out = 24'(15272);
			9462: out = 24'(15236);
			9463: out = 24'(15152);
			9464: out = 24'(15168);
			9465: out = 24'(15088);
			9466: out = 24'(15148);
			9467: out = 24'(15092);
			9468: out = 24'(15164);
			9469: out = 24'(15168);
			9470: out = 24'(15128);
			9471: out = 24'(15212);
			9472: out = 24'(15092);
			9473: out = 24'(15116);
			9474: out = 24'(15116);
			9475: out = 24'(15176);
			9476: out = 24'(15060);
			9477: out = 24'(15104);
			9478: out = 24'(15088);
			9479: out = 24'(15132);
			9480: out = 24'(15100);
			9481: out = 24'(15100);
			9482: out = 24'(15068);
			9483: out = 24'(15108);
			9484: out = 24'(15108);
			9485: out = 24'(15044);
			9486: out = 24'(15020);
			9487: out = 24'(15048);
			9488: out = 24'(15028);
			9489: out = 24'(14936);
			9490: out = 24'(14992);
			9491: out = 24'(14952);
			9492: out = 24'(15024);
			9493: out = 24'(14976);
			9494: out = 24'(15032);
			9495: out = 24'(14968);
			9496: out = 24'(14980);
			9497: out = 24'(14928);
			9498: out = 24'(14932);
			9499: out = 24'(14988);
			9500: out = 24'(14912);
			9501: out = 24'(14900);
			9502: out = 24'(14980);
			9503: out = 24'(14900);
			9504: out = 24'(14980);
			9505: out = 24'(14820);
			9506: out = 24'(14848);
			9507: out = 24'(14884);
			9508: out = 24'(14944);
			9509: out = 24'(14796);
			9510: out = 24'(14892);
			9511: out = 24'(14876);
			9512: out = 24'(14916);
			9513: out = 24'(14836);
			9514: out = 24'(14792);
			9515: out = 24'(14824);
			9516: out = 24'(14832);
			9517: out = 24'(14828);
			9518: out = 24'(14664);
			9519: out = 24'(14780);
			9520: out = 24'(14744);
			9521: out = 24'(14752);
			9522: out = 24'(14656);
			9523: out = 24'(14668);
			9524: out = 24'(14660);
			9525: out = 24'(14616);
			9526: out = 24'(14696);
			9527: out = 24'(14668);
			9528: out = 24'(14700);
			9529: out = 24'(14564);
			9530: out = 24'(14592);
			9531: out = 24'(14440);
			9532: out = 24'(14428);
			9533: out = 24'(14480);
			9534: out = 24'(14396);
			9535: out = 24'(14316);
			9536: out = 24'(14276);
			9537: out = 24'(14308);
			9538: out = 24'(14176);
			9539: out = 24'(14236);
			9540: out = 24'(14116);
			9541: out = 24'(14084);
			9542: out = 24'(14064);
			9543: out = 24'(13964);
			9544: out = 24'(13980);
			9545: out = 24'(13884);
			9546: out = 24'(13856);
			9547: out = 24'(13844);
			9548: out = 24'(13768);
			9549: out = 24'(13652);
			9550: out = 24'(13580);
			9551: out = 24'(13456);
			9552: out = 24'(13388);
			9553: out = 24'(13332);
			9554: out = 24'(13264);
			9555: out = 24'(13168);
			9556: out = 24'(13096);
			9557: out = 24'(13052);
			9558: out = 24'(12960);
			9559: out = 24'(12900);
			9560: out = 24'(12804);
			9561: out = 24'(12760);
			9562: out = 24'(12640);
			9563: out = 24'(12580);
			9564: out = 24'(12468);
			9565: out = 24'(12312);
			9566: out = 24'(12284);
			9567: out = 24'(12216);
			9568: out = 24'(12128);
			9569: out = 24'(12000);
			9570: out = 24'(11932);
			9571: out = 24'(11816);
			9572: out = 24'(11716);
			9573: out = 24'(11600);
			9574: out = 24'(11476);
			9575: out = 24'(11444);
			9576: out = 24'(11292);
			9577: out = 24'(11224);
			9578: out = 24'(11136);
			9579: out = 24'(11032);
			9580: out = 24'(11004);
			9581: out = 24'(10816);
			9582: out = 24'(10756);
			9583: out = 24'(10616);
			9584: out = 24'(10596);
			9585: out = 24'(10428);
			9586: out = 24'(10352);
			9587: out = 24'(10236);
			9588: out = 24'(10156);
			9589: out = 24'(10004);
			9590: out = 24'(9924);
			9591: out = 24'(9884);
			9592: out = 24'(9784);
			9593: out = 24'(9632);
			9594: out = 24'(9588);
			9595: out = 24'(9440);
			9596: out = 24'(9400);
			9597: out = 24'(9284);
			9598: out = 24'(9188);
			9599: out = 24'(9116);
			9600: out = 24'(9048);
			9601: out = 24'(8856);
			9602: out = 24'(8780);
			9603: out = 24'(8744);
			9604: out = 24'(8548);
			9605: out = 24'(8496);
			9606: out = 24'(8408);
			9607: out = 24'(8324);
			9608: out = 24'(8204);
			9609: out = 24'(8200);
			9610: out = 24'(7964);
			9611: out = 24'(7976);
			9612: out = 24'(7868);
			9613: out = 24'(7776);
			9614: out = 24'(7724);
			9615: out = 24'(7544);
			9616: out = 24'(7516);
			9617: out = 24'(7368);
			9618: out = 24'(7356);
			9619: out = 24'(7228);
			9620: out = 24'(7168);
			9621: out = 24'(7020);
			9622: out = 24'(7028);
			9623: out = 24'(6880);
			9624: out = 24'(6788);
			9625: out = 24'(6740);
			9626: out = 24'(6708);
			9627: out = 24'(6572);
			9628: out = 24'(6428);
			9629: out = 24'(6408);
			9630: out = 24'(6288);
			9631: out = 24'(6228);
			9632: out = 24'(6196);
			9633: out = 24'(6080);
			9634: out = 24'(6040);
			9635: out = 24'(5936);
			9636: out = 24'(5860);
			9637: out = 24'(5848);
			9638: out = 24'(5732);
			9639: out = 24'(5616);
			9640: out = 24'(5608);
			9641: out = 24'(5516);
			9642: out = 24'(5452);
			9643: out = 24'(5404);
			9644: out = 24'(5248);
			9645: out = 24'(5240);
			9646: out = 24'(5200);
			9647: out = 24'(5136);
			9648: out = 24'(5024);
			9649: out = 24'(5020);
			9650: out = 24'(4960);
			9651: out = 24'(4856);
			9652: out = 24'(4840);
			9653: out = 24'(4744);
			9654: out = 24'(4720);
			9655: out = 24'(4620);
			9656: out = 24'(4540);
			9657: out = 24'(4524);
			9658: out = 24'(4388);
			9659: out = 24'(4388);
			9660: out = 24'(4344);
			9661: out = 24'(4264);
			9662: out = 24'(4196);
			9663: out = 24'(4104);
			9664: out = 24'(4140);
			9665: out = 24'(4032);
			9666: out = 24'(3952);
			9667: out = 24'(3972);
			9668: out = 24'(3896);
			9669: out = 24'(3788);
			9670: out = 24'(3752);
			9671: out = 24'(3732);
			9672: out = 24'(3664);
			9673: out = 24'(3556);
			9674: out = 24'(3564);
			9675: out = 24'(3480);
			9676: out = 24'(3448);
			9677: out = 24'(3384);
			9678: out = 24'(3396);
			9679: out = 24'(3308);
			9680: out = 24'(3268);
			9681: out = 24'(3220);
			9682: out = 24'(3120);
			9683: out = 24'(3116);
			9684: out = 24'(3112);
			9685: out = 24'(2952);
			9686: out = 24'(2956);
			9687: out = 24'(2936);
			9688: out = 24'(2860);
			9689: out = 24'(2844);
			9690: out = 24'(2788);
			9691: out = 24'(2668);
			9692: out = 24'(2584);
			9693: out = 24'(2448);
			9694: out = 24'(2320);
			9695: out = 24'(2236);
			9696: out = 24'(2076);
			9697: out = 24'(1968);
			9698: out = 24'(1876);
			9699: out = 24'(1740);
			9700: out = 24'(1636);
			9701: out = 24'(1544);
			9702: out = 24'(1456);
			9703: out = 24'(1328);
			9704: out = 24'(1272);
			9705: out = 24'(1148);
			9706: out = 24'(1056);
			9707: out = 24'(904);
			9708: out = 24'(888);
			9709: out = 24'(728);
			9710: out = 24'(644);
			9711: out = 24'(548);
			9712: out = 24'(484);
			9713: out = 24'(364);
			9714: out = 24'(256);
			9715: out = 24'(176);
			9716: out = 24'(64);
			9717: out = 24'(24);
			9718: out = 24'(-76);
			9719: out = 24'(-168);
			9720: out = 24'(-248);
			9721: out = 24'(-352);
			9722: out = 24'(-448);
			9723: out = 24'(-508);
			9724: out = 24'(-548);
			9725: out = 24'(-712);
			9726: out = 24'(-764);
			9727: out = 24'(-844);
			9728: out = 24'(-948);
			9729: out = 24'(-1012);
			9730: out = 24'(-1036);
			9731: out = 24'(-1152);
			9732: out = 24'(-1204);
			9733: out = 24'(-1320);
			9734: out = 24'(-1388);
			9735: out = 24'(-1424);
			9736: out = 24'(-1536);
			9737: out = 24'(-1604);
			9738: out = 24'(-1700);
			9739: out = 24'(-1740);
			9740: out = 24'(-1824);
			9741: out = 24'(-1864);
			9742: out = 24'(-1964);
			9743: out = 24'(-2008);
			9744: out = 24'(-2088);
			9745: out = 24'(-2168);
			9746: out = 24'(-2216);
			9747: out = 24'(-2304);
			9748: out = 24'(-2368);
			9749: out = 24'(-2468);
			9750: out = 24'(-2516);
			9751: out = 24'(-2572);
			9752: out = 24'(-2656);
			9753: out = 24'(-2704);
			9754: out = 24'(-2752);
			9755: out = 24'(-2892);
			9756: out = 24'(-2888);
			9757: out = 24'(-3016);
			9758: out = 24'(-3036);
			9759: out = 24'(-3128);
			9760: out = 24'(-3172);
			9761: out = 24'(-3280);
			9762: out = 24'(-3336);
			9763: out = 24'(-3436);
			9764: out = 24'(-3436);
			9765: out = 24'(-3528);
			9766: out = 24'(-3628);
			9767: out = 24'(-3680);
			9768: out = 24'(-3752);
			9769: out = 24'(-3808);
			9770: out = 24'(-3848);
			9771: out = 24'(-3948);
			9772: out = 24'(-4072);
			9773: out = 24'(-4092);
			9774: out = 24'(-4196);
			9775: out = 24'(-4280);
			9776: out = 24'(-4340);
			9777: out = 24'(-4396);
			9778: out = 24'(-4484);
			9779: out = 24'(-4576);
			9780: out = 24'(-4664);
			9781: out = 24'(-4728);
			9782: out = 24'(-4788);
			9783: out = 24'(-4900);
			9784: out = 24'(-4936);
			9785: out = 24'(-4992);
			9786: out = 24'(-5168);
			9787: out = 24'(-5180);
			9788: out = 24'(-5352);
			9789: out = 24'(-5432);
			9790: out = 24'(-5568);
			9791: out = 24'(-5616);
			9792: out = 24'(-5700);
			9793: out = 24'(-5864);
			9794: out = 24'(-5888);
			9795: out = 24'(-5988);
			9796: out = 24'(-6100);
			9797: out = 24'(-6232);
			9798: out = 24'(-6316);
			9799: out = 24'(-6440);
			9800: out = 24'(-6548);
			9801: out = 24'(-6648);
			9802: out = 24'(-6776);
			9803: out = 24'(-6868);
			9804: out = 24'(-6992);
			9805: out = 24'(-7116);
			9806: out = 24'(-7216);
			9807: out = 24'(-7316);
			9808: out = 24'(-7488);
			9809: out = 24'(-7584);
			9810: out = 24'(-7696);
			9811: out = 24'(-7840);
			9812: out = 24'(-7968);
			9813: out = 24'(-8100);
			9814: out = 24'(-8228);
			9815: out = 24'(-8352);
			9816: out = 24'(-8440);
			9817: out = 24'(-8684);
			9818: out = 24'(-8720);
			9819: out = 24'(-8904);
			9820: out = 24'(-9032);
			9821: out = 24'(-9148);
			9822: out = 24'(-9296);
			9823: out = 24'(-9412);
			9824: out = 24'(-9600);
			9825: out = 24'(-9724);
			9826: out = 24'(-9872);
			9827: out = 24'(-9976);
			9828: out = 24'(-10164);
			9829: out = 24'(-10220);
			9830: out = 24'(-10404);
			9831: out = 24'(-10524);
			9832: out = 24'(-10632);
			9833: out = 24'(-10796);
			9834: out = 24'(-10900);
			9835: out = 24'(-11032);
			9836: out = 24'(-11160);
			9837: out = 24'(-11304);
			9838: out = 24'(-11416);
			9839: out = 24'(-11508);
			9840: out = 24'(-11628);
			9841: out = 24'(-11768);
			9842: out = 24'(-11820);
			9843: out = 24'(-11992);
			9844: out = 24'(-12064);
			9845: out = 24'(-12172);
			9846: out = 24'(-12308);
			9847: out = 24'(-12388);
			9848: out = 24'(-12492);
			9849: out = 24'(-12592);
			9850: out = 24'(-12660);
			9851: out = 24'(-12792);
			9852: out = 24'(-12852);
			9853: out = 24'(-12944);
			9854: out = 24'(-13052);
			9855: out = 24'(-13104);
			9856: out = 24'(-13192);
			9857: out = 24'(-13324);
			9858: out = 24'(-13332);
			9859: out = 24'(-13432);
			9860: out = 24'(-13484);
			9861: out = 24'(-13580);
			9862: out = 24'(-13684);
			9863: out = 24'(-13664);
			9864: out = 24'(-13792);
			9865: out = 24'(-13880);
			9866: out = 24'(-13884);
			9867: out = 24'(-13956);
			9868: out = 24'(-13980);
			9869: out = 24'(-14028);
			9870: out = 24'(-14148);
			9871: out = 24'(-14144);
			9872: out = 24'(-14236);
			9873: out = 24'(-14296);
			9874: out = 24'(-14348);
			9875: out = 24'(-14348);
			9876: out = 24'(-14444);
			9877: out = 24'(-14424);
			9878: out = 24'(-14512);
			9879: out = 24'(-14520);
			9880: out = 24'(-14560);
			9881: out = 24'(-14620);
			9882: out = 24'(-14628);
			9883: out = 24'(-14660);
			9884: out = 24'(-14724);
			9885: out = 24'(-14708);
			9886: out = 24'(-14780);
			9887: out = 24'(-14788);
			9888: out = 24'(-14792);
			9889: out = 24'(-14824);
			9890: out = 24'(-14832);
			9891: out = 24'(-14888);
			9892: out = 24'(-14876);
			9893: out = 24'(-14920);
			9894: out = 24'(-14896);
			9895: out = 24'(-14928);
			9896: out = 24'(-14936);
			9897: out = 24'(-14960);
			9898: out = 24'(-14964);
			9899: out = 24'(-14944);
			9900: out = 24'(-14944);
			9901: out = 24'(-14988);
			9902: out = 24'(-14984);
			9903: out = 24'(-14992);
			9904: out = 24'(-14988);
			9905: out = 24'(-15016);
			9906: out = 24'(-15012);
			9907: out = 24'(-14968);
			9908: out = 24'(-14984);
			9909: out = 24'(-15008);
			9910: out = 24'(-14988);
			9911: out = 24'(-14992);
			9912: out = 24'(-14964);
			9913: out = 24'(-14996);
			9914: out = 24'(-15020);
			9915: out = 24'(-14976);
			9916: out = 24'(-14984);
			9917: out = 24'(-14948);
			9918: out = 24'(-14932);
			9919: out = 24'(-14976);
			9920: out = 24'(-14924);
			9921: out = 24'(-14912);
			9922: out = 24'(-14940);
			9923: out = 24'(-14888);
			9924: out = 24'(-14880);
			9925: out = 24'(-14844);
			9926: out = 24'(-14900);
			9927: out = 24'(-14844);
			9928: out = 24'(-14828);
			9929: out = 24'(-14808);
			9930: out = 24'(-14784);
			9931: out = 24'(-14760);
			9932: out = 24'(-14788);
			9933: out = 24'(-14696);
			9934: out = 24'(-14744);
			9935: out = 24'(-14676);
			9936: out = 24'(-14664);
			9937: out = 24'(-14684);
			9938: out = 24'(-14616);
			9939: out = 24'(-14600);
			9940: out = 24'(-14608);
			9941: out = 24'(-14548);
			9942: out = 24'(-14540);
			9943: out = 24'(-14492);
			9944: out = 24'(-14544);
			9945: out = 24'(-14460);
			9946: out = 24'(-14424);
			9947: out = 24'(-14404);
			9948: out = 24'(-14352);
			9949: out = 24'(-14396);
			9950: out = 24'(-14312);
			9951: out = 24'(-14280);
			9952: out = 24'(-14272);
			9953: out = 24'(-14228);
			9954: out = 24'(-14196);
			9955: out = 24'(-14160);
			9956: out = 24'(-14176);
			9957: out = 24'(-14112);
			9958: out = 24'(-14068);
			9959: out = 24'(-14080);
			9960: out = 24'(-14004);
			9961: out = 24'(-14000);
			9962: out = 24'(-13980);
			9963: out = 24'(-13928);
			9964: out = 24'(-13908);
			9965: out = 24'(-13860);
			9966: out = 24'(-13852);
			9967: out = 24'(-13732);
			9968: out = 24'(-13740);
			9969: out = 24'(-13740);
			9970: out = 24'(-13652);
			9971: out = 24'(-13612);
			9972: out = 24'(-13588);
			9973: out = 24'(-13576);
			9974: out = 24'(-13496);
			9975: out = 24'(-13500);
			9976: out = 24'(-13408);
			9977: out = 24'(-13400);
			9978: out = 24'(-13332);
			9979: out = 24'(-13324);
			9980: out = 24'(-13232);
			9981: out = 24'(-13248);
			9982: out = 24'(-13152);
			9983: out = 24'(-13096);
			9984: out = 24'(-13112);
			9985: out = 24'(-12988);
			9986: out = 24'(-13020);
			9987: out = 24'(-12900);
			9988: out = 24'(-12892);
			9989: out = 24'(-12788);
			9990: out = 24'(-12796);
			9991: out = 24'(-12748);
			9992: out = 24'(-12640);
			9993: out = 24'(-12612);
			9994: out = 24'(-12528);
			9995: out = 24'(-12488);
			9996: out = 24'(-12384);
			9997: out = 24'(-12376);
			9998: out = 24'(-12244);
			9999: out = 24'(-12236);
			10000: out = 24'(-12120);
			10001: out = 24'(-12100);
			10002: out = 24'(-12000);
			10003: out = 24'(-11952);
			10004: out = 24'(-11876);
			10005: out = 24'(-11800);
			10006: out = 24'(-11684);
			10007: out = 24'(-11624);
			10008: out = 24'(-11528);
			10009: out = 24'(-11456);
			10010: out = 24'(-11372);
			10011: out = 24'(-11288);
			10012: out = 24'(-11180);
			10013: out = 24'(-11132);
			10014: out = 24'(-11004);
			10015: out = 24'(-10920);
			10016: out = 24'(-10840);
			10017: out = 24'(-10672);
			10018: out = 24'(-10672);
			10019: out = 24'(-10524);
			10020: out = 24'(-10424);
			10021: out = 24'(-10308);
			10022: out = 24'(-10240);
			10023: out = 24'(-10112);
			10024: out = 24'(-10028);
			10025: out = 24'(-9896);
			10026: out = 24'(-9828);
			10027: out = 24'(-9736);
			10028: out = 24'(-9544);
			10029: out = 24'(-9516);
			10030: out = 24'(-9420);
			10031: out = 24'(-9268);
			10032: out = 24'(-9176);
			10033: out = 24'(-9084);
			10034: out = 24'(-8952);
			10035: out = 24'(-8876);
			10036: out = 24'(-8772);
			10037: out = 24'(-8664);
			10038: out = 24'(-8524);
			10039: out = 24'(-8484);
			10040: out = 24'(-8340);
			10041: out = 24'(-8220);
			10042: out = 24'(-8160);
			10043: out = 24'(-8012);
			10044: out = 24'(-7944);
			10045: out = 24'(-7860);
			10046: out = 24'(-7688);
			10047: out = 24'(-7604);
			10048: out = 24'(-7496);
			10049: out = 24'(-7432);
			10050: out = 24'(-7324);
			10051: out = 24'(-7236);
			10052: out = 24'(-7156);
			10053: out = 24'(-7012);
			10054: out = 24'(-6960);
			10055: out = 24'(-6848);
			10056: out = 24'(-6760);
			10057: out = 24'(-6696);
			10058: out = 24'(-6556);
			10059: out = 24'(-6472);
			10060: out = 24'(-6416);
			10061: out = 24'(-6284);
			10062: out = 24'(-6196);
			10063: out = 24'(-6136);
			10064: out = 24'(-6020);
			10065: out = 24'(-5948);
			10066: out = 24'(-5860);
			10067: out = 24'(-5784);
			10068: out = 24'(-5664);
			10069: out = 24'(-5636);
			10070: out = 24'(-5476);
			10071: out = 24'(-5452);
			10072: out = 24'(-5376);
			10073: out = 24'(-5276);
			10074: out = 24'(-5176);
			10075: out = 24'(-5072);
			10076: out = 24'(-5080);
			10077: out = 24'(-4948);
			10078: out = 24'(-4876);
			10079: out = 24'(-4796);
			10080: out = 24'(-4752);
			10081: out = 24'(-4652);
			10082: out = 24'(-4604);
			10083: out = 24'(-4492);
			10084: out = 24'(-4428);
			10085: out = 24'(-4384);
			10086: out = 24'(-4272);
			10087: out = 24'(-4236);
			10088: out = 24'(-4152);
			10089: out = 24'(-4108);
			10090: out = 24'(-4024);
			10091: out = 24'(-3964);
			10092: out = 24'(-3872);
			10093: out = 24'(-3816);
			10094: out = 24'(-3768);
			10095: out = 24'(-3672);
			10096: out = 24'(-3668);
			10097: out = 24'(-3532);
			10098: out = 24'(-3556);
			10099: out = 24'(-3440);
			10100: out = 24'(-3416);
			10101: out = 24'(-3308);
			10102: out = 24'(-3288);
			10103: out = 24'(-3232);
			10104: out = 24'(-3156);
			10105: out = 24'(-3100);
			10106: out = 24'(-3056);
			10107: out = 24'(-3036);
			10108: out = 24'(-2940);
			10109: out = 24'(-2852);
			10110: out = 24'(-2820);
			10111: out = 24'(-2824);
			10112: out = 24'(-2728);
			10113: out = 24'(-2688);
			10114: out = 24'(-2616);
			10115: out = 24'(-2568);
			10116: out = 24'(-2432);
			10117: out = 24'(-2404);
			10118: out = 24'(-2280);
			10119: out = 24'(-2160);
			10120: out = 24'(-2124);
			10121: out = 24'(-2012);
			10122: out = 24'(-1960);
			10123: out = 24'(-1836);
			10124: out = 24'(-1828);
			10125: out = 24'(-1692);
			10126: out = 24'(-1644);
			10127: out = 24'(-1532);
			10128: out = 24'(-1492);
			10129: out = 24'(-1396);
			10130: out = 24'(-1352);
			10131: out = 24'(-1208);
			10132: out = 24'(-1212);
			10133: out = 24'(-1144);
			10134: out = 24'(-1048);
			10135: out = 24'(-960);
			10136: out = 24'(-932);
			10137: out = 24'(-844);
			10138: out = 24'(-768);
			10139: out = 24'(-752);
			10140: out = 24'(-664);
			10141: out = 24'(-540);
			10142: out = 24'(-584);
			10143: out = 24'(-440);
			10144: out = 24'(-416);
			10145: out = 24'(-320);
			10146: out = 24'(-304);
			10147: out = 24'(-240);
			10148: out = 24'(-228);
			10149: out = 24'(-104);
			10150: out = 24'(-56);
			10151: out = 24'(4);
			10152: out = 24'(72);
			10153: out = 24'(80);
			10154: out = 24'(152);
			10155: out = 24'(228);
			10156: out = 24'(288);
			10157: out = 24'(332);
			10158: out = 24'(348);
			10159: out = 24'(448);
			10160: out = 24'(496);
			10161: out = 24'(544);
			10162: out = 24'(564);
			10163: out = 24'(664);
			10164: out = 24'(672);
			10165: out = 24'(740);
			10166: out = 24'(796);
			10167: out = 24'(836);
			10168: out = 24'(868);
			10169: out = 24'(976);
			10170: out = 24'(956);
			10171: out = 24'(1052);
			10172: out = 24'(1068);
			10173: out = 24'(1144);
			10174: out = 24'(1204);
			10175: out = 24'(1212);
			10176: out = 24'(1284);
			10177: out = 24'(1344);
			10178: out = 24'(1396);
			10179: out = 24'(1428);
			10180: out = 24'(1484);
			10181: out = 24'(1544);
			10182: out = 24'(1564);
			10183: out = 24'(1624);
			10184: out = 24'(1664);
			10185: out = 24'(1768);
			10186: out = 24'(1728);
			10187: out = 24'(1836);
			10188: out = 24'(1880);
			10189: out = 24'(1920);
			10190: out = 24'(2000);
			10191: out = 24'(2044);
			10192: out = 24'(2124);
			10193: out = 24'(2120);
			10194: out = 24'(2204);
			10195: out = 24'(2240);
			10196: out = 24'(2308);
			10197: out = 24'(2368);
			10198: out = 24'(2376);
			10199: out = 24'(2468);
			10200: out = 24'(2560);
			10201: out = 24'(2564);
			10202: out = 24'(2656);
			10203: out = 24'(2712);
			10204: out = 24'(2768);
			10205: out = 24'(2800);
			10206: out = 24'(2896);
			10207: out = 24'(2952);
			10208: out = 24'(2988);
			10209: out = 24'(3112);
			10210: out = 24'(3100);
			10211: out = 24'(3228);
			10212: out = 24'(3296);
			10213: out = 24'(3356);
			10214: out = 24'(3460);
			10215: out = 24'(3456);
			10216: out = 24'(3616);
			10217: out = 24'(3640);
			10218: out = 24'(3728);
			10219: out = 24'(3780);
			10220: out = 24'(3944);
			10221: out = 24'(3924);
			10222: out = 24'(4048);
			10223: out = 24'(4148);
			10224: out = 24'(4228);
			10225: out = 24'(4300);
			10226: out = 24'(4392);
			10227: out = 24'(4516);
			10228: out = 24'(4528);
			10229: out = 24'(4696);
			10230: out = 24'(4748);
			10231: out = 24'(4824);
			10232: out = 24'(4964);
			10233: out = 24'(5032);
			10234: out = 24'(5168);
			10235: out = 24'(5200);
			10236: out = 24'(5308);
			10237: out = 24'(5380);
			10238: out = 24'(5544);
			10239: out = 24'(5580);
			10240: out = 24'(5704);
			10241: out = 24'(5776);
			10242: out = 24'(5876);
			10243: out = 24'(5968);
			10244: out = 24'(6012);
			10245: out = 24'(6148);
			10246: out = 24'(6236);
			10247: out = 24'(6324);
			10248: out = 24'(6432);
			10249: out = 24'(6512);
			10250: out = 24'(6656);
			10251: out = 24'(6668);
			10252: out = 24'(6784);
			10253: out = 24'(6880);
			10254: out = 24'(6992);
			10255: out = 24'(7036);
			10256: out = 24'(7176);
			10257: out = 24'(7228);
			10258: out = 24'(7352);
			10259: out = 24'(7376);
			10260: out = 24'(7484);
			10261: out = 24'(7600);
			10262: out = 24'(7660);
			10263: out = 24'(7732);
			10264: out = 24'(7816);
			10265: out = 24'(7936);
			10266: out = 24'(7928);
			10267: out = 24'(8096);
			10268: out = 24'(8120);
			10269: out = 24'(8212);
			10270: out = 24'(8308);
			10271: out = 24'(8336);
			10272: out = 24'(8408);
			10273: out = 24'(8532);
			10274: out = 24'(8600);
			10275: out = 24'(8684);
			10276: out = 24'(8700);
			10277: out = 24'(8812);
			10278: out = 24'(8892);
			10279: out = 24'(8892);
			10280: out = 24'(9028);
			10281: out = 24'(9044);
			10282: out = 24'(9148);
			10283: out = 24'(9200);
			10284: out = 24'(9260);
			10285: out = 24'(9376);
			10286: out = 24'(9396);
			10287: out = 24'(9460);
			10288: out = 24'(9544);
			10289: out = 24'(9600);
			10290: out = 24'(9640);
			10291: out = 24'(9724);
			10292: out = 24'(9784);
			10293: out = 24'(9812);
			10294: out = 24'(9876);
			10295: out = 24'(9924);
			10296: out = 24'(10008);
			10297: out = 24'(10056);
			10298: out = 24'(10156);
			10299: out = 24'(10168);
			10300: out = 24'(10216);
			10301: out = 24'(10276);
			10302: out = 24'(10348);
			10303: out = 24'(10380);
			10304: out = 24'(10456);
			10305: out = 24'(10472);
			10306: out = 24'(10544);
			10307: out = 24'(10632);
			10308: out = 24'(10584);
			10309: out = 24'(10716);
			10310: out = 24'(10756);
			10311: out = 24'(10824);
			10312: out = 24'(10840);
			10313: out = 24'(10880);
			10314: out = 24'(10960);
			10315: out = 24'(11012);
			10316: out = 24'(11000);
			10317: out = 24'(11060);
			10318: out = 24'(11112);
			10319: out = 24'(11140);
			10320: out = 24'(11260);
			10321: out = 24'(11248);
			10322: out = 24'(11328);
			10323: out = 24'(11368);
			10324: out = 24'(11384);
			10325: out = 24'(11508);
			10326: out = 24'(11432);
			10327: out = 24'(11552);
			10328: out = 24'(11568);
			10329: out = 24'(11620);
			10330: out = 24'(11668);
			10331: out = 24'(11676);
			10332: out = 24'(11744);
			10333: out = 24'(11772);
			10334: out = 24'(11812);
			10335: out = 24'(11836);
			10336: out = 24'(11932);
			10337: out = 24'(11916);
			10338: out = 24'(12012);
			10339: out = 24'(12008);
			10340: out = 24'(12036);
			10341: out = 24'(12108);
			10342: out = 24'(12120);
			10343: out = 24'(12196);
			10344: out = 24'(12188);
			10345: out = 24'(12236);
			10346: out = 24'(12248);
			10347: out = 24'(12328);
			10348: out = 24'(12300);
			10349: out = 24'(12360);
			10350: out = 24'(12340);
			10351: out = 24'(12376);
			10352: out = 24'(12380);
			10353: out = 24'(12376);
			10354: out = 24'(12328);
			10355: out = 24'(12292);
			10356: out = 24'(12276);
			10357: out = 24'(12292);
			10358: out = 24'(12296);
			10359: out = 24'(12300);
			10360: out = 24'(12316);
			10361: out = 24'(12288);
			10362: out = 24'(12272);
			10363: out = 24'(12276);
			10364: out = 24'(12216);
			10365: out = 24'(12268);
			10366: out = 24'(12340);
			10367: out = 24'(12252);
			10368: out = 24'(12208);
			10369: out = 24'(12180);
			10370: out = 24'(12124);
			10371: out = 24'(12196);
			10372: out = 24'(12188);
			10373: out = 24'(12152);
			10374: out = 24'(12172);
			10375: out = 24'(12204);
			10376: out = 24'(12152);
			10377: out = 24'(12252);
			10378: out = 24'(12188);
			10379: out = 24'(12196);
			10380: out = 24'(12200);
			10381: out = 24'(12224);
			10382: out = 24'(12228);
			10383: out = 24'(12188);
			10384: out = 24'(12216);
			10385: out = 24'(12192);
			10386: out = 24'(12112);
			10387: out = 24'(12184);
			10388: out = 24'(12176);
			10389: out = 24'(12176);
			10390: out = 24'(12184);
			10391: out = 24'(12124);
			10392: out = 24'(12208);
			10393: out = 24'(12196);
			10394: out = 24'(12188);
			10395: out = 24'(12200);
			10396: out = 24'(12208);
			10397: out = 24'(12084);
			10398: out = 24'(12076);
			10399: out = 24'(12148);
			10400: out = 24'(12052);
			10401: out = 24'(12072);
			10402: out = 24'(12152);
			10403: out = 24'(12028);
			10404: out = 24'(12152);
			10405: out = 24'(12056);
			10406: out = 24'(12056);
			10407: out = 24'(12100);
			10408: out = 24'(12016);
			10409: out = 24'(12056);
			10410: out = 24'(12056);
			10411: out = 24'(12040);
			10412: out = 24'(12104);
			10413: out = 24'(12064);
			10414: out = 24'(11984);
			10415: out = 24'(12024);
			10416: out = 24'(11888);
			10417: out = 24'(11948);
			10418: out = 24'(11932);
			10419: out = 24'(11860);
			10420: out = 24'(11804);
			10421: out = 24'(11864);
			10422: out = 24'(11764);
			10423: out = 24'(11836);
			10424: out = 24'(11752);
			10425: out = 24'(11800);
			10426: out = 24'(11716);
			10427: out = 24'(11764);
			10428: out = 24'(11692);
			10429: out = 24'(11680);
			10430: out = 24'(11600);
			10431: out = 24'(11612);
			10432: out = 24'(11468);
			10433: out = 24'(11432);
			10434: out = 24'(11400);
			10435: out = 24'(11388);
			10436: out = 24'(11292);
			10437: out = 24'(11324);
			10438: out = 24'(11140);
			10439: out = 24'(11212);
			10440: out = 24'(11052);
			10441: out = 24'(11000);
			10442: out = 24'(11004);
			10443: out = 24'(10916);
			10444: out = 24'(10860);
			10445: out = 24'(10860);
			10446: out = 24'(10788);
			10447: out = 24'(10664);
			10448: out = 24'(10640);
			10449: out = 24'(10536);
			10450: out = 24'(10448);
			10451: out = 24'(10400);
			10452: out = 24'(10324);
			10453: out = 24'(10256);
			10454: out = 24'(10228);
			10455: out = 24'(10124);
			10456: out = 24'(10064);
			10457: out = 24'(9956);
			10458: out = 24'(9924);
			10459: out = 24'(9824);
			10460: out = 24'(9720);
			10461: out = 24'(9724);
			10462: out = 24'(9544);
			10463: out = 24'(9532);
			10464: out = 24'(9400);
			10465: out = 24'(9352);
			10466: out = 24'(9248);
			10467: out = 24'(9240);
			10468: out = 24'(9056);
			10469: out = 24'(9016);
			10470: out = 24'(8952);
			10471: out = 24'(8872);
			10472: out = 24'(8792);
			10473: out = 24'(8680);
			10474: out = 24'(8664);
			10475: out = 24'(8568);
			10476: out = 24'(8476);
			10477: out = 24'(8388);
			10478: out = 24'(8320);
			10479: out = 24'(8172);
			10480: out = 24'(8136);
			10481: out = 24'(8064);
			10482: out = 24'(8016);
			10483: out = 24'(7884);
			10484: out = 24'(7840);
			10485: out = 24'(7768);
			10486: out = 24'(7584);
			10487: out = 24'(7584);
			10488: out = 24'(7532);
			10489: out = 24'(7392);
			10490: out = 24'(7332);
			10491: out = 24'(7248);
			10492: out = 24'(7208);
			10493: out = 24'(7096);
			10494: out = 24'(7028);
			10495: out = 24'(6948);
			10496: out = 24'(6888);
			10497: out = 24'(6808);
			10498: out = 24'(6728);
			10499: out = 24'(6640);
			10500: out = 24'(6556);
			10501: out = 24'(6468);
			10502: out = 24'(6440);
			10503: out = 24'(6412);
			10504: out = 24'(6308);
			10505: out = 24'(6232);
			10506: out = 24'(6168);
			10507: out = 24'(6096);
			10508: out = 24'(5972);
			10509: out = 24'(5976);
			10510: out = 24'(5792);
			10511: out = 24'(5792);
			10512: out = 24'(5732);
			10513: out = 24'(5640);
			10514: out = 24'(5612);
			10515: out = 24'(5516);
			10516: out = 24'(5444);
			10517: out = 24'(5392);
			10518: out = 24'(5364);
			10519: out = 24'(5280);
			10520: out = 24'(5176);
			10521: out = 24'(5120);
			10522: out = 24'(5076);
			10523: out = 24'(5032);
			10524: out = 24'(5000);
			10525: out = 24'(4856);
			10526: out = 24'(4824);
			10527: out = 24'(4816);
			10528: out = 24'(4632);
			10529: out = 24'(4672);
			10530: out = 24'(4612);
			10531: out = 24'(4472);
			10532: out = 24'(4460);
			10533: out = 24'(4468);
			10534: out = 24'(4376);
			10535: out = 24'(4324);
			10536: out = 24'(4232);
			10537: out = 24'(4220);
			10538: out = 24'(4108);
			10539: out = 24'(4088);
			10540: out = 24'(4040);
			10541: out = 24'(3984);
			10542: out = 24'(3932);
			10543: out = 24'(3864);
			10544: out = 24'(3820);
			10545: out = 24'(3812);
			10546: out = 24'(3724);
			10547: out = 24'(3656);
			10548: out = 24'(3616);
			10549: out = 24'(3624);
			10550: out = 24'(3484);
			10551: out = 24'(3468);
			10552: out = 24'(3472);
			10553: out = 24'(3344);
			10554: out = 24'(3336);
			10555: out = 24'(3272);
			10556: out = 24'(3280);
			10557: out = 24'(3160);
			10558: out = 24'(3192);
			10559: out = 24'(3068);
			10560: out = 24'(3084);
			10561: out = 24'(3056);
			10562: out = 24'(2916);
			10563: out = 24'(2952);
			10564: out = 24'(2944);
			10565: out = 24'(2824);
			10566: out = 24'(2828);
			10567: out = 24'(2724);
			10568: out = 24'(2756);
			10569: out = 24'(2676);
			10570: out = 24'(2632);
			10571: out = 24'(2616);
			10572: out = 24'(2568);
			10573: out = 24'(2536);
			10574: out = 24'(2492);
			10575: out = 24'(2496);
			10576: out = 24'(2400);
			10577: out = 24'(2404);
			10578: out = 24'(2308);
			10579: out = 24'(2308);
			10580: out = 24'(2268);
			10581: out = 24'(2212);
			10582: out = 24'(2100);
			10583: out = 24'(2044);
			10584: out = 24'(1920);
			10585: out = 24'(1824);
			10586: out = 24'(1728);
			10587: out = 24'(1648);
			10588: out = 24'(1540);
			10589: out = 24'(1428);
			10590: out = 24'(1380);
			10591: out = 24'(1280);
			10592: out = 24'(1160);
			10593: out = 24'(1120);
			10594: out = 24'(1044);
			10595: out = 24'(864);
			10596: out = 24'(880);
			10597: out = 24'(736);
			10598: out = 24'(684);
			10599: out = 24'(592);
			10600: out = 24'(512);
			10601: out = 24'(432);
			10602: out = 24'(336);
			10603: out = 24'(308);
			10604: out = 24'(168);
			10605: out = 24'(68);
			10606: out = 24'(24);
			10607: out = 24'(-4);
			10608: out = 24'(-172);
			10609: out = 24'(-156);
			10610: out = 24'(-272);
			10611: out = 24'(-312);
			10612: out = 24'(-400);
			10613: out = 24'(-444);
			10614: out = 24'(-488);
			10615: out = 24'(-584);
			10616: out = 24'(-644);
			10617: out = 24'(-684);
			10618: out = 24'(-808);
			10619: out = 24'(-876);
			10620: out = 24'(-908);
			10621: out = 24'(-960);
			10622: out = 24'(-1004);
			10623: out = 24'(-1096);
			10624: out = 24'(-1120);
			10625: out = 24'(-1236);
			10626: out = 24'(-1216);
			10627: out = 24'(-1340);
			10628: out = 24'(-1356);
			10629: out = 24'(-1428);
			10630: out = 24'(-1516);
			10631: out = 24'(-1532);
			10632: out = 24'(-1596);
			10633: out = 24'(-1688);
			10634: out = 24'(-1696);
			10635: out = 24'(-1792);
			10636: out = 24'(-1792);
			10637: out = 24'(-1924);
			10638: out = 24'(-1920);
			10639: out = 24'(-1992);
			10640: out = 24'(-2076);
			10641: out = 24'(-2100);
			10642: out = 24'(-2164);
			10643: out = 24'(-2208);
			10644: out = 24'(-2312);
			10645: out = 24'(-2368);
			10646: out = 24'(-2400);
			10647: out = 24'(-2492);
			10648: out = 24'(-2504);
			10649: out = 24'(-2564);
			10650: out = 24'(-2640);
			10651: out = 24'(-2680);
			10652: out = 24'(-2768);
			10653: out = 24'(-2768);
			10654: out = 24'(-2864);
			10655: out = 24'(-2908);
			10656: out = 24'(-2964);
			10657: out = 24'(-3024);
			10658: out = 24'(-3112);
			10659: out = 24'(-3116);
			10660: out = 24'(-3188);
			10661: out = 24'(-3268);
			10662: out = 24'(-3272);
			10663: out = 24'(-3380);
			10664: out = 24'(-3488);
			10665: out = 24'(-3412);
			10666: out = 24'(-3584);
			10667: out = 24'(-3616);
			10668: out = 24'(-3708);
			10669: out = 24'(-3732);
			10670: out = 24'(-3792);
			10671: out = 24'(-3872);
			10672: out = 24'(-3952);
			10673: out = 24'(-3996);
			10674: out = 24'(-4048);
			10675: out = 24'(-4176);
			10676: out = 24'(-4204);
			10677: out = 24'(-4268);
			10678: out = 24'(-4348);
			10679: out = 24'(-4460);
			10680: out = 24'(-4536);
			10681: out = 24'(-4540);
			10682: out = 24'(-4652);
			10683: out = 24'(-4760);
			10684: out = 24'(-4788);
			10685: out = 24'(-4908);
			10686: out = 24'(-4976);
			10687: out = 24'(-5076);
			10688: out = 24'(-5116);
			10689: out = 24'(-5232);
			10690: out = 24'(-5284);
			10691: out = 24'(-5388);
			10692: out = 24'(-5496);
			10693: out = 24'(-5588);
			10694: out = 24'(-5712);
			10695: out = 24'(-5840);
			10696: out = 24'(-5864);
			10697: out = 24'(-6036);
			10698: out = 24'(-6108);
			10699: out = 24'(-6176);
			10700: out = 24'(-6296);
			10701: out = 24'(-6416);
			10702: out = 24'(-6448);
			10703: out = 24'(-6580);
			10704: out = 24'(-6752);
			10705: out = 24'(-6808);
			10706: out = 24'(-6928);
			10707: out = 24'(-7060);
			10708: out = 24'(-7196);
			10709: out = 24'(-7236);
			10710: out = 24'(-7408);
			10711: out = 24'(-7460);
			10712: out = 24'(-7588);
			10713: out = 24'(-7740);
			10714: out = 24'(-7812);
			10715: out = 24'(-7936);
			10716: out = 24'(-8036);
			10717: out = 24'(-8192);
			10718: out = 24'(-8276);
			10719: out = 24'(-8392);
			10720: out = 24'(-8500);
			10721: out = 24'(-8596);
			10722: out = 24'(-8716);
			10723: out = 24'(-8788);
			10724: out = 24'(-8932);
			10725: out = 24'(-8988);
			10726: out = 24'(-9128);
			10727: out = 24'(-9236);
			10728: out = 24'(-9248);
			10729: out = 24'(-9472);
			10730: out = 24'(-9496);
			10731: out = 24'(-9604);
			10732: out = 24'(-9676);
			10733: out = 24'(-9780);
			10734: out = 24'(-9872);
			10735: out = 24'(-9928);
			10736: out = 24'(-10068);
			10737: out = 24'(-10132);
			10738: out = 24'(-10212);
			10739: out = 24'(-10324);
			10740: out = 24'(-10328);
			10741: out = 24'(-10484);
			10742: out = 24'(-10516);
			10743: out = 24'(-10636);
			10744: out = 24'(-10644);
			10745: out = 24'(-10780);
			10746: out = 24'(-10772);
			10747: out = 24'(-10880);
			10748: out = 24'(-10928);
			10749: out = 24'(-11000);
			10750: out = 24'(-11052);
			10751: out = 24'(-11096);
			10752: out = 24'(-11184);
			10753: out = 24'(-11192);
			10754: out = 24'(-11300);
			10755: out = 24'(-11344);
			10756: out = 24'(-11396);
			10757: out = 24'(-11444);
			10758: out = 24'(-11456);
			10759: out = 24'(-11576);
			10760: out = 24'(-11540);
			10761: out = 24'(-11616);
			10762: out = 24'(-11612);
			10763: out = 24'(-11716);
			10764: out = 24'(-11704);
			10765: out = 24'(-11772);
			10766: out = 24'(-11800);
			10767: out = 24'(-11820);
			10768: out = 24'(-11876);
			10769: out = 24'(-11872);
			10770: out = 24'(-11936);
			10771: out = 24'(-11920);
			10772: out = 24'(-12008);
			10773: out = 24'(-11976);
			10774: out = 24'(-12024);
			10775: out = 24'(-12016);
			10776: out = 24'(-12036);
			10777: out = 24'(-12136);
			10778: out = 24'(-12076);
			10779: out = 24'(-12148);
			10780: out = 24'(-12112);
			10781: out = 24'(-12204);
			10782: out = 24'(-12180);
			10783: out = 24'(-12224);
			10784: out = 24'(-12184);
			10785: out = 24'(-12228);
			10786: out = 24'(-12252);
			10787: out = 24'(-12240);
			10788: out = 24'(-12208);
			10789: out = 24'(-12296);
			10790: out = 24'(-12252);
			10791: out = 24'(-12240);
			10792: out = 24'(-12288);
			10793: out = 24'(-12300);
			10794: out = 24'(-12260);
			10795: out = 24'(-12272);
			10796: out = 24'(-12332);
			10797: out = 24'(-12244);
			10798: out = 24'(-12288);
			10799: out = 24'(-12252);
			10800: out = 24'(-12272);
			10801: out = 24'(-12300);
			10802: out = 24'(-12272);
			10803: out = 24'(-12240);
			10804: out = 24'(-12264);
			10805: out = 24'(-12260);
			10806: out = 24'(-12272);
			10807: out = 24'(-12216);
			10808: out = 24'(-12252);
			10809: out = 24'(-12244);
			10810: out = 24'(-12200);
			10811: out = 24'(-12184);
			10812: out = 24'(-12204);
			10813: out = 24'(-12172);
			10814: out = 24'(-12184);
			10815: out = 24'(-12144);
			10816: out = 24'(-12132);
			10817: out = 24'(-12188);
			10818: out = 24'(-12132);
			10819: out = 24'(-12084);
			10820: out = 24'(-12104);
			10821: out = 24'(-12052);
			10822: out = 24'(-12092);
			10823: out = 24'(-12000);
			10824: out = 24'(-12036);
			10825: out = 24'(-12032);
			10826: out = 24'(-11976);
			10827: out = 24'(-11948);
			10828: out = 24'(-11996);
			10829: out = 24'(-11920);
			10830: out = 24'(-11932);
			10831: out = 24'(-11872);
			10832: out = 24'(-11912);
			10833: out = 24'(-11836);
			10834: out = 24'(-11808);
			10835: out = 24'(-11812);
			10836: out = 24'(-11788);
			10837: out = 24'(-11756);
			10838: out = 24'(-11728);
			10839: out = 24'(-11696);
			10840: out = 24'(-11692);
			10841: out = 24'(-11684);
			10842: out = 24'(-11668);
			10843: out = 24'(-11560);
			10844: out = 24'(-11640);
			10845: out = 24'(-11568);
			10846: out = 24'(-11520);
			10847: out = 24'(-11544);
			10848: out = 24'(-11472);
			10849: out = 24'(-11456);
			10850: out = 24'(-11460);
			10851: out = 24'(-11392);
			10852: out = 24'(-11372);
			10853: out = 24'(-11376);
			10854: out = 24'(-11328);
			10855: out = 24'(-11280);
			10856: out = 24'(-11288);
			10857: out = 24'(-11220);
			10858: out = 24'(-11220);
			10859: out = 24'(-11188);
			10860: out = 24'(-11128);
			10861: out = 24'(-11140);
			10862: out = 24'(-11084);
			10863: out = 24'(-11064);
			10864: out = 24'(-11040);
			10865: out = 24'(-10984);
			10866: out = 24'(-10992);
			10867: out = 24'(-10900);
			10868: out = 24'(-10956);
			10869: out = 24'(-10864);
			10870: out = 24'(-10824);
			10871: out = 24'(-10800);
			10872: out = 24'(-10776);
			10873: out = 24'(-10676);
			10874: out = 24'(-10692);
			10875: out = 24'(-10616);
			10876: out = 24'(-10612);
			10877: out = 24'(-10540);
			10878: out = 24'(-10504);
			10879: out = 24'(-10476);
			10880: out = 24'(-10396);
			10881: out = 24'(-10400);
			10882: out = 24'(-10340);
			10883: out = 24'(-10292);
			10884: out = 24'(-10228);
			10885: out = 24'(-10180);
			10886: out = 24'(-10120);
			10887: out = 24'(-10096);
			10888: out = 24'(-10024);
			10889: out = 24'(-9992);
			10890: out = 24'(-9888);
			10891: out = 24'(-9864);
			10892: out = 24'(-9820);
			10893: out = 24'(-9760);
			10894: out = 24'(-9660);
			10895: out = 24'(-9632);
			10896: out = 24'(-9556);
			10897: out = 24'(-9468);
			10898: out = 24'(-9436);
			10899: out = 24'(-9332);
			10900: out = 24'(-9316);
			10901: out = 24'(-9224);
			10902: out = 24'(-9136);
			10903: out = 24'(-9072);
			10904: out = 24'(-8972);
			10905: out = 24'(-8936);
			10906: out = 24'(-8832);
			10907: out = 24'(-8760);
			10908: out = 24'(-8700);
			10909: out = 24'(-8608);
			10910: out = 24'(-8532);
			10911: out = 24'(-8428);
			10912: out = 24'(-8356);
			10913: out = 24'(-8304);
			10914: out = 24'(-8132);
			10915: out = 24'(-8136);
			10916: out = 24'(-8060);
			10917: out = 24'(-7928);
			10918: out = 24'(-7864);
			10919: out = 24'(-7776);
			10920: out = 24'(-7684);
			10921: out = 24'(-7600);
			10922: out = 24'(-7500);
			10923: out = 24'(-7408);
			10924: out = 24'(-7360);
			10925: out = 24'(-7256);
			10926: out = 24'(-7172);
			10927: out = 24'(-7076);
			10928: out = 24'(-7016);
			10929: out = 24'(-6896);
			10930: out = 24'(-6856);
			10931: out = 24'(-6744);
			10932: out = 24'(-6664);
			10933: out = 24'(-6568);
			10934: out = 24'(-6508);
			10935: out = 24'(-6424);
			10936: out = 24'(-6300);
			10937: out = 24'(-6280);
			10938: out = 24'(-6160);
			10939: out = 24'(-6084);
			10940: out = 24'(-6028);
			10941: out = 24'(-5948);
			10942: out = 24'(-5828);
			10943: out = 24'(-5792);
			10944: out = 24'(-5688);
			10945: out = 24'(-5604);
			10946: out = 24'(-5564);
			10947: out = 24'(-5484);
			10948: out = 24'(-5400);
			10949: out = 24'(-5268);
			10950: out = 24'(-5312);
			10951: out = 24'(-5184);
			10952: out = 24'(-5056);
			10953: out = 24'(-5024);
			10954: out = 24'(-4936);
			10955: out = 24'(-4912);
			10956: out = 24'(-4776);
			10957: out = 24'(-4756);
			10958: out = 24'(-4676);
			10959: out = 24'(-4600);
			10960: out = 24'(-4584);
			10961: out = 24'(-4460);
			10962: out = 24'(-4396);
			10963: out = 24'(-4376);
			10964: out = 24'(-4268);
			10965: out = 24'(-4220);
			10966: out = 24'(-4156);
			10967: out = 24'(-4084);
			10968: out = 24'(-4052);
			10969: out = 24'(-3980);
			10970: out = 24'(-3896);
			10971: out = 24'(-3856);
			10972: out = 24'(-3772);
			10973: out = 24'(-3712);
			10974: out = 24'(-3680);
			10975: out = 24'(-3592);
			10976: out = 24'(-3568);
			10977: out = 24'(-3524);
			10978: out = 24'(-3440);
			10979: out = 24'(-3380);
			10980: out = 24'(-3356);
			10981: out = 24'(-3276);
			10982: out = 24'(-3240);
			10983: out = 24'(-3152);
			10984: out = 24'(-3120);
			10985: out = 24'(-3088);
			10986: out = 24'(-3016);
			10987: out = 24'(-2952);
			10988: out = 24'(-2936);
			10989: out = 24'(-2836);
			10990: out = 24'(-2820);
			10991: out = 24'(-2824);
			10992: out = 24'(-2692);
			10993: out = 24'(-2712);
			10994: out = 24'(-2632);
			10995: out = 24'(-2572);
			10996: out = 24'(-2560);
			10997: out = 24'(-2476);
			10998: out = 24'(-2472);
			10999: out = 24'(-2396);
			11000: out = 24'(-2356);
			11001: out = 24'(-2348);
			11002: out = 24'(-2276);
			11003: out = 24'(-2248);
			11004: out = 24'(-2208);
			11005: out = 24'(-2144);
			11006: out = 24'(-2084);
			11007: out = 24'(-1992);
			11008: out = 24'(-1912);
			11009: out = 24'(-1864);
			11010: out = 24'(-1808);
			11011: out = 24'(-1708);
			11012: out = 24'(-1632);
			11013: out = 24'(-1592);
			11014: out = 24'(-1544);
			11015: out = 24'(-1448);
			11016: out = 24'(-1412);
			11017: out = 24'(-1304);
			11018: out = 24'(-1308);
			11019: out = 24'(-1196);
			11020: out = 24'(-1108);
			11021: out = 24'(-1112);
			11022: out = 24'(-1056);
			11023: out = 24'(-920);
			11024: out = 24'(-920);
			11025: out = 24'(-900);
			11026: out = 24'(-776);
			11027: out = 24'(-732);
			11028: out = 24'(-724);
			11029: out = 24'(-628);
			11030: out = 24'(-572);
			11031: out = 24'(-588);
			11032: out = 24'(-440);
			11033: out = 24'(-444);
			11034: out = 24'(-404);
			11035: out = 24'(-336);
			11036: out = 24'(-316);
			11037: out = 24'(-232);
			11038: out = 24'(-176);
			11039: out = 24'(-176);
			11040: out = 24'(-104);
			11041: out = 24'(-64);
			11042: out = 24'(24);
			11043: out = 24'(16);
			11044: out = 24'(48);
			11045: out = 24'(148);
			11046: out = 24'(184);
			11047: out = 24'(204);
			11048: out = 24'(224);
			11049: out = 24'(312);
			11050: out = 24'(288);
			11051: out = 24'(448);
			11052: out = 24'(332);
			11053: out = 24'(456);
			11054: out = 24'(468);
			11055: out = 24'(576);
			11056: out = 24'(560);
			11057: out = 24'(592);
			11058: out = 24'(676);
			11059: out = 24'(728);
			11060: out = 24'(752);
			11061: out = 24'(776);
			11062: out = 24'(836);
			11063: out = 24'(880);
			11064: out = 24'(888);
			11065: out = 24'(964);
			11066: out = 24'(960);
			11067: out = 24'(1036);
			11068: out = 24'(1072);
			11069: out = 24'(1096);
			11070: out = 24'(1164);
			11071: out = 24'(1176);
			11072: out = 24'(1236);
			11073: out = 24'(1272);
			11074: out = 24'(1320);
			11075: out = 24'(1368);
			11076: out = 24'(1384);
			11077: out = 24'(1440);
			11078: out = 24'(1436);
			11079: out = 24'(1520);
			11080: out = 24'(1552);
			11081: out = 24'(1592);
			11082: out = 24'(1612);
			11083: out = 24'(1668);
			11084: out = 24'(1744);
			11085: out = 24'(1752);
			11086: out = 24'(1812);
			11087: out = 24'(1836);
			11088: out = 24'(1900);
			11089: out = 24'(1928);
			11090: out = 24'(1984);
			11091: out = 24'(2040);
			11092: out = 24'(2072);
			11093: out = 24'(2148);
			11094: out = 24'(2180);
			11095: out = 24'(2212);
			11096: out = 24'(2264);
			11097: out = 24'(2356);
			11098: out = 24'(2376);
			11099: out = 24'(2440);
			11100: out = 24'(2504);
			11101: out = 24'(2544);
			11102: out = 24'(2628);
			11103: out = 24'(2644);
			11104: out = 24'(2728);
			11105: out = 24'(2756);
			11106: out = 24'(2872);
			11107: out = 24'(2888);
			11108: out = 24'(2976);
			11109: out = 24'(3020);
			11110: out = 24'(3112);
			11111: out = 24'(3156);
			11112: out = 24'(3208);
			11113: out = 24'(3308);
			11114: out = 24'(3352);
			11115: out = 24'(3424);
			11116: out = 24'(3552);
			11117: out = 24'(3580);
			11118: out = 24'(3700);
			11119: out = 24'(3724);
			11120: out = 24'(3792);
			11121: out = 24'(3904);
			11122: out = 24'(3980);
			11123: out = 24'(3972);
			11124: out = 24'(4152);
			11125: out = 24'(4148);
			11126: out = 24'(4292);
			11127: out = 24'(4328);
			11128: out = 24'(4404);
			11129: out = 24'(4488);
			11130: out = 24'(4548);
			11131: out = 24'(4676);
			11132: out = 24'(4728);
			11133: out = 24'(4804);
			11134: out = 24'(4880);
			11135: out = 24'(4976);
			11136: out = 24'(5004);
			11137: out = 24'(5132);
			11138: out = 24'(5212);
			11139: out = 24'(5216);
			11140: out = 24'(5376);
			11141: out = 24'(5412);
			11142: out = 24'(5512);
			11143: out = 24'(5548);
			11144: out = 24'(5604);
			11145: out = 24'(5728);
			11146: out = 24'(5740);
			11147: out = 24'(5828);
			11148: out = 24'(5904);
			11149: out = 24'(5988);
			11150: out = 24'(6060);
			11151: out = 24'(6136);
			11152: out = 24'(6168);
			11153: out = 24'(6264);
			11154: out = 24'(6308);
			11155: out = 24'(6344);
			11156: out = 24'(6444);
			11157: out = 24'(6552);
			11158: out = 24'(6584);
			11159: out = 24'(6648);
			11160: out = 24'(6700);
			11161: out = 24'(6780);
			11162: out = 24'(6848);
			11163: out = 24'(6836);
			11164: out = 24'(6952);
			11165: out = 24'(6988);
			11166: out = 24'(7068);
			11167: out = 24'(7120);
			11168: out = 24'(7208);
			11169: out = 24'(7188);
			11170: out = 24'(7328);
			11171: out = 24'(7348);
			11172: out = 24'(7376);
			11173: out = 24'(7492);
			11174: out = 24'(7500);
			11175: out = 24'(7472);
			11176: out = 24'(7660);
			11177: out = 24'(7656);
			11178: out = 24'(7736);
			11179: out = 24'(7748);
			11180: out = 24'(7820);
			11181: out = 24'(7852);
			11182: out = 24'(7900);
			11183: out = 24'(7984);
			11184: out = 24'(7964);
			11185: out = 24'(8096);
			11186: out = 24'(8056);
			11187: out = 24'(8168);
			11188: out = 24'(8164);
			11189: out = 24'(8232);
			11190: out = 24'(8316);
			11191: out = 24'(8300);
			11192: out = 24'(8356);
			11193: out = 24'(8428);
			11194: out = 24'(8440);
			11195: out = 24'(8536);
			11196: out = 24'(8496);
			11197: out = 24'(8584);
			11198: out = 24'(8624);
			11199: out = 24'(8676);
			11200: out = 24'(8688);
			11201: out = 24'(8772);
			11202: out = 24'(8812);
			11203: out = 24'(8820);
			11204: out = 24'(8864);
			11205: out = 24'(8908);
			11206: out = 24'(8932);
			11207: out = 24'(8976);
			11208: out = 24'(9016);
			11209: out = 24'(9072);
			11210: out = 24'(9084);
			11211: out = 24'(9124);
			11212: out = 24'(9204);
			11213: out = 24'(9208);
			11214: out = 24'(9224);
			11215: out = 24'(9292);
			11216: out = 24'(9332);
			11217: out = 24'(9328);
			11218: out = 24'(9396);
			11219: out = 24'(9412);
			11220: out = 24'(9452);
			11221: out = 24'(9472);
			11222: out = 24'(9532);
			11223: out = 24'(9548);
			11224: out = 24'(9604);
			11225: out = 24'(9616);
			11226: out = 24'(9648);
			11227: out = 24'(9708);
			11228: out = 24'(9680);
			11229: out = 24'(9764);
			11230: out = 24'(9760);
			11231: out = 24'(9792);
			11232: out = 24'(9808);
			11233: out = 24'(9884);
			11234: out = 24'(9868);
			11235: out = 24'(9920);
			11236: out = 24'(9948);
			11237: out = 24'(9952);
			11238: out = 24'(9968);
			11239: out = 24'(9992);
			11240: out = 24'(9968);
			11241: out = 24'(10024);
			11242: out = 24'(10004);
			11243: out = 24'(9980);
			11244: out = 24'(10028);
			11245: out = 24'(9996);
			11246: out = 24'(9988);
			11247: out = 24'(10024);
			11248: out = 24'(9932);
			11249: out = 24'(9980);
			11250: out = 24'(9928);
			11251: out = 24'(9936);
			11252: out = 24'(9964);
			11253: out = 24'(9964);
			11254: out = 24'(9952);
			11255: out = 24'(9960);
			11256: out = 24'(9960);
			11257: out = 24'(9988);
			11258: out = 24'(9964);
			11259: out = 24'(9964);
			11260: out = 24'(9976);
			11261: out = 24'(9912);
			11262: out = 24'(9960);
			11263: out = 24'(9856);
			11264: out = 24'(9876);
			11265: out = 24'(9900);
			11266: out = 24'(9944);
			11267: out = 24'(9856);
			11268: out = 24'(9920);
			11269: out = 24'(9876);
			11270: out = 24'(9912);
			11271: out = 24'(9936);
			11272: out = 24'(9836);
			11273: out = 24'(9904);
			11274: out = 24'(9896);
			11275: out = 24'(9960);
			11276: out = 24'(9920);
			11277: out = 24'(9868);
			11278: out = 24'(9928);
			11279: out = 24'(9920);
			11280: out = 24'(9964);
			11281: out = 24'(9908);
			11282: out = 24'(9932);
			11283: out = 24'(9936);
			11284: out = 24'(9964);
			11285: out = 24'(9884);
			11286: out = 24'(9908);
			11287: out = 24'(9884);
			11288: out = 24'(9908);
			11289: out = 24'(9852);
			11290: out = 24'(9848);
			11291: out = 24'(9880);
			11292: out = 24'(9932);
			11293: out = 24'(9792);
			11294: out = 24'(9820);
			11295: out = 24'(9816);
			11296: out = 24'(9744);
			11297: out = 24'(9768);
			11298: out = 24'(9816);
			11299: out = 24'(9772);
			11300: out = 24'(9720);
			11301: out = 24'(9788);
			11302: out = 24'(9696);
			11303: out = 24'(9680);
			11304: out = 24'(9760);
			11305: out = 24'(9732);
			11306: out = 24'(9660);
			11307: out = 24'(9644);
			11308: out = 24'(9640);
			11309: out = 24'(9660);
			11310: out = 24'(9640);
			11311: out = 24'(9584);
			11312: out = 24'(9600);
			11313: out = 24'(9584);
			11314: out = 24'(9540);
			11315: out = 24'(9556);
			11316: out = 24'(9408);
			11317: out = 24'(9424);
			11318: out = 24'(9376);
			11319: out = 24'(9428);
			11320: out = 24'(9356);
			11321: out = 24'(9300);
			11322: out = 24'(9320);
			11323: out = 24'(9260);
			11324: out = 24'(9256);
			11325: out = 24'(9240);
			11326: out = 24'(9168);
			11327: out = 24'(9140);
			11328: out = 24'(9116);
			11329: out = 24'(9048);
			11330: out = 24'(8960);
			11331: out = 24'(8984);
			11332: out = 24'(8860);
			11333: out = 24'(8868);
			11334: out = 24'(8800);
			11335: out = 24'(8776);
			11336: out = 24'(8700);
			11337: out = 24'(8692);
			11338: out = 24'(8588);
			11339: out = 24'(8584);
			11340: out = 24'(8548);
			11341: out = 24'(8480);
			11342: out = 24'(8432);
			11343: out = 24'(8312);
			11344: out = 24'(8316);
			11345: out = 24'(8212);
			11346: out = 24'(8160);
			11347: out = 24'(8124);
			11348: out = 24'(8020);
			11349: out = 24'(7968);
			11350: out = 24'(7920);
			11351: out = 24'(7884);
			11352: out = 24'(7752);
			11353: out = 24'(7720);
			11354: out = 24'(7696);
			11355: out = 24'(7616);
			11356: out = 24'(7532);
			11357: out = 24'(7484);
			11358: out = 24'(7404);
			11359: out = 24'(7396);
			11360: out = 24'(7276);
			11361: out = 24'(7176);
			11362: out = 24'(7180);
			11363: out = 24'(7108);
			11364: out = 24'(7000);
			11365: out = 24'(6972);
			11366: out = 24'(6872);
			11367: out = 24'(6776);
			11368: out = 24'(6772);
			11369: out = 24'(6680);
			11370: out = 24'(6676);
			11371: out = 24'(6492);
			11372: out = 24'(6500);
			11373: out = 24'(6448);
			11374: out = 24'(6344);
			11375: out = 24'(6284);
			11376: out = 24'(6260);
			11377: out = 24'(6144);
			11378: out = 24'(6148);
			11379: out = 24'(6020);
			11380: out = 24'(5968);
			11381: out = 24'(5928);
			11382: out = 24'(5884);
			11383: out = 24'(5748);
			11384: out = 24'(5688);
			11385: out = 24'(5704);
			11386: out = 24'(5556);
			11387: out = 24'(5540);
			11388: out = 24'(5476);
			11389: out = 24'(5408);
			11390: out = 24'(5384);
			11391: out = 24'(5280);
			11392: out = 24'(5244);
			11393: out = 24'(5188);
			11394: out = 24'(5116);
			11395: out = 24'(5048);
			11396: out = 24'(4992);
			11397: out = 24'(4948);
			11398: out = 24'(4944);
			11399: out = 24'(4844);
			11400: out = 24'(4772);
			11401: out = 24'(4784);
			11402: out = 24'(4708);
			11403: out = 24'(4620);
			11404: out = 24'(4536);
			11405: out = 24'(4512);
			11406: out = 24'(4508);
			11407: out = 24'(4336);
			11408: out = 24'(4332);
			11409: out = 24'(4328);
			11410: out = 24'(4224);
			11411: out = 24'(4192);
			11412: out = 24'(4124);
			11413: out = 24'(4112);
			11414: out = 24'(4024);
			11415: out = 24'(3992);
			11416: out = 24'(3948);
			11417: out = 24'(3860);
			11418: out = 24'(3828);
			11419: out = 24'(3776);
			11420: out = 24'(3744);
			11421: out = 24'(3660);
			11422: out = 24'(3616);
			11423: out = 24'(3608);
			11424: out = 24'(3572);
			11425: out = 24'(3484);
			11426: out = 24'(3472);
			11427: out = 24'(3416);
			11428: out = 24'(3352);
			11429: out = 24'(3284);
			11430: out = 24'(3308);
			11431: out = 24'(3188);
			11432: out = 24'(3188);
			11433: out = 24'(3128);
			11434: out = 24'(3080);
			11435: out = 24'(3068);
			11436: out = 24'(3004);
			11437: out = 24'(3004);
			11438: out = 24'(2904);
			11439: out = 24'(2900);
			11440: out = 24'(2844);
			11441: out = 24'(2812);
			11442: out = 24'(2808);
			11443: out = 24'(2720);
			11444: out = 24'(2684);
			11445: out = 24'(2660);
			11446: out = 24'(2612);
			11447: out = 24'(2580);
			11448: out = 24'(2548);
			11449: out = 24'(2512);
			11450: out = 24'(2436);
			11451: out = 24'(2444);
			11452: out = 24'(2388);
			11453: out = 24'(2368);
			11454: out = 24'(2300);
			11455: out = 24'(2324);
			11456: out = 24'(2268);
			11457: out = 24'(2200);
			11458: out = 24'(2228);
			11459: out = 24'(2140);
			11460: out = 24'(2124);
			11461: out = 24'(2140);
			11462: out = 24'(1992);
			11463: out = 24'(2064);
			11464: out = 24'(2000);
			11465: out = 24'(1956);
			11466: out = 24'(1964);
			11467: out = 24'(1896);
			11468: out = 24'(1864);
			11469: out = 24'(1872);
			11470: out = 24'(1836);
			11471: out = 24'(1780);
			11472: out = 24'(1764);
			11473: out = 24'(1596);
			11474: out = 24'(1536);
			11475: out = 24'(1520);
			11476: out = 24'(1380);
			11477: out = 24'(1316);
			11478: out = 24'(1260);
			11479: out = 24'(1140);
			11480: out = 24'(1092);
			11481: out = 24'(1024);
			11482: out = 24'(924);
			11483: out = 24'(872);
			11484: out = 24'(788);
			11485: out = 24'(744);
			11486: out = 24'(648);
			11487: out = 24'(580);
			11488: out = 24'(532);
			11489: out = 24'(440);
			11490: out = 24'(408);
			11491: out = 24'(316);
			11492: out = 24'(268);
			11493: out = 24'(212);
			11494: out = 24'(148);
			11495: out = 24'(88);
			11496: out = 24'(16);
			11497: out = 24'(-56);
			11498: out = 24'(-72);
			11499: out = 24'(-148);
			11500: out = 24'(-184);
			11501: out = 24'(-308);
			11502: out = 24'(-344);
			11503: out = 24'(-388);
			11504: out = 24'(-464);
			11505: out = 24'(-480);
			11506: out = 24'(-512);
			11507: out = 24'(-604);
			11508: out = 24'(-616);
			11509: out = 24'(-680);
			11510: out = 24'(-736);
			11511: out = 24'(-784);
			11512: out = 24'(-832);
			11513: out = 24'(-920);
			11514: out = 24'(-968);
			11515: out = 24'(-960);
			11516: out = 24'(-1048);
			11517: out = 24'(-1076);
			11518: out = 24'(-1128);
			11519: out = 24'(-1204);
			11520: out = 24'(-1216);
			11521: out = 24'(-1264);
			11522: out = 24'(-1360);
			11523: out = 24'(-1360);
			11524: out = 24'(-1440);
			11525: out = 24'(-1468);
			11526: out = 24'(-1508);
			11527: out = 24'(-1564);
			11528: out = 24'(-1604);
			11529: out = 24'(-1644);
			11530: out = 24'(-1672);
			11531: out = 24'(-1760);
			11532: out = 24'(-1772);
			11533: out = 24'(-1872);
			11534: out = 24'(-1856);
			11535: out = 24'(-1932);
			11536: out = 24'(-1956);
			11537: out = 24'(-2024);
			11538: out = 24'(-2068);
			11539: out = 24'(-2064);
			11540: out = 24'(-2192);
			11541: out = 24'(-2156);
			11542: out = 24'(-2252);
			11543: out = 24'(-2320);
			11544: out = 24'(-2300);
			11545: out = 24'(-2352);
			11546: out = 24'(-2428);
			11547: out = 24'(-2432);
			11548: out = 24'(-2540);
			11549: out = 24'(-2536);
			11550: out = 24'(-2644);
			11551: out = 24'(-2612);
			11552: out = 24'(-2688);
			11553: out = 24'(-2772);
			11554: out = 24'(-2804);
			11555: out = 24'(-2828);
			11556: out = 24'(-2912);
			11557: out = 24'(-2956);
			11558: out = 24'(-2976);
			11559: out = 24'(-3052);
			11560: out = 24'(-3116);
			11561: out = 24'(-3128);
			11562: out = 24'(-3192);
			11563: out = 24'(-3292);
			11564: out = 24'(-3300);
			11565: out = 24'(-3352);
			11566: out = 24'(-3428);
			11567: out = 24'(-3460);
			11568: out = 24'(-3536);
			11569: out = 24'(-3592);
			11570: out = 24'(-3632);
			11571: out = 24'(-3728);
			11572: out = 24'(-3844);
			11573: out = 24'(-3808);
			11574: out = 24'(-3936);
			11575: out = 24'(-3924);
			11576: out = 24'(-4048);
			11577: out = 24'(-4108);
			11578: out = 24'(-4192);
			11579: out = 24'(-4236);
			11580: out = 24'(-4292);
			11581: out = 24'(-4396);
			11582: out = 24'(-4472);
			11583: out = 24'(-4508);
			11584: out = 24'(-4668);
			11585: out = 24'(-4696);
			11586: out = 24'(-4744);
			11587: out = 24'(-4840);
			11588: out = 24'(-4888);
			11589: out = 24'(-5032);
			11590: out = 24'(-5060);
			11591: out = 24'(-5184);
			11592: out = 24'(-5264);
			11593: out = 24'(-5404);
			11594: out = 24'(-5428);
			11595: out = 24'(-5548);
			11596: out = 24'(-5596);
			11597: out = 24'(-5732);
			11598: out = 24'(-5764);
			11599: out = 24'(-5884);
			11600: out = 24'(-5988);
			11601: out = 24'(-6072);
			11602: out = 24'(-6136);
			11603: out = 24'(-6256);
			11604: out = 24'(-6328);
			11605: out = 24'(-6420);
			11606: out = 24'(-6540);
			11607: out = 24'(-6580);
			11608: out = 24'(-6700);
			11609: out = 24'(-6756);
			11610: out = 24'(-6892);
			11611: out = 24'(-6924);
			11612: out = 24'(-7072);
			11613: out = 24'(-7132);
			11614: out = 24'(-7212);
			11615: out = 24'(-7332);
			11616: out = 24'(-7372);
			11617: out = 24'(-7472);
			11618: out = 24'(-7536);
			11619: out = 24'(-7592);
			11620: out = 24'(-7740);
			11621: out = 24'(-7780);
			11622: out = 24'(-7844);
			11623: out = 24'(-7968);
			11624: out = 24'(-8032);
			11625: out = 24'(-8076);
			11626: out = 24'(-8152);
			11627: out = 24'(-8212);
			11628: out = 24'(-8304);
			11629: out = 24'(-8364);
			11630: out = 24'(-8440);
			11631: out = 24'(-8480);
			11632: out = 24'(-8528);
			11633: out = 24'(-8620);
			11634: out = 24'(-8652);
			11635: out = 24'(-8724);
			11636: out = 24'(-8776);
			11637: out = 24'(-8832);
			11638: out = 24'(-8876);
			11639: out = 24'(-8940);
			11640: out = 24'(-8980);
			11641: out = 24'(-9044);
			11642: out = 24'(-9092);
			11643: out = 24'(-9080);
			11644: out = 24'(-9160);
			11645: out = 24'(-9244);
			11646: out = 24'(-9236);
			11647: out = 24'(-9288);
			11648: out = 24'(-9332);
			11649: out = 24'(-9376);
			11650: out = 24'(-9392);
			11651: out = 24'(-9432);
			11652: out = 24'(-9488);
			11653: out = 24'(-9476);
			11654: out = 24'(-9536);
			11655: out = 24'(-9556);
			11656: out = 24'(-9572);
			11657: out = 24'(-9616);
			11658: out = 24'(-9664);
			11659: out = 24'(-9668);
			11660: out = 24'(-9712);
			11661: out = 24'(-9732);
			11662: out = 24'(-9728);
			11663: out = 24'(-9760);
			11664: out = 24'(-9768);
			11665: out = 24'(-9848);
			11666: out = 24'(-9788);
			11667: out = 24'(-9836);
			11668: out = 24'(-9896);
			11669: out = 24'(-9896);
			11670: out = 24'(-9880);
			11671: out = 24'(-9868);
			11672: out = 24'(-9920);
			11673: out = 24'(-9916);
			11674: out = 24'(-9960);
			11675: out = 24'(-9980);
			11676: out = 24'(-9928);
			11677: out = 24'(-9980);
			11678: out = 24'(-10020);
			11679: out = 24'(-9968);
			11680: out = 24'(-9996);
			11681: out = 24'(-9988);
			11682: out = 24'(-10036);
			11683: out = 24'(-10016);
			11684: out = 24'(-9988);
			11685: out = 24'(-10036);
			11686: out = 24'(-10028);
			11687: out = 24'(-9988);
			11688: out = 24'(-10044);
			11689: out = 24'(-9996);
			11690: out = 24'(-10028);
			11691: out = 24'(-10016);
			11692: out = 24'(-9996);
			11693: out = 24'(-9980);
			11694: out = 24'(-10040);
			11695: out = 24'(-10008);
			11696: out = 24'(-9964);
			11697: out = 24'(-10012);
			11698: out = 24'(-9980);
			11699: out = 24'(-10000);
			11700: out = 24'(-9944);
			11701: out = 24'(-9976);
			11702: out = 24'(-9944);
			11703: out = 24'(-9968);
			11704: out = 24'(-9924);
			11705: out = 24'(-9952);
			11706: out = 24'(-9924);
			11707: out = 24'(-9904);
			11708: out = 24'(-9904);
			11709: out = 24'(-9884);
			11710: out = 24'(-9904);
			11711: out = 24'(-9864);
			11712: out = 24'(-9856);
			11713: out = 24'(-9856);
			11714: out = 24'(-9816);
			11715: out = 24'(-9836);
			11716: out = 24'(-9784);
			11717: out = 24'(-9832);
			11718: out = 24'(-9788);
			11719: out = 24'(-9764);
			11720: out = 24'(-9736);
			11721: out = 24'(-9728);
			11722: out = 24'(-9744);
			11723: out = 24'(-9708);
			11724: out = 24'(-9676);
			11725: out = 24'(-9636);
			11726: out = 24'(-9684);
			11727: out = 24'(-9636);
			11728: out = 24'(-9620);
			11729: out = 24'(-9548);
			11730: out = 24'(-9616);
			11731: out = 24'(-9548);
			11732: out = 24'(-9536);
			11733: out = 24'(-9488);
			11734: out = 24'(-9540);
			11735: out = 24'(-9472);
			11736: out = 24'(-9436);
			11737: out = 24'(-9452);
			11738: out = 24'(-9440);
			11739: out = 24'(-9368);
			11740: out = 24'(-9388);
			11741: out = 24'(-9380);
			11742: out = 24'(-9292);
			11743: out = 24'(-9300);
			11744: out = 24'(-9320);
			11745: out = 24'(-9240);
			11746: out = 24'(-9240);
			11747: out = 24'(-9240);
			11748: out = 24'(-9172);
			11749: out = 24'(-9188);
			11750: out = 24'(-9128);
			11751: out = 24'(-9128);
			11752: out = 24'(-9080);
			11753: out = 24'(-9044);
			11754: out = 24'(-9024);
			11755: out = 24'(-9032);
			11756: out = 24'(-8996);
			11757: out = 24'(-8920);
			11758: out = 24'(-8912);
			11759: out = 24'(-8908);
			11760: out = 24'(-8872);
			11761: out = 24'(-8856);
			11762: out = 24'(-8792);
			11763: out = 24'(-8792);
			11764: out = 24'(-8744);
			11765: out = 24'(-8752);
			11766: out = 24'(-8672);
			11767: out = 24'(-8676);
			11768: out = 24'(-8624);
			11769: out = 24'(-8568);
			11770: out = 24'(-8580);
			11771: out = 24'(-8512);
			11772: out = 24'(-8460);
			11773: out = 24'(-8428);
			11774: out = 24'(-8392);
			11775: out = 24'(-8360);
			11776: out = 24'(-8332);
			11777: out = 24'(-8272);
			11778: out = 24'(-8192);
			11779: out = 24'(-8200);
			11780: out = 24'(-8172);
			11781: out = 24'(-8068);
			11782: out = 24'(-8048);
			11783: out = 24'(-8004);
			11784: out = 24'(-7936);
			11785: out = 24'(-7916);
			11786: out = 24'(-7860);
			11787: out = 24'(-7804);
			11788: out = 24'(-7720);
			11789: out = 24'(-7696);
			11790: out = 24'(-7600);
			11791: out = 24'(-7580);
			11792: out = 24'(-7504);
			11793: out = 24'(-7424);
			11794: out = 24'(-7416);
			11795: out = 24'(-7308);
			11796: out = 24'(-7264);
			11797: out = 24'(-7180);
			11798: out = 24'(-7188);
			11799: out = 24'(-7028);
			11800: out = 24'(-7016);
			11801: out = 24'(-6928);
			11802: out = 24'(-6856);
			11803: out = 24'(-6828);
			11804: out = 24'(-6740);
			11805: out = 24'(-6632);
			11806: out = 24'(-6620);
			11807: out = 24'(-6516);
			11808: out = 24'(-6472);
			11809: out = 24'(-6396);
			11810: out = 24'(-6324);
			11811: out = 24'(-6244);
			11812: out = 24'(-6180);
			11813: out = 24'(-6124);
			11814: out = 24'(-6044);
			11815: out = 24'(-5968);
			11816: out = 24'(-5900);
			11817: out = 24'(-5864);
			11818: out = 24'(-5792);
			11819: out = 24'(-5696);
			11820: out = 24'(-5616);
			11821: out = 24'(-5564);
			11822: out = 24'(-5524);
			11823: out = 24'(-5416);
			11824: out = 24'(-5352);
			11825: out = 24'(-5332);
			11826: out = 24'(-5184);
			11827: out = 24'(-5220);
			11828: out = 24'(-5096);
			11829: out = 24'(-5012);
			11830: out = 24'(-4948);
			11831: out = 24'(-4908);
			11832: out = 24'(-4840);
			11833: out = 24'(-4756);
			11834: out = 24'(-4724);
			11835: out = 24'(-4624);
			11836: out = 24'(-4568);
			11837: out = 24'(-4596);
			11838: out = 24'(-4416);
			11839: out = 24'(-4396);
			11840: out = 24'(-4328);
			11841: out = 24'(-4252);
			11842: out = 24'(-4264);
			11843: out = 24'(-4144);
			11844: out = 24'(-4100);
			11845: out = 24'(-4012);
			11846: out = 24'(-3972);
			11847: out = 24'(-3948);
			11848: out = 24'(-3860);
			11849: out = 24'(-3768);
			11850: out = 24'(-3772);
			11851: out = 24'(-3684);
			11852: out = 24'(-3640);
			11853: out = 24'(-3572);
			11854: out = 24'(-3540);
			11855: out = 24'(-3472);
			11856: out = 24'(-3396);
			11857: out = 24'(-3432);
			11858: out = 24'(-3304);
			11859: out = 24'(-3268);
			11860: out = 24'(-3240);
			11861: out = 24'(-3152);
			11862: out = 24'(-3136);
			11863: out = 24'(-3068);
			11864: out = 24'(-3044);
			11865: out = 24'(-3016);
			11866: out = 24'(-2948);
			11867: out = 24'(-2864);
			11868: out = 24'(-2864);
			11869: out = 24'(-2788);
			11870: out = 24'(-2752);
			11871: out = 24'(-2724);
			11872: out = 24'(-2640);
			11873: out = 24'(-2668);
			11874: out = 24'(-2576);
			11875: out = 24'(-2532);
			11876: out = 24'(-2520);
			11877: out = 24'(-2424);
			11878: out = 24'(-2436);
			11879: out = 24'(-2360);
			11880: out = 24'(-2368);
			11881: out = 24'(-2280);
			11882: out = 24'(-2276);
			11883: out = 24'(-2240);
			11884: out = 24'(-2168);
			11885: out = 24'(-2156);
			11886: out = 24'(-2136);
			11887: out = 24'(-2072);
			11888: out = 24'(-2040);
			11889: out = 24'(-2004);
			11890: out = 24'(-2020);
			11891: out = 24'(-1920);
			11892: out = 24'(-1908);
			11893: out = 24'(-1856);
			11894: out = 24'(-1864);
			11895: out = 24'(-1808);
			11896: out = 24'(-1744);
			11897: out = 24'(-1712);
			11898: out = 24'(-1616);
			11899: out = 24'(-1600);
			11900: out = 24'(-1520);
			11901: out = 24'(-1452);
			11902: out = 24'(-1396);
			11903: out = 24'(-1388);
			11904: out = 24'(-1284);
			11905: out = 24'(-1248);
			11906: out = 24'(-1232);
			11907: out = 24'(-1144);
			11908: out = 24'(-1108);
			11909: out = 24'(-1012);
			11910: out = 24'(-1016);
			11911: out = 24'(-928);
			11912: out = 24'(-904);
			11913: out = 24'(-840);
			11914: out = 24'(-792);
			11915: out = 24'(-768);
			11916: out = 24'(-724);
			11917: out = 24'(-680);
			11918: out = 24'(-620);
			11919: out = 24'(-584);
			11920: out = 24'(-556);
			11921: out = 24'(-496);
			11922: out = 24'(-432);
			11923: out = 24'(-404);
			11924: out = 24'(-408);
			11925: out = 24'(-312);
			11926: out = 24'(-312);
			11927: out = 24'(-196);
			11928: out = 24'(-276);
			11929: out = 24'(-184);
			11930: out = 24'(-144);
			11931: out = 24'(-104);
			11932: out = 24'(-60);
			11933: out = 24'(-24);
			11934: out = 24'(8);
			11935: out = 24'(80);
			11936: out = 24'(60);
			11937: out = 24'(108);
			11938: out = 24'(168);
			11939: out = 24'(184);
			11940: out = 24'(184);
			11941: out = 24'(264);
			11942: out = 24'(308);
			11943: out = 24'(300);
			11944: out = 24'(360);
			11945: out = 24'(408);
			11946: out = 24'(404);
			11947: out = 24'(432);
			11948: out = 24'(516);
			11949: out = 24'(544);
			11950: out = 24'(524);
			11951: out = 24'(596);
			11952: out = 24'(604);
			11953: out = 24'(628);
			11954: out = 24'(720);
			11955: out = 24'(688);
			11956: out = 24'(764);
			11957: out = 24'(800);
			11958: out = 24'(784);
			11959: out = 24'(848);
			11960: out = 24'(892);
			11961: out = 24'(932);
			11962: out = 24'(940);
			11963: out = 24'(972);
			11964: out = 24'(1012);
			11965: out = 24'(1012);
			11966: out = 24'(1096);
			11967: out = 24'(1080);
			11968: out = 24'(1128);
			11969: out = 24'(1168);
			11970: out = 24'(1196);
			11971: out = 24'(1248);
			11972: out = 24'(1272);
			11973: out = 24'(1316);
			11974: out = 24'(1328);
			11975: out = 24'(1396);
			11976: out = 24'(1436);
			11977: out = 24'(1444);
			11978: out = 24'(1476);
			11979: out = 24'(1536);
			11980: out = 24'(1552);
			11981: out = 24'(1556);
			11982: out = 24'(1636);
			11983: out = 24'(1672);
			11984: out = 24'(1716);
			11985: out = 24'(1736);
			11986: out = 24'(1816);
			11987: out = 24'(1836);
			11988: out = 24'(1868);
			11989: out = 24'(1920);
			11990: out = 24'(1948);
			11991: out = 24'(2008);
			11992: out = 24'(2040);
			11993: out = 24'(2096);
			11994: out = 24'(2156);
			11995: out = 24'(2172);
			11996: out = 24'(2248);
			11997: out = 24'(2268);
			11998: out = 24'(2348);
			11999: out = 24'(2356);
			12000: out = 24'(2452);
			12001: out = 24'(2480);
			12002: out = 24'(2560);
			12003: out = 24'(2564);
			12004: out = 24'(2664);
			12005: out = 24'(2700);
			12006: out = 24'(2740);
			12007: out = 24'(2812);
			12008: out = 24'(2896);
			12009: out = 24'(2920);
			12010: out = 24'(2988);
			12011: out = 24'(3068);
			12012: out = 24'(3120);
			12013: out = 24'(3192);
			12014: out = 24'(3212);
			12015: out = 24'(3296);
			12016: out = 24'(3344);
			12017: out = 24'(3436);
			12018: out = 24'(3456);
			12019: out = 24'(3568);
			12020: out = 24'(3604);
			12021: out = 24'(3676);
			12022: out = 24'(3732);
			12023: out = 24'(3804);
			12024: out = 24'(3840);
			12025: out = 24'(3936);
			12026: out = 24'(3984);
			12027: out = 24'(4036);
			12028: out = 24'(4096);
			12029: out = 24'(4176);
			12030: out = 24'(4220);
			12031: out = 24'(4316);
			12032: out = 24'(4324);
			12033: out = 24'(4356);
			12034: out = 24'(4480);
			12035: out = 24'(4532);
			12036: out = 24'(4624);
			12037: out = 24'(4616);
			12038: out = 24'(4704);
			12039: out = 24'(4768);
			12040: out = 24'(4800);
			12041: out = 24'(4836);
			12042: out = 24'(4904);
			12043: out = 24'(4952);
			12044: out = 24'(5044);
			12045: out = 24'(5088);
			12046: out = 24'(5116);
			12047: out = 24'(5184);
			12048: out = 24'(5248);
			12049: out = 24'(5304);
			12050: out = 24'(5336);
			12051: out = 24'(5340);
			12052: out = 24'(5464);
			12053: out = 24'(5500);
			12054: out = 24'(5556);
			12055: out = 24'(5572);
			12056: out = 24'(5620);
			12057: out = 24'(5692);
			12058: out = 24'(5732);
			12059: out = 24'(5776);
			12060: out = 24'(5808);
			12061: out = 24'(5860);
			12062: out = 24'(5904);
			12063: out = 24'(5980);
			12064: out = 24'(6000);
			12065: out = 24'(6044);
			12066: out = 24'(6064);
			12067: out = 24'(6172);
			12068: out = 24'(6108);
			12069: out = 24'(6208);
			12070: out = 24'(6240);
			12071: out = 24'(6304);
			12072: out = 24'(6344);
			12073: out = 24'(6332);
			12074: out = 24'(6432);
			12075: out = 24'(6452);
			12076: out = 24'(6500);
			12077: out = 24'(6476);
			12078: out = 24'(6564);
			12079: out = 24'(6604);
			12080: out = 24'(6644);
			12081: out = 24'(6636);
			12082: out = 24'(6752);
			12083: out = 24'(6736);
			12084: out = 24'(6760);
			12085: out = 24'(6812);
			12086: out = 24'(6876);
			12087: out = 24'(6852);
			12088: out = 24'(6936);
			12089: out = 24'(6968);
			12090: out = 24'(6980);
			12091: out = 24'(7000);
			12092: out = 24'(7072);
			12093: out = 24'(7076);
			12094: out = 24'(7112);
			12095: out = 24'(7184);
			12096: out = 24'(7164);
			12097: out = 24'(7252);
			12098: out = 24'(7212);
			12099: out = 24'(7296);
			12100: out = 24'(7312);
			12101: out = 24'(7344);
			12102: out = 24'(7396);
			12103: out = 24'(7376);
			12104: out = 24'(7424);
			12105: out = 24'(7484);
			12106: out = 24'(7492);
			12107: out = 24'(7488);
			12108: out = 24'(7544);
			12109: out = 24'(7564);
			12110: out = 24'(7608);
			12111: out = 24'(7656);
			12112: out = 24'(7648);
			12113: out = 24'(7664);
			12114: out = 24'(7740);
			12115: out = 24'(7716);
			12116: out = 24'(7748);
			12117: out = 24'(7796);
			12118: out = 24'(7840);
			12119: out = 24'(7812);
			12120: out = 24'(7908);
			12121: out = 24'(7920);
			12122: out = 24'(7924);
			12123: out = 24'(7964);
			12124: out = 24'(7964);
			12125: out = 24'(8000);
			12126: out = 24'(8040);
			12127: out = 24'(8036);
			12128: out = 24'(8028);
			12129: out = 24'(8096);
			12130: out = 24'(8108);
			12131: out = 24'(8136);
			12132: out = 24'(8108);
			12133: out = 24'(8104);
			12134: out = 24'(8144);
			12135: out = 24'(8108);
			12136: out = 24'(8104);
			12137: out = 24'(8104);
			12138: out = 24'(8052);
			12139: out = 24'(8104);
			12140: out = 24'(8088);
			12141: out = 24'(8064);
			12142: out = 24'(8096);
			12143: out = 24'(8112);
			12144: out = 24'(8068);
			12145: out = 24'(8064);
			12146: out = 24'(8048);
			12147: out = 24'(8052);
			12148: out = 24'(8052);
			12149: out = 24'(8028);
			12150: out = 24'(8004);
			12151: out = 24'(8060);
			12152: out = 24'(8032);
			12153: out = 24'(8060);
			12154: out = 24'(8004);
			12155: out = 24'(8032);
			12156: out = 24'(8036);
			12157: out = 24'(8008);
			12158: out = 24'(8036);
			12159: out = 24'(8024);
			12160: out = 24'(8008);
			12161: out = 24'(8012);
			12162: out = 24'(8016);
			12163: out = 24'(7984);
			12164: out = 24'(8036);
			12165: out = 24'(8012);
			12166: out = 24'(8024);
			12167: out = 24'(8048);
			12168: out = 24'(8036);
			12169: out = 24'(8020);
			12170: out = 24'(7992);
			12171: out = 24'(8000);
			12172: out = 24'(8000);
			12173: out = 24'(7964);
			12174: out = 24'(8000);
			12175: out = 24'(7928);
			12176: out = 24'(7940);
			12177: out = 24'(8012);
			12178: out = 24'(7956);
			12179: out = 24'(7988);
			12180: out = 24'(7944);
			12181: out = 24'(7988);
			12182: out = 24'(7932);
			12183: out = 24'(7944);
			12184: out = 24'(7976);
			12185: out = 24'(7932);
			12186: out = 24'(7928);
			12187: out = 24'(7912);
			12188: out = 24'(7920);
			12189: out = 24'(7868);
			12190: out = 24'(7872);
			12191: out = 24'(7944);
			12192: out = 24'(7876);
			12193: out = 24'(7864);
			12194: out = 24'(7880);
			12195: out = 24'(7848);
			12196: out = 24'(7832);
			12197: out = 24'(7876);
			12198: out = 24'(7832);
			12199: out = 24'(7836);
			12200: out = 24'(7768);
			12201: out = 24'(7768);
			12202: out = 24'(7764);
			12203: out = 24'(7736);
			12204: out = 24'(7696);
			12205: out = 24'(7776);
			12206: out = 24'(7700);
			12207: out = 24'(7688);
			12208: out = 24'(7636);
			12209: out = 24'(7612);
			12210: out = 24'(7644);
			12211: out = 24'(7508);
			12212: out = 24'(7560);
			12213: out = 24'(7520);
			12214: out = 24'(7460);
			12215: out = 24'(7432);
			12216: out = 24'(7424);
			12217: out = 24'(7376);
			12218: out = 24'(7380);
			12219: out = 24'(7320);
			12220: out = 24'(7328);
			12221: out = 24'(7292);
			12222: out = 24'(7236);
			12223: out = 24'(7224);
			12224: out = 24'(7200);
			12225: out = 24'(7124);
			12226: out = 24'(7136);
			12227: out = 24'(7064);
			12228: out = 24'(6980);
			12229: out = 24'(6972);
			12230: out = 24'(6960);
			12231: out = 24'(6892);
			12232: out = 24'(6804);
			12233: out = 24'(6764);
			12234: out = 24'(6772);
			12235: out = 24'(6644);
			12236: out = 24'(6656);
			12237: out = 24'(6612);
			12238: out = 24'(6568);
			12239: out = 24'(6460);
			12240: out = 24'(6452);
			12241: out = 24'(6404);
			12242: out = 24'(6380);
			12243: out = 24'(6264);
			12244: out = 24'(6264);
			12245: out = 24'(6204);
			12246: out = 24'(6136);
			12247: out = 24'(6088);
			12248: out = 24'(6052);
			12249: out = 24'(6036);
			12250: out = 24'(5880);
			12251: out = 24'(5860);
			12252: out = 24'(5848);
			12253: out = 24'(5764);
			12254: out = 24'(5732);
			12255: out = 24'(5656);
			12256: out = 24'(5580);
			12257: out = 24'(5572);
			12258: out = 24'(5496);
			12259: out = 24'(5464);
			12260: out = 24'(5412);
			12261: out = 24'(5332);
			12262: out = 24'(5316);
			12263: out = 24'(5200);
			12264: out = 24'(5196);
			12265: out = 24'(5120);
			12266: out = 24'(5068);
			12267: out = 24'(5028);
			12268: out = 24'(4988);
			12269: out = 24'(4896);
			12270: out = 24'(4908);
			12271: out = 24'(4840);
			12272: out = 24'(4736);
			12273: out = 24'(4744);
			12274: out = 24'(4672);
			12275: out = 24'(4628);
			12276: out = 24'(4568);
			12277: out = 24'(4524);
			12278: out = 24'(4432);
			12279: out = 24'(4404);
			12280: out = 24'(4420);
			12281: out = 24'(4296);
			12282: out = 24'(4272);
			12283: out = 24'(4264);
			12284: out = 24'(4192);
			12285: out = 24'(4148);
			12286: out = 24'(4092);
			12287: out = 24'(4044);
			12288: out = 24'(3996);
			12289: out = 24'(3968);
			12290: out = 24'(3932);
			12291: out = 24'(3856);
			12292: out = 24'(3776);
			12293: out = 24'(3804);
			12294: out = 24'(3708);
			12295: out = 24'(3668);
			12296: out = 24'(3636);
			12297: out = 24'(3604);
			12298: out = 24'(3600);
			12299: out = 24'(3540);
			12300: out = 24'(3488);
			12301: out = 24'(3440);
			12302: out = 24'(3376);
			12303: out = 24'(3364);
			12304: out = 24'(3320);
			12305: out = 24'(3240);
			12306: out = 24'(3212);
			12307: out = 24'(3212);
			12308: out = 24'(3136);
			12309: out = 24'(3112);
			12310: out = 24'(3000);
			12311: out = 24'(3084);
			12312: out = 24'(2964);
			12313: out = 24'(2908);
			12314: out = 24'(2916);
			12315: out = 24'(2916);
			12316: out = 24'(2824);
			12317: out = 24'(2808);
			12318: out = 24'(2780);
			12319: out = 24'(2704);
			12320: out = 24'(2688);
			12321: out = 24'(2668);
			12322: out = 24'(2572);
			12323: out = 24'(2596);
			12324: out = 24'(2568);
			12325: out = 24'(2512);
			12326: out = 24'(2476);
			12327: out = 24'(2436);
			12328: out = 24'(2420);
			12329: out = 24'(2360);
			12330: out = 24'(2400);
			12331: out = 24'(2256);
			12332: out = 24'(2288);
			12333: out = 24'(2260);
			12334: out = 24'(2188);
			12335: out = 24'(2200);
			12336: out = 24'(2116);
			12337: out = 24'(2124);
			12338: out = 24'(2088);
			12339: out = 24'(2044);
			12340: out = 24'(2060);
			12341: out = 24'(2004);
			12342: out = 24'(1956);
			12343: out = 24'(1924);
			12344: out = 24'(1924);
			12345: out = 24'(1884);
			12346: out = 24'(1860);
			12347: out = 24'(1792);
			12348: out = 24'(1852);
			12349: out = 24'(1740);
			12350: out = 24'(1744);
			12351: out = 24'(1716);
			12352: out = 24'(1768);
			12353: out = 24'(1644);
			12354: out = 24'(1620);
			12355: out = 24'(1628);
			12356: out = 24'(1572);
			12357: out = 24'(1556);
			12358: out = 24'(1540);
			12359: out = 24'(1504);
			12360: out = 24'(1476);
			12361: out = 24'(1484);
			12362: out = 24'(1440);
			12363: out = 24'(1388);
			12364: out = 24'(1328);
			12365: out = 24'(1244);
			12366: out = 24'(1188);
			12367: out = 24'(1140);
			12368: out = 24'(1048);
			12369: out = 24'(988);
			12370: out = 24'(928);
			12371: out = 24'(892);
			12372: out = 24'(796);
			12373: out = 24'(728);
			12374: out = 24'(720);
			12375: out = 24'(628);
			12376: out = 24'(624);
			12377: out = 24'(468);
			12378: out = 24'(480);
			12379: out = 24'(404);
			12380: out = 24'(356);
			12381: out = 24'(340);
			12382: out = 24'(240);
			12383: out = 24'(216);
			12384: out = 24'(196);
			12385: out = 24'(60);
			12386: out = 24'(72);
			12387: out = 24'(28);
			12388: out = 24'(-60);
			12389: out = 24'(-88);
			12390: out = 24'(-116);
			12391: out = 24'(-180);
			12392: out = 24'(-208);
			12393: out = 24'(-276);
			12394: out = 24'(-332);
			12395: out = 24'(-384);
			12396: out = 24'(-356);
			12397: out = 24'(-456);
			12398: out = 24'(-512);
			12399: out = 24'(-544);
			12400: out = 24'(-588);
			12401: out = 24'(-632);
			12402: out = 24'(-676);
			12403: out = 24'(-700);
			12404: out = 24'(-768);
			12405: out = 24'(-744);
			12406: out = 24'(-840);
			12407: out = 24'(-864);
			12408: out = 24'(-872);
			12409: out = 24'(-988);
			12410: out = 24'(-976);
			12411: out = 24'(-1016);
			12412: out = 24'(-1052);
			12413: out = 24'(-1112);
			12414: out = 24'(-1164);
			12415: out = 24'(-1176);
			12416: out = 24'(-1196);
			12417: out = 24'(-1284);
			12418: out = 24'(-1284);
			12419: out = 24'(-1348);
			12420: out = 24'(-1344);
			12421: out = 24'(-1408);
			12422: out = 24'(-1440);
			12423: out = 24'(-1480);
			12424: out = 24'(-1516);
			12425: out = 24'(-1568);
			12426: out = 24'(-1600);
			12427: out = 24'(-1628);
			12428: out = 24'(-1668);
			12429: out = 24'(-1708);
			12430: out = 24'(-1772);
			12431: out = 24'(-1756);
			12432: out = 24'(-1852);
			12433: out = 24'(-1840);
			12434: out = 24'(-1860);
			12435: out = 24'(-1928);
			12436: out = 24'(-2008);
			12437: out = 24'(-1960);
			12438: out = 24'(-2060);
			12439: out = 24'(-2092);
			12440: out = 24'(-2104);
			12441: out = 24'(-2152);
			12442: out = 24'(-2228);
			12443: out = 24'(-2204);
			12444: out = 24'(-2288);
			12445: out = 24'(-2308);
			12446: out = 24'(-2336);
			12447: out = 24'(-2420);
			12448: out = 24'(-2440);
			12449: out = 24'(-2488);
			12450: out = 24'(-2520);
			12451: out = 24'(-2544);
			12452: out = 24'(-2620);
			12453: out = 24'(-2672);
			12454: out = 24'(-2680);
			12455: out = 24'(-2752);
			12456: out = 24'(-2776);
			12457: out = 24'(-2824);
			12458: out = 24'(-2900);
			12459: out = 24'(-2948);
			12460: out = 24'(-2992);
			12461: out = 24'(-3036);
			12462: out = 24'(-3048);
			12463: out = 24'(-3136);
			12464: out = 24'(-3180);
			12465: out = 24'(-3204);
			12466: out = 24'(-3320);
			12467: out = 24'(-3336);
			12468: out = 24'(-3380);
			12469: out = 24'(-3456);
			12470: out = 24'(-3524);
			12471: out = 24'(-3528);
			12472: out = 24'(-3668);
			12473: out = 24'(-3648);
			12474: out = 24'(-3756);
			12475: out = 24'(-3792);
			12476: out = 24'(-3912);
			12477: out = 24'(-3916);
			12478: out = 24'(-3992);
			12479: out = 24'(-4080);
			12480: out = 24'(-4132);
			12481: out = 24'(-4224);
			12482: out = 24'(-4248);
			12483: out = 24'(-4340);
			12484: out = 24'(-4360);
			12485: out = 24'(-4468);
			12486: out = 24'(-4520);
			12487: out = 24'(-4580);
			12488: out = 24'(-4752);
			12489: out = 24'(-4736);
			12490: out = 24'(-4864);
			12491: out = 24'(-4900);
			12492: out = 24'(-5008);
			12493: out = 24'(-5048);
			12494: out = 24'(-5136);
			12495: out = 24'(-5184);
			12496: out = 24'(-5248);
			12497: out = 24'(-5368);
			12498: out = 24'(-5400);
			12499: out = 24'(-5504);
			12500: out = 24'(-5556);
			12501: out = 24'(-5660);
			12502: out = 24'(-5696);
			12503: out = 24'(-5796);
			12504: out = 24'(-5836);
			12505: out = 24'(-5940);
			12506: out = 24'(-5972);
			12507: out = 24'(-6048);
			12508: out = 24'(-6116);
			12509: out = 24'(-6188);
			12510: out = 24'(-6256);
			12511: out = 24'(-6280);
			12512: out = 24'(-6396);
			12513: out = 24'(-6428);
			12514: out = 24'(-6468);
			12515: out = 24'(-6612);
			12516: out = 24'(-6616);
			12517: out = 24'(-6648);
			12518: out = 24'(-6748);
			12519: out = 24'(-6788);
			12520: out = 24'(-6836);
			12521: out = 24'(-6844);
			12522: out = 24'(-6928);
			12523: out = 24'(-7028);
			12524: out = 24'(-7044);
			12525: out = 24'(-7056);
			12526: out = 24'(-7172);
			12527: out = 24'(-7196);
			12528: out = 24'(-7208);
			12529: out = 24'(-7272);
			12530: out = 24'(-7300);
			12531: out = 24'(-7360);
			12532: out = 24'(-7340);
			12533: out = 24'(-7448);
			12534: out = 24'(-7460);
			12535: out = 24'(-7496);
			12536: out = 24'(-7520);
			12537: out = 24'(-7540);
			12538: out = 24'(-7632);
			12539: out = 24'(-7616);
			12540: out = 24'(-7640);
			12541: out = 24'(-7664);
			12542: out = 24'(-7732);
			12543: out = 24'(-7728);
			12544: out = 24'(-7780);
			12545: out = 24'(-7752);
			12546: out = 24'(-7844);
			12547: out = 24'(-7844);
			12548: out = 24'(-7840);
			12549: out = 24'(-7896);
			12550: out = 24'(-7908);
			12551: out = 24'(-7908);
			12552: out = 24'(-7976);
			12553: out = 24'(-7936);
			12554: out = 24'(-7980);
			12555: out = 24'(-8008);
			12556: out = 24'(-7968);
			12557: out = 24'(-8056);
			12558: out = 24'(-8036);
			12559: out = 24'(-8048);
			12560: out = 24'(-8068);
			12561: out = 24'(-8080);
			12562: out = 24'(-8072);
			12563: out = 24'(-8120);
			12564: out = 24'(-8088);
			12565: out = 24'(-8116);
			12566: out = 24'(-8100);
			12567: out = 24'(-8164);
			12568: out = 24'(-8096);
			12569: out = 24'(-8176);
			12570: out = 24'(-8088);
			12571: out = 24'(-8164);
			12572: out = 24'(-8164);
			12573: out = 24'(-8128);
			12574: out = 24'(-8148);
			12575: out = 24'(-8184);
			12576: out = 24'(-8160);
			12577: out = 24'(-8156);
			12578: out = 24'(-8156);
			12579: out = 24'(-8196);
			12580: out = 24'(-8164);
			12581: out = 24'(-8160);
			12582: out = 24'(-8152);
			12583: out = 24'(-8172);
			12584: out = 24'(-8156);
			12585: out = 24'(-8156);
			12586: out = 24'(-8100);
			12587: out = 24'(-8176);
			12588: out = 24'(-8124);
			12589: out = 24'(-8112);
			12590: out = 24'(-8132);
			12591: out = 24'(-8112);
			12592: out = 24'(-8124);
			12593: out = 24'(-8100);
			12594: out = 24'(-8116);
			12595: out = 24'(-8068);
			12596: out = 24'(-8084);
			12597: out = 24'(-8060);
			12598: out = 24'(-8072);
			12599: out = 24'(-8012);
			12600: out = 24'(-8100);
			12601: out = 24'(-8012);
			12602: out = 24'(-8024);
			12603: out = 24'(-8024);
			12604: out = 24'(-7980);
			12605: out = 24'(-8012);
			12606: out = 24'(-7984);
			12607: out = 24'(-7948);
			12608: out = 24'(-7964);
			12609: out = 24'(-7896);
			12610: out = 24'(-7956);
			12611: out = 24'(-7900);
			12612: out = 24'(-7932);
			12613: out = 24'(-7888);
			12614: out = 24'(-7860);
			12615: out = 24'(-7872);
			12616: out = 24'(-7852);
			12617: out = 24'(-7844);
			12618: out = 24'(-7796);
			12619: out = 24'(-7824);
			12620: out = 24'(-7784);
			12621: out = 24'(-7764);
			12622: out = 24'(-7764);
			12623: out = 24'(-7736);
			12624: out = 24'(-7744);
			12625: out = 24'(-7728);
			12626: out = 24'(-7684);
			12627: out = 24'(-7692);
			12628: out = 24'(-7660);
			12629: out = 24'(-7656);
			12630: out = 24'(-7636);
			12631: out = 24'(-7584);
			12632: out = 24'(-7592);
			12633: out = 24'(-7600);
			12634: out = 24'(-7544);
			12635: out = 24'(-7516);
			12636: out = 24'(-7540);
			12637: out = 24'(-7508);
			12638: out = 24'(-7456);
			12639: out = 24'(-7492);
			12640: out = 24'(-7444);
			12641: out = 24'(-7372);
			12642: out = 24'(-7448);
			12643: out = 24'(-7364);
			12644: out = 24'(-7388);
			12645: out = 24'(-7300);
			12646: out = 24'(-7344);
			12647: out = 24'(-7292);
			12648: out = 24'(-7276);
			12649: out = 24'(-7228);
			12650: out = 24'(-7260);
			12651: out = 24'(-7172);
			12652: out = 24'(-7180);
			12653: out = 24'(-7168);
			12654: out = 24'(-7112);
			12655: out = 24'(-7108);
			12656: out = 24'(-7072);
			12657: out = 24'(-7064);
			12658: out = 24'(-7000);
			12659: out = 24'(-7008);
			12660: out = 24'(-6992);
			12661: out = 24'(-6932);
			12662: out = 24'(-6884);
			12663: out = 24'(-6892);
			12664: out = 24'(-6864);
			12665: out = 24'(-6836);
			12666: out = 24'(-6772);
			12667: out = 24'(-6776);
			12668: out = 24'(-6716);
			12669: out = 24'(-6712);
			12670: out = 24'(-6648);
			12671: out = 24'(-6640);
			12672: out = 24'(-6568);
			12673: out = 24'(-6560);
			12674: out = 24'(-6500);
			12675: out = 24'(-6456);
			12676: out = 24'(-6432);
			12677: out = 24'(-6380);
			12678: out = 24'(-6348);
			12679: out = 24'(-6272);
			12680: out = 24'(-6252);
			12681: out = 24'(-6196);
			12682: out = 24'(-6156);
			12683: out = 24'(-6096);
			12684: out = 24'(-6052);
			12685: out = 24'(-5992);
			12686: out = 24'(-5976);
			12687: out = 24'(-5892);
			12688: out = 24'(-5884);
			12689: out = 24'(-5776);
			12690: out = 24'(-5736);
			12691: out = 24'(-5732);
			12692: out = 24'(-5624);
			12693: out = 24'(-5596);
			12694: out = 24'(-5548);
			12695: out = 24'(-5520);
			12696: out = 24'(-5404);
			12697: out = 24'(-5372);
			12698: out = 24'(-5356);
			12699: out = 24'(-5268);
			12700: out = 24'(-5196);
			12701: out = 24'(-5164);
			12702: out = 24'(-5100);
			12703: out = 24'(-5028);
			12704: out = 24'(-4984);
			12705: out = 24'(-4900);
			12706: out = 24'(-4884);
			12707: out = 24'(-4852);
			12708: out = 24'(-4748);
			12709: out = 24'(-4676);
			12710: out = 24'(-4660);
			12711: out = 24'(-4600);
			12712: out = 24'(-4532);
			12713: out = 24'(-4452);
			12714: out = 24'(-4436);
			12715: out = 24'(-4376);
			12716: out = 24'(-4324);
			12717: out = 24'(-4252);
			12718: out = 24'(-4224);
			12719: out = 24'(-4128);
			12720: out = 24'(-4084);
			12721: out = 24'(-4080);
			12722: out = 24'(-3956);
			12723: out = 24'(-3960);
			12724: out = 24'(-3892);
			12725: out = 24'(-3856);
			12726: out = 24'(-3748);
			12727: out = 24'(-3792);
			12728: out = 24'(-3668);
			12729: out = 24'(-3632);
			12730: out = 24'(-3580);
			12731: out = 24'(-3508);
			12732: out = 24'(-3520);
			12733: out = 24'(-3432);
			12734: out = 24'(-3424);
			12735: out = 24'(-3332);
			12736: out = 24'(-3300);
			12737: out = 24'(-3268);
			12738: out = 24'(-3208);
			12739: out = 24'(-3128);
			12740: out = 24'(-3136);
			12741: out = 24'(-3068);
			12742: out = 24'(-3008);
			12743: out = 24'(-2972);
			12744: out = 24'(-2952);
			12745: out = 24'(-2912);
			12746: out = 24'(-2832);
			12747: out = 24'(-2800);
			12748: out = 24'(-2796);
			12749: out = 24'(-2716);
			12750: out = 24'(-2676);
			12751: out = 24'(-2664);
			12752: out = 24'(-2624);
			12753: out = 24'(-2532);
			12754: out = 24'(-2536);
			12755: out = 24'(-2484);
			12756: out = 24'(-2424);
			12757: out = 24'(-2356);
			12758: out = 24'(-2416);
			12759: out = 24'(-2304);
			12760: out = 24'(-2348);
			12761: out = 24'(-2208);
			12762: out = 24'(-2256);
			12763: out = 24'(-2220);
			12764: out = 24'(-2136);
			12765: out = 24'(-2124);
			12766: out = 24'(-2088);
			12767: out = 24'(-2084);
			12768: out = 24'(-2008);
			12769: out = 24'(-1992);
			12770: out = 24'(-1936);
			12771: out = 24'(-1932);
			12772: out = 24'(-1872);
			12773: out = 24'(-1888);
			12774: out = 24'(-1828);
			12775: out = 24'(-1800);
			12776: out = 24'(-1760);
			12777: out = 24'(-1764);
			12778: out = 24'(-1680);
			12779: out = 24'(-1696);
			12780: out = 24'(-1652);
			12781: out = 24'(-1596);
			12782: out = 24'(-1620);
			12783: out = 24'(-1600);
			12784: out = 24'(-1496);
			12785: out = 24'(-1524);
			12786: out = 24'(-1492);
			12787: out = 24'(-1432);
			12788: out = 24'(-1396);
			12789: out = 24'(-1360);
			12790: out = 24'(-1320);
			12791: out = 24'(-1200);
			12792: out = 24'(-1240);
			12793: out = 24'(-1152);
			12794: out = 24'(-1108);
			12795: out = 24'(-1068);
			12796: out = 24'(-1052);
			12797: out = 24'(-984);
			12798: out = 24'(-964);
			12799: out = 24'(-932);
			12800: out = 24'(-884);
			12801: out = 24'(-796);
			12802: out = 24'(-792);
			12803: out = 24'(-764);
			12804: out = 24'(-732);
			12805: out = 24'(-644);
			12806: out = 24'(-652);
			12807: out = 24'(-596);
			12808: out = 24'(-564);
			12809: out = 24'(-552);
			12810: out = 24'(-524);
			12811: out = 24'(-448);
			12812: out = 24'(-440);
			12813: out = 24'(-368);
			12814: out = 24'(-380);
			12815: out = 24'(-336);
			12816: out = 24'(-276);
			12817: out = 24'(-288);
			12818: out = 24'(-212);
			12819: out = 24'(-216);
			12820: out = 24'(-176);
			12821: out = 24'(-164);
			12822: out = 24'(-80);
			12823: out = 24'(-76);
			12824: out = 24'(-60);
			12825: out = 24'(-12);
			12826: out = 24'(4);
			12827: out = 24'(12);
			12828: out = 24'(76);
			12829: out = 24'(104);
			12830: out = 24'(124);
			12831: out = 24'(160);
			12832: out = 24'(144);
			12833: out = 24'(248);
			12834: out = 24'(216);
			12835: out = 24'(264);
			12836: out = 24'(304);
			12837: out = 24'(292);
			12838: out = 24'(332);
			12839: out = 24'(396);
			12840: out = 24'(404);
			12841: out = 24'(432);
			12842: out = 24'(456);
			12843: out = 24'(476);
			12844: out = 24'(480);
			12845: out = 24'(552);
			12846: out = 24'(508);
			12847: out = 24'(592);
			12848: out = 24'(592);
			12849: out = 24'(620);
			12850: out = 24'(672);
			12851: out = 24'(672);
			12852: out = 24'(736);
			12853: out = 24'(700);
			12854: out = 24'(792);
			12855: out = 24'(748);
			12856: out = 24'(816);
			12857: out = 24'(816);
			12858: out = 24'(868);
			12859: out = 24'(880);
			12860: out = 24'(956);
			12861: out = 24'(920);
			12862: out = 24'(996);
			12863: out = 24'(996);
			12864: out = 24'(1028);
			12865: out = 24'(1076);
			12866: out = 24'(1092);
			12867: out = 24'(1096);
			12868: out = 24'(1132);
			12869: out = 24'(1216);
			12870: out = 24'(1176);
			12871: out = 24'(1220);
			12872: out = 24'(1264);
			12873: out = 24'(1320);
			12874: out = 24'(1300);
			12875: out = 24'(1364);
			12876: out = 24'(1396);
			12877: out = 24'(1448);
			12878: out = 24'(1472);
			12879: out = 24'(1460);
			12880: out = 24'(1524);
			12881: out = 24'(1564);
			12882: out = 24'(1632);
			12883: out = 24'(1632);
			12884: out = 24'(1632);
			12885: out = 24'(1724);
			12886: out = 24'(1736);
			12887: out = 24'(1824);
			12888: out = 24'(1776);
			12889: out = 24'(1868);
			12890: out = 24'(1920);
			12891: out = 24'(1996);
			12892: out = 24'(1972);
			12893: out = 24'(2060);
			12894: out = 24'(2088);
			12895: out = 24'(2140);
			12896: out = 24'(2152);
			12897: out = 24'(2228);
			12898: out = 24'(2232);
			12899: out = 24'(2340);
			12900: out = 24'(2356);
			12901: out = 24'(2408);
			12902: out = 24'(2472);
			12903: out = 24'(2492);
			12904: out = 24'(2576);
			12905: out = 24'(2580);
			12906: out = 24'(2668);
			12907: out = 24'(2684);
			12908: out = 24'(2736);
			12909: out = 24'(2788);
			12910: out = 24'(2888);
			12911: out = 24'(2904);
			12912: out = 24'(2936);
			12913: out = 24'(3012);
			12914: out = 24'(3056);
			12915: out = 24'(3084);
			12916: out = 24'(3172);
			12917: out = 24'(3192);
			12918: out = 24'(3240);
			12919: out = 24'(3332);
			12920: out = 24'(3324);
			12921: out = 24'(3416);
			12922: out = 24'(3416);
			12923: out = 24'(3512);
			12924: out = 24'(3576);
			12925: out = 24'(3576);
			12926: out = 24'(3636);
			12927: out = 24'(3700);
			12928: out = 24'(3772);
			12929: out = 24'(3760);
			12930: out = 24'(3840);
			12931: out = 24'(3856);
			12932: out = 24'(3972);
			12933: out = 24'(3912);
			12934: out = 24'(4028);
			12935: out = 24'(4048);
			12936: out = 24'(4112);
			12937: out = 24'(4132);
			12938: out = 24'(4204);
			12939: out = 24'(4236);
			12940: out = 24'(4284);
			12941: out = 24'(4332);
			12942: out = 24'(4316);
			12943: out = 24'(4432);
			12944: out = 24'(4384);
			12945: out = 24'(4484);
			12946: out = 24'(4480);
			12947: out = 24'(4548);
			12948: out = 24'(4576);
			12949: out = 24'(4584);
			12950: out = 24'(4676);
			12951: out = 24'(4664);
			12952: out = 24'(4752);
			12953: out = 24'(4736);
			12954: out = 24'(4808);
			12955: out = 24'(4840);
			12956: out = 24'(4876);
			12957: out = 24'(4876);
			12958: out = 24'(4944);
			12959: out = 24'(4956);
			12960: out = 24'(4996);
			12961: out = 24'(5028);
			12962: out = 24'(5096);
			12963: out = 24'(5068);
			12964: out = 24'(5136);
			12965: out = 24'(5176);
			12966: out = 24'(5172);
			12967: out = 24'(5256);
			12968: out = 24'(5236);
			12969: out = 24'(5308);
			12970: out = 24'(5304);
			12971: out = 24'(5320);
			12972: out = 24'(5392);
			12973: out = 24'(5408);
			12974: out = 24'(5432);
			12975: out = 24'(5464);
			12976: out = 24'(5504);
			12977: out = 24'(5480);
			12978: out = 24'(5596);
			12979: out = 24'(5564);
			12980: out = 24'(5612);
			12981: out = 24'(5620);
			12982: out = 24'(5664);
			12983: out = 24'(5700);
			12984: out = 24'(5688);
			12985: out = 24'(5764);
			12986: out = 24'(5736);
			12987: out = 24'(5800);
			12988: out = 24'(5796);
			12989: out = 24'(5848);
			12990: out = 24'(5876);
			12991: out = 24'(5856);
			12992: out = 24'(5924);
			12993: out = 24'(5924);
			12994: out = 24'(5968);
			12995: out = 24'(5972);
			12996: out = 24'(6012);
			12997: out = 24'(6020);
			12998: out = 24'(6084);
			12999: out = 24'(6068);
			13000: out = 24'(6080);
			13001: out = 24'(6120);
			13002: out = 24'(6176);
			13003: out = 24'(6156);
			13004: out = 24'(6172);
			13005: out = 24'(6252);
			13006: out = 24'(6220);
			13007: out = 24'(6232);
			13008: out = 24'(6300);
			13009: out = 24'(6280);
			13010: out = 24'(6328);
			13011: out = 24'(6336);
			13012: out = 24'(6364);
			13013: out = 24'(6392);
			13014: out = 24'(6404);
			13015: out = 24'(6396);
			13016: out = 24'(6456);
			13017: out = 24'(6464);
			13018: out = 24'(6492);
			13019: out = 24'(6496);
			13020: out = 24'(6480);
			13021: out = 24'(6512);
			13022: out = 24'(6512);
			13023: out = 24'(6520);
			13024: out = 24'(6512);
			13025: out = 24'(6524);
			13026: out = 24'(6512);
			13027: out = 24'(6504);
			13028: out = 24'(6508);
			13029: out = 24'(6520);
			13030: out = 24'(6512);
			13031: out = 24'(6548);
			13032: out = 24'(6536);
			13033: out = 24'(6492);
			13034: out = 24'(6472);
			13035: out = 24'(6528);
			13036: out = 24'(6416);
			13037: out = 24'(6464);
			13038: out = 24'(6496);
			13039: out = 24'(6468);
			13040: out = 24'(6472);
			13041: out = 24'(6452);
			13042: out = 24'(6448);
			13043: out = 24'(6476);
			13044: out = 24'(6480);
			13045: out = 24'(6444);
			13046: out = 24'(6460);
			13047: out = 24'(6408);
			13048: out = 24'(6488);
			13049: out = 24'(6496);
			13050: out = 24'(6404);
			13051: out = 24'(6488);
			13052: out = 24'(6492);
			13053: out = 24'(6504);
			13054: out = 24'(6412);
			13055: out = 24'(6424);
			13056: out = 24'(6448);
			13057: out = 24'(6448);
			13058: out = 24'(6428);
			13059: out = 24'(6428);
			13060: out = 24'(6472);
			13061: out = 24'(6500);
			13062: out = 24'(6496);
			13063: out = 24'(6460);
			13064: out = 24'(6472);
			13065: out = 24'(6464);
			13066: out = 24'(6356);
			13067: out = 24'(6400);
			13068: out = 24'(6444);
			13069: out = 24'(6392);
			13070: out = 24'(6372);
			13071: out = 24'(6420);
			13072: out = 24'(6428);
			13073: out = 24'(6400);
			13074: out = 24'(6420);
			13075: out = 24'(6440);
			13076: out = 24'(6396);
			13077: out = 24'(6400);
			13078: out = 24'(6404);
			13079: out = 24'(6348);
			13080: out = 24'(6428);
			13081: out = 24'(6352);
			13082: out = 24'(6372);
			13083: out = 24'(6368);
			13084: out = 24'(6304);
			13085: out = 24'(6380);
			13086: out = 24'(6324);
			13087: out = 24'(6344);
			13088: out = 24'(6324);
			13089: out = 24'(6324);
			13090: out = 24'(6304);
			13091: out = 24'(6296);
			13092: out = 24'(6280);
			13093: out = 24'(6268);
			13094: out = 24'(6220);
			13095: out = 24'(6244);
			13096: out = 24'(6264);
			13097: out = 24'(6216);
			13098: out = 24'(6216);
			13099: out = 24'(6160);
			13100: out = 24'(6192);
			13101: out = 24'(6164);
			13102: out = 24'(6092);
			13103: out = 24'(6088);
			13104: out = 24'(6072);
			13105: out = 24'(6060);
			13106: out = 24'(6052);
			13107: out = 24'(5968);
			13108: out = 24'(6000);
			13109: out = 24'(5936);
			13110: out = 24'(5920);
			13111: out = 24'(5920);
			13112: out = 24'(5912);
			13113: out = 24'(5816);
			13114: out = 24'(5832);
			13115: out = 24'(5804);
			13116: out = 24'(5740);
			13117: out = 24'(5740);
			13118: out = 24'(5688);
			13119: out = 24'(5620);
			13120: out = 24'(5640);
			13121: out = 24'(5576);
			13122: out = 24'(5548);
			13123: out = 24'(5540);
			13124: out = 24'(5456);
			13125: out = 24'(5456);
			13126: out = 24'(5376);
			13127: out = 24'(5388);
			13128: out = 24'(5328);
			13129: out = 24'(5280);
			13130: out = 24'(5212);
			13131: out = 24'(5192);
			13132: out = 24'(5176);
			13133: out = 24'(5096);
			13134: out = 24'(5052);
			13135: out = 24'(5056);
			13136: out = 24'(4976);
			13137: out = 24'(4948);
			13138: out = 24'(4896);
			13139: out = 24'(4848);
			13140: out = 24'(4816);
			13141: out = 24'(4756);
			13142: out = 24'(4708);
			13143: out = 24'(4692);
			13144: out = 24'(4628);
			13145: out = 24'(4628);
			13146: out = 24'(4524);
			13147: out = 24'(4472);
			13148: out = 24'(4476);
			13149: out = 24'(4388);
			13150: out = 24'(4376);
			13151: out = 24'(4364);
			13152: out = 24'(4236);
			13153: out = 24'(4268);
			13154: out = 24'(4188);
			13155: out = 24'(4152);
			13156: out = 24'(4092);
			13157: out = 24'(4072);
			13158: out = 24'(4036);
			13159: out = 24'(3952);
			13160: out = 24'(3956);
			13161: out = 24'(3900);
			13162: out = 24'(3852);
			13163: out = 24'(3812);
			13164: out = 24'(3812);
			13165: out = 24'(3724);
			13166: out = 24'(3684);
			13167: out = 24'(3636);
			13168: out = 24'(3560);
			13169: out = 24'(3588);
			13170: out = 24'(3508);
			13171: out = 24'(3432);
			13172: out = 24'(3448);
			13173: out = 24'(3392);
			13174: out = 24'(3392);
			13175: out = 24'(3272);
			13176: out = 24'(3304);
			13177: out = 24'(3212);
			13178: out = 24'(3220);
			13179: out = 24'(3156);
			13180: out = 24'(3128);
			13181: out = 24'(3096);
			13182: out = 24'(3016);
			13183: out = 24'(3052);
			13184: out = 24'(2952);
			13185: out = 24'(2972);
			13186: out = 24'(2876);
			13187: out = 24'(2920);
			13188: out = 24'(2800);
			13189: out = 24'(2812);
			13190: out = 24'(2768);
			13191: out = 24'(2732);
			13192: out = 24'(2704);
			13193: out = 24'(2664);
			13194: out = 24'(2620);
			13195: out = 24'(2620);
			13196: out = 24'(2536);
			13197: out = 24'(2572);
			13198: out = 24'(2492);
			13199: out = 24'(2468);
			13200: out = 24'(2444);
			13201: out = 24'(2400);
			13202: out = 24'(2348);
			13203: out = 24'(2368);
			13204: out = 24'(2360);
			13205: out = 24'(2268);
			13206: out = 24'(2236);
			13207: out = 24'(2216);
			13208: out = 24'(2208);
			13209: out = 24'(2148);
			13210: out = 24'(2104);
			13211: out = 24'(2092);
			13212: out = 24'(2084);
			13213: out = 24'(2072);
			13214: out = 24'(1984);
			13215: out = 24'(1956);
			13216: out = 24'(1960);
			13217: out = 24'(1904);
			13218: out = 24'(1936);
			13219: out = 24'(1812);
			13220: out = 24'(1832);
			13221: out = 24'(1840);
			13222: out = 24'(1800);
			13223: out = 24'(1764);
			13224: out = 24'(1740);
			13225: out = 24'(1732);
			13226: out = 24'(1688);
			13227: out = 24'(1644);
			13228: out = 24'(1644);
			13229: out = 24'(1612);
			13230: out = 24'(1540);
			13231: out = 24'(1576);
			13232: out = 24'(1568);
			13233: out = 24'(1548);
			13234: out = 24'(1468);
			13235: out = 24'(1496);
			13236: out = 24'(1456);
			13237: out = 24'(1424);
			13238: out = 24'(1424);
			13239: out = 24'(1380);
			13240: out = 24'(1308);
			13241: out = 24'(1392);
			13242: out = 24'(1292);
			13243: out = 24'(1316);
			13244: out = 24'(1236);
			13245: out = 24'(1256);
			13246: out = 24'(1260);
			13247: out = 24'(1184);
			13248: out = 24'(1220);
			13249: out = 24'(1200);
			13250: out = 24'(1152);
			13251: out = 24'(1148);
			13252: out = 24'(1148);
			13253: out = 24'(1060);
			13254: out = 24'(1064);
			13255: out = 24'(1068);
			13256: out = 24'(904);
			13257: out = 24'(884);
			13258: out = 24'(876);
			13259: out = 24'(784);
			13260: out = 24'(768);
			13261: out = 24'(680);
			13262: out = 24'(648);
			13263: out = 24'(592);
			13264: out = 24'(596);
			13265: out = 24'(456);
			13266: out = 24'(480);
			13267: out = 24'(412);
			13268: out = 24'(348);
			13269: out = 24'(324);
			13270: out = 24'(288);
			13271: out = 24'(208);
			13272: out = 24'(248);
			13273: out = 24'(136);
			13274: out = 24'(132);
			13275: out = 24'(68);
			13276: out = 24'(20);
			13277: out = 24'(16);
			13278: out = 24'(-76);
			13279: out = 24'(-76);
			13280: out = 24'(-112);
			13281: out = 24'(-204);
			13282: out = 24'(-160);
			13283: out = 24'(-256);
			13284: out = 24'(-256);
			13285: out = 24'(-304);
			13286: out = 24'(-360);
			13287: out = 24'(-384);
			13288: out = 24'(-452);
			13289: out = 24'(-452);
			13290: out = 24'(-468);
			13291: out = 24'(-556);
			13292: out = 24'(-552);
			13293: out = 24'(-604);
			13294: out = 24'(-608);
			13295: out = 24'(-668);
			13296: out = 24'(-676);
			13297: out = 24'(-740);
			13298: out = 24'(-744);
			13299: out = 24'(-792);
			13300: out = 24'(-824);
			13301: out = 24'(-824);
			13302: out = 24'(-892);
			13303: out = 24'(-912);
			13304: out = 24'(-956);
			13305: out = 24'(-1000);
			13306: out = 24'(-1004);
			13307: out = 24'(-1036);
			13308: out = 24'(-1080);
			13309: out = 24'(-1072);
			13310: out = 24'(-1148);
			13311: out = 24'(-1144);
			13312: out = 24'(-1196);
			13313: out = 24'(-1232);
			13314: out = 24'(-1236);
			13315: out = 24'(-1248);
			13316: out = 24'(-1320);
			13317: out = 24'(-1340);
			13318: out = 24'(-1316);
			13319: out = 24'(-1392);
			13320: out = 24'(-1404);
			13321: out = 24'(-1472);
			13322: out = 24'(-1484);
			13323: out = 24'(-1508);
			13324: out = 24'(-1564);
			13325: out = 24'(-1564);
			13326: out = 24'(-1592);
			13327: out = 24'(-1628);
			13328: out = 24'(-1660);
			13329: out = 24'(-1664);
			13330: out = 24'(-1708);
			13331: out = 24'(-1728);
			13332: out = 24'(-1780);
			13333: out = 24'(-1800);
			13334: out = 24'(-1872);
			13335: out = 24'(-1864);
			13336: out = 24'(-1884);
			13337: out = 24'(-1968);
			13338: out = 24'(-1968);
			13339: out = 24'(-1992);
			13340: out = 24'(-2024);
			13341: out = 24'(-2088);
			13342: out = 24'(-2052);
			13343: out = 24'(-2120);
			13344: out = 24'(-2212);
			13345: out = 24'(-2196);
			13346: out = 24'(-2236);
			13347: out = 24'(-2308);
			13348: out = 24'(-2308);
			13349: out = 24'(-2388);
			13350: out = 24'(-2360);
			13351: out = 24'(-2440);
			13352: out = 24'(-2472);
			13353: out = 24'(-2516);
			13354: out = 24'(-2548);
			13355: out = 24'(-2588);
			13356: out = 24'(-2652);
			13357: out = 24'(-2708);
			13358: out = 24'(-2724);
			13359: out = 24'(-2740);
			13360: out = 24'(-2828);
			13361: out = 24'(-2868);
			13362: out = 24'(-2920);
			13363: out = 24'(-2944);
			13364: out = 24'(-3020);
			13365: out = 24'(-3040);
			13366: out = 24'(-3116);
			13367: out = 24'(-3152);
			13368: out = 24'(-3180);
			13369: out = 24'(-3288);
			13370: out = 24'(-3308);
			13371: out = 24'(-3384);
			13372: out = 24'(-3356);
			13373: out = 24'(-3524);
			13374: out = 24'(-3544);
			13375: out = 24'(-3560);
			13376: out = 24'(-3640);
			13377: out = 24'(-3676);
			13378: out = 24'(-3792);
			13379: out = 24'(-3800);
			13380: out = 24'(-3884);
			13381: out = 24'(-3888);
			13382: out = 24'(-4012);
			13383: out = 24'(-4040);
			13384: out = 24'(-4140);
			13385: out = 24'(-4132);
			13386: out = 24'(-4232);
			13387: out = 24'(-4312);
			13388: out = 24'(-4340);
			13389: out = 24'(-4408);
			13390: out = 24'(-4408);
			13391: out = 24'(-4572);
			13392: out = 24'(-4536);
			13393: out = 24'(-4632);
			13394: out = 24'(-4700);
			13395: out = 24'(-4756);
			13396: out = 24'(-4788);
			13397: out = 24'(-4848);
			13398: out = 24'(-4952);
			13399: out = 24'(-4976);
			13400: out = 24'(-4980);
			13401: out = 24'(-5116);
			13402: out = 24'(-5092);
			13403: out = 24'(-5184);
			13404: out = 24'(-5224);
			13405: out = 24'(-5264);
			13406: out = 24'(-5364);
			13407: out = 24'(-5296);
			13408: out = 24'(-5432);
			13409: out = 24'(-5448);
			13410: out = 24'(-5508);
			13411: out = 24'(-5496);
			13412: out = 24'(-5580);
			13413: out = 24'(-5640);
			13414: out = 24'(-5656);
			13415: out = 24'(-5676);
			13416: out = 24'(-5752);
			13417: out = 24'(-5804);
			13418: out = 24'(-5800);
			13419: out = 24'(-5860);
			13420: out = 24'(-5852);
			13421: out = 24'(-5952);
			13422: out = 24'(-5912);
			13423: out = 24'(-5984);
			13424: out = 24'(-6016);
			13425: out = 24'(-6020);
			13426: out = 24'(-6076);
			13427: out = 24'(-6092);
			13428: out = 24'(-6128);
			13429: out = 24'(-6156);
			13430: out = 24'(-6164);
			13431: out = 24'(-6216);
			13432: out = 24'(-6204);
			13433: out = 24'(-6252);
			13434: out = 24'(-6284);
			13435: out = 24'(-6284);
			13436: out = 24'(-6308);
			13437: out = 24'(-6320);
			13438: out = 24'(-6376);
			13439: out = 24'(-6364);
			13440: out = 24'(-6368);
			13441: out = 24'(-6408);
			13442: out = 24'(-6408);
			13443: out = 24'(-6448);
			13444: out = 24'(-6432);
			13445: out = 24'(-6452);
			13446: out = 24'(-6504);
			13447: out = 24'(-6452);
			13448: out = 24'(-6520);
			13449: out = 24'(-6508);
			13450: out = 24'(-6496);
			13451: out = 24'(-6560);
			13452: out = 24'(-6552);
			13453: out = 24'(-6508);
			13454: out = 24'(-6548);
			13455: out = 24'(-6580);
			13456: out = 24'(-6548);
			13457: out = 24'(-6560);
			13458: out = 24'(-6600);
			13459: out = 24'(-6592);
			13460: out = 24'(-6572);
			13461: out = 24'(-6616);
			13462: out = 24'(-6592);
			13463: out = 24'(-6604);
			13464: out = 24'(-6616);
			13465: out = 24'(-6600);
			13466: out = 24'(-6616);
			13467: out = 24'(-6608);
			13468: out = 24'(-6588);
			13469: out = 24'(-6656);
			13470: out = 24'(-6604);
			13471: out = 24'(-6612);
			13472: out = 24'(-6592);
			13473: out = 24'(-6592);
			13474: out = 24'(-6600);
			13475: out = 24'(-6604);
			13476: out = 24'(-6612);
			13477: out = 24'(-6592);
			13478: out = 24'(-6608);
			13479: out = 24'(-6628);
			13480: out = 24'(-6600);
			13481: out = 24'(-6588);
			13482: out = 24'(-6568);
			13483: out = 24'(-6608);
			13484: out = 24'(-6548);
			13485: out = 24'(-6580);
			13486: out = 24'(-6580);
			13487: out = 24'(-6528);
			13488: out = 24'(-6552);
			13489: out = 24'(-6556);
			13490: out = 24'(-6536);
			13491: out = 24'(-6544);
			13492: out = 24'(-6496);
			13493: out = 24'(-6536);
			13494: out = 24'(-6528);
			13495: out = 24'(-6480);
			13496: out = 24'(-6460);
			13497: out = 24'(-6500);
			13498: out = 24'(-6444);
			13499: out = 24'(-6452);
			13500: out = 24'(-6472);
			13501: out = 24'(-6428);
			13502: out = 24'(-6428);
			13503: out = 24'(-6476);
			13504: out = 24'(-6412);
			13505: out = 24'(-6380);
			13506: out = 24'(-6368);
			13507: out = 24'(-6412);
			13508: out = 24'(-6360);
			13509: out = 24'(-6332);
			13510: out = 24'(-6368);
			13511: out = 24'(-6320);
			13512: out = 24'(-6296);
			13513: out = 24'(-6320);
			13514: out = 24'(-6276);
			13515: out = 24'(-6284);
			13516: out = 24'(-6268);
			13517: out = 24'(-6244);
			13518: out = 24'(-6232);
			13519: out = 24'(-6228);
			13520: out = 24'(-6240);
			13521: out = 24'(-6148);
			13522: out = 24'(-6196);
			13523: out = 24'(-6180);
			13524: out = 24'(-6140);
			13525: out = 24'(-6128);
			13526: out = 24'(-6112);
			13527: out = 24'(-6156);
			13528: out = 24'(-6052);
			13529: out = 24'(-6108);
			13530: out = 24'(-6052);
			13531: out = 24'(-6076);
			13532: out = 24'(-6016);
			13533: out = 24'(-6012);
			13534: out = 24'(-6000);
			13535: out = 24'(-5984);
			13536: out = 24'(-5944);
			13537: out = 24'(-5944);
			13538: out = 24'(-5944);
			13539: out = 24'(-5928);
			13540: out = 24'(-5876);
			13541: out = 24'(-5892);
			13542: out = 24'(-5848);
			13543: out = 24'(-5848);
			13544: out = 24'(-5816);
			13545: out = 24'(-5788);
			13546: out = 24'(-5796);
			13547: out = 24'(-5740);
			13548: out = 24'(-5748);
			13549: out = 24'(-5716);
			13550: out = 24'(-5700);
			13551: out = 24'(-5652);
			13552: out = 24'(-5660);
			13553: out = 24'(-5600);
			13554: out = 24'(-5600);
			13555: out = 24'(-5552);
			13556: out = 24'(-5564);
			13557: out = 24'(-5496);
			13558: out = 24'(-5524);
			13559: out = 24'(-5468);
			13560: out = 24'(-5416);
			13561: out = 24'(-5420);
			13562: out = 24'(-5324);
			13563: out = 24'(-5364);
			13564: out = 24'(-5316);
			13565: out = 24'(-5268);
			13566: out = 24'(-5260);
			13567: out = 24'(-5196);
			13568: out = 24'(-5192);
			13569: out = 24'(-5140);
			13570: out = 24'(-5116);
			13571: out = 24'(-5060);
			13572: out = 24'(-5052);
			13573: out = 24'(-4964);
			13574: out = 24'(-4984);
			13575: out = 24'(-4952);
			13576: out = 24'(-4864);
			13577: out = 24'(-4832);
			13578: out = 24'(-4832);
			13579: out = 24'(-4724);
			13580: out = 24'(-4728);
			13581: out = 24'(-4696);
			13582: out = 24'(-4608);
			13583: out = 24'(-4596);
			13584: out = 24'(-4572);
			13585: out = 24'(-4504);
			13586: out = 24'(-4456);
			13587: out = 24'(-4388);
			13588: out = 24'(-4396);
			13589: out = 24'(-4308);
			13590: out = 24'(-4284);
			13591: out = 24'(-4240);
			13592: out = 24'(-4184);
			13593: out = 24'(-4148);
			13594: out = 24'(-4076);
			13595: out = 24'(-4060);
			13596: out = 24'(-4012);
			13597: out = 24'(-3956);
			13598: out = 24'(-3932);
			13599: out = 24'(-3860);
			13600: out = 24'(-3848);
			13601: out = 24'(-3760);
			13602: out = 24'(-3732);
			13603: out = 24'(-3720);
			13604: out = 24'(-3616);
			13605: out = 24'(-3612);
			13606: out = 24'(-3524);
			13607: out = 24'(-3528);
			13608: out = 24'(-3472);
			13609: out = 24'(-3432);
			13610: out = 24'(-3412);
			13611: out = 24'(-3332);
			13612: out = 24'(-3276);
			13613: out = 24'(-3280);
			13614: out = 24'(-3240);
			13615: out = 24'(-3152);
			13616: out = 24'(-3112);
			13617: out = 24'(-3084);
			13618: out = 24'(-3052);
			13619: out = 24'(-3016);
			13620: out = 24'(-2972);
			13621: out = 24'(-2912);
			13622: out = 24'(-2876);
			13623: out = 24'(-2856);
			13624: out = 24'(-2780);
			13625: out = 24'(-2796);
			13626: out = 24'(-2708);
			13627: out = 24'(-2708);
			13628: out = 24'(-2660);
			13629: out = 24'(-2620);
			13630: out = 24'(-2592);
			13631: out = 24'(-2512);
			13632: out = 24'(-2536);
			13633: out = 24'(-2468);
			13634: out = 24'(-2416);
			13635: out = 24'(-2416);
			13636: out = 24'(-2380);
			13637: out = 24'(-2328);
			13638: out = 24'(-2296);
			13639: out = 24'(-2288);
			13640: out = 24'(-2220);
			13641: out = 24'(-2180);
			13642: out = 24'(-2160);
			13643: out = 24'(-2156);
			13644: out = 24'(-2068);
			13645: out = 24'(-2104);
			13646: out = 24'(-2056);
			13647: out = 24'(-1980);
			13648: out = 24'(-1996);
			13649: out = 24'(-1948);
			13650: out = 24'(-1920);
			13651: out = 24'(-1904);
			13652: out = 24'(-1816);
			13653: out = 24'(-1832);
			13654: out = 24'(-1792);
			13655: out = 24'(-1784);
			13656: out = 24'(-1752);
			13657: out = 24'(-1684);
			13658: out = 24'(-1696);
			13659: out = 24'(-1660);
			13660: out = 24'(-1684);
			13661: out = 24'(-1592);
			13662: out = 24'(-1600);
			13663: out = 24'(-1580);
			13664: out = 24'(-1544);
			13665: out = 24'(-1508);
			13666: out = 24'(-1460);
			13667: out = 24'(-1500);
			13668: out = 24'(-1404);
			13669: out = 24'(-1416);
			13670: out = 24'(-1404);
			13671: out = 24'(-1368);
			13672: out = 24'(-1336);
			13673: out = 24'(-1356);
			13674: out = 24'(-1272);
			13675: out = 24'(-1328);
			13676: out = 24'(-1216);
			13677: out = 24'(-1268);
			13678: out = 24'(-1212);
			13679: out = 24'(-1164);
			13680: out = 24'(-1124);
			13681: out = 24'(-1116);
			13682: out = 24'(-1056);
			13683: out = 24'(-996);
			13684: out = 24'(-988);
			13685: out = 24'(-960);
			13686: out = 24'(-924);
			13687: out = 24'(-868);
			13688: out = 24'(-836);
			13689: out = 24'(-832);
			13690: out = 24'(-800);
			13691: out = 24'(-744);
			13692: out = 24'(-712);
			13693: out = 24'(-656);
			13694: out = 24'(-684);
			13695: out = 24'(-588);
			13696: out = 24'(-584);
			13697: out = 24'(-580);
			13698: out = 24'(-536);
			13699: out = 24'(-476);
			13700: out = 24'(-456);
			13701: out = 24'(-448);
			13702: out = 24'(-436);
			13703: out = 24'(-380);
			13704: out = 24'(-356);
			13705: out = 24'(-320);
			13706: out = 24'(-344);
			13707: out = 24'(-276);
			13708: out = 24'(-224);
			13709: out = 24'(-216);
			13710: out = 24'(-208);
			13711: out = 24'(-156);
			13712: out = 24'(-168);
			13713: out = 24'(-128);
			13714: out = 24'(-68);
			13715: out = 24'(-108);
			13716: out = 24'(-40);
			13717: out = 24'(-20);
			13718: out = 24'(0);
			13719: out = 24'(28);
			13720: out = 24'(-20);
			13721: out = 24'(104);
			13722: out = 24'(96);
			13723: out = 24'(100);
			13724: out = 24'(108);
			13725: out = 24'(196);
			13726: out = 24'(152);
			13727: out = 24'(212);
			13728: out = 24'(228);
			13729: out = 24'(232);
			13730: out = 24'(280);
			13731: out = 24'(288);
			13732: out = 24'(296);
			13733: out = 24'(344);
			13734: out = 24'(356);
			13735: out = 24'(380);
			13736: out = 24'(400);
			13737: out = 24'(396);
			13738: out = 24'(464);
			13739: out = 24'(468);
			13740: out = 24'(452);
			13741: out = 24'(492);
			13742: out = 24'(536);
			13743: out = 24'(544);
			13744: out = 24'(556);
			13745: out = 24'(564);
			13746: out = 24'(680);
			13747: out = 24'(588);
			13748: out = 24'(656);
			13749: out = 24'(688);
			13750: out = 24'(704);
			13751: out = 24'(688);
			13752: out = 24'(776);
			13753: out = 24'(736);
			13754: out = 24'(800);
			13755: out = 24'(780);
			13756: out = 24'(824);
			13757: out = 24'(844);
			13758: out = 24'(872);
			13759: out = 24'(888);
			13760: out = 24'(920);
			13761: out = 24'(956);
			13762: out = 24'(952);
			13763: out = 24'(1016);
			13764: out = 24'(1028);
			13765: out = 24'(1020);
			13766: out = 24'(1084);
			13767: out = 24'(1116);
			13768: out = 24'(1056);
			13769: out = 24'(1200);
			13770: out = 24'(1152);
			13771: out = 24'(1248);
			13772: out = 24'(1224);
			13773: out = 24'(1256);
			13774: out = 24'(1312);
			13775: out = 24'(1300);
			13776: out = 24'(1392);
			13777: out = 24'(1380);
			13778: out = 24'(1412);
			13779: out = 24'(1468);
			13780: out = 24'(1500);
			13781: out = 24'(1500);
			13782: out = 24'(1556);
			13783: out = 24'(1596);
			13784: out = 24'(1640);
			13785: out = 24'(1640);
			13786: out = 24'(1692);
			13787: out = 24'(1752);
			13788: out = 24'(1768);
			13789: out = 24'(1800);
			13790: out = 24'(1816);
			13791: out = 24'(1916);
			13792: out = 24'(1888);
			13793: out = 24'(1956);
			13794: out = 24'(2016);
			13795: out = 24'(2040);
			13796: out = 24'(2068);
			13797: out = 24'(2116);
			13798: out = 24'(2172);
			13799: out = 24'(2196);
			13800: out = 24'(2228);
			13801: out = 24'(2252);
			13802: out = 24'(2332);
			13803: out = 24'(2356);
			13804: out = 24'(2380);
			13805: out = 24'(2440);
			13806: out = 24'(2480);
			13807: out = 24'(2536);
			13808: out = 24'(2560);
			13809: out = 24'(2572);
			13810: out = 24'(2652);
			13811: out = 24'(2692);
			13812: out = 24'(2720);
			13813: out = 24'(2772);
			13814: out = 24'(2780);
			13815: out = 24'(2828);
			13816: out = 24'(2904);
			13817: out = 24'(2868);
			13818: out = 24'(2976);
			13819: out = 24'(2992);
			13820: out = 24'(3008);
			13821: out = 24'(3080);
			13822: out = 24'(3092);
			13823: out = 24'(3160);
			13824: out = 24'(3144);
			13825: out = 24'(3196);
			13826: out = 24'(3256);
			13827: out = 24'(3280);
			13828: out = 24'(3276);
			13829: out = 24'(3356);
			13830: out = 24'(3388);
			13831: out = 24'(3428);
			13832: out = 24'(3440);
			13833: out = 24'(3448);
			13834: out = 24'(3528);
			13835: out = 24'(3540);
			13836: out = 24'(3560);
			13837: out = 24'(3604);
			13838: out = 24'(3660);
			13839: out = 24'(3620);
			13840: out = 24'(3752);
			13841: out = 24'(3716);
			13842: out = 24'(3752);
			13843: out = 24'(3792);
			13844: out = 24'(3836);
			13845: out = 24'(3812);
			13846: out = 24'(3868);
			13847: out = 24'(3900);
			13848: out = 24'(3904);
			13849: out = 24'(4000);
			13850: out = 24'(3960);
			13851: out = 24'(4000);
			13852: out = 24'(4040);
			13853: out = 24'(4092);
			13854: out = 24'(4048);
			13855: out = 24'(4132);
			13856: out = 24'(4140);
			13857: out = 24'(4160);
			13858: out = 24'(4188);
			13859: out = 24'(4224);
			13860: out = 24'(4236);
			13861: out = 24'(4248);
			13862: out = 24'(4328);
			13863: out = 24'(4276);
			13864: out = 24'(4340);
			13865: out = 24'(4360);
			13866: out = 24'(4372);
			13867: out = 24'(4420);
			13868: out = 24'(4404);
			13869: out = 24'(4476);
			13870: out = 24'(4468);
			13871: out = 24'(4484);
			13872: out = 24'(4520);
			13873: out = 24'(4520);
			13874: out = 24'(4540);
			13875: out = 24'(4596);
			13876: out = 24'(4600);
			13877: out = 24'(4604);
			13878: out = 24'(4620);
			13879: out = 24'(4708);
			13880: out = 24'(4672);
			13881: out = 24'(4688);
			13882: out = 24'(4748);
			13883: out = 24'(4716);
			13884: out = 24'(4792);
			13885: out = 24'(4752);
			13886: out = 24'(4832);
			13887: out = 24'(4808);
			13888: out = 24'(4844);
			13889: out = 24'(4844);
			13890: out = 24'(4876);
			13891: out = 24'(4904);
			13892: out = 24'(4900);
			13893: out = 24'(4948);
			13894: out = 24'(4972);
			13895: out = 24'(4948);
			13896: out = 24'(4984);
			13897: out = 24'(5008);
			13898: out = 24'(5024);
			13899: out = 24'(5052);
			13900: out = 24'(4988);
			13901: out = 24'(5084);
			13902: out = 24'(5096);
			13903: out = 24'(5088);
			13904: out = 24'(5144);
			13905: out = 24'(5120);
			13906: out = 24'(5152);
			13907: out = 24'(5192);
			13908: out = 24'(5132);
			13909: out = 24'(5220);
			13910: out = 24'(5184);
			13911: out = 24'(5192);
			13912: out = 24'(5244);
			13913: out = 24'(5200);
			13914: out = 24'(5240);
			13915: out = 24'(5224);
			13916: out = 24'(5260);
			13917: out = 24'(5200);
			13918: out = 24'(5196);
			13919: out = 24'(5232);
			13920: out = 24'(5220);
			13921: out = 24'(5232);
			13922: out = 24'(5180);
			13923: out = 24'(5216);
			13924: out = 24'(5244);
			13925: out = 24'(5200);
			13926: out = 24'(5180);
			13927: out = 24'(5176);
			13928: out = 24'(5232);
			13929: out = 24'(5200);
			13930: out = 24'(5164);
			13931: out = 24'(5148);
			13932: out = 24'(5168);
			13933: out = 24'(5132);
			13934: out = 24'(5144);
			13935: out = 24'(5168);
			13936: out = 24'(5168);
			13937: out = 24'(5120);
			13938: out = 24'(5192);
			13939: out = 24'(5152);
			13940: out = 24'(5188);
			13941: out = 24'(5128);
			13942: out = 24'(5180);
			13943: out = 24'(5172);
			13944: out = 24'(5136);
			13945: out = 24'(5180);
			13946: out = 24'(5160);
			13947: out = 24'(5080);
			13948: out = 24'(5192);
			13949: out = 24'(5116);
			13950: out = 24'(5104);
			13951: out = 24'(5152);
			13952: out = 24'(5116);
			13953: out = 24'(5152);
			13954: out = 24'(5080);
			13955: out = 24'(5132);
			13956: out = 24'(5152);
			13957: out = 24'(5124);
			13958: out = 24'(5108);
			13959: out = 24'(5116);
			13960: out = 24'(5144);
			13961: out = 24'(5124);
			13962: out = 24'(5076);
			13963: out = 24'(5124);
			13964: out = 24'(5140);
			13965: out = 24'(5080);
			13966: out = 24'(5124);
			13967: out = 24'(5128);
			13968: out = 24'(5104);
			13969: out = 24'(5116);
			13970: out = 24'(5056);
			13971: out = 24'(5072);
			13972: out = 24'(5096);
			13973: out = 24'(5088);
			13974: out = 24'(5040);
			13975: out = 24'(5072);
			13976: out = 24'(4996);
			13977: out = 24'(5096);
			13978: out = 24'(5020);
			13979: out = 24'(5040);
			13980: out = 24'(5012);
			13981: out = 24'(5080);
			13982: out = 24'(5044);
			13983: out = 24'(5012);
			13984: out = 24'(4988);
			13985: out = 24'(5020);
			13986: out = 24'(4960);
			13987: out = 24'(4916);
			13988: out = 24'(4972);
			13989: out = 24'(4924);
			13990: out = 24'(4908);
			13991: out = 24'(4912);
			13992: out = 24'(4856);
			13993: out = 24'(4852);
			13994: out = 24'(4860);
			13995: out = 24'(4832);
			13996: out = 24'(4776);
			13997: out = 24'(4824);
			13998: out = 24'(4760);
			13999: out = 24'(4764);
			14000: out = 24'(4760);
			14001: out = 24'(4672);
			14002: out = 24'(4700);
			14003: out = 24'(4668);
			14004: out = 24'(4680);
			14005: out = 24'(4552);
			14006: out = 24'(4644);
			14007: out = 24'(4568);
			14008: out = 24'(4596);
			14009: out = 24'(4512);
			14010: out = 24'(4480);
			14011: out = 24'(4472);
			14012: out = 24'(4468);
			14013: out = 24'(4404);
			14014: out = 24'(4356);
			14015: out = 24'(4340);
			14016: out = 24'(4332);
			14017: out = 24'(4276);
			14018: out = 24'(4240);
			14019: out = 24'(4216);
			14020: out = 24'(4188);
			14021: out = 24'(4140);
			14022: out = 24'(4104);
			14023: out = 24'(4072);
			14024: out = 24'(4084);
			14025: out = 24'(4000);
			14026: out = 24'(3992);
			14027: out = 24'(3968);
			14028: out = 24'(3896);
			14029: out = 24'(3912);
			14030: out = 24'(3828);
			14031: out = 24'(3812);
			14032: out = 24'(3780);
			14033: out = 24'(3744);
			14034: out = 24'(3744);
			14035: out = 24'(3660);
			14036: out = 24'(3648);
			14037: out = 24'(3632);
			14038: out = 24'(3604);
			14039: out = 24'(3540);
			14040: out = 24'(3520);
			14041: out = 24'(3472);
			14042: out = 24'(3448);
			14043: out = 24'(3400);
			14044: out = 24'(3352);
			14045: out = 24'(3372);
			14046: out = 24'(3260);
			14047: out = 24'(3268);
			14048: out = 24'(3272);
			14049: out = 24'(3228);
			14050: out = 24'(3156);
			14051: out = 24'(3120);
			14052: out = 24'(3088);
			14053: out = 24'(3064);
			14054: out = 24'(3032);
			14055: out = 24'(2984);
			14056: out = 24'(2912);
			14057: out = 24'(2956);
			14058: out = 24'(2908);
			14059: out = 24'(2892);
			14060: out = 24'(2808);
			14061: out = 24'(2828);
			14062: out = 24'(2804);
			14063: out = 24'(2712);
			14064: out = 24'(2724);
			14065: out = 24'(2708);
			14066: out = 24'(2616);
			14067: out = 24'(2660);
			14068: out = 24'(2568);
			14069: out = 24'(2564);
			14070: out = 24'(2524);
			14071: out = 24'(2492);
			14072: out = 24'(2472);
			14073: out = 24'(2444);
			14074: out = 24'(2392);
			14075: out = 24'(2368);
			14076: out = 24'(2388);
			14077: out = 24'(2300);
			14078: out = 24'(2288);
			14079: out = 24'(2264);
			14080: out = 24'(2240);
			14081: out = 24'(2196);
			14082: out = 24'(2164);
			14083: out = 24'(2164);
			14084: out = 24'(2132);
			14085: out = 24'(2068);
			14086: out = 24'(2072);
			14087: out = 24'(2028);
			14088: out = 24'(2016);
			14089: out = 24'(1996);
			14090: out = 24'(1984);
			14091: out = 24'(1928);
			14092: out = 24'(1916);
			14093: out = 24'(1896);
			14094: out = 24'(1820);
			14095: out = 24'(1856);
			14096: out = 24'(1768);
			14097: out = 24'(1768);
			14098: out = 24'(1776);
			14099: out = 24'(1720);
			14100: out = 24'(1720);
			14101: out = 24'(1736);
			14102: out = 24'(1688);
			14103: out = 24'(1628);
			14104: out = 24'(1640);
			14105: out = 24'(1620);
			14106: out = 24'(1556);
			14107: out = 24'(1564);
			14108: out = 24'(1500);
			14109: out = 24'(1504);
			14110: out = 24'(1492);
			14111: out = 24'(1440);
			14112: out = 24'(1432);
			14113: out = 24'(1428);
			14114: out = 24'(1436);
			14115: out = 24'(1348);
			14116: out = 24'(1360);
			14117: out = 24'(1328);
			14118: out = 24'(1312);
			14119: out = 24'(1292);
			14120: out = 24'(1272);
			14121: out = 24'(1224);
			14122: out = 24'(1236);
			14123: out = 24'(1220);
			14124: out = 24'(1212);
			14125: out = 24'(1184);
			14126: out = 24'(1156);
			14127: out = 24'(1100);
			14128: out = 24'(1148);
			14129: out = 24'(1104);
			14130: out = 24'(1036);
			14131: out = 24'(1068);
			14132: out = 24'(1068);
			14133: out = 24'(1036);
			14134: out = 24'(1008);
			14135: out = 24'(1008);
			14136: out = 24'(980);
			14137: out = 24'(976);
			14138: out = 24'(936);
			14139: out = 24'(932);
			14140: out = 24'(912);
			14141: out = 24'(908);
			14142: out = 24'(892);
			14143: out = 24'(876);
			14144: out = 24'(832);
			14145: out = 24'(820);
			14146: out = 24'(764);
			14147: out = 24'(712);
			14148: out = 24'(696);
			14149: out = 24'(640);
			14150: out = 24'(596);
			14151: out = 24'(572);
			14152: out = 24'(512);
			14153: out = 24'(476);
			14154: out = 24'(440);
			14155: out = 24'(408);
			14156: out = 24'(352);
			14157: out = 24'(364);
			14158: out = 24'(260);
			14159: out = 24'(304);
			14160: out = 24'(184);
			14161: out = 24'(212);
			14162: out = 24'(120);
			14163: out = 24'(152);
			14164: out = 24'(68);
			14165: out = 24'(68);
			14166: out = 24'(28);
			14167: out = 24'(-8);
			14168: out = 24'(-52);
			14169: out = 24'(-76);
			14170: out = 24'(-96);
			14171: out = 24'(-160);
			14172: out = 24'(-164);
			14173: out = 24'(-204);
			14174: out = 24'(-204);
			14175: out = 24'(-264);
			14176: out = 24'(-288);
			14177: out = 24'(-296);
			14178: out = 24'(-348);
			14179: out = 24'(-380);
			14180: out = 24'(-372);
			14181: out = 24'(-436);
			14182: out = 24'(-460);
			14183: out = 24'(-508);
			14184: out = 24'(-504);
			14185: out = 24'(-544);
			14186: out = 24'(-548);
			14187: out = 24'(-552);
			14188: out = 24'(-664);
			14189: out = 24'(-608);
			14190: out = 24'(-648);
			14191: out = 24'(-688);
			14192: out = 24'(-696);
			14193: out = 24'(-780);
			14194: out = 24'(-768);
			14195: out = 24'(-808);
			14196: out = 24'(-824);
			14197: out = 24'(-824);
			14198: out = 24'(-876);
			14199: out = 24'(-884);
			14200: out = 24'(-908);
			14201: out = 24'(-912);
			14202: out = 24'(-1008);
			14203: out = 24'(-996);
			14204: out = 24'(-1008);
			14205: out = 24'(-1116);
			14206: out = 24'(-1036);
			14207: out = 24'(-1076);
			14208: out = 24'(-1120);
			14209: out = 24'(-1104);
			14210: out = 24'(-1168);
			14211: out = 24'(-1176);
			14212: out = 24'(-1216);
			14213: out = 24'(-1196);
			14214: out = 24'(-1280);
			14215: out = 24'(-1232);
			14216: out = 24'(-1336);
			14217: out = 24'(-1308);
			14218: out = 24'(-1308);
			14219: out = 24'(-1408);
			14220: out = 24'(-1364);
			14221: out = 24'(-1412);
			14222: out = 24'(-1456);
			14223: out = 24'(-1472);
			14224: out = 24'(-1492);
			14225: out = 24'(-1520);
			14226: out = 24'(-1536);
			14227: out = 24'(-1552);
			14228: out = 24'(-1640);
			14229: out = 24'(-1592);
			14230: out = 24'(-1672);
			14231: out = 24'(-1688);
			14232: out = 24'(-1680);
			14233: out = 24'(-1772);
			14234: out = 24'(-1764);
			14235: out = 24'(-1784);
			14236: out = 24'(-1812);
			14237: out = 24'(-1856);
			14238: out = 24'(-1868);
			14239: out = 24'(-1920);
			14240: out = 24'(-1920);
			14241: out = 24'(-1968);
			14242: out = 24'(-2028);
			14243: out = 24'(-2044);
			14244: out = 24'(-2036);
			14245: out = 24'(-2112);
			14246: out = 24'(-2152);
			14247: out = 24'(-2144);
			14248: out = 24'(-2208);
			14249: out = 24'(-2256);
			14250: out = 24'(-2232);
			14251: out = 24'(-2340);
			14252: out = 24'(-2340);
			14253: out = 24'(-2424);
			14254: out = 24'(-2408);
			14255: out = 24'(-2428);
			14256: out = 24'(-2528);
			14257: out = 24'(-2572);
			14258: out = 24'(-2568);
			14259: out = 24'(-2608);
			14260: out = 24'(-2684);
			14261: out = 24'(-2676);
			14262: out = 24'(-2764);
			14263: out = 24'(-2780);
			14264: out = 24'(-2868);
			14265: out = 24'(-2864);
			14266: out = 24'(-2912);
			14267: out = 24'(-3008);
			14268: out = 24'(-3044);
			14269: out = 24'(-3052);
			14270: out = 24'(-3128);
			14271: out = 24'(-3160);
			14272: out = 24'(-3256);
			14273: out = 24'(-3224);
			14274: out = 24'(-3316);
			14275: out = 24'(-3336);
			14276: out = 24'(-3424);
			14277: out = 24'(-3480);
			14278: out = 24'(-3484);
			14279: out = 24'(-3552);
			14280: out = 24'(-3608);
			14281: out = 24'(-3640);
			14282: out = 24'(-3716);
			14283: out = 24'(-3704);
			14284: out = 24'(-3808);
			14285: out = 24'(-3820);
			14286: out = 24'(-3856);
			14287: out = 24'(-3904);
			14288: out = 24'(-3964);
			14289: out = 24'(-3952);
			14290: out = 24'(-4052);
			14291: out = 24'(-4056);
			14292: out = 24'(-4152);
			14293: out = 24'(-4184);
			14294: out = 24'(-4216);
			14295: out = 24'(-4252);
			14296: out = 24'(-4296);
			14297: out = 24'(-4324);
			14298: out = 24'(-4344);
			14299: out = 24'(-4420);
			14300: out = 24'(-4420);
			14301: out = 24'(-4480);
			14302: out = 24'(-4500);
			14303: out = 24'(-4540);
			14304: out = 24'(-4584);
			14305: out = 24'(-4600);
			14306: out = 24'(-4624);
			14307: out = 24'(-4660);
			14308: out = 24'(-4708);
			14309: out = 24'(-4736);
			14310: out = 24'(-4724);
			14311: out = 24'(-4768);
			14312: out = 24'(-4788);
			14313: out = 24'(-4852);
			14314: out = 24'(-4816);
			14315: out = 24'(-4884);
			14316: out = 24'(-4908);
			14317: out = 24'(-4916);
			14318: out = 24'(-4944);
			14319: out = 24'(-4980);
			14320: out = 24'(-4964);
			14321: out = 24'(-5024);
			14322: out = 24'(-5032);
			14323: out = 24'(-5040);
			14324: out = 24'(-5044);
			14325: out = 24'(-5092);
			14326: out = 24'(-5100);
			14327: out = 24'(-5120);
			14328: out = 24'(-5080);
			14329: out = 24'(-5152);
			14330: out = 24'(-5172);
			14331: out = 24'(-5168);
			14332: out = 24'(-5152);
			14333: out = 24'(-5192);
			14334: out = 24'(-5236);
			14335: out = 24'(-5208);
			14336: out = 24'(-5216);
			14337: out = 24'(-5260);
			14338: out = 24'(-5244);
			14339: out = 24'(-5260);
			14340: out = 24'(-5264);
			14341: out = 24'(-5312);
			14342: out = 24'(-5228);
			14343: out = 24'(-5328);
			14344: out = 24'(-5324);
			14345: out = 24'(-5280);
			14346: out = 24'(-5324);
			14347: out = 24'(-5292);
			14348: out = 24'(-5364);
			14349: out = 24'(-5312);
			14350: out = 24'(-5352);
			14351: out = 24'(-5320);
			14352: out = 24'(-5344);
			14353: out = 24'(-5352);
			14354: out = 24'(-5324);
			14355: out = 24'(-5332);
			14356: out = 24'(-5368);
			14357: out = 24'(-5340);
			14358: out = 24'(-5316);
			14359: out = 24'(-5364);
			14360: out = 24'(-5372);
			14361: out = 24'(-5308);
			14362: out = 24'(-5344);
			14363: out = 24'(-5380);
			14364: out = 24'(-5316);
			14365: out = 24'(-5336);
			14366: out = 24'(-5360);
			14367: out = 24'(-5344);
			14368: out = 24'(-5324);
			14369: out = 24'(-5316);
			14370: out = 24'(-5364);
			14371: out = 24'(-5284);
			14372: out = 24'(-5308);
			14373: out = 24'(-5316);
			14374: out = 24'(-5332);
			14375: out = 24'(-5316);
			14376: out = 24'(-5280);
			14377: out = 24'(-5296);
			14378: out = 24'(-5288);
			14379: out = 24'(-5276);
			14380: out = 24'(-5276);
			14381: out = 24'(-5292);
			14382: out = 24'(-5240);
			14383: out = 24'(-5288);
			14384: out = 24'(-5284);
			14385: out = 24'(-5240);
			14386: out = 24'(-5264);
			14387: out = 24'(-5248);
			14388: out = 24'(-5232);
			14389: out = 24'(-5236);
			14390: out = 24'(-5196);
			14391: out = 24'(-5200);
			14392: out = 24'(-5212);
			14393: out = 24'(-5188);
			14394: out = 24'(-5200);
			14395: out = 24'(-5152);
			14396: out = 24'(-5176);
			14397: out = 24'(-5180);
			14398: out = 24'(-5136);
			14399: out = 24'(-5164);
			14400: out = 24'(-5084);
			14401: out = 24'(-5164);
			14402: out = 24'(-5108);
			14403: out = 24'(-5120);
			14404: out = 24'(-5052);
			14405: out = 24'(-5088);
			14406: out = 24'(-5076);
			14407: out = 24'(-5080);
			14408: out = 24'(-5020);
			14409: out = 24'(-5024);
			14410: out = 24'(-5052);
			14411: out = 24'(-5024);
			14412: out = 24'(-4988);
			14413: out = 24'(-4988);
			14414: out = 24'(-5036);
			14415: out = 24'(-4948);
			14416: out = 24'(-4956);
			14417: out = 24'(-5000);
			14418: out = 24'(-4928);
			14419: out = 24'(-4948);
			14420: out = 24'(-4904);
			14421: out = 24'(-4940);
			14422: out = 24'(-4884);
			14423: out = 24'(-4864);
			14424: out = 24'(-4876);
			14425: out = 24'(-4864);
			14426: out = 24'(-4832);
			14427: out = 24'(-4808);
			14428: out = 24'(-4804);
			14429: out = 24'(-4784);
			14430: out = 24'(-4808);
			14431: out = 24'(-4764);
			14432: out = 24'(-4716);
			14433: out = 24'(-4760);
			14434: out = 24'(-4720);
			14435: out = 24'(-4672);
			14436: out = 24'(-4664);
			14437: out = 24'(-4700);
			14438: out = 24'(-4656);
			14439: out = 24'(-4616);
			14440: out = 24'(-4628);
			14441: out = 24'(-4616);
			14442: out = 24'(-4552);
			14443: out = 24'(-4556);
			14444: out = 24'(-4548);
			14445: out = 24'(-4540);
			14446: out = 24'(-4484);
			14447: out = 24'(-4488);
			14448: out = 24'(-4472);
			14449: out = 24'(-4452);
			14450: out = 24'(-4432);
			14451: out = 24'(-4404);
			14452: out = 24'(-4344);
			14453: out = 24'(-4388);
			14454: out = 24'(-4308);
			14455: out = 24'(-4276);
			14456: out = 24'(-4296);
			14457: out = 24'(-4236);
			14458: out = 24'(-4216);
			14459: out = 24'(-4196);
			14460: out = 24'(-4176);
			14461: out = 24'(-4144);
			14462: out = 24'(-4100);
			14463: out = 24'(-4100);
			14464: out = 24'(-4044);
			14465: out = 24'(-4016);
			14466: out = 24'(-4036);
			14467: out = 24'(-3940);
			14468: out = 24'(-3932);
			14469: out = 24'(-3900);
			14470: out = 24'(-3836);
			14471: out = 24'(-3828);
			14472: out = 24'(-3808);
			14473: out = 24'(-3744);
			14474: out = 24'(-3704);
			14475: out = 24'(-3688);
			14476: out = 24'(-3676);
			14477: out = 24'(-3580);
			14478: out = 24'(-3576);
			14479: out = 24'(-3528);
			14480: out = 24'(-3504);
			14481: out = 24'(-3424);
			14482: out = 24'(-3444);
			14483: out = 24'(-3388);
			14484: out = 24'(-3356);
			14485: out = 24'(-3336);
			14486: out = 24'(-3240);
			14487: out = 24'(-3300);
			14488: out = 24'(-3208);
			14489: out = 24'(-3160);
			14490: out = 24'(-3136);
			14491: out = 24'(-3084);
			14492: out = 24'(-3068);
			14493: out = 24'(-3016);
			14494: out = 24'(-2968);
			14495: out = 24'(-2960);
			14496: out = 24'(-2912);
			14497: out = 24'(-2888);
			14498: out = 24'(-2852);
			14499: out = 24'(-2788);
			14500: out = 24'(-2816);
			14501: out = 24'(-2720);
			14502: out = 24'(-2716);
			14503: out = 24'(-2652);
			14504: out = 24'(-2668);
			14505: out = 24'(-2576);
			14506: out = 24'(-2592);
			14507: out = 24'(-2500);
			14508: out = 24'(-2540);
			14509: out = 24'(-2444);
			14510: out = 24'(-2440);
			14511: out = 24'(-2400);
			14512: out = 24'(-2392);
			14513: out = 24'(-2312);
			14514: out = 24'(-2332);
			14515: out = 24'(-2304);
			14516: out = 24'(-2184);
			14517: out = 24'(-2236);
			14518: out = 24'(-2200);
			14519: out = 24'(-2152);
			14520: out = 24'(-2112);
			14521: out = 24'(-2112);
			14522: out = 24'(-2024);
			14523: out = 24'(-2056);
			14524: out = 24'(-2016);
			14525: out = 24'(-1960);
			14526: out = 24'(-1948);
			14527: out = 24'(-1920);
			14528: out = 24'(-1888);
			14529: out = 24'(-1852);
			14530: out = 24'(-1824);
			14531: out = 24'(-1840);
			14532: out = 24'(-1752);
			14533: out = 24'(-1732);
			14534: out = 24'(-1776);
			14535: out = 24'(-1708);
			14536: out = 24'(-1648);
			14537: out = 24'(-1664);
			14538: out = 24'(-1668);
			14539: out = 24'(-1568);
			14540: out = 24'(-1592);
			14541: out = 24'(-1568);
			14542: out = 24'(-1528);
			14543: out = 24'(-1524);
			14544: out = 24'(-1484);
			14545: out = 24'(-1448);
			14546: out = 24'(-1472);
			14547: out = 24'(-1428);
			14548: out = 24'(-1368);
			14549: out = 24'(-1416);
			14550: out = 24'(-1352);
			14551: out = 24'(-1292);
			14552: out = 24'(-1340);
			14553: out = 24'(-1252);
			14554: out = 24'(-1300);
			14555: out = 24'(-1240);
			14556: out = 24'(-1220);
			14557: out = 24'(-1232);
			14558: out = 24'(-1204);
			14559: out = 24'(-1188);
			14560: out = 24'(-1124);
			14561: out = 24'(-1160);
			14562: out = 24'(-1104);
			14563: out = 24'(-1108);
			14564: out = 24'(-1092);
			14565: out = 24'(-1084);
			14566: out = 24'(-1016);
			14567: out = 24'(-1016);
			14568: out = 24'(-1012);
			14569: out = 24'(-988);
			14570: out = 24'(-936);
			14571: out = 24'(-928);
			14572: out = 24'(-892);
			14573: out = 24'(-904);
			14574: out = 24'(-832);
			14575: out = 24'(-780);
			14576: out = 24'(-828);
			14577: out = 24'(-692);
			14578: out = 24'(-764);
			14579: out = 24'(-680);
			14580: out = 24'(-676);
			14581: out = 24'(-640);
			14582: out = 24'(-636);
			14583: out = 24'(-564);
			14584: out = 24'(-576);
			14585: out = 24'(-540);
			14586: out = 24'(-528);
			14587: out = 24'(-496);
			14588: out = 24'(-456);
			14589: out = 24'(-444);
			14590: out = 24'(-404);
			14591: out = 24'(-408);
			14592: out = 24'(-380);
			14593: out = 24'(-336);
			14594: out = 24'(-348);
			14595: out = 24'(-316);
			14596: out = 24'(-276);
			14597: out = 24'(-280);
			14598: out = 24'(-220);
			14599: out = 24'(-228);
			14600: out = 24'(-180);
			14601: out = 24'(-172);
			14602: out = 24'(-180);
			14603: out = 24'(-116);
			14604: out = 24'(-144);
			14605: out = 24'(-80);
			14606: out = 24'(-80);
			14607: out = 24'(-68);
			14608: out = 24'(-40);
			14609: out = 24'(-48);
			14610: out = 24'(4);
			14611: out = 24'(28);
			14612: out = 24'(-16);
			14613: out = 24'(80);
			14614: out = 24'(36);
			14615: out = 24'(84);
			14616: out = 24'(108);
			14617: out = 24'(108);
			14618: out = 24'(148);
			14619: out = 24'(144);
			14620: out = 24'(152);
			14621: out = 24'(168);
			14622: out = 24'(240);
			14623: out = 24'(208);
			14624: out = 24'(244);
			14625: out = 24'(272);
			14626: out = 24'(268);
			14627: out = 24'(256);
			14628: out = 24'(348);
			14629: out = 24'(304);
			14630: out = 24'(336);
			14631: out = 24'(364);
			14632: out = 24'(340);
			14633: out = 24'(388);
			14634: out = 24'(428);
			14635: out = 24'(400);
			14636: out = 24'(404);
			14637: out = 24'(496);
			14638: out = 24'(440);
			14639: out = 24'(532);
			14640: out = 24'(512);
			14641: out = 24'(456);
			14642: out = 24'(572);
			14643: out = 24'(552);
			14644: out = 24'(588);
			14645: out = 24'(584);
			14646: out = 24'(600);
			14647: out = 24'(616);
			14648: out = 24'(688);
			14649: out = 24'(664);
			14650: out = 24'(632);
			14651: out = 24'(688);
			14652: out = 24'(728);
			14653: out = 24'(752);
			14654: out = 24'(736);
			14655: out = 24'(780);
			14656: out = 24'(776);
			14657: out = 24'(880);
			14658: out = 24'(808);
			14659: out = 24'(880);
			14660: out = 24'(872);
			14661: out = 24'(924);
			14662: out = 24'(888);
			14663: out = 24'(960);
			14664: out = 24'(988);
			14665: out = 24'(968);
			14666: out = 24'(1028);
			14667: out = 24'(1036);
			14668: out = 24'(1056);
			14669: out = 24'(1116);
			14670: out = 24'(1092);
			14671: out = 24'(1144);
			14672: out = 24'(1156);
			14673: out = 24'(1188);
			14674: out = 24'(1232);
			14675: out = 24'(1240);
			14676: out = 24'(1284);
			14677: out = 24'(1300);
			14678: out = 24'(1360);
			14679: out = 24'(1368);
			14680: out = 24'(1384);
			14681: out = 24'(1432);
			14682: out = 24'(1432);
			14683: out = 24'(1468);
			14684: out = 24'(1564);
			14685: out = 24'(1536);
			14686: out = 24'(1572);
			14687: out = 24'(1620);
			14688: out = 24'(1672);
			14689: out = 24'(1676);
			14690: out = 24'(1716);
			14691: out = 24'(1760);
			14692: out = 24'(1760);
			14693: out = 24'(1816);
			14694: out = 24'(1852);
			14695: out = 24'(1864);
			14696: out = 24'(1876);
			14697: out = 24'(1980);
			14698: out = 24'(1948);
			14699: out = 24'(2028);
			14700: out = 24'(2040);
			14701: out = 24'(2076);
			14702: out = 24'(2100);
			14703: out = 24'(2172);
			14704: out = 24'(2144);
			14705: out = 24'(2208);
			14706: out = 24'(2220);
			14707: out = 24'(2264);
			14708: out = 24'(2264);
			14709: out = 24'(2336);
			14710: out = 24'(2336);
			14711: out = 24'(2376);
			14712: out = 24'(2440);
			14713: out = 24'(2416);
			14714: out = 24'(2512);
			14715: out = 24'(2496);
			14716: out = 24'(2500);
			14717: out = 24'(2568);
			14718: out = 24'(2588);
			14719: out = 24'(2620);
			14720: out = 24'(2644);
			14721: out = 24'(2644);
			14722: out = 24'(2708);
			14723: out = 24'(2728);
			14724: out = 24'(2724);
			14725: out = 24'(2764);
			14726: out = 24'(2800);
			14727: out = 24'(2832);
			14728: out = 24'(2864);
			14729: out = 24'(2876);
			14730: out = 24'(2876);
			14731: out = 24'(2920);
			14732: out = 24'(2960);
			14733: out = 24'(3000);
			14734: out = 24'(2956);
			14735: out = 24'(3016);
			14736: out = 24'(3084);
			14737: out = 24'(3084);
			14738: out = 24'(3084);
			14739: out = 24'(3104);
			14740: out = 24'(3148);
			14741: out = 24'(3184);
			14742: out = 24'(3140);
			14743: out = 24'(3204);
			14744: out = 24'(3224);
			14745: out = 24'(3224);
			14746: out = 24'(3272);
			14747: out = 24'(3272);
			14748: out = 24'(3316);
			14749: out = 24'(3288);
			14750: out = 24'(3388);
			14751: out = 24'(3320);
			14752: out = 24'(3396);
			14753: out = 24'(3368);
			14754: out = 24'(3404);
			14755: out = 24'(3448);
			14756: out = 24'(3420);
			14757: out = 24'(3480);
			14758: out = 24'(3464);
			14759: out = 24'(3536);
			14760: out = 24'(3512);
			14761: out = 24'(3560);
			14762: out = 24'(3544);
			14763: out = 24'(3584);
			14764: out = 24'(3588);
			14765: out = 24'(3592);
			14766: out = 24'(3632);
			14767: out = 24'(3640);
			14768: out = 24'(3652);
			14769: out = 24'(3688);
			14770: out = 24'(3672);
			14771: out = 24'(3724);
			14772: out = 24'(3700);
			14773: out = 24'(3768);
			14774: out = 24'(3740);
			14775: out = 24'(3780);
			14776: out = 24'(3776);
			14777: out = 24'(3844);
			14778: out = 24'(3764);
			14779: out = 24'(3864);
			14780: out = 24'(3856);
			14781: out = 24'(3824);
			14782: out = 24'(3872);
			14783: out = 24'(3888);
			14784: out = 24'(3892);
			14785: out = 24'(3912);
			14786: out = 24'(3932);
			14787: out = 24'(3984);
			14788: out = 24'(3936);
			14789: out = 24'(3980);
			14790: out = 24'(3996);
			14791: out = 24'(4012);
			14792: out = 24'(3980);
			14793: out = 24'(4064);
			14794: out = 24'(4052);
			14795: out = 24'(4040);
			14796: out = 24'(4080);
			14797: out = 24'(4120);
			14798: out = 24'(4076);
			14799: out = 24'(4100);
			14800: out = 24'(4156);
			14801: out = 24'(4132);
			14802: out = 24'(4152);
			14803: out = 24'(4144);
			14804: out = 24'(4152);
			14805: out = 24'(4128);
			14806: out = 24'(4204);
			14807: out = 24'(4140);
			14808: out = 24'(4180);
			14809: out = 24'(4140);
			14810: out = 24'(4184);
			14811: out = 24'(4128);
			14812: out = 24'(4152);
			14813: out = 24'(4188);
			14814: out = 24'(4128);
			14815: out = 24'(4144);
			14816: out = 24'(4160);
			14817: out = 24'(4156);
			14818: out = 24'(4112);
			14819: out = 24'(4140);
			14820: out = 24'(4140);
			14821: out = 24'(4096);
			14822: out = 24'(4124);
			14823: out = 24'(4124);
			14824: out = 24'(4140);
			14825: out = 24'(4096);
			14826: out = 24'(4092);
			14827: out = 24'(4108);
			14828: out = 24'(4072);
			14829: out = 24'(4120);
			14830: out = 24'(4084);
			14831: out = 24'(4064);
			14832: out = 24'(4124);
			14833: out = 24'(4140);
			14834: out = 24'(4048);
			14835: out = 24'(4136);
			14836: out = 24'(4076);
			14837: out = 24'(4144);
			14838: out = 24'(4056);
			14839: out = 24'(4088);
			14840: out = 24'(4128);
			14841: out = 24'(4064);
			14842: out = 24'(4080);
			14843: out = 24'(4144);
			14844: out = 24'(4072);
			14845: out = 24'(4100);
			14846: out = 24'(4120);
			14847: out = 24'(4108);
			14848: out = 24'(4092);
			14849: out = 24'(4096);
			14850: out = 24'(4080);
			14851: out = 24'(4076);
			14852: out = 24'(4104);
			14853: out = 24'(4060);
			14854: out = 24'(4028);
			14855: out = 24'(4064);
			14856: out = 24'(4060);
			14857: out = 24'(4040);
			14858: out = 24'(4048);
			14859: out = 24'(4064);
			14860: out = 24'(4088);
			14861: out = 24'(4036);
			14862: out = 24'(4060);
			14863: out = 24'(4064);
			14864: out = 24'(4028);
			14865: out = 24'(4008);
			14866: out = 24'(4024);
			14867: out = 24'(3996);
			14868: out = 24'(4008);
			14869: out = 24'(4012);
			14870: out = 24'(4004);
			14871: out = 24'(4044);
			14872: out = 24'(4008);
			14873: out = 24'(4016);
			14874: out = 24'(3992);
			14875: out = 24'(3996);
			14876: out = 24'(3956);
			14877: out = 24'(3968);
			14878: out = 24'(3912);
			14879: out = 24'(3924);
			14880: out = 24'(3948);
			14881: out = 24'(3912);
			14882: out = 24'(3912);
			14883: out = 24'(3900);
			14884: out = 24'(3916);
			14885: out = 24'(3820);
			14886: out = 24'(3808);
			14887: out = 24'(3884);
			14888: out = 24'(3800);
			14889: out = 24'(3788);
			14890: out = 24'(3792);
			14891: out = 24'(3748);
			14892: out = 24'(3788);
			14893: out = 24'(3704);
			14894: out = 24'(3720);
			14895: out = 24'(3688);
			14896: out = 24'(3708);
			14897: out = 24'(3700);
			14898: out = 24'(3656);
			14899: out = 24'(3624);
			14900: out = 24'(3616);
			14901: out = 24'(3588);
			14902: out = 24'(3496);
			14903: out = 24'(3552);
			14904: out = 24'(3512);
			14905: out = 24'(3440);
			14906: out = 24'(3464);
			14907: out = 24'(3448);
			14908: out = 24'(3400);
			14909: out = 24'(3376);
			14910: out = 24'(3400);
			14911: out = 24'(3296);
			14912: out = 24'(3324);
			14913: out = 24'(3288);
			14914: out = 24'(3200);
			14915: out = 24'(3220);
			14916: out = 24'(3184);
			14917: out = 24'(3144);
			14918: out = 24'(3160);
			14919: out = 24'(3136);
			14920: out = 24'(3096);
			14921: out = 24'(3104);
			14922: out = 24'(3016);
			14923: out = 24'(3024);
			14924: out = 24'(2976);
			14925: out = 24'(2944);
			14926: out = 24'(2940);
			14927: out = 24'(2880);
			14928: out = 24'(2880);
			14929: out = 24'(2860);
			14930: out = 24'(2836);
			14931: out = 24'(2780);
			14932: out = 24'(2796);
			14933: out = 24'(2740);
			14934: out = 24'(2704);
			14935: out = 24'(2660);
			14936: out = 24'(2620);
			14937: out = 24'(2660);
			14938: out = 24'(2536);
			14939: out = 24'(2584);
			14940: out = 24'(2520);
			14941: out = 24'(2536);
			14942: out = 24'(2488);
			14943: out = 24'(2424);
			14944: out = 24'(2456);
			14945: out = 24'(2408);
			14946: out = 24'(2344);
			14947: out = 24'(2368);
			14948: out = 24'(2304);
			14949: out = 24'(2304);
			14950: out = 24'(2300);
			14951: out = 24'(2216);
			14952: out = 24'(2200);
			14953: out = 24'(2232);
			14954: out = 24'(2136);
			14955: out = 24'(2136);
			14956: out = 24'(2148);
			14957: out = 24'(2072);
			14958: out = 24'(2064);
			14959: out = 24'(2056);
			14960: out = 24'(2008);
			14961: out = 24'(1968);
			14962: out = 24'(1968);
			14963: out = 24'(1972);
			14964: out = 24'(1824);
			14965: out = 24'(1952);
			14966: out = 24'(1816);
			14967: out = 24'(1864);
			14968: out = 24'(1836);
			14969: out = 24'(1756);
			14970: out = 24'(1812);
			14971: out = 24'(1744);
			14972: out = 24'(1736);
			14973: out = 24'(1712);
			14974: out = 24'(1688);
			14975: out = 24'(1684);
			14976: out = 24'(1648);
			14977: out = 24'(1556);
			14978: out = 24'(1648);
			14979: out = 24'(1568);
			14980: out = 24'(1516);
			14981: out = 24'(1536);
			14982: out = 24'(1540);
			14983: out = 24'(1484);
			14984: out = 24'(1452);
			14985: out = 24'(1468);
			14986: out = 24'(1428);
			14987: out = 24'(1400);
			14988: out = 24'(1396);
			14989: out = 24'(1328);
			14990: out = 24'(1384);
			14991: out = 24'(1308);
			14992: out = 24'(1320);
			14993: out = 24'(1308);
			14994: out = 24'(1244);
			14995: out = 24'(1252);
			14996: out = 24'(1264);
			14997: out = 24'(1224);
			14998: out = 24'(1224);
			14999: out = 24'(1224);
			15000: out = 24'(1156);
			15001: out = 24'(1168);
			15002: out = 24'(1124);
			15003: out = 24'(1112);
			15004: out = 24'(1076);
			15005: out = 24'(1080);
			15006: out = 24'(1048);
			15007: out = 24'(1056);
			15008: out = 24'(1036);
			15009: out = 24'(988);
			15010: out = 24'(1036);
			15011: out = 24'(964);
			15012: out = 24'(968);
			15013: out = 24'(932);
			15014: out = 24'(920);
			15015: out = 24'(972);
			15016: out = 24'(876);
			15017: out = 24'(904);
			15018: out = 24'(892);
			15019: out = 24'(888);
			15020: out = 24'(840);
			15021: out = 24'(840);
			15022: out = 24'(864);
			15023: out = 24'(772);
			15024: out = 24'(792);
			15025: out = 24'(784);
			15026: out = 24'(788);
			15027: out = 24'(732);
			15028: out = 24'(744);
			15029: out = 24'(752);
			15030: out = 24'(720);
			15031: out = 24'(728);
			15032: out = 24'(668);
			15033: out = 24'(684);
			15034: out = 24'(676);
			15035: out = 24'(620);
			15036: out = 24'(628);
			15037: out = 24'(616);
			15038: out = 24'(576);
			15039: out = 24'(500);
			15040: out = 24'(512);
			15041: out = 24'(468);
			15042: out = 24'(388);
			15043: out = 24'(408);
			15044: out = 24'(352);
			15045: out = 24'(336);
			15046: out = 24'(256);
			15047: out = 24'(300);
			15048: out = 24'(252);
			15049: out = 24'(156);
			15050: out = 24'(196);
			15051: out = 24'(152);
			15052: out = 24'(152);
			15053: out = 24'(64);
			15054: out = 24'(96);
			15055: out = 24'(4);
			15056: out = 24'(36);
			15057: out = 24'(-16);
			15058: out = 24'(-28);
			15059: out = 24'(-76);
			15060: out = 24'(-72);
			15061: out = 24'(-80);
			15062: out = 24'(-196);
			15063: out = 24'(-116);
			15064: out = 24'(-228);
			15065: out = 24'(-172);
			15066: out = 24'(-244);
			15067: out = 24'(-240);
			15068: out = 24'(-260);
			15069: out = 24'(-320);
			15070: out = 24'(-304);
			15071: out = 24'(-340);
			15072: out = 24'(-396);
			15073: out = 24'(-388);
			15074: out = 24'(-404);
			15075: out = 24'(-440);
			15076: out = 24'(-460);
			15077: out = 24'(-496);
			15078: out = 24'(-480);
			15079: out = 24'(-500);
			15080: out = 24'(-560);
			15081: out = 24'(-584);
			15082: out = 24'(-560);
			15083: out = 24'(-600);
			15084: out = 24'(-648);
			15085: out = 24'(-636);
			15086: out = 24'(-636);
			15087: out = 24'(-692);
			15088: out = 24'(-696);
			15089: out = 24'(-724);
			15090: out = 24'(-740);
			15091: out = 24'(-772);
			15092: out = 24'(-824);
			15093: out = 24'(-772);
			15094: out = 24'(-828);
			15095: out = 24'(-844);
			15096: out = 24'(-836);
			15097: out = 24'(-888);
			15098: out = 24'(-848);
			15099: out = 24'(-960);
			15100: out = 24'(-952);
			15101: out = 24'(-936);
			15102: out = 24'(-976);
			15103: out = 24'(-1012);
			15104: out = 24'(-956);
			15105: out = 24'(-1056);
			15106: out = 24'(-1036);
			15107: out = 24'(-1068);
			15108: out = 24'(-1076);
			15109: out = 24'(-1108);
			15110: out = 24'(-1140);
			15111: out = 24'(-1152);
			15112: out = 24'(-1164);
			15113: out = 24'(-1184);
			15114: out = 24'(-1200);
			15115: out = 24'(-1256);
			15116: out = 24'(-1220);
			15117: out = 24'(-1288);
			15118: out = 24'(-1264);
			15119: out = 24'(-1340);
			15120: out = 24'(-1308);
			15121: out = 24'(-1400);
			15122: out = 24'(-1344);
			15123: out = 24'(-1408);
			15124: out = 24'(-1424);
			15125: out = 24'(-1444);
			15126: out = 24'(-1484);
			15127: out = 24'(-1488);
			15128: out = 24'(-1520);
			15129: out = 24'(-1528);
			15130: out = 24'(-1552);
			15131: out = 24'(-1568);
			15132: out = 24'(-1640);
			15133: out = 24'(-1612);
			15134: out = 24'(-1672);
			15135: out = 24'(-1716);
			15136: out = 24'(-1696);
			15137: out = 24'(-1732);
			15138: out = 24'(-1760);
			15139: out = 24'(-1808);
			15140: out = 24'(-1788);
			15141: out = 24'(-1880);
			15142: out = 24'(-1872);
			15143: out = 24'(-1888);
			15144: out = 24'(-1968);
			15145: out = 24'(-1976);
			15146: out = 24'(-1984);
			15147: out = 24'(-2012);
			15148: out = 24'(-2064);
			15149: out = 24'(-2140);
			15150: out = 24'(-2104);
			15151: out = 24'(-2192);
			15152: out = 24'(-2188);
			15153: out = 24'(-2232);
			15154: out = 24'(-2292);
			15155: out = 24'(-2320);
			15156: out = 24'(-2332);
			15157: out = 24'(-2384);
			15158: out = 24'(-2428);
			15159: out = 24'(-2456);
			15160: out = 24'(-2484);
			15161: out = 24'(-2528);
			15162: out = 24'(-2560);
			15163: out = 24'(-2592);
			15164: out = 24'(-2692);
			15165: out = 24'(-2652);
			15166: out = 24'(-2720);
			15167: out = 24'(-2732);
			15168: out = 24'(-2804);
			15169: out = 24'(-2820);
			15170: out = 24'(-2876);
			15171: out = 24'(-2868);
			15172: out = 24'(-3008);
			15173: out = 24'(-2940);
			15174: out = 24'(-2996);
			15175: out = 24'(-3084);
			15176: out = 24'(-3080);
			15177: out = 24'(-3068);
			15178: out = 24'(-3164);
			15179: out = 24'(-3192);
			15180: out = 24'(-3220);
			15181: out = 24'(-3256);
			15182: out = 24'(-3300);
			15183: out = 24'(-3332);
			15184: out = 24'(-3352);
			15185: out = 24'(-3400);
			15186: out = 24'(-3384);
			15187: out = 24'(-3468);
			15188: out = 24'(-3464);
			15189: out = 24'(-3492);
			15190: out = 24'(-3556);
			15191: out = 24'(-3584);
			15192: out = 24'(-3584);
			15193: out = 24'(-3624);
			15194: out = 24'(-3652);
			15195: out = 24'(-3688);
			15196: out = 24'(-3708);
			15197: out = 24'(-3712);
			15198: out = 24'(-3772);
			15199: out = 24'(-3772);
			15200: out = 24'(-3792);
			15201: out = 24'(-3804);
			15202: out = 24'(-3864);
			15203: out = 24'(-3828);
			15204: out = 24'(-3876);
			15205: out = 24'(-3924);
			15206: out = 24'(-3900);
			15207: out = 24'(-3956);
			15208: out = 24'(-3980);
			15209: out = 24'(-3956);
			15210: out = 24'(-3992);
			15211: out = 24'(-3992);
			15212: out = 24'(-4064);
			15213: out = 24'(-4016);
			15214: out = 24'(-4060);
			15215: out = 24'(-4080);
			15216: out = 24'(-4040);
			15217: out = 24'(-4144);
			15218: out = 24'(-4096);
			15219: out = 24'(-4104);
			15220: out = 24'(-4176);
			15221: out = 24'(-4112);
			15222: out = 24'(-4184);
			15223: out = 24'(-4160);
			15224: out = 24'(-4160);
			15225: out = 24'(-4220);
			15226: out = 24'(-4184);
			15227: out = 24'(-4224);
			15228: out = 24'(-4200);
			15229: out = 24'(-4220);
			15230: out = 24'(-4228);
			15231: out = 24'(-4248);
			15232: out = 24'(-4224);
			15233: out = 24'(-4248);
			15234: out = 24'(-4268);
			15235: out = 24'(-4240);
			15236: out = 24'(-4288);
			15237: out = 24'(-4292);
			15238: out = 24'(-4252);
			15239: out = 24'(-4268);
			15240: out = 24'(-4300);
			15241: out = 24'(-4268);
			15242: out = 24'(-4296);
			15243: out = 24'(-4292);
			15244: out = 24'(-4300);
			15245: out = 24'(-4268);
			15246: out = 24'(-4364);
			15247: out = 24'(-4264);
			15248: out = 24'(-4296);
			15249: out = 24'(-4300);
			15250: out = 24'(-4284);
			15251: out = 24'(-4296);
			15252: out = 24'(-4308);
			15253: out = 24'(-4300);
			15254: out = 24'(-4284);
			15255: out = 24'(-4252);
			15256: out = 24'(-4288);
			15257: out = 24'(-4316);
			15258: out = 24'(-4312);
			15259: out = 24'(-4264);
			15260: out = 24'(-4332);
			15261: out = 24'(-4264);
			15262: out = 24'(-4292);
			15263: out = 24'(-4296);
			15264: out = 24'(-4268);
			15265: out = 24'(-4280);
			15266: out = 24'(-4264);
			15267: out = 24'(-4264);
			15268: out = 24'(-4264);
			15269: out = 24'(-4244);
			15270: out = 24'(-4248);
			15271: out = 24'(-4244);
			15272: out = 24'(-4252);
			15273: out = 24'(-4220);
			15274: out = 24'(-4252);
			15275: out = 24'(-4236);
			15276: out = 24'(-4244);
			15277: out = 24'(-4232);
			15278: out = 24'(-4232);
			15279: out = 24'(-4220);
			15280: out = 24'(-4176);
			15281: out = 24'(-4256);
			15282: out = 24'(-4172);
			15283: out = 24'(-4208);
			15284: out = 24'(-4180);
			15285: out = 24'(-4168);
			15286: out = 24'(-4196);
			15287: out = 24'(-4184);
			15288: out = 24'(-4132);
			15289: out = 24'(-4176);
			15290: out = 24'(-4124);
			15291: out = 24'(-4136);
			15292: out = 24'(-4128);
			15293: out = 24'(-4120);
			15294: out = 24'(-4100);
			15295: out = 24'(-4088);
			15296: out = 24'(-4076);
			15297: out = 24'(-4112);
			15298: out = 24'(-4064);
			15299: out = 24'(-4072);
			15300: out = 24'(-4076);
			15301: out = 24'(-4048);
			15302: out = 24'(-4044);
			15303: out = 24'(-4028);
			15304: out = 24'(-4052);
			15305: out = 24'(-4008);
			15306: out = 24'(-4000);
			15307: out = 24'(-4032);
			15308: out = 24'(-3984);
			15309: out = 24'(-3968);
			15310: out = 24'(-3980);
			15311: out = 24'(-3952);
			15312: out = 24'(-3964);
			15313: out = 24'(-3948);
			15314: out = 24'(-3960);
			15315: out = 24'(-3864);
			15316: out = 24'(-3916);
			15317: out = 24'(-3916);
			15318: out = 24'(-3892);
			15319: out = 24'(-3848);
			15320: out = 24'(-3896);
			15321: out = 24'(-3812);
			15322: out = 24'(-3856);
			15323: out = 24'(-3828);
			15324: out = 24'(-3776);
			15325: out = 24'(-3836);
			15326: out = 24'(-3760);
			15327: out = 24'(-3780);
			15328: out = 24'(-3780);
			15329: out = 24'(-3724);
			15330: out = 24'(-3752);
			15331: out = 24'(-3716);
			15332: out = 24'(-3720);
			15333: out = 24'(-3664);
			15334: out = 24'(-3716);
			15335: out = 24'(-3640);
			15336: out = 24'(-3652);
			15337: out = 24'(-3616);
			15338: out = 24'(-3588);
			15339: out = 24'(-3636);
			15340: out = 24'(-3592);
			15341: out = 24'(-3528);
			15342: out = 24'(-3552);
			15343: out = 24'(-3524);
			15344: out = 24'(-3524);
			15345: out = 24'(-3436);
			15346: out = 24'(-3464);
			15347: out = 24'(-3480);
			15348: out = 24'(-3404);
			15349: out = 24'(-3432);
			15350: out = 24'(-3412);
			15351: out = 24'(-3352);
			15352: out = 24'(-3344);
			15353: out = 24'(-3296);
			15354: out = 24'(-3296);
			15355: out = 24'(-3284);
			15356: out = 24'(-3204);
			15357: out = 24'(-3212);
			15358: out = 24'(-3212);
			15359: out = 24'(-3156);
			15360: out = 24'(-3116);
			15361: out = 24'(-3132);
			15362: out = 24'(-3088);
			15363: out = 24'(-3056);
			15364: out = 24'(-3052);
			15365: out = 24'(-3008);
			15366: out = 24'(-2936);
			15367: out = 24'(-3008);
			15368: out = 24'(-2880);
			15369: out = 24'(-2912);
			15370: out = 24'(-2856);
			15371: out = 24'(-2816);
			15372: out = 24'(-2844);
			15373: out = 24'(-2776);
			15374: out = 24'(-2724);
			15375: out = 24'(-2700);
			15376: out = 24'(-2700);
			15377: out = 24'(-2640);
			15378: out = 24'(-2632);
			15379: out = 24'(-2604);
			15380: out = 24'(-2588);
			15381: out = 24'(-2532);
			15382: out = 24'(-2540);
			15383: out = 24'(-2496);
			15384: out = 24'(-2448);
			15385: out = 24'(-2440);
			15386: out = 24'(-2380);
			15387: out = 24'(-2388);
			15388: out = 24'(-2352);
			15389: out = 24'(-2300);
			15390: out = 24'(-2284);
			15391: out = 24'(-2268);
			15392: out = 24'(-2248);
			15393: out = 24'(-2204);
			15394: out = 24'(-2192);
			15395: out = 24'(-2124);
			15396: out = 24'(-2124);
			15397: out = 24'(-2116);
			15398: out = 24'(-2052);
			15399: out = 24'(-2044);
			15400: out = 24'(-1996);
			15401: out = 24'(-2000);
			15402: out = 24'(-1976);
			15403: out = 24'(-1932);
			15404: out = 24'(-1888);
			15405: out = 24'(-1908);
			15406: out = 24'(-1852);
			15407: out = 24'(-1832);
			15408: out = 24'(-1792);
			15409: out = 24'(-1820);
			15410: out = 24'(-1764);
			15411: out = 24'(-1756);
			15412: out = 24'(-1736);
			15413: out = 24'(-1684);
			15414: out = 24'(-1692);
			15415: out = 24'(-1644);
			15416: out = 24'(-1644);
			15417: out = 24'(-1604);
			15418: out = 24'(-1588);
			15419: out = 24'(-1536);
			15420: out = 24'(-1544);
			15421: out = 24'(-1568);
			15422: out = 24'(-1468);
			15423: out = 24'(-1476);
			15424: out = 24'(-1428);
			15425: out = 24'(-1448);
			15426: out = 24'(-1444);
			15427: out = 24'(-1388);
			15428: out = 24'(-1356);
			15429: out = 24'(-1360);
			15430: out = 24'(-1352);
			15431: out = 24'(-1316);
			15432: out = 24'(-1288);
			15433: out = 24'(-1268);
			15434: out = 24'(-1248);
			15435: out = 24'(-1236);
			15436: out = 24'(-1192);
			15437: out = 24'(-1204);
			15438: out = 24'(-1208);
			15439: out = 24'(-1156);
			15440: out = 24'(-1144);
			15441: out = 24'(-1160);
			15442: out = 24'(-1128);
			15443: out = 24'(-1092);
			15444: out = 24'(-1080);
			15445: out = 24'(-1084);
			15446: out = 24'(-1032);
			15447: out = 24'(-1020);
			15448: out = 24'(-1028);
			15449: out = 24'(-996);
			15450: out = 24'(-968);
			15451: out = 24'(-1024);
			15452: out = 24'(-936);
			15453: out = 24'(-948);
			15454: out = 24'(-952);
			15455: out = 24'(-920);
			15456: out = 24'(-888);
			15457: out = 24'(-880);
			15458: out = 24'(-872);
			15459: out = 24'(-816);
			15460: out = 24'(-836);
			15461: out = 24'(-792);
			15462: out = 24'(-816);
			15463: out = 24'(-704);
			15464: out = 24'(-760);
			15465: out = 24'(-724);
			15466: out = 24'(-668);
			15467: out = 24'(-640);
			15468: out = 24'(-652);
			15469: out = 24'(-592);
			15470: out = 24'(-580);
			15471: out = 24'(-576);
			15472: out = 24'(-524);
			15473: out = 24'(-552);
			15474: out = 24'(-544);
			15475: out = 24'(-476);
			15476: out = 24'(-444);
			15477: out = 24'(-464);
			15478: out = 24'(-440);
			15479: out = 24'(-400);
			15480: out = 24'(-388);
			15481: out = 24'(-388);
			15482: out = 24'(-360);
			15483: out = 24'(-324);
			15484: out = 24'(-340);
			15485: out = 24'(-276);
			15486: out = 24'(-276);
			15487: out = 24'(-240);
			15488: out = 24'(-296);
			15489: out = 24'(-208);
			15490: out = 24'(-216);
			15491: out = 24'(-216);
			15492: out = 24'(-164);
			15493: out = 24'(-172);
			15494: out = 24'(-124);
			15495: out = 24'(-148);
			15496: out = 24'(-80);
			15497: out = 24'(-108);
			15498: out = 24'(-48);
			15499: out = 24'(-76);
			15500: out = 24'(-64);
			15501: out = 24'(-28);
			15502: out = 24'(-20);
			15503: out = 24'(-4);
			15504: out = 24'(28);
			15505: out = 24'(16);
			15506: out = 24'(28);
			15507: out = 24'(56);
			15508: out = 24'(80);
			15509: out = 24'(68);
			15510: out = 24'(116);
			15511: out = 24'(84);
			15512: out = 24'(108);
			15513: out = 24'(160);
			15514: out = 24'(144);
			15515: out = 24'(164);
			15516: out = 24'(164);
			15517: out = 24'(184);
			15518: out = 24'(204);
			15519: out = 24'(228);
			15520: out = 24'(216);
			15521: out = 24'(260);
			15522: out = 24'(232);
			15523: out = 24'(320);
			15524: out = 24'(272);
			15525: out = 24'(252);
			15526: out = 24'(332);
			15527: out = 24'(340);
			15528: out = 24'(348);
			15529: out = 24'(332);
			15530: out = 24'(372);
			15531: out = 24'(392);
			15532: out = 24'(412);
			15533: out = 24'(400);
			15534: out = 24'(444);
			15535: out = 24'(436);
			15536: out = 24'(468);
			15537: out = 24'(484);
			15538: out = 24'(492);
			15539: out = 24'(512);
			15540: out = 24'(512);
			15541: out = 24'(528);
			15542: out = 24'(548);
			15543: out = 24'(580);
			15544: out = 24'(544);
			15545: out = 24'(596);
			15546: out = 24'(640);
			15547: out = 24'(580);
			15548: out = 24'(684);
			15549: out = 24'(620);
			15550: out = 24'(684);
			15551: out = 24'(652);
			15552: out = 24'(752);
			15553: out = 24'(696);
			15554: out = 24'(748);
			15555: out = 24'(744);
			15556: out = 24'(832);
			15557: out = 24'(772);
			15558: out = 24'(848);
			15559: out = 24'(844);
			15560: out = 24'(880);
			15561: out = 24'(884);
			15562: out = 24'(888);
			15563: out = 24'(936);
			15564: out = 24'(948);
			15565: out = 24'(948);
			15566: out = 24'(1016);
			15567: out = 24'(1000);
			15568: out = 24'(1044);
			15569: out = 24'(1076);
			15570: out = 24'(1072);
			15571: out = 24'(1120);
			15572: out = 24'(1124);
			15573: out = 24'(1168);
			15574: out = 24'(1188);
			15575: out = 24'(1232);
			15576: out = 24'(1192);
			15577: out = 24'(1304);
			15578: out = 24'(1244);
			15579: out = 24'(1344);
			15580: out = 24'(1328);
			15581: out = 24'(1340);
			15582: out = 24'(1376);
			15583: out = 24'(1412);
			15584: out = 24'(1488);
			15585: out = 24'(1412);
			15586: out = 24'(1524);
			15587: out = 24'(1484);
			15588: out = 24'(1588);
			15589: out = 24'(1552);
			15590: out = 24'(1592);
			15591: out = 24'(1616);
			15592: out = 24'(1680);
			15593: out = 24'(1664);
			15594: out = 24'(1728);
			15595: out = 24'(1720);
			15596: out = 24'(1772);
			15597: out = 24'(1776);
			15598: out = 24'(1780);
			15599: out = 24'(1808);
			15600: out = 24'(1836);
			15601: out = 24'(1888);
			15602: out = 24'(1872);
			15603: out = 24'(1904);
			15604: out = 24'(1960);
			15605: out = 24'(1972);
			15606: out = 24'(1968);
			15607: out = 24'(1984);
			15608: out = 24'(2068);
			15609: out = 24'(2056);
			15610: out = 24'(2072);
			15611: out = 24'(2084);
			15612: out = 24'(2116);
			15613: out = 24'(2140);
			15614: out = 24'(2192);
			15615: out = 24'(2164);
			15616: out = 24'(2180);
			15617: out = 24'(2240);
			15618: out = 24'(2236);
			15619: out = 24'(2308);
			15620: out = 24'(2240);
			15621: out = 24'(2292);
			15622: out = 24'(2328);
			15623: out = 24'(2388);
			15624: out = 24'(2356);
			15625: out = 24'(2372);
			15626: out = 24'(2396);
			15627: out = 24'(2436);
			15628: out = 24'(2436);
			15629: out = 24'(2432);
			15630: out = 24'(2468);
			15631: out = 24'(2480);
			15632: out = 24'(2524);
			15633: out = 24'(2500);
			15634: out = 24'(2544);
			15635: out = 24'(2564);
			15636: out = 24'(2568);
			15637: out = 24'(2580);
			15638: out = 24'(2624);
			15639: out = 24'(2616);
			15640: out = 24'(2620);
			15641: out = 24'(2636);
			15642: out = 24'(2680);
			15643: out = 24'(2688);
			15644: out = 24'(2668);
			15645: out = 24'(2712);
			15646: out = 24'(2732);
			15647: out = 24'(2776);
			15648: out = 24'(2736);
			15649: out = 24'(2780);
			15650: out = 24'(2772);
			15651: out = 24'(2804);
			15652: out = 24'(2848);
			15653: out = 24'(2820);
			15654: out = 24'(2820);
			15655: out = 24'(2852);
			15656: out = 24'(2908);
			15657: out = 24'(2848);
			15658: out = 24'(2924);
			15659: out = 24'(2900);
			15660: out = 24'(2916);
			15661: out = 24'(2940);
			15662: out = 24'(2940);
			15663: out = 24'(2984);
			15664: out = 24'(2976);
			15665: out = 24'(2968);
			15666: out = 24'(3008);
			15667: out = 24'(3008);
			15668: out = 24'(3048);
			15669: out = 24'(2984);
			15670: out = 24'(3060);
			15671: out = 24'(3048);
			15672: out = 24'(3056);
			15673: out = 24'(3104);
			15674: out = 24'(3060);
			15675: out = 24'(3108);
			15676: out = 24'(3112);
			15677: out = 24'(3132);
			15678: out = 24'(3128);
			15679: out = 24'(3132);
			15680: out = 24'(3156);
			15681: out = 24'(3180);
			15682: out = 24'(3184);
			15683: out = 24'(3156);
			15684: out = 24'(3228);
			15685: out = 24'(3200);
			15686: out = 24'(3220);
			15687: out = 24'(3212);
			15688: out = 24'(3252);
			15689: out = 24'(3268);
			15690: out = 24'(3252);
			15691: out = 24'(3256);
			15692: out = 24'(3276);
			15693: out = 24'(3276);
			15694: out = 24'(3288);
			15695: out = 24'(3276);
			15696: out = 24'(3244);
			15697: out = 24'(3296);
			15698: out = 24'(3276);
			15699: out = 24'(3288);
			15700: out = 24'(3240);
			15701: out = 24'(3288);
			15702: out = 24'(3272);
			15703: out = 24'(3276);
			15704: out = 24'(3228);
			15705: out = 24'(3296);
			15706: out = 24'(3248);
			15707: out = 24'(3284);
			15708: out = 24'(3252);
			15709: out = 24'(3188);
			15710: out = 24'(3272);
			15711: out = 24'(3204);
			15712: out = 24'(3272);
			15713: out = 24'(3244);
			15714: out = 24'(3240);
			15715: out = 24'(3252);
			15716: out = 24'(3248);
			15717: out = 24'(3248);
			15718: out = 24'(3288);
			15719: out = 24'(3244);
			15720: out = 24'(3220);
			15721: out = 24'(3252);
			15722: out = 24'(3256);
			15723: out = 24'(3252);
			15724: out = 24'(3204);
			15725: out = 24'(3196);
			15726: out = 24'(3244);
			15727: out = 24'(3164);
			15728: out = 24'(3220);
			15729: out = 24'(3228);
			15730: out = 24'(3172);
			15731: out = 24'(3240);
			15732: out = 24'(3244);
			15733: out = 24'(3200);
			15734: out = 24'(3196);
			15735: out = 24'(3196);
			15736: out = 24'(3204);
			15737: out = 24'(3152);
			15738: out = 24'(3232);
			15739: out = 24'(3184);
			15740: out = 24'(3172);
			15741: out = 24'(3220);
			15742: out = 24'(3196);
			15743: out = 24'(3220);
			15744: out = 24'(3156);
			15745: out = 24'(3192);
			15746: out = 24'(3232);
			15747: out = 24'(3172);
			15748: out = 24'(3188);
			15749: out = 24'(3228);
			15750: out = 24'(3204);
			15751: out = 24'(3184);
			15752: out = 24'(3184);
			15753: out = 24'(3140);
			15754: out = 24'(3224);
			15755: out = 24'(3152);
			15756: out = 24'(3128);
			15757: out = 24'(3144);
			15758: out = 24'(3200);
			15759: out = 24'(3128);
			15760: out = 24'(3112);
			15761: out = 24'(3156);
			15762: out = 24'(3120);
			15763: out = 24'(3112);
			15764: out = 24'(3140);
			15765: out = 24'(3100);
			15766: out = 24'(3136);
			15767: out = 24'(3092);
			15768: out = 24'(3096);
			15769: out = 24'(3108);
			15770: out = 24'(3084);
			15771: out = 24'(3048);
			15772: out = 24'(3080);
			15773: out = 24'(3084);
			15774: out = 24'(3012);
			15775: out = 24'(3064);
			15776: out = 24'(2996);
			15777: out = 24'(3040);
			15778: out = 24'(2964);
			15779: out = 24'(2996);
			15780: out = 24'(2988);
			15781: out = 24'(2960);
			15782: out = 24'(2944);
			15783: out = 24'(2928);
			15784: out = 24'(2936);
			15785: out = 24'(2876);
			15786: out = 24'(2924);
			15787: out = 24'(2828);
			15788: out = 24'(2856);
			15789: out = 24'(2864);
			15790: out = 24'(2828);
			15791: out = 24'(2816);
			15792: out = 24'(2772);
			15793: out = 24'(2808);
			15794: out = 24'(2784);
			15795: out = 24'(2736);
			15796: out = 24'(2716);
			15797: out = 24'(2712);
			15798: out = 24'(2676);
			15799: out = 24'(2668);
			15800: out = 24'(2672);
			15801: out = 24'(2580);
			15802: out = 24'(2624);
			15803: out = 24'(2532);
			15804: out = 24'(2536);
			15805: out = 24'(2548);
			15806: out = 24'(2480);
			15807: out = 24'(2496);
			15808: out = 24'(2468);
			15809: out = 24'(2464);
			15810: out = 24'(2416);
			15811: out = 24'(2428);
			15812: out = 24'(2384);
			15813: out = 24'(2388);
			15814: out = 24'(2328);
			15815: out = 24'(2320);
			15816: out = 24'(2288);
			15817: out = 24'(2260);
			15818: out = 24'(2252);
			15819: out = 24'(2236);
			15820: out = 24'(2168);
			15821: out = 24'(2172);
			15822: out = 24'(2152);
			15823: out = 24'(2152);
			15824: out = 24'(2124);
			15825: out = 24'(2056);
			15826: out = 24'(2104);
			15827: out = 24'(2044);
			15828: out = 24'(2060);
			15829: out = 24'(1992);
			15830: out = 24'(2000);
			15831: out = 24'(1964);
			15832: out = 24'(1960);
			15833: out = 24'(1876);
			15834: out = 24'(1924);
			15835: out = 24'(1888);
			15836: out = 24'(1864);
			15837: out = 24'(1840);
			15838: out = 24'(1816);
			15839: out = 24'(1824);
			15840: out = 24'(1764);
			15841: out = 24'(1744);
			15842: out = 24'(1724);
			15843: out = 24'(1676);
			15844: out = 24'(1720);
			15845: out = 24'(1644);
			15846: out = 24'(1632);
			15847: out = 24'(1660);
			15848: out = 24'(1596);
			15849: out = 24'(1624);
			15850: out = 24'(1544);
			15851: out = 24'(1568);
			15852: out = 24'(1544);
			15853: out = 24'(1492);
			15854: out = 24'(1504);
			15855: out = 24'(1452);
			15856: out = 24'(1452);
			15857: out = 24'(1440);
			15858: out = 24'(1396);
			15859: out = 24'(1396);
			15860: out = 24'(1380);
			15861: out = 24'(1364);
			15862: out = 24'(1312);
			15863: out = 24'(1332);
			15864: out = 24'(1308);
			15865: out = 24'(1296);
			15866: out = 24'(1248);
			15867: out = 24'(1260);
			15868: out = 24'(1224);
			15869: out = 24'(1236);
			15870: out = 24'(1188);
			15871: out = 24'(1216);
			15872: out = 24'(1140);
			15873: out = 24'(1176);
			15874: out = 24'(1144);
			15875: out = 24'(1108);
			15876: out = 24'(1068);
			15877: out = 24'(1104);
			15878: out = 24'(1096);
			15879: out = 24'(1004);
			15880: out = 24'(1028);
			15881: out = 24'(1064);
			15882: out = 24'(1000);
			15883: out = 24'(968);
			15884: out = 24'(1000);
			15885: out = 24'(968);
			15886: out = 24'(928);
			15887: out = 24'(952);
			15888: out = 24'(908);
			15889: out = 24'(868);
			15890: out = 24'(912);
			15891: out = 24'(836);
			15892: out = 24'(832);
			15893: out = 24'(864);
			15894: out = 24'(796);
			15895: out = 24'(816);
			15896: out = 24'(836);
			15897: out = 24'(764);
			15898: out = 24'(796);
			15899: out = 24'(748);
			15900: out = 24'(748);
			15901: out = 24'(752);
			15902: out = 24'(712);
			15903: out = 24'(712);
			15904: out = 24'(720);
			15905: out = 24'(704);
			15906: out = 24'(688);
			15907: out = 24'(676);
			15908: out = 24'(656);
			15909: out = 24'(656);
			15910: out = 24'(632);
			15911: out = 24'(596);
			15912: out = 24'(640);
			15913: out = 24'(556);
			15914: out = 24'(608);
			15915: out = 24'(588);
			15916: out = 24'(532);
			15917: out = 24'(560);
			15918: out = 24'(532);
			15919: out = 24'(564);
			15920: out = 24'(512);
			15921: out = 24'(500);
			15922: out = 24'(492);
			15923: out = 24'(512);
			15924: out = 24'(516);
			15925: out = 24'(432);
			15926: out = 24'(452);
			15927: out = 24'(444);
			15928: out = 24'(416);
			15929: out = 24'(340);
			15930: out = 24'(372);
			15931: out = 24'(312);
			15932: out = 24'(296);
			15933: out = 24'(272);
			15934: out = 24'(260);
			15935: out = 24'(220);
			15936: out = 24'(204);
			15937: out = 24'(172);
			15938: out = 24'(128);
			15939: out = 24'(132);
			15940: out = 24'(120);
			15941: out = 24'(76);
			15942: out = 24'(32);
			15943: out = 24'(48);
			15944: out = 24'(60);
			15945: out = 24'(-36);
			15946: out = 24'(-4);
			15947: out = 24'(-28);
			15948: out = 24'(-36);
			15949: out = 24'(-100);
			15950: out = 24'(-96);
			15951: out = 24'(-100);
			15952: out = 24'(-128);
			15953: out = 24'(-152);
			15954: out = 24'(-208);
			15955: out = 24'(-196);
			15956: out = 24'(-200);
			15957: out = 24'(-240);
			15958: out = 24'(-252);
			15959: out = 24'(-276);
			15960: out = 24'(-272);
			15961: out = 24'(-316);
			15962: out = 24'(-292);
			15963: out = 24'(-364);
			15964: out = 24'(-324);
			15965: out = 24'(-388);
			15966: out = 24'(-412);
			15967: out = 24'(-432);
			15968: out = 24'(-388);
			15969: out = 24'(-432);
			15970: out = 24'(-468);
			15971: out = 24'(-476);
			15972: out = 24'(-452);
			15973: out = 24'(-524);
			15974: out = 24'(-500);
			15975: out = 24'(-532);
			15976: out = 24'(-560);
			15977: out = 24'(-552);
			15978: out = 24'(-584);
			15979: out = 24'(-576);
			15980: out = 24'(-616);
			15981: out = 24'(-624);
			15982: out = 24'(-628);
			15983: out = 24'(-632);
			15984: out = 24'(-668);
			15985: out = 24'(-684);
			15986: out = 24'(-668);
			15987: out = 24'(-716);
			15988: out = 24'(-716);
			15989: out = 24'(-740);
			15990: out = 24'(-780);
			15991: out = 24'(-764);
			15992: out = 24'(-768);
			15993: out = 24'(-844);
			15994: out = 24'(-780);
			15995: out = 24'(-868);
			15996: out = 24'(-820);
			15997: out = 24'(-868);
			15998: out = 24'(-876);
			15999: out = 24'(-912);
			16000: out = 24'(-884);
			16001: out = 24'(-940);
			16002: out = 24'(-964);
			16003: out = 24'(-952);
			16004: out = 24'(-984);
			16005: out = 24'(-1008);
			16006: out = 24'(-1028);
			16007: out = 24'(-996);
			16008: out = 24'(-1072);
			16009: out = 24'(-1032);
			16010: out = 24'(-1096);
			16011: out = 24'(-1084);
			16012: out = 24'(-1112);
			16013: out = 24'(-1148);
			16014: out = 24'(-1132);
			16015: out = 24'(-1144);
			16016: out = 24'(-1204);
			16017: out = 24'(-1188);
			16018: out = 24'(-1216);
			16019: out = 24'(-1212);
			16020: out = 24'(-1272);
			16021: out = 24'(-1248);
			16022: out = 24'(-1292);
			16023: out = 24'(-1300);
			16024: out = 24'(-1344);
			16025: out = 24'(-1348);
			16026: out = 24'(-1368);
			16027: out = 24'(-1400);
			16028: out = 24'(-1392);
			16029: out = 24'(-1460);
			16030: out = 24'(-1476);
			16031: out = 24'(-1468);
			16032: out = 24'(-1480);
			16033: out = 24'(-1536);
			16034: out = 24'(-1544);
			16035: out = 24'(-1572);
			16036: out = 24'(-1620);
			16037: out = 24'(-1620);
			16038: out = 24'(-1632);
			16039: out = 24'(-1684);
			16040: out = 24'(-1696);
			16041: out = 24'(-1732);
			16042: out = 24'(-1724);
			16043: out = 24'(-1792);
			16044: out = 24'(-1808);
			16045: out = 24'(-1852);
			16046: out = 24'(-1864);
			16047: out = 24'(-1904);
			16048: out = 24'(-1924);
			16049: out = 24'(-1908);
			16050: out = 24'(-2020);
			16051: out = 24'(-2008);
			16052: out = 24'(-2028);
			16053: out = 24'(-2092);
			16054: out = 24'(-2100);
			16055: out = 24'(-2140);
			16056: out = 24'(-2156);
			16057: out = 24'(-2168);
			16058: out = 24'(-2204);
			16059: out = 24'(-2240);
			16060: out = 24'(-2324);
			16061: out = 24'(-2284);
			16062: out = 24'(-2340);
			16063: out = 24'(-2344);
			16064: out = 24'(-2436);
			16065: out = 24'(-2440);
			16066: out = 24'(-2456);
			16067: out = 24'(-2452);
			16068: out = 24'(-2528);
			16069: out = 24'(-2548);
			16070: out = 24'(-2588);
			16071: out = 24'(-2548);
			16072: out = 24'(-2640);
			16073: out = 24'(-2652);
			16074: out = 24'(-2676);
			16075: out = 24'(-2688);
			16076: out = 24'(-2732);
			16077: out = 24'(-2780);
			16078: out = 24'(-2768);
			16079: out = 24'(-2776);
			16080: out = 24'(-2824);
			16081: out = 24'(-2880);
			16082: out = 24'(-2848);
			16083: out = 24'(-2908);
			16084: out = 24'(-2892);
			16085: out = 24'(-2968);
			16086: out = 24'(-2960);
			16087: out = 24'(-2988);
			16088: out = 24'(-2992);
			16089: out = 24'(-3012);
			16090: out = 24'(-3040);
			16091: out = 24'(-3032);
			16092: out = 24'(-3096);
			16093: out = 24'(-3064);
			16094: out = 24'(-3112);
			16095: out = 24'(-3132);
			16096: out = 24'(-3144);
			16097: out = 24'(-3160);
			16098: out = 24'(-3148);
			16099: out = 24'(-3180);
			16100: out = 24'(-3176);
			16101: out = 24'(-3244);
			16102: out = 24'(-3176);
			16103: out = 24'(-3248);
			16104: out = 24'(-3276);
			16105: out = 24'(-3224);
			16106: out = 24'(-3296);
			16107: out = 24'(-3252);
			16108: out = 24'(-3304);
			16109: out = 24'(-3284);
			16110: out = 24'(-3332);
			16111: out = 24'(-3292);
			16112: out = 24'(-3348);
			16113: out = 24'(-3340);
			16114: out = 24'(-3336);
			16115: out = 24'(-3368);
			16116: out = 24'(-3344);
			16117: out = 24'(-3372);
			16118: out = 24'(-3388);
			16119: out = 24'(-3352);
			16120: out = 24'(-3428);
			16121: out = 24'(-3352);
			16122: out = 24'(-3428);
			16123: out = 24'(-3400);
			16124: out = 24'(-3388);
			16125: out = 24'(-3436);
			16126: out = 24'(-3412);
			16127: out = 24'(-3428);
			16128: out = 24'(-3404);
			16129: out = 24'(-3460);
			16130: out = 24'(-3392);
			16131: out = 24'(-3464);
			16132: out = 24'(-3420);
			16133: out = 24'(-3480);
			16134: out = 24'(-3412);
			16135: out = 24'(-3456);
			16136: out = 24'(-3468);
			16137: out = 24'(-3448);
			16138: out = 24'(-3432);
			16139: out = 24'(-3444);
			16140: out = 24'(-3468);
			16141: out = 24'(-3468);
			16142: out = 24'(-3428);
			16143: out = 24'(-3460);
			16144: out = 24'(-3468);
			16145: out = 24'(-3436);
			16146: out = 24'(-3444);
			16147: out = 24'(-3460);
			16148: out = 24'(-3464);
			16149: out = 24'(-3432);
			16150: out = 24'(-3492);
			16151: out = 24'(-3412);
			16152: out = 24'(-3456);
			16153: out = 24'(-3460);
			16154: out = 24'(-3436);
			16155: out = 24'(-3448);
			16156: out = 24'(-3372);
			16157: out = 24'(-3516);
			16158: out = 24'(-3388);
			16159: out = 24'(-3436);
			16160: out = 24'(-3384);
			16161: out = 24'(-3460);
			16162: out = 24'(-3384);
			16163: out = 24'(-3412);
			16164: out = 24'(-3384);
			16165: out = 24'(-3388);
			16166: out = 24'(-3420);
			16167: out = 24'(-3372);
			16168: out = 24'(-3384);
			16169: out = 24'(-3356);
			16170: out = 24'(-3400);
			16171: out = 24'(-3392);
			16172: out = 24'(-3368);
			16173: out = 24'(-3376);
			16174: out = 24'(-3320);
			16175: out = 24'(-3392);
			16176: out = 24'(-3344);
			16177: out = 24'(-3356);
			16178: out = 24'(-3304);
			16179: out = 24'(-3328);
			16180: out = 24'(-3364);
			16181: out = 24'(-3332);
			16182: out = 24'(-3288);
			16183: out = 24'(-3292);
			16184: out = 24'(-3368);
			16185: out = 24'(-3272);
			16186: out = 24'(-3292);
			16187: out = 24'(-3256);
			16188: out = 24'(-3300);
			16189: out = 24'(-3284);
			16190: out = 24'(-3248);
			16191: out = 24'(-3272);
			16192: out = 24'(-3248);
			16193: out = 24'(-3276);
			16194: out = 24'(-3212);
			16195: out = 24'(-3248);
			16196: out = 24'(-3204);
			16197: out = 24'(-3232);
			16198: out = 24'(-3204);
			16199: out = 24'(-3200);
			16200: out = 24'(-3224);
			16201: out = 24'(-3176);
			16202: out = 24'(-3164);
			16203: out = 24'(-3188);
			16204: out = 24'(-3176);
			16205: out = 24'(-3140);
			16206: out = 24'(-3140);
			16207: out = 24'(-3160);
			16208: out = 24'(-3136);
			16209: out = 24'(-3116);
			16210: out = 24'(-3100);
			16211: out = 24'(-3128);
			16212: out = 24'(-3080);
			16213: out = 24'(-3092);
			16214: out = 24'(-3108);
			16215: out = 24'(-3044);
			16216: out = 24'(-3060);
			16217: out = 24'(-3052);
			16218: out = 24'(-3032);
			16219: out = 24'(-3032);
			16220: out = 24'(-2976);
			16221: out = 24'(-3016);
			16222: out = 24'(-3032);
			16223: out = 24'(-2968);
			16224: out = 24'(-2968);
			16225: out = 24'(-2964);
			16226: out = 24'(-2920);
			16227: out = 24'(-2960);
			16228: out = 24'(-2900);
			16229: out = 24'(-2916);
			16230: out = 24'(-2896);
			16231: out = 24'(-2864);
			16232: out = 24'(-2868);
			16233: out = 24'(-2836);
			16234: out = 24'(-2832);
			16235: out = 24'(-2844);
			16236: out = 24'(-2812);
			16237: out = 24'(-2776);
			16238: out = 24'(-2764);
			16239: out = 24'(-2800);
			16240: out = 24'(-2732);
			16241: out = 24'(-2720);
			16242: out = 24'(-2676);
			16243: out = 24'(-2724);
			16244: out = 24'(-2668);
			16245: out = 24'(-2652);
			16246: out = 24'(-2640);
			16247: out = 24'(-2604);
			16248: out = 24'(-2592);
			16249: out = 24'(-2580);
			16250: out = 24'(-2540);
			16251: out = 24'(-2520);
			16252: out = 24'(-2560);
			16253: out = 24'(-2452);
			16254: out = 24'(-2480);
			16255: out = 24'(-2452);
			16256: out = 24'(-2396);
			16257: out = 24'(-2444);
			16258: out = 24'(-2360);
			16259: out = 24'(-2356);
			16260: out = 24'(-2336);
			16261: out = 24'(-2280);
			16262: out = 24'(-2320);
			16263: out = 24'(-2268);
			16264: out = 24'(-2228);
			16265: out = 24'(-2192);
			16266: out = 24'(-2200);
			16267: out = 24'(-2196);
			16268: out = 24'(-2108);
			16269: out = 24'(-2136);
			16270: out = 24'(-2072);
			16271: out = 24'(-2100);
			16272: out = 24'(-2060);
			16273: out = 24'(-2000);
			16274: out = 24'(-2012);
			16275: out = 24'(-1992);
			16276: out = 24'(-1932);
			16277: out = 24'(-1952);
			16278: out = 24'(-1904);
			16279: out = 24'(-1896);
			16280: out = 24'(-1840);
			16281: out = 24'(-1832);
			16282: out = 24'(-1832);
			16283: out = 24'(-1792);
			16284: out = 24'(-1772);
			16285: out = 24'(-1764);
			16286: out = 24'(-1752);
			16287: out = 24'(-1724);
			16288: out = 24'(-1672);
			16289: out = 24'(-1684);
			16290: out = 24'(-1664);
			16291: out = 24'(-1616);
			16292: out = 24'(-1604);
			16293: out = 24'(-1604);
			16294: out = 24'(-1564);
			16295: out = 24'(-1544);
			16296: out = 24'(-1544);
			16297: out = 24'(-1504);
			16298: out = 24'(-1496);
			16299: out = 24'(-1444);
			16300: out = 24'(-1460);
			16301: out = 24'(-1440);
			16302: out = 24'(-1416);
			16303: out = 24'(-1356);
			16304: out = 24'(-1388);
			16305: out = 24'(-1356);
			16306: out = 24'(-1308);
			16307: out = 24'(-1340);
			16308: out = 24'(-1268);
			16309: out = 24'(-1320);
			16310: out = 24'(-1224);
			16311: out = 24'(-1280);
			16312: out = 24'(-1208);
			16313: out = 24'(-1208);
			16314: out = 24'(-1200);
			16315: out = 24'(-1152);
			16316: out = 24'(-1192);
			16317: out = 24'(-1128);
			16318: out = 24'(-1112);
			16319: out = 24'(-1084);
			16320: out = 24'(-1120);
			16321: out = 24'(-1048);
			16322: out = 24'(-1056);
			16323: out = 24'(-1068);
			16324: out = 24'(-1020);
			16325: out = 24'(-1004);
			16326: out = 24'(-1060);
			16327: out = 24'(-956);
			16328: out = 24'(-988);
			16329: out = 24'(-980);
			16330: out = 24'(-968);
			16331: out = 24'(-904);
			16332: out = 24'(-952);
			16333: out = 24'(-924);
			16334: out = 24'(-884);
			16335: out = 24'(-908);
			16336: out = 24'(-840);
			16337: out = 24'(-848);
			16338: out = 24'(-904);
			16339: out = 24'(-828);
			16340: out = 24'(-812);
			16341: out = 24'(-796);
			16342: out = 24'(-772);
			16343: out = 24'(-816);
			16344: out = 24'(-736);
			16345: out = 24'(-760);
			16346: out = 24'(-740);
			16347: out = 24'(-736);
			16348: out = 24'(-724);
			16349: out = 24'(-720);
			16350: out = 24'(-692);
			16351: out = 24'(-688);
			16352: out = 24'(-648);
			16353: out = 24'(-644);
			16354: out = 24'(-616);
			16355: out = 24'(-588);
			16356: out = 24'(-588);
			16357: out = 24'(-556);
			16358: out = 24'(-552);
			16359: out = 24'(-532);
			16360: out = 24'(-532);
			16361: out = 24'(-504);
			16362: out = 24'(-452);
			16363: out = 24'(-456);
			16364: out = 24'(-432);
			16365: out = 24'(-440);
			16366: out = 24'(-392);
			16367: out = 24'(-372);
			16368: out = 24'(-380);
			16369: out = 24'(-404);
			16370: out = 24'(-344);
			16371: out = 24'(-312);
			16372: out = 24'(-296);
			16373: out = 24'(-332);
			16374: out = 24'(-272);
			16375: out = 24'(-256);
			16376: out = 24'(-268);
			16377: out = 24'(-260);
			16378: out = 24'(-224);
			16379: out = 24'(-244);
			16380: out = 24'(-204);
			16381: out = 24'(-196);
			16382: out = 24'(-180);
			16383: out = 24'(-180);
			16384: out = 24'(-152);
			16385: out = 24'(-164);
			16386: out = 24'(-116);
			16387: out = 24'(-136);
			16388: out = 24'(-96);
			16389: out = 24'(-84);
			16390: out = 24'(-68);
			16391: out = 24'(-60);
			16392: out = 24'(-64);
			16393: out = 24'(-32);
			16394: out = 24'(-12);
			16395: out = 24'(-48);
			16396: out = 24'(-16);
			16397: out = 24'(0);
			16398: out = 24'(0);
			16399: out = 24'(28);
			16400: out = 24'(36);
			16401: out = 24'(12);
			16402: out = 24'(80);
			16403: out = 24'(40);
			16404: out = 24'(80);
			16405: out = 24'(64);
			16406: out = 24'(96);
			16407: out = 24'(124);
			16408: out = 24'(128);
			16409: out = 24'(128);
			16410: out = 24'(132);
			16411: out = 24'(180);
			16412: out = 24'(152);
			16413: out = 24'(156);
			16414: out = 24'(180);
			16415: out = 24'(176);
			16416: out = 24'(228);
			16417: out = 24'(200);
			16418: out = 24'(224);
			16419: out = 24'(240);
			16420: out = 24'(280);
			16421: out = 24'(248);
			16422: out = 24'(272);
			16423: out = 24'(288);
			16424: out = 24'(340);
			16425: out = 24'(276);
			16426: out = 24'(308);
			16427: out = 24'(344);
			16428: out = 24'(356);
			16429: out = 24'(316);
			16430: out = 24'(408);
			16431: out = 24'(360);
			16432: out = 24'(404);
			16433: out = 24'(404);
			16434: out = 24'(404);
			16435: out = 24'(452);
			16436: out = 24'(444);
			16437: out = 24'(436);
			16438: out = 24'(476);
			16439: out = 24'(488);
			16440: out = 24'(508);
			16441: out = 24'(464);
			16442: out = 24'(532);
			16443: out = 24'(528);
			16444: out = 24'(524);
			16445: out = 24'(588);
			16446: out = 24'(532);
			16447: out = 24'(616);
			16448: out = 24'(572);
			16449: out = 24'(664);
			16450: out = 24'(628);
			16451: out = 24'(644);
			16452: out = 24'(688);
			16453: out = 24'(720);
			16454: out = 24'(704);
			16455: out = 24'(720);
			16456: out = 24'(760);
			16457: out = 24'(764);
			16458: out = 24'(764);
			16459: out = 24'(784);
			16460: out = 24'(876);
			16461: out = 24'(812);
			16462: out = 24'(848);
			16463: out = 24'(876);
			16464: out = 24'(916);
			16465: out = 24'(900);
			16466: out = 24'(960);
			16467: out = 24'(980);
			16468: out = 24'(968);
			16469: out = 24'(1008);
			16470: out = 24'(1020);
			16471: out = 24'(1036);
			16472: out = 24'(1056);
			16473: out = 24'(1080);
			16474: out = 24'(1120);
			16475: out = 24'(1092);
			16476: out = 24'(1128);
			16477: out = 24'(1172);
			16478: out = 24'(1188);
			16479: out = 24'(1168);
			16480: out = 24'(1236);
			16481: out = 24'(1252);
			16482: out = 24'(1272);
			16483: out = 24'(1280);
			16484: out = 24'(1312);
			16485: out = 24'(1308);
			16486: out = 24'(1376);
			16487: out = 24'(1360);
			16488: out = 24'(1368);
			16489: out = 24'(1412);
			16490: out = 24'(1412);
			16491: out = 24'(1428);
			16492: out = 24'(1468);
			16493: out = 24'(1472);
			16494: out = 24'(1520);
			16495: out = 24'(1496);
			16496: out = 24'(1588);
			16497: out = 24'(1532);
			16498: out = 24'(1532);
			16499: out = 24'(1604);
			16500: out = 24'(1616);
			16501: out = 24'(1628);
			16502: out = 24'(1668);
			16503: out = 24'(1600);
			16504: out = 24'(1728);
			16505: out = 24'(1680);
			16506: out = 24'(1688);
			16507: out = 24'(1776);
			16508: out = 24'(1716);
			16509: out = 24'(1712);
			16510: out = 24'(1808);
			16511: out = 24'(1804);
			16512: out = 24'(1824);
			16513: out = 24'(1784);
			16514: out = 24'(1840);
			16515: out = 24'(1868);
			16516: out = 24'(1828);
			16517: out = 24'(1872);
			16518: out = 24'(1860);
			16519: out = 24'(1936);
			16520: out = 24'(1896);
			16521: out = 24'(1952);
			16522: out = 24'(1932);
			16523: out = 24'(1980);
			16524: out = 24'(1980);
			16525: out = 24'(1968);
			16526: out = 24'(2008);
			16527: out = 24'(1992);
			16528: out = 24'(2028);
			16529: out = 24'(2024);
			16530: out = 24'(2056);
			16531: out = 24'(2056);
			16532: out = 24'(2120);
			16533: out = 24'(2064);
			16534: out = 24'(2084);
			16535: out = 24'(2132);
			16536: out = 24'(2116);
			16537: out = 24'(2116);
			16538: out = 24'(2124);
			16539: out = 24'(2160);
			16540: out = 24'(2188);
			16541: out = 24'(2124);
			16542: out = 24'(2208);
			16543: out = 24'(2184);
			16544: out = 24'(2228);
			16545: out = 24'(2192);
			16546: out = 24'(2244);
			16547: out = 24'(2252);
			16548: out = 24'(2244);
			16549: out = 24'(2256);
			16550: out = 24'(2276);
			16551: out = 24'(2268);
			16552: out = 24'(2288);
			16553: out = 24'(2264);
			16554: out = 24'(2332);
			16555: out = 24'(2300);
			16556: out = 24'(2324);
			16557: out = 24'(2340);
			16558: out = 24'(2368);
			16559: out = 24'(2332);
			16560: out = 24'(2348);
			16561: out = 24'(2392);
			16562: out = 24'(2416);
			16563: out = 24'(2348);
			16564: out = 24'(2420);
			16565: out = 24'(2420);
			16566: out = 24'(2404);
			16567: out = 24'(2452);
			16568: out = 24'(2408);
			16569: out = 24'(2468);
			16570: out = 24'(2444);
			16571: out = 24'(2476);
			16572: out = 24'(2480);
			16573: out = 24'(2500);
			16574: out = 24'(2480);
			16575: out = 24'(2520);
			16576: out = 24'(2480);
			16577: out = 24'(2548);
			16578: out = 24'(2484);
			16579: out = 24'(2504);
			16580: out = 24'(2532);
			16581: out = 24'(2520);
			16582: out = 24'(2588);
			16583: out = 24'(2500);
			16584: out = 24'(2584);
			16585: out = 24'(2532);
			16586: out = 24'(2584);
			16587: out = 24'(2540);
			16588: out = 24'(2584);
			16589: out = 24'(2560);
			16590: out = 24'(2596);
			16591: out = 24'(2528);
			16592: out = 24'(2560);
			16593: out = 24'(2552);
			16594: out = 24'(2564);
			16595: out = 24'(2488);
			16596: out = 24'(2536);
			16597: out = 24'(2520);
			16598: out = 24'(2500);
			16599: out = 24'(2576);
			16600: out = 24'(2492);
			16601: out = 24'(2548);
			16602: out = 24'(2524);
			16603: out = 24'(2552);
			16604: out = 24'(2528);
			16605: out = 24'(2504);
			16606: out = 24'(2552);
			16607: out = 24'(2512);
			16608: out = 24'(2536);
			16609: out = 24'(2492);
			16610: out = 24'(2568);
			16611: out = 24'(2524);
			16612: out = 24'(2552);
			16613: out = 24'(2488);
			16614: out = 24'(2552);
			16615: out = 24'(2536);
			16616: out = 24'(2500);
			16617: out = 24'(2512);
			16618: out = 24'(2500);
			16619: out = 24'(2528);
			16620: out = 24'(2532);
			16621: out = 24'(2484);
			16622: out = 24'(2528);
			16623: out = 24'(2488);
			16624: out = 24'(2492);
			16625: out = 24'(2488);
			16626: out = 24'(2504);
			16627: out = 24'(2488);
			16628: out = 24'(2492);
			16629: out = 24'(2512);
			16630: out = 24'(2476);
			16631: out = 24'(2476);
			16632: out = 24'(2524);
			16633: out = 24'(2472);
			16634: out = 24'(2456);
			16635: out = 24'(2516);
			16636: out = 24'(2456);
			16637: out = 24'(2540);
			16638: out = 24'(2464);
			16639: out = 24'(2480);
			16640: out = 24'(2456);
			16641: out = 24'(2544);
			16642: out = 24'(2444);
			16643: out = 24'(2476);
			16644: out = 24'(2476);
			16645: out = 24'(2512);
			16646: out = 24'(2420);
			16647: out = 24'(2488);
			16648: out = 24'(2440);
			16649: out = 24'(2472);
			16650: out = 24'(2464);
			16651: out = 24'(2428);
			16652: out = 24'(2476);
			16653: out = 24'(2444);
			16654: out = 24'(2456);
			16655: out = 24'(2404);
			16656: out = 24'(2440);
			16657: out = 24'(2428);
			16658: out = 24'(2400);
			16659: out = 24'(2384);
			16660: out = 24'(2408);
			16661: out = 24'(2408);
			16662: out = 24'(2372);
			16663: out = 24'(2368);
			16664: out = 24'(2392);
			16665: out = 24'(2384);
			16666: out = 24'(2360);
			16667: out = 24'(2300);
			16668: out = 24'(2392);
			16669: out = 24'(2324);
			16670: out = 24'(2320);
			16671: out = 24'(2292);
			16672: out = 24'(2332);
			16673: out = 24'(2268);
			16674: out = 24'(2276);
			16675: out = 24'(2260);
			16676: out = 24'(2232);
			16677: out = 24'(2292);
			16678: out = 24'(2180);
			16679: out = 24'(2228);
			16680: out = 24'(2196);
			16681: out = 24'(2212);
			16682: out = 24'(2188);
			16683: out = 24'(2096);
			16684: out = 24'(2172);
			16685: out = 24'(2132);
			16686: out = 24'(2132);
			16687: out = 24'(2088);
			16688: out = 24'(2104);
			16689: out = 24'(2068);
			16690: out = 24'(2068);
			16691: out = 24'(2048);
			16692: out = 24'(2020);
			16693: out = 24'(1996);
			16694: out = 24'(2016);
			16695: out = 24'(1968);
			16696: out = 24'(1908);
			16697: out = 24'(1972);
			16698: out = 24'(1908);
			16699: out = 24'(1864);
			16700: out = 24'(1908);
			16701: out = 24'(1872);
			16702: out = 24'(1836);
			16703: out = 24'(1836);
			16704: out = 24'(1816);
			16705: out = 24'(1804);
			16706: out = 24'(1756);
			16707: out = 24'(1768);
			16708: out = 24'(1780);
			16709: out = 24'(1696);
			16710: out = 24'(1724);
			16711: out = 24'(1688);
			16712: out = 24'(1700);
			16713: out = 24'(1648);
			16714: out = 24'(1628);
			16715: out = 24'(1632);
			16716: out = 24'(1616);
			16717: out = 24'(1604);
			16718: out = 24'(1580);
			16719: out = 24'(1556);
			16720: out = 24'(1568);
			16721: out = 24'(1484);
			16722: out = 24'(1508);
			16723: out = 24'(1516);
			16724: out = 24'(1452);
			16725: out = 24'(1432);
			16726: out = 24'(1440);
			16727: out = 24'(1416);
			16728: out = 24'(1388);
			16729: out = 24'(1396);
			16730: out = 24'(1356);
			16731: out = 24'(1380);
			16732: out = 24'(1332);
			16733: out = 24'(1316);
			16734: out = 24'(1308);
			16735: out = 24'(1296);
			16736: out = 24'(1248);
			16737: out = 24'(1240);
			16738: out = 24'(1244);
			16739: out = 24'(1196);
			16740: out = 24'(1256);
			16741: out = 24'(1168);
			16742: out = 24'(1172);
			16743: out = 24'(1156);
			16744: out = 24'(1184);
			16745: out = 24'(1128);
			16746: out = 24'(1104);
			16747: out = 24'(1120);
			16748: out = 24'(1068);
			16749: out = 24'(1048);
			16750: out = 24'(1056);
			16751: out = 24'(1064);
			16752: out = 24'(1020);
			16753: out = 24'(1044);
			16754: out = 24'(980);
			16755: out = 24'(1004);
			16756: out = 24'(980);
			16757: out = 24'(952);
			16758: out = 24'(924);
			16759: out = 24'(912);
			16760: out = 24'(924);
			16761: out = 24'(920);
			16762: out = 24'(880);
			16763: out = 24'(888);
			16764: out = 24'(880);
			16765: out = 24'(828);
			16766: out = 24'(872);
			16767: out = 24'(808);
			16768: out = 24'(808);
			16769: out = 24'(812);
			16770: out = 24'(764);
			16771: out = 24'(808);
			16772: out = 24'(740);
			16773: out = 24'(764);
			16774: out = 24'(740);
			16775: out = 24'(744);
			16776: out = 24'(704);
			16777: out = 24'(700);
			16778: out = 24'(696);
			16779: out = 24'(672);
			16780: out = 24'(692);
			16781: out = 24'(640);
			16782: out = 24'(636);
			16783: out = 24'(644);
			16784: out = 24'(644);
			16785: out = 24'(608);
			16786: out = 24'(592);
			16787: out = 24'(596);
			16788: out = 24'(640);
			16789: out = 24'(544);
			16790: out = 24'(580);
			16791: out = 24'(584);
			16792: out = 24'(536);
			16793: out = 24'(496);
			16794: out = 24'(548);
			16795: out = 24'(532);
			16796: out = 24'(496);
			16797: out = 24'(492);
			16798: out = 24'(516);
			16799: out = 24'(476);
			16800: out = 24'(484);
			16801: out = 24'(448);
			16802: out = 24'(456);
			16803: out = 24'(448);
			16804: out = 24'(440);
			16805: out = 24'(456);
			16806: out = 24'(408);
			16807: out = 24'(444);
			16808: out = 24'(368);
			16809: out = 24'(444);
			16810: out = 24'(388);
			16811: out = 24'(396);
			16812: out = 24'(388);
			16813: out = 24'(384);
			16814: out = 24'(340);
			16815: out = 24'(384);
			16816: out = 24'(352);
			16817: out = 24'(256);
			16818: out = 24'(344);
			16819: out = 24'(256);
			16820: out = 24'(268);
			16821: out = 24'(240);
			16822: out = 24'(216);
			16823: out = 24'(192);
			16824: out = 24'(200);
			16825: out = 24'(164);
			16826: out = 24'(132);
			16827: out = 24'(120);
			16828: out = 24'(124);
			16829: out = 24'(40);
			16830: out = 24'(52);
			16831: out = 24'(60);
			16832: out = 24'(12);
			16833: out = 24'(20);
			16834: out = 24'(-28);
			16835: out = 24'(-16);
			16836: out = 24'(-28);
			16837: out = 24'(-64);
			16838: out = 24'(-72);
			16839: out = 24'(-128);
			16840: out = 24'(-64);
			16841: out = 24'(-148);
			16842: out = 24'(-124);
			16843: out = 24'(-168);
			16844: out = 24'(-152);
			16845: out = 24'(-220);
			16846: out = 24'(-160);
			16847: out = 24'(-244);
			16848: out = 24'(-212);
			16849: out = 24'(-248);
			16850: out = 24'(-260);
			16851: out = 24'(-252);
			16852: out = 24'(-300);
			16853: out = 24'(-296);
			16854: out = 24'(-292);
			16855: out = 24'(-340);
			16856: out = 24'(-340);
			16857: out = 24'(-348);
			16858: out = 24'(-360);
			16859: out = 24'(-384);
			16860: out = 24'(-408);
			16861: out = 24'(-388);
			16862: out = 24'(-444);
			16863: out = 24'(-420);
			16864: out = 24'(-492);
			16865: out = 24'(-412);
			16866: out = 24'(-492);
			16867: out = 24'(-480);
			16868: out = 24'(-508);
			16869: out = 24'(-500);
			16870: out = 24'(-500);
			16871: out = 24'(-552);
			16872: out = 24'(-528);
			16873: out = 24'(-564);
			16874: out = 24'(-576);
			16875: out = 24'(-580);
			16876: out = 24'(-592);
			16877: out = 24'(-640);
			16878: out = 24'(-624);
			16879: out = 24'(-596);
			16880: out = 24'(-692);
			16881: out = 24'(-656);
			16882: out = 24'(-680);
			16883: out = 24'(-644);
			16884: out = 24'(-724);
			16885: out = 24'(-704);
			16886: out = 24'(-712);
			16887: out = 24'(-732);
			16888: out = 24'(-724);
			16889: out = 24'(-772);
			16890: out = 24'(-744);
			16891: out = 24'(-764);
			16892: out = 24'(-796);
			16893: out = 24'(-764);
			16894: out = 24'(-848);
			16895: out = 24'(-832);
			16896: out = 24'(-820);
			16897: out = 24'(-868);
			16898: out = 24'(-844);
			16899: out = 24'(-916);
			16900: out = 24'(-840);
			16901: out = 24'(-908);
			16902: out = 24'(-900);
			16903: out = 24'(-940);
			16904: out = 24'(-940);
			16905: out = 24'(-936);
			16906: out = 24'(-972);
			16907: out = 24'(-972);
			16908: out = 24'(-996);
			16909: out = 24'(-996);
			16910: out = 24'(-1044);
			16911: out = 24'(-1064);
			16912: out = 24'(-1044);
			16913: out = 24'(-1080);
			16914: out = 24'(-1100);
			16915: out = 24'(-1100);
			16916: out = 24'(-1132);
			16917: out = 24'(-1120);
			16918: out = 24'(-1144);
			16919: out = 24'(-1220);
			16920: out = 24'(-1168);
			16921: out = 24'(-1192);
			16922: out = 24'(-1248);
			16923: out = 24'(-1208);
			16924: out = 24'(-1280);
			16925: out = 24'(-1264);
			16926: out = 24'(-1304);
			16927: out = 24'(-1292);
			16928: out = 24'(-1348);
			16929: out = 24'(-1360);
			16930: out = 24'(-1356);
			16931: out = 24'(-1396);
			16932: out = 24'(-1436);
			16933: out = 24'(-1416);
			16934: out = 24'(-1428);
			16935: out = 24'(-1492);
			16936: out = 24'(-1516);
			16937: out = 24'(-1472);
			16938: out = 24'(-1564);
			16939: out = 24'(-1556);
			16940: out = 24'(-1584);
			16941: out = 24'(-1648);
			16942: out = 24'(-1628);
			16943: out = 24'(-1648);
			16944: out = 24'(-1660);
			16945: out = 24'(-1740);
			16946: out = 24'(-1720);
			16947: out = 24'(-1752);
			16948: out = 24'(-1760);
			16949: out = 24'(-1828);
			16950: out = 24'(-1816);
			16951: out = 24'(-1840);
			16952: out = 24'(-1832);
			16953: out = 24'(-1868);
			16954: out = 24'(-1924);
			16955: out = 24'(-1932);
			16956: out = 24'(-1936);
			16957: out = 24'(-1976);
			16958: out = 24'(-2016);
			16959: out = 24'(-2024);
			16960: out = 24'(-2072);
			16961: out = 24'(-2020);
			16962: out = 24'(-2100);
			16963: out = 24'(-2108);
			16964: out = 24'(-2108);
			16965: out = 24'(-2168);
			16966: out = 24'(-2124);
			16967: out = 24'(-2212);
			16968: out = 24'(-2216);
			16969: out = 24'(-2240);
			16970: out = 24'(-2240);
			16971: out = 24'(-2268);
			16972: out = 24'(-2236);
			16973: out = 24'(-2308);
			16974: out = 24'(-2300);
			16975: out = 24'(-2324);
			16976: out = 24'(-2360);
			16977: out = 24'(-2380);
			16978: out = 24'(-2360);
			16979: out = 24'(-2408);
			16980: out = 24'(-2420);
			16981: out = 24'(-2392);
			16982: out = 24'(-2484);
			16983: out = 24'(-2408);
			16984: out = 24'(-2472);
			16985: out = 24'(-2500);
			16986: out = 24'(-2496);
			16987: out = 24'(-2492);
			16988: out = 24'(-2516);
			16989: out = 24'(-2528);
			16990: out = 24'(-2532);
			16991: out = 24'(-2544);
			16992: out = 24'(-2568);
			16993: out = 24'(-2564);
			16994: out = 24'(-2608);
			16995: out = 24'(-2568);
			16996: out = 24'(-2580);
			16997: out = 24'(-2636);
			16998: out = 24'(-2584);
			16999: out = 24'(-2616);
			17000: out = 24'(-2632);
			17001: out = 24'(-2604);
			17002: out = 24'(-2668);
			17003: out = 24'(-2624);
			17004: out = 24'(-2660);
			17005: out = 24'(-2640);
			17006: out = 24'(-2672);
			17007: out = 24'(-2664);
			17008: out = 24'(-2700);
			17009: out = 24'(-2704);
			17010: out = 24'(-2656);
			17011: out = 24'(-2688);
			17012: out = 24'(-2708);
			17013: out = 24'(-2668);
			17014: out = 24'(-2740);
			17015: out = 24'(-2676);
			17016: out = 24'(-2724);
			17017: out = 24'(-2748);
			17018: out = 24'(-2716);
			17019: out = 24'(-2720);
			17020: out = 24'(-2724);
			17021: out = 24'(-2712);
			17022: out = 24'(-2756);
			17023: out = 24'(-2684);
			17024: out = 24'(-2752);
			17025: out = 24'(-2732);
			17026: out = 24'(-2748);
			17027: out = 24'(-2732);
			17028: out = 24'(-2760);
			17029: out = 24'(-2732);
			17030: out = 24'(-2764);
			17031: out = 24'(-2724);
			17032: out = 24'(-2752);
			17033: out = 24'(-2764);
			17034: out = 24'(-2728);
			17035: out = 24'(-2756);
			17036: out = 24'(-2748);
			17037: out = 24'(-2748);
			17038: out = 24'(-2740);
			17039: out = 24'(-2740);
			17040: out = 24'(-2736);
			17041: out = 24'(-2780);
			17042: out = 24'(-2716);
			17043: out = 24'(-2736);
			17044: out = 24'(-2736);
			17045: out = 24'(-2732);
			17046: out = 24'(-2728);
			17047: out = 24'(-2720);
			17048: out = 24'(-2724);
			17049: out = 24'(-2736);
			17050: out = 24'(-2712);
			17051: out = 24'(-2764);
			17052: out = 24'(-2716);
			17053: out = 24'(-2684);
			17054: out = 24'(-2748);
			17055: out = 24'(-2708);
			17056: out = 24'(-2716);
			17057: out = 24'(-2688);
			17058: out = 24'(-2716);
			17059: out = 24'(-2716);
			17060: out = 24'(-2652);
			17061: out = 24'(-2732);
			17062: out = 24'(-2656);
			17063: out = 24'(-2712);
			17064: out = 24'(-2680);
			17065: out = 24'(-2688);
			17066: out = 24'(-2636);
			17067: out = 24'(-2692);
			17068: out = 24'(-2664);
			17069: out = 24'(-2640);
			17070: out = 24'(-2676);
			17071: out = 24'(-2608);
			17072: out = 24'(-2672);
			17073: out = 24'(-2636);
			17074: out = 24'(-2624);
			17075: out = 24'(-2660);
			17076: out = 24'(-2624);
			17077: out = 24'(-2616);
			17078: out = 24'(-2628);
			17079: out = 24'(-2608);
			17080: out = 24'(-2624);
			17081: out = 24'(-2584);
			17082: out = 24'(-2572);
			17083: out = 24'(-2596);
			17084: out = 24'(-2580);
			17085: out = 24'(-2572);
			17086: out = 24'(-2564);
			17087: out = 24'(-2568);
			17088: out = 24'(-2584);
			17089: out = 24'(-2552);
			17090: out = 24'(-2564);
			17091: out = 24'(-2564);
			17092: out = 24'(-2532);
			17093: out = 24'(-2544);
			17094: out = 24'(-2532);
			17095: out = 24'(-2516);
			17096: out = 24'(-2516);
			17097: out = 24'(-2516);
			17098: out = 24'(-2492);
			17099: out = 24'(-2524);
			17100: out = 24'(-2440);
			17101: out = 24'(-2520);
			17102: out = 24'(-2488);
			17103: out = 24'(-2440);
			17104: out = 24'(-2468);
			17105: out = 24'(-2452);
			17106: out = 24'(-2420);
			17107: out = 24'(-2440);
			17108: out = 24'(-2440);
			17109: out = 24'(-2396);
			17110: out = 24'(-2416);
			17111: out = 24'(-2380);
			17112: out = 24'(-2408);
			17113: out = 24'(-2376);
			17114: out = 24'(-2352);
			17115: out = 24'(-2388);
			17116: out = 24'(-2332);
			17117: out = 24'(-2348);
			17118: out = 24'(-2356);
			17119: out = 24'(-2328);
			17120: out = 24'(-2304);
			17121: out = 24'(-2304);
			17122: out = 24'(-2292);
			17123: out = 24'(-2304);
			17124: out = 24'(-2240);
			17125: out = 24'(-2268);
			17126: out = 24'(-2256);
			17127: out = 24'(-2228);
			17128: out = 24'(-2192);
			17129: out = 24'(-2208);
			17130: out = 24'(-2184);
			17131: out = 24'(-2196);
			17132: out = 24'(-2160);
			17133: out = 24'(-2132);
			17134: out = 24'(-2140);
			17135: out = 24'(-2188);
			17136: out = 24'(-2064);
			17137: out = 24'(-2120);
			17138: out = 24'(-2052);
			17139: out = 24'(-2096);
			17140: out = 24'(-2036);
			17141: out = 24'(-2040);
			17142: out = 24'(-2008);
			17143: out = 24'(-2000);
			17144: out = 24'(-1976);
			17145: out = 24'(-1960);
			17146: out = 24'(-1956);
			17147: out = 24'(-1916);
			17148: out = 24'(-1904);
			17149: out = 24'(-1872);
			17150: out = 24'(-1920);
			17151: out = 24'(-1840);
			17152: out = 24'(-1852);
			17153: out = 24'(-1820);
			17154: out = 24'(-1800);
			17155: out = 24'(-1812);
			17156: out = 24'(-1752);
			17157: out = 24'(-1744);
			17158: out = 24'(-1712);
			17159: out = 24'(-1716);
			17160: out = 24'(-1728);
			17161: out = 24'(-1616);
			17162: out = 24'(-1680);
			17163: out = 24'(-1664);
			17164: out = 24'(-1588);
			17165: out = 24'(-1588);
			17166: out = 24'(-1580);
			17167: out = 24'(-1580);
			17168: out = 24'(-1524);
			17169: out = 24'(-1524);
			17170: out = 24'(-1516);
			17171: out = 24'(-1496);
			17172: out = 24'(-1476);
			17173: out = 24'(-1468);
			17174: out = 24'(-1424);
			17175: out = 24'(-1428);
			17176: out = 24'(-1424);
			17177: out = 24'(-1380);
			17178: out = 24'(-1360);
			17179: out = 24'(-1400);
			17180: out = 24'(-1320);
			17181: out = 24'(-1376);
			17182: out = 24'(-1304);
			17183: out = 24'(-1288);
			17184: out = 24'(-1308);
			17185: out = 24'(-1244);
			17186: out = 24'(-1280);
			17187: out = 24'(-1220);
			17188: out = 24'(-1232);
			17189: out = 24'(-1176);
			17190: out = 24'(-1212);
			17191: out = 24'(-1144);
			17192: out = 24'(-1176);
			17193: out = 24'(-1120);
			17194: out = 24'(-1108);
			17195: out = 24'(-1128);
			17196: out = 24'(-1104);
			17197: out = 24'(-1060);
			17198: out = 24'(-1076);
			17199: out = 24'(-1064);
			17200: out = 24'(-1048);
			17201: out = 24'(-1032);
			17202: out = 24'(-1000);
			17203: out = 24'(-1060);
			17204: out = 24'(-928);
			17205: out = 24'(-1016);
			17206: out = 24'(-940);
			17207: out = 24'(-936);
			17208: out = 24'(-956);
			17209: out = 24'(-928);
			17210: out = 24'(-920);
			17211: out = 24'(-876);
			17212: out = 24'(-876);
			17213: out = 24'(-884);
			17214: out = 24'(-856);
			17215: out = 24'(-868);
			17216: out = 24'(-832);
			17217: out = 24'(-824);
			17218: out = 24'(-820);
			17219: out = 24'(-832);
			17220: out = 24'(-772);
			17221: out = 24'(-784);
			17222: out = 24'(-780);
			17223: out = 24'(-772);
			17224: out = 24'(-720);
			17225: out = 24'(-796);
			17226: out = 24'(-712);
			17227: out = 24'(-720);
			17228: out = 24'(-736);
			17229: out = 24'(-680);
			17230: out = 24'(-724);
			17231: out = 24'(-688);
			17232: out = 24'(-680);
			17233: out = 24'(-656);
			17234: out = 24'(-640);
			17235: out = 24'(-684);
			17236: out = 24'(-616);
			17237: out = 24'(-616);
			17238: out = 24'(-656);
			17239: out = 24'(-608);
			17240: out = 24'(-588);
			17241: out = 24'(-592);
			17242: out = 24'(-580);
			17243: out = 24'(-552);
			17244: out = 24'(-524);
			17245: out = 24'(-512);
			17246: out = 24'(-516);
			17247: out = 24'(-444);
			17248: out = 24'(-512);
			17249: out = 24'(-460);
			17250: out = 24'(-416);
			17251: out = 24'(-460);
			17252: out = 24'(-420);
			17253: out = 24'(-400);
			17254: out = 24'(-392);
			17255: out = 24'(-380);
			17256: out = 24'(-380);
			17257: out = 24'(-356);
			17258: out = 24'(-356);
			17259: out = 24'(-308);
			17260: out = 24'(-304);
			17261: out = 24'(-332);
			17262: out = 24'(-304);
			17263: out = 24'(-232);
			17264: out = 24'(-312);
			17265: out = 24'(-244);
			17266: out = 24'(-268);
			17267: out = 24'(-200);
			17268: out = 24'(-212);
			17269: out = 24'(-216);
			17270: out = 24'(-208);
			17271: out = 24'(-176);
			17272: out = 24'(-160);
			17273: out = 24'(-176);
			17274: out = 24'(-160);
			17275: out = 24'(-160);
			17276: out = 24'(-164);
			17277: out = 24'(-96);
			17278: out = 24'(-132);
			17279: out = 24'(-144);
			17280: out = 24'(-84);
			17281: out = 24'(-84);
			17282: out = 24'(-60);
			17283: out = 24'(-64);
			17284: out = 24'(-88);
			17285: out = 24'(-60);
			17286: out = 24'(-36);
			17287: out = 24'(-32);
			17288: out = 24'(-32);
			17289: out = 24'(-20);
			17290: out = 24'(-20);
			17291: out = 24'(24);
			17292: out = 24'(-24);
			17293: out = 24'(16);
			17294: out = 24'(24);
			17295: out = 24'(68);
			17296: out = 24'(52);
			17297: out = 24'(8);
			17298: out = 24'(80);
			17299: out = 24'(84);
			17300: out = 24'(84);
			17301: out = 24'(84);
			17302: out = 24'(80);
			17303: out = 24'(104);
			17304: out = 24'(136);
			17305: out = 24'(112);
			17306: out = 24'(136);
			17307: out = 24'(144);
			17308: out = 24'(152);
			17309: out = 24'(180);
			17310: out = 24'(164);
			17311: out = 24'(164);
			17312: out = 24'(216);
			17313: out = 24'(172);
			17314: out = 24'(180);
			17315: out = 24'(212);
			17316: out = 24'(224);
			17317: out = 24'(208);
			17318: out = 24'(248);
			17319: out = 24'(232);
			17320: out = 24'(268);
			17321: out = 24'(216);
			17322: out = 24'(300);
			17323: out = 24'(268);
			17324: out = 24'(268);
			17325: out = 24'(332);
			17326: out = 24'(256);
			17327: out = 24'(340);
			17328: out = 24'(316);
			17329: out = 24'(340);
			17330: out = 24'(372);
			17331: out = 24'(348);
			17332: out = 24'(384);
			17333: out = 24'(404);
			17334: out = 24'(412);
			17335: out = 24'(408);
			17336: out = 24'(412);
			17337: out = 24'(428);
			17338: out = 24'(484);
			17339: out = 24'(440);
			17340: out = 24'(452);
			17341: out = 24'(488);
			17342: out = 24'(532);
			17343: out = 24'(504);
			17344: out = 24'(500);
			17345: out = 24'(576);
			17346: out = 24'(552);
			17347: out = 24'(572);
			17348: out = 24'(536);
			17349: out = 24'(620);
			17350: out = 24'(588);
			17351: out = 24'(608);
			17352: out = 24'(632);
			17353: out = 24'(644);
			17354: out = 24'(680);
			17355: out = 24'(668);
			17356: out = 24'(704);
			17357: out = 24'(716);
			17358: out = 24'(704);
			17359: out = 24'(732);
			17360: out = 24'(776);
			17361: out = 24'(740);
			17362: out = 24'(824);
			17363: out = 24'(796);
			17364: out = 24'(808);
			17365: out = 24'(864);
			17366: out = 24'(840);
			17367: out = 24'(848);
			17368: out = 24'(884);
			17369: out = 24'(932);
			17370: out = 24'(936);
			17371: out = 24'(952);
			17372: out = 24'(912);
			17373: out = 24'(1016);
			17374: out = 24'(980);
			17375: out = 24'(1004);
			17376: out = 24'(1020);
			17377: out = 24'(1028);
			17378: out = 24'(1048);
			17379: out = 24'(1064);
			17380: out = 24'(1104);
			17381: out = 24'(1076);
			17382: out = 24'(1140);
			17383: out = 24'(1116);
			17384: out = 24'(1112);
			17385: out = 24'(1184);
			17386: out = 24'(1164);
			17387: out = 24'(1148);
			17388: out = 24'(1224);
			17389: out = 24'(1188);
			17390: out = 24'(1252);
			17391: out = 24'(1236);
			17392: out = 24'(1260);
			17393: out = 24'(1264);
			17394: out = 24'(1316);
			17395: out = 24'(1260);
			17396: out = 24'(1304);
			17397: out = 24'(1336);
			17398: out = 24'(1316);
			17399: out = 24'(1364);
			17400: out = 24'(1332);
			17401: out = 24'(1360);
			17402: out = 24'(1360);
			17403: out = 24'(1400);
			17404: out = 24'(1360);
			17405: out = 24'(1432);
			17406: out = 24'(1408);
			17407: out = 24'(1444);
			17408: out = 24'(1456);
			17409: out = 24'(1456);
			17410: out = 24'(1500);
			17411: out = 24'(1488);
			17412: out = 24'(1492);
			17413: out = 24'(1496);
			17414: out = 24'(1532);
			17415: out = 24'(1520);
			17416: out = 24'(1536);
			17417: out = 24'(1524);
			17418: out = 24'(1588);
			17419: out = 24'(1572);
			17420: out = 24'(1544);
			17421: out = 24'(1604);
			17422: out = 24'(1612);
			17423: out = 24'(1612);
			17424: out = 24'(1600);
			17425: out = 24'(1596);
			17426: out = 24'(1652);
			17427: out = 24'(1668);
			17428: out = 24'(1652);
			17429: out = 24'(1636);
			17430: out = 24'(1680);
			17431: out = 24'(1720);
			17432: out = 24'(1672);
			17433: out = 24'(1688);
			17434: out = 24'(1720);
			17435: out = 24'(1752);
			17436: out = 24'(1688);
			17437: out = 24'(1728);
			17438: out = 24'(1756);
			17439: out = 24'(1712);
			17440: out = 24'(1776);
			17441: out = 24'(1764);
			17442: out = 24'(1776);
			17443: out = 24'(1764);
			17444: out = 24'(1800);
			17445: out = 24'(1824);
			17446: out = 24'(1768);
			17447: out = 24'(1824);
			17448: out = 24'(1800);
			17449: out = 24'(1820);
			17450: out = 24'(1860);
			17451: out = 24'(1824);
			17452: out = 24'(1896);
			17453: out = 24'(1820);
			17454: out = 24'(1872);
			17455: out = 24'(1860);
			17456: out = 24'(1868);
			17457: out = 24'(1908);
			17458: out = 24'(1876);
			17459: out = 24'(1880);
			17460: out = 24'(1944);
			17461: out = 24'(1876);
			17462: out = 24'(1952);
			17463: out = 24'(1912);
			17464: out = 24'(1932);
			17465: out = 24'(1944);
			17466: out = 24'(1956);
			17467: out = 24'(1952);
			17468: out = 24'(1956);
			17469: out = 24'(1952);
			17470: out = 24'(1948);
			17471: out = 24'(1960);
			17472: out = 24'(1956);
			17473: out = 24'(1964);
			17474: out = 24'(1968);
			17475: out = 24'(1980);
			17476: out = 24'(1928);
			17477: out = 24'(2000);
			17478: out = 24'(1964);
			17479: out = 24'(1956);
			17480: out = 24'(1972);
			17481: out = 24'(1976);
			17482: out = 24'(1956);
			17483: out = 24'(1968);
			17484: out = 24'(2000);
			17485: out = 24'(1920);
			17486: out = 24'(2000);
			17487: out = 24'(1912);
			17488: out = 24'(2004);
			17489: out = 24'(1924);
			17490: out = 24'(1948);
			17491: out = 24'(2000);
			17492: out = 24'(1972);
			17493: out = 24'(1956);
			17494: out = 24'(1972);
			17495: out = 24'(1992);
			17496: out = 24'(1944);
			17497: out = 24'(1972);
			17498: out = 24'(1936);
			17499: out = 24'(1928);
			17500: out = 24'(1960);
			17501: out = 24'(1948);
			17502: out = 24'(1896);
			17503: out = 24'(1956);
			17504: out = 24'(1928);
			17505: out = 24'(1920);
			17506: out = 24'(1924);
			17507: out = 24'(1932);
			17508: out = 24'(1928);
			17509: out = 24'(1932);
			17510: out = 24'(1920);
			17511: out = 24'(1960);
			17512: out = 24'(1900);
			17513: out = 24'(1936);
			17514: out = 24'(1948);
			17515: out = 24'(1948);
			17516: out = 24'(1904);
			17517: out = 24'(1952);
			17518: out = 24'(1916);
			17519: out = 24'(1948);
			17520: out = 24'(1880);
			17521: out = 24'(1920);
			17522: out = 24'(1896);
			17523: out = 24'(1928);
			17524: out = 24'(1872);
			17525: out = 24'(1932);
			17526: out = 24'(1920);
			17527: out = 24'(1908);
			17528: out = 24'(1916);
			17529: out = 24'(1880);
			17530: out = 24'(1936);
			17531: out = 24'(1896);
			17532: out = 24'(1848);
			17533: out = 24'(1932);
			17534: out = 24'(1888);
			17535: out = 24'(1880);
			17536: out = 24'(1928);
			17537: out = 24'(1884);
			17538: out = 24'(1908);
			17539: out = 24'(1896);
			17540: out = 24'(1888);
			17541: out = 24'(1868);
			17542: out = 24'(1872);
			17543: out = 24'(1884);
			17544: out = 24'(1860);
			17545: out = 24'(1848);
			17546: out = 24'(1880);
			17547: out = 24'(1856);
			17548: out = 24'(1852);
			17549: out = 24'(1876);
			17550: out = 24'(1824);
			17551: out = 24'(1868);
			17552: out = 24'(1832);
			17553: out = 24'(1852);
			17554: out = 24'(1832);
			17555: out = 24'(1804);
			17556: out = 24'(1788);
			17557: out = 24'(1820);
			17558: out = 24'(1776);
			17559: out = 24'(1740);
			17560: out = 24'(1776);
			17561: out = 24'(1760);
			17562: out = 24'(1768);
			17563: out = 24'(1724);
			17564: out = 24'(1744);
			17565: out = 24'(1716);
			17566: out = 24'(1736);
			17567: out = 24'(1720);
			17568: out = 24'(1668);
			17569: out = 24'(1692);
			17570: out = 24'(1668);
			17571: out = 24'(1712);
			17572: out = 24'(1644);
			17573: out = 24'(1632);
			17574: out = 24'(1644);
			17575: out = 24'(1668);
			17576: out = 24'(1620);
			17577: out = 24'(1612);
			17578: out = 24'(1576);
			17579: out = 24'(1620);
			17580: out = 24'(1564);
			17581: out = 24'(1556);
			17582: out = 24'(1584);
			17583: out = 24'(1516);
			17584: out = 24'(1508);
			17585: out = 24'(1548);
			17586: out = 24'(1456);
			17587: out = 24'(1488);
			17588: out = 24'(1448);
			17589: out = 24'(1480);
			17590: out = 24'(1400);
			17591: out = 24'(1436);
			17592: out = 24'(1408);
			17593: out = 24'(1396);
			17594: out = 24'(1364);
			17595: out = 24'(1360);
			17596: out = 24'(1364);
			17597: out = 24'(1332);
			17598: out = 24'(1332);
			17599: out = 24'(1312);
			17600: out = 24'(1308);
			17601: out = 24'(1280);
			17602: out = 24'(1268);
			17603: out = 24'(1296);
			17604: out = 24'(1220);
			17605: out = 24'(1216);
			17606: out = 24'(1236);
			17607: out = 24'(1220);
			17608: out = 24'(1156);
			17609: out = 24'(1164);
			17610: out = 24'(1176);
			17611: out = 24'(1144);
			17612: out = 24'(1144);
			17613: out = 24'(1132);
			17614: out = 24'(1116);
			17615: out = 24'(1080);
			17616: out = 24'(1108);
			17617: out = 24'(1032);
			17618: out = 24'(1068);
			17619: out = 24'(1032);
			17620: out = 24'(1012);
			17621: out = 24'(1048);
			17622: out = 24'(972);
			17623: out = 24'(1024);
			17624: out = 24'(964);
			17625: out = 24'(952);
			17626: out = 24'(980);
			17627: out = 24'(948);
			17628: out = 24'(892);
			17629: out = 24'(936);
			17630: out = 24'(920);
			17631: out = 24'(860);
			17632: out = 24'(880);
			17633: out = 24'(856);
			17634: out = 24'(864);
			17635: out = 24'(844);
			17636: out = 24'(788);
			17637: out = 24'(832);
			17638: out = 24'(812);
			17639: out = 24'(784);
			17640: out = 24'(772);
			17641: out = 24'(768);
			17642: out = 24'(740);
			17643: out = 24'(736);
			17644: out = 24'(744);
			17645: out = 24'(716);
			17646: out = 24'(684);
			17647: out = 24'(704);
			17648: out = 24'(680);
			17649: out = 24'(676);
			17650: out = 24'(684);
			17651: out = 24'(656);
			17652: out = 24'(644);
			17653: out = 24'(656);
			17654: out = 24'(624);
			17655: out = 24'(620);
			17656: out = 24'(596);
			17657: out = 24'(600);
			17658: out = 24'(592);
			17659: out = 24'(588);
			17660: out = 24'(556);
			17661: out = 24'(540);
			17662: out = 24'(576);
			17663: out = 24'(552);
			17664: out = 24'(480);
			17665: out = 24'(556);
			17666: out = 24'(476);
			17667: out = 24'(512);
			17668: out = 24'(496);
			17669: out = 24'(500);
			17670: out = 24'(488);
			17671: out = 24'(444);
			17672: out = 24'(476);
			17673: out = 24'(452);
			17674: out = 24'(460);
			17675: out = 24'(444);
			17676: out = 24'(372);
			17677: out = 24'(416);
			17678: out = 24'(448);
			17679: out = 24'(392);
			17680: out = 24'(392);
			17681: out = 24'(364);
			17682: out = 24'(404);
			17683: out = 24'(384);
			17684: out = 24'(352);
			17685: out = 24'(368);
			17686: out = 24'(352);
			17687: out = 24'(324);
			17688: out = 24'(320);
			17689: out = 24'(336);
			17690: out = 24'(296);
			17691: out = 24'(324);
			17692: out = 24'(296);
			17693: out = 24'(308);
			17694: out = 24'(292);
			17695: out = 24'(292);
			17696: out = 24'(260);
			17697: out = 24'(264);
			17698: out = 24'(308);
			17699: out = 24'(220);
			17700: out = 24'(212);
			17701: out = 24'(272);
			17702: out = 24'(256);
			17703: out = 24'(224);
			17704: out = 24'(204);
			17705: out = 24'(244);
			17706: out = 24'(216);
			17707: out = 24'(200);
			17708: out = 24'(176);
			17709: out = 24'(200);
			17710: out = 24'(124);
			17711: out = 24'(156);
			17712: out = 24'(144);
			17713: out = 24'(88);
			17714: out = 24'(100);
			17715: out = 24'(88);
			17716: out = 24'(56);
			17717: out = 24'(68);
			17718: out = 24'(20);
			17719: out = 24'(16);
			17720: out = 24'(20);
			17721: out = 24'(-12);
			17722: out = 24'(-24);
			17723: out = 24'(-52);
			17724: out = 24'(-20);
			17725: out = 24'(-88);
			17726: out = 24'(-24);
			17727: out = 24'(-120);
			17728: out = 24'(-84);
			17729: out = 24'(-104);
			17730: out = 24'(-116);
			17731: out = 24'(-152);
			17732: out = 24'(-128);
			17733: out = 24'(-168);
			17734: out = 24'(-128);
			17735: out = 24'(-196);
			17736: out = 24'(-192);
			17737: out = 24'(-176);
			17738: out = 24'(-228);
			17739: out = 24'(-228);
			17740: out = 24'(-240);
			17741: out = 24'(-228);
			17742: out = 24'(-256);
			17743: out = 24'(-276);
			17744: out = 24'(-252);
			17745: out = 24'(-288);
			17746: out = 24'(-332);
			17747: out = 24'(-292);
			17748: out = 24'(-304);
			17749: out = 24'(-296);
			17750: out = 24'(-372);
			17751: out = 24'(-364);
			17752: out = 24'(-324);
			17753: out = 24'(-380);
			17754: out = 24'(-388);
			17755: out = 24'(-388);
			17756: out = 24'(-388);
			17757: out = 24'(-408);
			17758: out = 24'(-412);
			17759: out = 24'(-432);
			17760: out = 24'(-416);
			17761: out = 24'(-440);
			17762: out = 24'(-448);
			17763: out = 24'(-496);
			17764: out = 24'(-444);
			17765: out = 24'(-456);
			17766: out = 24'(-544);
			17767: out = 24'(-492);
			17768: out = 24'(-524);
			17769: out = 24'(-488);
			17770: out = 24'(-556);
			17771: out = 24'(-548);
			17772: out = 24'(-532);
			17773: out = 24'(-584);
			17774: out = 24'(-540);
			17775: out = 24'(-580);
			17776: out = 24'(-620);
			17777: out = 24'(-564);
			17778: out = 24'(-600);
			17779: out = 24'(-604);
			17780: out = 24'(-624);
			17781: out = 24'(-608);
			17782: out = 24'(-680);
			17783: out = 24'(-616);
			17784: out = 24'(-676);
			17785: out = 24'(-676);
			17786: out = 24'(-636);
			17787: out = 24'(-736);
			17788: out = 24'(-728);
			17789: out = 24'(-672);
			17790: out = 24'(-716);
			17791: out = 24'(-732);
			17792: out = 24'(-732);
			17793: out = 24'(-772);
			17794: out = 24'(-732);
			17795: out = 24'(-780);
			17796: out = 24'(-784);
			17797: out = 24'(-836);
			17798: out = 24'(-776);
			17799: out = 24'(-820);
			17800: out = 24'(-824);
			17801: out = 24'(-816);
			17802: out = 24'(-844);
			17803: out = 24'(-864);
			17804: out = 24'(-856);
			17805: out = 24'(-872);
			17806: out = 24'(-884);
			17807: out = 24'(-928);
			17808: out = 24'(-916);
			17809: out = 24'(-940);
			17810: out = 24'(-940);
			17811: out = 24'(-952);
			17812: out = 24'(-988);
			17813: out = 24'(-980);
			17814: out = 24'(-984);
			17815: out = 24'(-1016);
			17816: out = 24'(-1020);
			17817: out = 24'(-1012);
			17818: out = 24'(-1100);
			17819: out = 24'(-1084);
			17820: out = 24'(-1044);
			17821: out = 24'(-1128);
			17822: out = 24'(-1108);
			17823: out = 24'(-1116);
			17824: out = 24'(-1192);
			17825: out = 24'(-1188);
			17826: out = 24'(-1176);
			17827: out = 24'(-1188);
			17828: out = 24'(-1240);
			17829: out = 24'(-1244);
			17830: out = 24'(-1240);
			17831: out = 24'(-1272);
			17832: out = 24'(-1256);
			17833: out = 24'(-1356);
			17834: out = 24'(-1352);
			17835: out = 24'(-1300);
			17836: out = 24'(-1392);
			17837: out = 24'(-1368);
			17838: out = 24'(-1400);
			17839: out = 24'(-1392);
			17840: out = 24'(-1460);
			17841: out = 24'(-1444);
			17842: out = 24'(-1448);
			17843: out = 24'(-1492);
			17844: out = 24'(-1516);
			17845: out = 24'(-1528);
			17846: out = 24'(-1564);
			17847: out = 24'(-1564);
			17848: out = 24'(-1564);
			17849: out = 24'(-1600);
			17850: out = 24'(-1640);
			17851: out = 24'(-1620);
			17852: out = 24'(-1640);
			17853: out = 24'(-1660);
			17854: out = 24'(-1644);
			17855: out = 24'(-1756);
			17856: out = 24'(-1696);
			17857: out = 24'(-1712);
			17858: out = 24'(-1736);
			17859: out = 24'(-1736);
			17860: out = 24'(-1780);
			17861: out = 24'(-1804);
			17862: out = 24'(-1804);
			17863: out = 24'(-1768);
			17864: out = 24'(-1872);
			17865: out = 24'(-1848);
			17866: out = 24'(-1856);
			17867: out = 24'(-1848);
			17868: out = 24'(-1848);
			17869: out = 24'(-1936);
			17870: out = 24'(-1868);
			17871: out = 24'(-1908);
			17872: out = 24'(-1888);
			17873: out = 24'(-1964);
			17874: out = 24'(-1952);
			17875: out = 24'(-1932);
			17876: out = 24'(-1932);
			17877: out = 24'(-2004);
			17878: out = 24'(-1960);
			17879: out = 24'(-1972);
			17880: out = 24'(-2012);
			17881: out = 24'(-1984);
			17882: out = 24'(-2024);
			17883: out = 24'(-2028);
			17884: out = 24'(-2020);
			17885: out = 24'(-2064);
			17886: out = 24'(-2040);
			17887: out = 24'(-2044);
			17888: out = 24'(-2072);
			17889: out = 24'(-2088);
			17890: out = 24'(-2052);
			17891: out = 24'(-2088);
			17892: out = 24'(-2104);
			17893: out = 24'(-2084);
			17894: out = 24'(-2072);
			17895: out = 24'(-2140);
			17896: out = 24'(-2104);
			17897: out = 24'(-2116);
			17898: out = 24'(-2120);
			17899: out = 24'(-2132);
			17900: out = 24'(-2160);
			17901: out = 24'(-2076);
			17902: out = 24'(-2124);
			17903: out = 24'(-2136);
			17904: out = 24'(-2124);
			17905: out = 24'(-2100);
			17906: out = 24'(-2140);
			17907: out = 24'(-2148);
			17908: out = 24'(-2152);
			17909: out = 24'(-2148);
			17910: out = 24'(-2132);
			17911: out = 24'(-2168);
			17912: out = 24'(-2160);
			17913: out = 24'(-2124);
			17914: out = 24'(-2156);
			17915: out = 24'(-2156);
			17916: out = 24'(-2172);
			17917: out = 24'(-2124);
			17918: out = 24'(-2164);
			17919: out = 24'(-2168);
			17920: out = 24'(-2132);
			17921: out = 24'(-2184);
			17922: out = 24'(-2204);
			17923: out = 24'(-2100);
			17924: out = 24'(-2212);
			17925: out = 24'(-2136);
			17926: out = 24'(-2188);
			17927: out = 24'(-2160);
			17928: out = 24'(-2156);
			17929: out = 24'(-2184);
			17930: out = 24'(-2136);
			17931: out = 24'(-2160);
			17932: out = 24'(-2160);
			17933: out = 24'(-2148);
			17934: out = 24'(-2148);
			17935: out = 24'(-2156);
			17936: out = 24'(-2180);
			17937: out = 24'(-2148);
			17938: out = 24'(-2148);
			17939: out = 24'(-2188);
			17940: out = 24'(-2148);
			17941: out = 24'(-2168);
			17942: out = 24'(-2112);
			17943: out = 24'(-2184);
			17944: out = 24'(-2152);
			17945: out = 24'(-2140);
			17946: out = 24'(-2156);
			17947: out = 24'(-2124);
			17948: out = 24'(-2136);
			17949: out = 24'(-2192);
			17950: out = 24'(-2112);
			17951: out = 24'(-2116);
			17952: out = 24'(-2124);
			17953: out = 24'(-2148);
			17954: out = 24'(-2120);
			17955: out = 24'(-2112);
			17956: out = 24'(-2112);
			17957: out = 24'(-2120);
			17958: out = 24'(-2112);
			17959: out = 24'(-2100);
			17960: out = 24'(-2076);
			17961: out = 24'(-2088);
			17962: out = 24'(-2144);
			17963: out = 24'(-2064);
			17964: out = 24'(-2072);
			17965: out = 24'(-2100);
			17966: out = 24'(-2124);
			17967: out = 24'(-2028);
			17968: out = 24'(-2108);
			17969: out = 24'(-2040);
			17970: out = 24'(-2096);
			17971: out = 24'(-2040);
			17972: out = 24'(-2064);
			17973: out = 24'(-2056);
			17974: out = 24'(-2040);
			17975: out = 24'(-2052);
			17976: out = 24'(-2028);
			17977: out = 24'(-2068);
			17978: out = 24'(-2024);
			17979: out = 24'(-2012);
			17980: out = 24'(-2060);
			17981: out = 24'(-2008);
			17982: out = 24'(-2044);
			17983: out = 24'(-1980);
			17984: out = 24'(-2076);
			17985: out = 24'(-1960);
			17986: out = 24'(-2016);
			17987: out = 24'(-1992);
			17988: out = 24'(-2004);
			17989: out = 24'(-1992);
			17990: out = 24'(-1952);
			17991: out = 24'(-1972);
			17992: out = 24'(-1984);
			17993: out = 24'(-1952);
			17994: out = 24'(-1916);
			17995: out = 24'(-1964);
			17996: out = 24'(-1948);
			17997: out = 24'(-1912);
			17998: out = 24'(-1968);
			17999: out = 24'(-1904);
			18000: out = 24'(-1944);
			18001: out = 24'(-1908);
			18002: out = 24'(-1920);
			18003: out = 24'(-1904);
			18004: out = 24'(-1880);
			18005: out = 24'(-1920);
			18006: out = 24'(-1876);
			18007: out = 24'(-1872);
			18008: out = 24'(-1868);
			18009: out = 24'(-1880);
			18010: out = 24'(-1820);
			18011: out = 24'(-1872);
			18012: out = 24'(-1840);
			18013: out = 24'(-1816);
			18014: out = 24'(-1832);
			18015: out = 24'(-1816);
			18016: out = 24'(-1816);
			18017: out = 24'(-1764);
			18018: out = 24'(-1776);
			18019: out = 24'(-1776);
			18020: out = 24'(-1732);
			18021: out = 24'(-1752);
			18022: out = 24'(-1752);
			18023: out = 24'(-1708);
			18024: out = 24'(-1728);
			18025: out = 24'(-1676);
			18026: out = 24'(-1728);
			18027: out = 24'(-1696);
			18028: out = 24'(-1652);
			18029: out = 24'(-1664);
			18030: out = 24'(-1620);
			18031: out = 24'(-1628);
			18032: out = 24'(-1588);
			18033: out = 24'(-1632);
			18034: out = 24'(-1596);
			18035: out = 24'(-1536);
			18036: out = 24'(-1596);
			18037: out = 24'(-1552);
			18038: out = 24'(-1492);
			18039: out = 24'(-1548);
			18040: out = 24'(-1476);
			18041: out = 24'(-1508);
			18042: out = 24'(-1460);
			18043: out = 24'(-1452);
			18044: out = 24'(-1476);
			18045: out = 24'(-1436);
			18046: out = 24'(-1412);
			18047: out = 24'(-1416);
			18048: out = 24'(-1400);
			18049: out = 24'(-1352);
			18050: out = 24'(-1388);
			18051: out = 24'(-1356);
			18052: out = 24'(-1328);
			18053: out = 24'(-1340);
			18054: out = 24'(-1344);
			18055: out = 24'(-1288);
			18056: out = 24'(-1316);
			18057: out = 24'(-1256);
			18058: out = 24'(-1252);
			18059: out = 24'(-1272);
			18060: out = 24'(-1192);
			18061: out = 24'(-1216);
			18062: out = 24'(-1216);
			18063: out = 24'(-1164);
			18064: out = 24'(-1188);
			18065: out = 24'(-1152);
			18066: out = 24'(-1128);
			18067: out = 24'(-1128);
			18068: out = 24'(-1100);
			18069: out = 24'(-1112);
			18070: out = 24'(-1072);
			18071: out = 24'(-1064);
			18072: out = 24'(-1076);
			18073: out = 24'(-1068);
			18074: out = 24'(-1028);
			18075: out = 24'(-996);
			18076: out = 24'(-988);
			18077: out = 24'(-1036);
			18078: out = 24'(-972);
			18079: out = 24'(-952);
			18080: out = 24'(-964);
			18081: out = 24'(-976);
			18082: out = 24'(-900);
			18083: out = 24'(-976);
			18084: out = 24'(-880);
			18085: out = 24'(-936);
			18086: out = 24'(-864);
			18087: out = 24'(-912);
			18088: out = 24'(-856);
			18089: out = 24'(-868);
			18090: out = 24'(-864);
			18091: out = 24'(-828);
			18092: out = 24'(-868);
			18093: out = 24'(-816);
			18094: out = 24'(-788);
			18095: out = 24'(-828);
			18096: out = 24'(-780);
			18097: out = 24'(-796);
			18098: out = 24'(-740);
			18099: out = 24'(-808);
			18100: out = 24'(-732);
			18101: out = 24'(-744);
			18102: out = 24'(-764);
			18103: out = 24'(-712);
			18104: out = 24'(-732);
			18105: out = 24'(-696);
			18106: out = 24'(-684);
			18107: out = 24'(-716);
			18108: out = 24'(-648);
			18109: out = 24'(-684);
			18110: out = 24'(-652);
			18111: out = 24'(-672);
			18112: out = 24'(-600);
			18113: out = 24'(-680);
			18114: out = 24'(-608);
			18115: out = 24'(-628);
			18116: out = 24'(-600);
			18117: out = 24'(-588);
			18118: out = 24'(-624);
			18119: out = 24'(-580);
			18120: out = 24'(-572);
			18121: out = 24'(-572);
			18122: out = 24'(-560);
			18123: out = 24'(-552);
			18124: out = 24'(-548);
			18125: out = 24'(-540);
			18126: out = 24'(-540);
			18127: out = 24'(-540);
			18128: out = 24'(-536);
			18129: out = 24'(-524);
			18130: out = 24'(-512);
			18131: out = 24'(-480);
			18132: out = 24'(-480);
			18133: out = 24'(-504);
			18134: out = 24'(-460);
			18135: out = 24'(-432);
			18136: out = 24'(-480);
			18137: out = 24'(-408);
			18138: out = 24'(-420);
			18139: out = 24'(-384);
			18140: out = 24'(-380);
			18141: out = 24'(-412);
			18142: out = 24'(-384);
			18143: out = 24'(-316);
			18144: out = 24'(-392);
			18145: out = 24'(-304);
			18146: out = 24'(-340);
			18147: out = 24'(-288);
			18148: out = 24'(-300);
			18149: out = 24'(-324);
			18150: out = 24'(-268);
			18151: out = 24'(-268);
			18152: out = 24'(-292);
			18153: out = 24'(-224);
			18154: out = 24'(-260);
			18155: out = 24'(-256);
			18156: out = 24'(-208);
			18157: out = 24'(-248);
			18158: out = 24'(-176);
			18159: out = 24'(-268);
			18160: out = 24'(-176);
			18161: out = 24'(-196);
			18162: out = 24'(-196);
			18163: out = 24'(-196);
			18164: out = 24'(-144);
			18165: out = 24'(-180);
			18166: out = 24'(-168);
			18167: out = 24'(-120);
			18168: out = 24'(-144);
			18169: out = 24'(-144);
			18170: out = 24'(-120);
			18171: out = 24'(-116);
			18172: out = 24'(-96);
			18173: out = 24'(-112);
			18174: out = 24'(-72);
			18175: out = 24'(-64);
			18176: out = 24'(-100);
			18177: out = 24'(-72);
			18178: out = 24'(-68);
			18179: out = 24'(-40);
			18180: out = 24'(-60);
			18181: out = 24'(-48);
			18182: out = 24'(-32);
			18183: out = 24'(-16);
			18184: out = 24'(-4);
			18185: out = 24'(-24);
			18186: out = 24'(4);
			18187: out = 24'(-16);
			18188: out = 24'(8);
			18189: out = 24'(24);
			18190: out = 24'(36);
			18191: out = 24'(36);
			18192: out = 24'(16);
			18193: out = 24'(68);
			18194: out = 24'(20);
			18195: out = 24'(68);
			18196: out = 24'(84);
			18197: out = 24'(8);
			18198: out = 24'(120);
			18199: out = 24'(100);
			18200: out = 24'(76);
			18201: out = 24'(120);
			18202: out = 24'(88);
			18203: out = 24'(148);
			18204: out = 24'(128);
			18205: out = 24'(76);
			18206: out = 24'(164);
			18207: out = 24'(136);
			18208: out = 24'(144);
			18209: out = 24'(180);
			18210: out = 24'(148);
			18211: out = 24'(196);
			18212: out = 24'(168);
			18213: out = 24'(192);
			18214: out = 24'(176);
			18215: out = 24'(224);
			18216: out = 24'(172);
			18217: out = 24'(212);
			18218: out = 24'(204);
			18219: out = 24'(260);
			18220: out = 24'(204);
			18221: out = 24'(264);
			18222: out = 24'(252);
			18223: out = 24'(272);
			18224: out = 24'(248);
			18225: out = 24'(288);
			18226: out = 24'(296);
			18227: out = 24'(288);
			18228: out = 24'(316);
			18229: out = 24'(320);
			18230: out = 24'(296);
			18231: out = 24'(360);
			18232: out = 24'(344);
			18233: out = 24'(324);
			18234: out = 24'(396);
			18235: out = 24'(336);
			18236: out = 24'(444);
			18237: out = 24'(364);
			18238: out = 24'(412);
			18239: out = 24'(408);
			18240: out = 24'(464);
			18241: out = 24'(436);
			18242: out = 24'(460);
			18243: out = 24'(476);
			18244: out = 24'(512);
			18245: out = 24'(504);
			18246: out = 24'(460);
			18247: out = 24'(544);
			18248: out = 24'(544);
			18249: out = 24'(516);
			18250: out = 24'(556);
			18251: out = 24'(576);
			18252: out = 24'(572);
			18253: out = 24'(580);
			18254: out = 24'(640);
			18255: out = 24'(600);
			18256: out = 24'(620);
			18257: out = 24'(668);
			18258: out = 24'(672);
			18259: out = 24'(672);
			18260: out = 24'(696);
			18261: out = 24'(640);
			18262: out = 24'(700);
			18263: out = 24'(744);
			18264: out = 24'(716);
			18265: out = 24'(748);
			18266: out = 24'(772);
			18267: out = 24'(764);
			18268: out = 24'(812);
			18269: out = 24'(772);
			18270: out = 24'(824);
			18271: out = 24'(828);
			18272: out = 24'(844);
			18273: out = 24'(824);
			18274: out = 24'(856);
			18275: out = 24'(836);
			18276: out = 24'(872);
			18277: out = 24'(888);
			18278: out = 24'(856);
			18279: out = 24'(892);
			18280: out = 24'(928);
			18281: out = 24'(920);
			18282: out = 24'(924);
			18283: out = 24'(952);
			18284: out = 24'(964);
			18285: out = 24'(964);
			18286: out = 24'(984);
			18287: out = 24'(972);
			18288: out = 24'(1012);
			18289: out = 24'(1004);
			18290: out = 24'(1024);
			18291: out = 24'(1004);
			18292: out = 24'(1048);
			18293: out = 24'(1060);
			18294: out = 24'(1080);
			18295: out = 24'(1048);
			18296: out = 24'(1108);
			18297: out = 24'(1096);
			18298: out = 24'(1068);
			18299: out = 24'(1112);
			18300: out = 24'(1132);
			18301: out = 24'(1060);
			18302: out = 24'(1128);
			18303: out = 24'(1132);
			18304: out = 24'(1132);
			18305: out = 24'(1128);
			18306: out = 24'(1152);
			18307: out = 24'(1172);
			18308: out = 24'(1176);
			18309: out = 24'(1164);
			18310: out = 24'(1192);
			18311: out = 24'(1176);
			18312: out = 24'(1164);
			18313: out = 24'(1248);
			18314: out = 24'(1212);
			18315: out = 24'(1208);
			18316: out = 24'(1224);
			18317: out = 24'(1252);
			18318: out = 24'(1236);
			18319: out = 24'(1260);
			18320: out = 24'(1248);
			18321: out = 24'(1224);
			18322: out = 24'(1272);
			18323: out = 24'(1288);
			18324: out = 24'(1288);
			18325: out = 24'(1256);
			18326: out = 24'(1344);
			18327: out = 24'(1280);
			18328: out = 24'(1288);
			18329: out = 24'(1308);
			18330: out = 24'(1340);
			18331: out = 24'(1320);
			18332: out = 24'(1308);
			18333: out = 24'(1320);
			18334: out = 24'(1368);
			18335: out = 24'(1336);
			18336: out = 24'(1360);
			18337: out = 24'(1340);
			18338: out = 24'(1376);
			18339: out = 24'(1384);
			18340: out = 24'(1352);
			18341: out = 24'(1388);
			18342: out = 24'(1428);
			18343: out = 24'(1356);
			18344: out = 24'(1388);
			18345: out = 24'(1428);
			18346: out = 24'(1384);
			18347: out = 24'(1424);
			18348: out = 24'(1392);
			18349: out = 24'(1440);
			18350: out = 24'(1408);
			18351: out = 24'(1396);
			18352: out = 24'(1444);
			18353: out = 24'(1456);
			18354: out = 24'(1448);
			18355: out = 24'(1408);
			18356: out = 24'(1468);
			18357: out = 24'(1468);
			18358: out = 24'(1476);
			18359: out = 24'(1456);
			18360: out = 24'(1476);
			18361: out = 24'(1484);
			18362: out = 24'(1468);
			18363: out = 24'(1492);
			18364: out = 24'(1520);
			18365: out = 24'(1444);
			18366: out = 24'(1496);
			18367: out = 24'(1488);
			18368: out = 24'(1520);
			18369: out = 24'(1472);
			18370: out = 24'(1496);
			18371: out = 24'(1504);
			18372: out = 24'(1456);
			18373: out = 24'(1476);
			18374: out = 24'(1492);
			18375: out = 24'(1500);
			18376: out = 24'(1468);
			18377: out = 24'(1468);
			18378: out = 24'(1468);
			18379: out = 24'(1500);
			18380: out = 24'(1452);
			18381: out = 24'(1444);
			18382: out = 24'(1472);
			18383: out = 24'(1468);
			18384: out = 24'(1496);
			18385: out = 24'(1452);
			18386: out = 24'(1444);
			18387: out = 24'(1504);
			18388: out = 24'(1488);
			18389: out = 24'(1452);
			18390: out = 24'(1468);
			18391: out = 24'(1452);
			18392: out = 24'(1496);
			18393: out = 24'(1428);
			18394: out = 24'(1452);
			18395: out = 24'(1456);
			18396: out = 24'(1492);
			18397: out = 24'(1436);
			18398: out = 24'(1404);
			18399: out = 24'(1504);
			18400: out = 24'(1392);
			18401: out = 24'(1476);
			18402: out = 24'(1444);
			18403: out = 24'(1432);
			18404: out = 24'(1432);
			18405: out = 24'(1492);
			18406: out = 24'(1440);
			18407: out = 24'(1448);
			18408: out = 24'(1436);
			18409: out = 24'(1456);
			18410: out = 24'(1424);
			18411: out = 24'(1428);
			18412: out = 24'(1456);
			18413: out = 24'(1412);
			18414: out = 24'(1460);
			18415: out = 24'(1440);
			18416: out = 24'(1452);
			18417: out = 24'(1416);
			18418: out = 24'(1468);
			18419: out = 24'(1432);
			18420: out = 24'(1408);
			18421: out = 24'(1440);
			18422: out = 24'(1404);
			18423: out = 24'(1416);
			18424: out = 24'(1444);
			18425: out = 24'(1404);
			18426: out = 24'(1428);
			18427: out = 24'(1400);
			18428: out = 24'(1444);
			18429: out = 24'(1416);
			18430: out = 24'(1424);
			18431: out = 24'(1428);
			18432: out = 24'(1404);
			18433: out = 24'(1428);
			18434: out = 24'(1424);
			18435: out = 24'(1376);
			18436: out = 24'(1428);
			18437: out = 24'(1356);
			18438: out = 24'(1380);
			18439: out = 24'(1404);
			18440: out = 24'(1368);
			18441: out = 24'(1392);
			18442: out = 24'(1384);
			18443: out = 24'(1368);
			18444: out = 24'(1364);
			18445: out = 24'(1376);
			18446: out = 24'(1340);
			18447: out = 24'(1316);
			18448: out = 24'(1320);
			18449: out = 24'(1380);
			18450: out = 24'(1272);
			18451: out = 24'(1316);
			18452: out = 24'(1332);
			18453: out = 24'(1284);
			18454: out = 24'(1316);
			18455: out = 24'(1300);
			18456: out = 24'(1268);
			18457: out = 24'(1280);
			18458: out = 24'(1268);
			18459: out = 24'(1296);
			18460: out = 24'(1244);
			18461: out = 24'(1216);
			18462: out = 24'(1260);
			18463: out = 24'(1236);
			18464: out = 24'(1232);
			18465: out = 24'(1208);
			18466: out = 24'(1236);
			18467: out = 24'(1216);
			18468: out = 24'(1224);
			18469: out = 24'(1164);
			18470: out = 24'(1208);
			18471: out = 24'(1168);
			18472: out = 24'(1124);
			18473: out = 24'(1160);
			18474: out = 24'(1148);
			18475: out = 24'(1060);
			18476: out = 24'(1152);
			18477: out = 24'(1084);
			18478: out = 24'(1104);
			18479: out = 24'(1052);
			18480: out = 24'(1076);
			18481: out = 24'(1068);
			18482: out = 24'(1032);
			18483: out = 24'(1060);
			18484: out = 24'(1024);
			18485: out = 24'(1028);
			18486: out = 24'(984);
			18487: out = 24'(1044);
			18488: out = 24'(940);
			18489: out = 24'(1020);
			18490: out = 24'(956);
			18491: out = 24'(972);
			18492: out = 24'(928);
			18493: out = 24'(948);
			18494: out = 24'(936);
			18495: out = 24'(920);
			18496: out = 24'(876);
			18497: out = 24'(900);
			18498: out = 24'(884);
			18499: out = 24'(880);
			18500: out = 24'(840);
			18501: out = 24'(856);
			18502: out = 24'(840);
			18503: out = 24'(860);
			18504: out = 24'(808);
			18505: out = 24'(828);
			18506: out = 24'(788);
			18507: out = 24'(808);
			18508: out = 24'(748);
			18509: out = 24'(780);
			18510: out = 24'(700);
			18511: out = 24'(796);
			18512: out = 24'(684);
			18513: out = 24'(748);
			18514: out = 24'(724);
			18515: out = 24'(688);
			18516: out = 24'(712);
			18517: out = 24'(688);
			18518: out = 24'(688);
			18519: out = 24'(672);
			18520: out = 24'(668);
			18521: out = 24'(644);
			18522: out = 24'(668);
			18523: out = 24'(640);
			18524: out = 24'(600);
			18525: out = 24'(584);
			18526: out = 24'(616);
			18527: out = 24'(592);
			18528: out = 24'(572);
			18529: out = 24'(564);
			18530: out = 24'(584);
			18531: out = 24'(556);
			18532: out = 24'(532);
			18533: out = 24'(560);
			18534: out = 24'(548);
			18535: out = 24'(504);
			18536: out = 24'(524);
			18537: out = 24'(508);
			18538: out = 24'(488);
			18539: out = 24'(496);
			18540: out = 24'(448);
			18541: out = 24'(488);
			18542: out = 24'(476);
			18543: out = 24'(456);
			18544: out = 24'(476);
			18545: out = 24'(440);
			18546: out = 24'(464);
			18547: out = 24'(408);
			18548: out = 24'(400);
			18549: out = 24'(432);
			18550: out = 24'(412);
			18551: out = 24'(392);
			18552: out = 24'(388);
			18553: out = 24'(412);
			18554: out = 24'(352);
			18555: out = 24'(400);
			18556: out = 24'(340);
			18557: out = 24'(360);
			18558: out = 24'(356);
			18559: out = 24'(348);
			18560: out = 24'(332);
			18561: out = 24'(292);
			18562: out = 24'(352);
			18563: out = 24'(296);
			18564: out = 24'(324);
			18565: out = 24'(268);
			18566: out = 24'(320);
			18567: out = 24'(272);
			18568: out = 24'(320);
			18569: out = 24'(252);
			18570: out = 24'(304);
			18571: out = 24'(268);
			18572: out = 24'(272);
			18573: out = 24'(248);
			18574: out = 24'(256);
			18575: out = 24'(228);
			18576: out = 24'(252);
			18577: out = 24'(200);
			18578: out = 24'(244);
			18579: out = 24'(200);
			18580: out = 24'(208);
			18581: out = 24'(208);
			18582: out = 24'(200);
			18583: out = 24'(192);
			18584: out = 24'(192);
			18585: out = 24'(184);
			18586: out = 24'(184);
			18587: out = 24'(176);
			18588: out = 24'(192);
			18589: out = 24'(148);
			18590: out = 24'(152);
			18591: out = 24'(172);
			18592: out = 24'(144);
			18593: out = 24'(136);
			18594: out = 24'(136);
			18595: out = 24'(144);
			18596: out = 24'(144);
			18597: out = 24'(128);
			18598: out = 24'(116);
			18599: out = 24'(112);
			18600: out = 24'(120);
			18601: out = 24'(80);
			18602: out = 24'(68);
			18603: out = 24'(56);
			18604: out = 24'(24);
			18605: out = 24'(56);
			18606: out = 24'(-4);
			18607: out = 24'(8);
			18608: out = 24'(8);
			18609: out = 24'(-16);
			18610: out = 24'(-40);
			18611: out = 24'(-36);
			18612: out = 24'(-20);
			18613: out = 24'(-116);
			18614: out = 24'(-40);
			18615: out = 24'(-76);
			18616: out = 24'(-64);
			18617: out = 24'(-124);
			18618: out = 24'(-96);
			18619: out = 24'(-124);
			18620: out = 24'(-96);
			18621: out = 24'(-156);
			18622: out = 24'(-108);
			18623: out = 24'(-152);
			18624: out = 24'(-168);
			18625: out = 24'(-172);
			18626: out = 24'(-196);
			18627: out = 24'(-180);
			18628: out = 24'(-216);
			18629: out = 24'(-216);
			18630: out = 24'(-216);
			18631: out = 24'(-220);
			18632: out = 24'(-220);
			18633: out = 24'(-244);
			18634: out = 24'(-240);
			18635: out = 24'(-256);
			18636: out = 24'(-268);
			18637: out = 24'(-272);
			18638: out = 24'(-276);
			18639: out = 24'(-296);
			18640: out = 24'(-332);
			18641: out = 24'(-304);
			18642: out = 24'(-296);
			18643: out = 24'(-336);
			18644: out = 24'(-332);
			18645: out = 24'(-348);
			18646: out = 24'(-320);
			18647: out = 24'(-340);
			18648: out = 24'(-344);
			18649: out = 24'(-380);
			18650: out = 24'(-356);
			18651: out = 24'(-352);
			18652: out = 24'(-436);
			18653: out = 24'(-408);
			18654: out = 24'(-364);
			18655: out = 24'(-428);
			18656: out = 24'(-436);
			18657: out = 24'(-400);
			18658: out = 24'(-416);
			18659: out = 24'(-436);
			18660: out = 24'(-464);
			18661: out = 24'(-412);
			18662: out = 24'(-488);
			18663: out = 24'(-480);
			18664: out = 24'(-440);
			18665: out = 24'(-528);
			18666: out = 24'(-464);
			18667: out = 24'(-496);
			18668: out = 24'(-512);
			18669: out = 24'(-496);
			18670: out = 24'(-516);
			18671: out = 24'(-528);
			18672: out = 24'(-536);
			18673: out = 24'(-528);
			18674: out = 24'(-536);
			18675: out = 24'(-540);
			18676: out = 24'(-604);
			18677: out = 24'(-532);
			18678: out = 24'(-564);
			18679: out = 24'(-632);
			18680: out = 24'(-576);
			18681: out = 24'(-592);
			18682: out = 24'(-600);
			18683: out = 24'(-608);
			18684: out = 24'(-636);
			18685: out = 24'(-592);
			18686: out = 24'(-652);
			18687: out = 24'(-628);
			18688: out = 24'(-664);
			18689: out = 24'(-672);
			18690: out = 24'(-656);
			18691: out = 24'(-684);
			18692: out = 24'(-664);
			18693: out = 24'(-696);
			18694: out = 24'(-704);
			18695: out = 24'(-688);
			18696: out = 24'(-732);
			18697: out = 24'(-728);
			18698: out = 24'(-716);
			18699: out = 24'(-744);
			18700: out = 24'(-768);
			18701: out = 24'(-760);
			18702: out = 24'(-760);
			18703: out = 24'(-788);
			18704: out = 24'(-784);
			18705: out = 24'(-832);
			18706: out = 24'(-816);
			18707: out = 24'(-868);
			18708: out = 24'(-812);
			18709: out = 24'(-884);
			18710: out = 24'(-812);
			18711: out = 24'(-920);
			18712: out = 24'(-868);
			18713: out = 24'(-900);
			18714: out = 24'(-916);
			18715: out = 24'(-928);
			18716: out = 24'(-936);
			18717: out = 24'(-968);
			18718: out = 24'(-948);
			18719: out = 24'(-968);
			18720: out = 24'(-996);
			18721: out = 24'(-984);
			18722: out = 24'(-1016);
			18723: out = 24'(-1024);
			18724: out = 24'(-1024);
			18725: out = 24'(-1064);
			18726: out = 24'(-1032);
			18727: out = 24'(-1112);
			18728: out = 24'(-1092);
			18729: out = 24'(-1092);
			18730: out = 24'(-1152);
			18731: out = 24'(-1160);
			18732: out = 24'(-1156);
			18733: out = 24'(-1144);
			18734: out = 24'(-1172);
			18735: out = 24'(-1200);
			18736: out = 24'(-1196);
			18737: out = 24'(-1204);
			18738: out = 24'(-1224);
			18739: out = 24'(-1232);
			18740: out = 24'(-1252);
			18741: out = 24'(-1284);
			18742: out = 24'(-1240);
			18743: out = 24'(-1308);
			18744: out = 24'(-1344);
			18745: out = 24'(-1292);
			18746: out = 24'(-1332);
			18747: out = 24'(-1336);
			18748: out = 24'(-1368);
			18749: out = 24'(-1356);
			18750: out = 24'(-1392);
			18751: out = 24'(-1360);
			18752: out = 24'(-1440);
			18753: out = 24'(-1392);
			18754: out = 24'(-1432);
			18755: out = 24'(-1448);
			18756: out = 24'(-1436);
			18757: out = 24'(-1444);
			18758: out = 24'(-1468);
			18759: out = 24'(-1480);
			18760: out = 24'(-1468);
			18761: out = 24'(-1496);
			18762: out = 24'(-1492);
			18763: out = 24'(-1496);
			18764: out = 24'(-1520);
			18765: out = 24'(-1536);
			18766: out = 24'(-1508);
			18767: out = 24'(-1524);
			18768: out = 24'(-1544);
			18769: out = 24'(-1544);
			18770: out = 24'(-1552);
			18771: out = 24'(-1568);
			18772: out = 24'(-1584);
			18773: out = 24'(-1528);
			18774: out = 24'(-1636);
			18775: out = 24'(-1544);
			18776: out = 24'(-1628);
			18777: out = 24'(-1540);
			18778: out = 24'(-1604);
			18779: out = 24'(-1632);
			18780: out = 24'(-1576);
			18781: out = 24'(-1616);
			18782: out = 24'(-1640);
			18783: out = 24'(-1624);
			18784: out = 24'(-1612);
			18785: out = 24'(-1632);
			18786: out = 24'(-1632);
			18787: out = 24'(-1668);
			18788: out = 24'(-1628);
			18789: out = 24'(-1652);
			18790: out = 24'(-1664);
			18791: out = 24'(-1632);
			18792: out = 24'(-1688);
			18793: out = 24'(-1680);
			18794: out = 24'(-1672);
			18795: out = 24'(-1676);
			18796: out = 24'(-1668);
			18797: out = 24'(-1700);
			18798: out = 24'(-1676);
			18799: out = 24'(-1688);
			18800: out = 24'(-1660);
			18801: out = 24'(-1712);
			18802: out = 24'(-1716);
			18803: out = 24'(-1676);
			18804: out = 24'(-1708);
			18805: out = 24'(-1684);
			18806: out = 24'(-1728);
			18807: out = 24'(-1680);
			18808: out = 24'(-1700);
			18809: out = 24'(-1680);
			18810: out = 24'(-1708);
			18811: out = 24'(-1672);
			18812: out = 24'(-1692);
			18813: out = 24'(-1680);
			18814: out = 24'(-1688);
			18815: out = 24'(-1716);
			18816: out = 24'(-1644);
			18817: out = 24'(-1720);
			18818: out = 24'(-1720);
			18819: out = 24'(-1692);
			18820: out = 24'(-1680);
			18821: out = 24'(-1692);
			18822: out = 24'(-1756);
			18823: out = 24'(-1668);
			18824: out = 24'(-1712);
			18825: out = 24'(-1688);
			18826: out = 24'(-1720);
			18827: out = 24'(-1672);
			18828: out = 24'(-1708);
			18829: out = 24'(-1676);
			18830: out = 24'(-1696);
			18831: out = 24'(-1688);
			18832: out = 24'(-1676);
			18833: out = 24'(-1668);
			18834: out = 24'(-1744);
			18835: out = 24'(-1672);
			18836: out = 24'(-1664);
			18837: out = 24'(-1700);
			18838: out = 24'(-1680);
			18839: out = 24'(-1692);
			18840: out = 24'(-1684);
			18841: out = 24'(-1676);
			18842: out = 24'(-1676);
			18843: out = 24'(-1652);
			18844: out = 24'(-1688);
			18845: out = 24'(-1652);
			18846: out = 24'(-1652);
			18847: out = 24'(-1700);
			18848: out = 24'(-1660);
			18849: out = 24'(-1680);
			18850: out = 24'(-1616);
			18851: out = 24'(-1672);
			18852: out = 24'(-1676);
			18853: out = 24'(-1628);
			18854: out = 24'(-1620);
			18855: out = 24'(-1668);
			18856: out = 24'(-1632);
			18857: out = 24'(-1620);
			18858: out = 24'(-1644);
			18859: out = 24'(-1600);
			18860: out = 24'(-1644);
			18861: out = 24'(-1624);
			18862: out = 24'(-1600);
			18863: out = 24'(-1616);
			18864: out = 24'(-1628);
			18865: out = 24'(-1628);
			18866: out = 24'(-1568);
			18867: out = 24'(-1644);
			18868: out = 24'(-1588);
			18869: out = 24'(-1600);
			18870: out = 24'(-1588);
			18871: out = 24'(-1592);
			18872: out = 24'(-1600);
			18873: out = 24'(-1572);
			18874: out = 24'(-1580);
			18875: out = 24'(-1564);
			18876: out = 24'(-1596);
			18877: out = 24'(-1604);
			18878: out = 24'(-1524);
			18879: out = 24'(-1604);
			18880: out = 24'(-1528);
			18881: out = 24'(-1572);
			18882: out = 24'(-1572);
			18883: out = 24'(-1520);
			18884: out = 24'(-1552);
			18885: out = 24'(-1516);
			18886: out = 24'(-1536);
			18887: out = 24'(-1504);
			18888: out = 24'(-1524);
			18889: out = 24'(-1492);
			18890: out = 24'(-1524);
			18891: out = 24'(-1520);
			18892: out = 24'(-1508);
			18893: out = 24'(-1484);
			18894: out = 24'(-1528);
			18895: out = 24'(-1484);
			18896: out = 24'(-1508);
			18897: out = 24'(-1476);
			18898: out = 24'(-1444);
			18899: out = 24'(-1480);
			18900: out = 24'(-1460);
			18901: out = 24'(-1456);
			18902: out = 24'(-1416);
			18903: out = 24'(-1448);
			18904: out = 24'(-1452);
			18905: out = 24'(-1440);
			18906: out = 24'(-1412);
			18907: out = 24'(-1412);
			18908: out = 24'(-1424);
			18909: out = 24'(-1404);
			18910: out = 24'(-1364);
			18911: out = 24'(-1352);
			18912: out = 24'(-1424);
			18913: out = 24'(-1348);
			18914: out = 24'(-1340);
			18915: out = 24'(-1380);
			18916: out = 24'(-1328);
			18917: out = 24'(-1308);
			18918: out = 24'(-1364);
			18919: out = 24'(-1320);
			18920: out = 24'(-1288);
			18921: out = 24'(-1280);
			18922: out = 24'(-1320);
			18923: out = 24'(-1264);
			18924: out = 24'(-1264);
			18925: out = 24'(-1272);
			18926: out = 24'(-1200);
			18927: out = 24'(-1296);
			18928: out = 24'(-1216);
			18929: out = 24'(-1208);
			18930: out = 24'(-1208);
			18931: out = 24'(-1184);
			18932: out = 24'(-1172);
			18933: out = 24'(-1172);
			18934: out = 24'(-1156);
			18935: out = 24'(-1172);
			18936: out = 24'(-1112);
			18937: out = 24'(-1108);
			18938: out = 24'(-1164);
			18939: out = 24'(-1084);
			18940: out = 24'(-1100);
			18941: out = 24'(-1060);
			18942: out = 24'(-1092);
			18943: out = 24'(-1076);
			18944: out = 24'(-1024);
			18945: out = 24'(-1060);
			18946: out = 24'(-1048);
			18947: out = 24'(-1008);
			18948: out = 24'(-1008);
			18949: out = 24'(-1032);
			18950: out = 24'(-964);
			18951: out = 24'(-996);
			18952: out = 24'(-1000);
			18953: out = 24'(-952);
			18954: out = 24'(-940);
			18955: out = 24'(-976);
			18956: out = 24'(-928);
			18957: out = 24'(-900);
			18958: out = 24'(-940);
			18959: out = 24'(-880);
			18960: out = 24'(-876);
			18961: out = 24'(-872);
			18962: out = 24'(-908);
			18963: out = 24'(-832);
			18964: out = 24'(-840);
			18965: out = 24'(-832);
			18966: out = 24'(-800);
			18967: out = 24'(-864);
			18968: out = 24'(-800);
			18969: out = 24'(-812);
			18970: out = 24'(-776);
			18971: out = 24'(-784);
			18972: out = 24'(-820);
			18973: out = 24'(-724);
			18974: out = 24'(-752);
			18975: out = 24'(-720);
			18976: out = 24'(-764);
			18977: out = 24'(-712);
			18978: out = 24'(-696);
			18979: out = 24'(-700);
			18980: out = 24'(-704);
			18981: out = 24'(-684);
			18982: out = 24'(-672);
			18983: out = 24'(-652);
			18984: out = 24'(-716);
			18985: out = 24'(-636);
			18986: out = 24'(-644);
			18987: out = 24'(-644);
			18988: out = 24'(-688);
			18989: out = 24'(-572);
			18990: out = 24'(-684);
			18991: out = 24'(-584);
			18992: out = 24'(-636);
			18993: out = 24'(-592);
			18994: out = 24'(-600);
			18995: out = 24'(-616);
			18996: out = 24'(-576);
			18997: out = 24'(-616);
			18998: out = 24'(-528);
			18999: out = 24'(-592);
			19000: out = 24'(-564);
			19001: out = 24'(-544);
			19002: out = 24'(-540);
			19003: out = 24'(-544);
			19004: out = 24'(-528);
			19005: out = 24'(-524);
			19006: out = 24'(-508);
			19007: out = 24'(-512);
			19008: out = 24'(-476);
			19009: out = 24'(-488);
			19010: out = 24'(-508);
			19011: out = 24'(-484);
			19012: out = 24'(-440);
			19013: out = 24'(-504);
			19014: out = 24'(-460);
			19015: out = 24'(-460);
			19016: out = 24'(-480);
			19017: out = 24'(-436);
			19018: out = 24'(-448);
			19019: out = 24'(-428);
			19020: out = 24'(-452);
			19021: out = 24'(-396);
			19022: out = 24'(-432);
			19023: out = 24'(-388);
			19024: out = 24'(-408);
			19025: out = 24'(-364);
			19026: out = 24'(-408);
			19027: out = 24'(-340);
			19028: out = 24'(-352);
			19029: out = 24'(-348);
			19030: out = 24'(-352);
			19031: out = 24'(-300);
			19032: out = 24'(-360);
			19033: out = 24'(-324);
			19034: out = 24'(-296);
			19035: out = 24'(-340);
			19036: out = 24'(-264);
			19037: out = 24'(-304);
			19038: out = 24'(-296);
			19039: out = 24'(-268);
			19040: out = 24'(-252);
			19041: out = 24'(-248);
			19042: out = 24'(-272);
			19043: out = 24'(-224);
			19044: out = 24'(-204);
			19045: out = 24'(-252);
			19046: out = 24'(-232);
			19047: out = 24'(-192);
			19048: out = 24'(-204);
			19049: out = 24'(-200);
			19050: out = 24'(-160);
			19051: out = 24'(-220);
			19052: out = 24'(-156);
			19053: out = 24'(-184);
			19054: out = 24'(-148);
			19055: out = 24'(-156);
			19056: out = 24'(-184);
			19057: out = 24'(-132);
			19058: out = 24'(-120);
			19059: out = 24'(-152);
			19060: out = 24'(-100);
			19061: out = 24'(-132);
			19062: out = 24'(-76);
			19063: out = 24'(-96);
			19064: out = 24'(-108);
			19065: out = 24'(-88);
			19066: out = 24'(-100);
			19067: out = 24'(-104);
			19068: out = 24'(-72);
			19069: out = 24'(-68);
			19070: out = 24'(-108);
			19071: out = 24'(-24);
			19072: out = 24'(-76);
			19073: out = 24'(-48);
			19074: out = 24'(-64);
			19075: out = 24'(-64);
			19076: out = 24'(-32);
			19077: out = 24'(-56);
			19078: out = 24'(-32);
			19079: out = 24'(-40);
			19080: out = 24'(4);
			19081: out = 24'(-28);
			19082: out = 24'(-4);
			19083: out = 24'(12);
			19084: out = 24'(-8);
			19085: out = 24'(0);
			19086: out = 24'(4);
			19087: out = 24'(28);
			19088: out = 24'(8);
			19089: out = 24'(28);
			19090: out = 24'(36);
			19091: out = 24'(48);
			19092: out = 24'(64);
			19093: out = 24'(12);
			19094: out = 24'(60);
			19095: out = 24'(68);
			19096: out = 24'(88);
			19097: out = 24'(52);
			19098: out = 24'(88);
			19099: out = 24'(56);
			19100: out = 24'(132);
			19101: out = 24'(64);
			19102: out = 24'(104);
			19103: out = 24'(104);
			19104: out = 24'(108);
			19105: out = 24'(96);
			19106: out = 24'(108);
			19107: out = 24'(156);
			19108: out = 24'(84);
			19109: out = 24'(156);
			19110: out = 24'(144);
			19111: out = 24'(112);
			19112: out = 24'(176);
			19113: out = 24'(136);
			19114: out = 24'(152);
			19115: out = 24'(184);
			19116: out = 24'(152);
			19117: out = 24'(196);
			19118: out = 24'(184);
			19119: out = 24'(204);
			19120: out = 24'(208);
			19121: out = 24'(184);
			19122: out = 24'(232);
			19123: out = 24'(276);
			19124: out = 24'(196);
			19125: out = 24'(264);
			19126: out = 24'(272);
			19127: out = 24'(260);
			19128: out = 24'(288);
			19129: out = 24'(272);
			19130: out = 24'(304);
			19131: out = 24'(288);
			19132: out = 24'(316);
			19133: out = 24'(300);
			19134: out = 24'(340);
			19135: out = 24'(356);
			19136: out = 24'(320);
			19137: out = 24'(392);
			19138: out = 24'(364);
			19139: out = 24'(400);
			19140: out = 24'(384);
			19141: out = 24'(364);
			19142: out = 24'(448);
			19143: out = 24'(388);
			19144: out = 24'(420);
			19145: out = 24'(412);
			19146: out = 24'(476);
			19147: out = 24'(460);
			19148: out = 24'(448);
			19149: out = 24'(484);
			19150: out = 24'(508);
			19151: out = 24'(492);
			19152: out = 24'(496);
			19153: out = 24'(512);
			19154: out = 24'(528);
			19155: out = 24'(544);
			19156: out = 24'(508);
			19157: out = 24'(548);
			19158: out = 24'(552);
			19159: out = 24'(584);
			19160: out = 24'(540);
			19161: out = 24'(624);
			19162: out = 24'(580);
			19163: out = 24'(580);
			19164: out = 24'(616);
			19165: out = 24'(652);
			19166: out = 24'(640);
			19167: out = 24'(616);
			19168: out = 24'(652);
			19169: out = 24'(664);
			19170: out = 24'(696);
			19171: out = 24'(664);
			19172: out = 24'(680);
			19173: out = 24'(672);
			19174: out = 24'(740);
			19175: out = 24'(704);
			19176: out = 24'(688);
			19177: out = 24'(744);
			19178: out = 24'(724);
			19179: out = 24'(736);
			19180: out = 24'(744);
			19181: out = 24'(740);
			19182: out = 24'(752);
			19183: out = 24'(796);
			19184: out = 24'(760);
			19185: out = 24'(800);
			19186: out = 24'(772);
			19187: out = 24'(788);
			19188: out = 24'(800);
			19189: out = 24'(812);
			19190: out = 24'(800);
			19191: out = 24'(820);
			19192: out = 24'(812);
			19193: out = 24'(824);
			19194: out = 24'(860);
			19195: out = 24'(876);
			19196: out = 24'(832);
			19197: out = 24'(840);
			19198: out = 24'(888);
			19199: out = 24'(868);
			19200: out = 24'(880);
			19201: out = 24'(876);
			19202: out = 24'(888);
			19203: out = 24'(900);
			19204: out = 24'(908);
			19205: out = 24'(904);
			19206: out = 24'(916);
			19207: out = 24'(956);
			19208: out = 24'(864);
			19209: out = 24'(920);
			19210: out = 24'(968);
			19211: out = 24'(920);
			19212: out = 24'(960);
			19213: out = 24'(936);
			19214: out = 24'(932);
			19215: out = 24'(972);
			19216: out = 24'(988);
			19217: out = 24'(936);
			19218: out = 24'(1004);
			19219: out = 24'(956);
			19220: out = 24'(1020);
			19221: out = 24'(980);
			19222: out = 24'(972);
			19223: out = 24'(980);
			19224: out = 24'(1024);
			19225: out = 24'(1020);
			19226: out = 24'(976);
			19227: out = 24'(1020);
			19228: out = 24'(1020);
			19229: out = 24'(1052);
			19230: out = 24'(976);
			19231: out = 24'(1044);
			19232: out = 24'(1008);
			19233: out = 24'(1032);
			19234: out = 24'(1060);
			19235: out = 24'(1008);
			19236: out = 24'(1076);
			19237: out = 24'(1032);
			19238: out = 24'(1056);
			19239: out = 24'(1048);
			19240: out = 24'(1052);
			19241: out = 24'(1096);
			19242: out = 24'(1028);
			19243: out = 24'(1072);
			19244: out = 24'(1092);
			19245: out = 24'(1068);
			19246: out = 24'(1104);
			19247: out = 24'(1060);
			19248: out = 24'(1092);
			19249: out = 24'(1100);
			19250: out = 24'(1108);
			19251: out = 24'(1080);
			19252: out = 24'(1080);
			19253: out = 24'(1124);
			19254: out = 24'(1072);
			19255: out = 24'(1100);
			19256: out = 24'(1100);
			19257: out = 24'(1072);
			19258: out = 24'(1148);
			19259: out = 24'(1048);
			19260: out = 24'(1128);
			19261: out = 24'(1080);
			19262: out = 24'(1104);
			19263: out = 24'(1076);
			19264: out = 24'(1112);
			19265: out = 24'(1092);
			19266: out = 24'(1140);
			19267: out = 24'(1084);
			19268: out = 24'(1100);
			19269: out = 24'(1084);
			19270: out = 24'(1072);
			19271: out = 24'(1128);
			19272: out = 24'(1020);
			19273: out = 24'(1064);
			19274: out = 24'(1084);
			19275: out = 24'(1084);
			19276: out = 24'(1068);
			19277: out = 24'(1036);
			19278: out = 24'(1104);
			19279: out = 24'(1064);
			19280: out = 24'(1068);
			19281: out = 24'(1092);
			19282: out = 24'(1048);
			19283: out = 24'(1076);
			19284: out = 24'(1096);
			19285: out = 24'(1060);
			19286: out = 24'(1092);
			19287: out = 24'(1064);
			19288: out = 24'(1048);
			19289: out = 24'(1064);
			19290: out = 24'(1084);
			19291: out = 24'(1028);
			19292: out = 24'(1044);
			19293: out = 24'(1068);
			19294: out = 24'(1052);
			19295: out = 24'(1084);
			19296: out = 24'(1016);
			19297: out = 24'(1100);
			19298: out = 24'(1032);
			19299: out = 24'(1064);
			19300: out = 24'(1068);
			19301: out = 24'(1036);
			19302: out = 24'(1068);
			19303: out = 24'(1076);
			19304: out = 24'(1024);
			19305: out = 24'(1096);
			19306: out = 24'(1032);
			19307: out = 24'(1056);
			19308: out = 24'(1072);
			19309: out = 24'(1020);
			19310: out = 24'(1056);
			19311: out = 24'(1068);
			19312: out = 24'(1012);
			19313: out = 24'(1076);
			19314: out = 24'(1016);
			19315: out = 24'(1036);
			19316: out = 24'(1044);
			19317: out = 24'(1016);
			19318: out = 24'(1020);
			19319: out = 24'(1044);
			19320: out = 24'(1004);
			19321: out = 24'(1016);
			19322: out = 24'(1032);
			19323: out = 24'(984);
			19324: out = 24'(1060);
			19325: out = 24'(956);
			19326: out = 24'(1020);
			19327: out = 24'(1008);
			19328: out = 24'(1000);
			19329: out = 24'(996);
			19330: out = 24'(1020);
			19331: out = 24'(996);
			19332: out = 24'(984);
			19333: out = 24'(1020);
			19334: out = 24'(960);
			19335: out = 24'(968);
			19336: out = 24'(1008);
			19337: out = 24'(956);
			19338: out = 24'(968);
			19339: out = 24'(980);
			19340: out = 24'(948);
			19341: out = 24'(980);
			19342: out = 24'(956);
			19343: out = 24'(932);
			19344: out = 24'(960);
			19345: out = 24'(956);
			19346: out = 24'(940);
			19347: out = 24'(936);
			19348: out = 24'(952);
			19349: out = 24'(900);
			19350: out = 24'(964);
			19351: out = 24'(864);
			19352: out = 24'(888);
			19353: out = 24'(912);
			19354: out = 24'(892);
			19355: out = 24'(872);
			19356: out = 24'(892);
			19357: out = 24'(856);
			19358: out = 24'(872);
			19359: out = 24'(872);
			19360: out = 24'(812);
			19361: out = 24'(836);
			19362: out = 24'(800);
			19363: out = 24'(848);
			19364: out = 24'(776);
			19365: out = 24'(848);
			19366: out = 24'(788);
			19367: out = 24'(760);
			19368: out = 24'(828);
			19369: out = 24'(760);
			19370: out = 24'(780);
			19371: out = 24'(760);
			19372: out = 24'(732);
			19373: out = 24'(800);
			19374: out = 24'(728);
			19375: out = 24'(724);
			19376: out = 24'(736);
			19377: out = 24'(732);
			19378: out = 24'(676);
			19379: out = 24'(724);
			19380: out = 24'(700);
			19381: out = 24'(680);
			19382: out = 24'(672);
			19383: out = 24'(668);
			19384: out = 24'(644);
			19385: out = 24'(664);
			19386: out = 24'(632);
			19387: out = 24'(632);
			19388: out = 24'(628);
			19389: out = 24'(628);
			19390: out = 24'(632);
			19391: out = 24'(572);
			19392: out = 24'(632);
			19393: out = 24'(576);
			19394: out = 24'(572);
			19395: out = 24'(576);
			19396: out = 24'(544);
			19397: out = 24'(588);
			19398: out = 24'(544);
			19399: out = 24'(516);
			19400: out = 24'(556);
			19401: out = 24'(528);
			19402: out = 24'(492);
			19403: out = 24'(504);
			19404: out = 24'(512);
			19405: out = 24'(456);
			19406: out = 24'(508);
			19407: out = 24'(476);
			19408: out = 24'(464);
			19409: out = 24'(476);
			19410: out = 24'(460);
			19411: out = 24'(404);
			19412: out = 24'(460);
			19413: out = 24'(416);
			19414: out = 24'(412);
			19415: out = 24'(416);
			19416: out = 24'(428);
			19417: out = 24'(364);
			19418: out = 24'(412);
			19419: out = 24'(396);
			19420: out = 24'(356);
			19421: out = 24'(400);
			19422: out = 24'(352);
			19423: out = 24'(384);
			19424: out = 24'(344);
			19425: out = 24'(380);
			19426: out = 24'(356);
			19427: out = 24'(356);
			19428: out = 24'(316);
			19429: out = 24'(340);
			19430: out = 24'(316);
			19431: out = 24'(332);
			19432: out = 24'(272);
			19433: out = 24'(312);
			19434: out = 24'(292);
			19435: out = 24'(296);
			19436: out = 24'(336);
			19437: out = 24'(212);
			19438: out = 24'(268);
			19439: out = 24'(248);
			19440: out = 24'(292);
			19441: out = 24'(228);
			19442: out = 24'(228);
			19443: out = 24'(244);
			19444: out = 24'(240);
			19445: out = 24'(204);
			19446: out = 24'(232);
			19447: out = 24'(212);
			19448: out = 24'(196);
			19449: out = 24'(204);
			19450: out = 24'(200);
			19451: out = 24'(224);
			19452: out = 24'(164);
			19453: out = 24'(196);
			19454: out = 24'(196);
			19455: out = 24'(184);
			19456: out = 24'(168);
			19457: out = 24'(164);
			19458: out = 24'(160);
			19459: out = 24'(156);
			19460: out = 24'(148);
			19461: out = 24'(148);
			19462: out = 24'(172);
			19463: out = 24'(116);
			19464: out = 24'(164);
			19465: out = 24'(124);
			19466: out = 24'(100);
			19467: out = 24'(148);
			19468: out = 24'(148);
			19469: out = 24'(84);
			19470: out = 24'(120);
			19471: out = 24'(88);
			19472: out = 24'(116);
			19473: out = 24'(96);
			19474: out = 24'(100);
			19475: out = 24'(84);
			19476: out = 24'(64);
			19477: out = 24'(112);
			19478: out = 24'(80);
			19479: out = 24'(68);
			19480: out = 24'(100);
			19481: out = 24'(52);
			19482: out = 24'(60);
			19483: out = 24'(32);
			19484: out = 24'(100);
			19485: out = 24'(36);
			19486: out = 24'(48);
			19487: out = 24'(20);
			19488: out = 24'(36);
			19489: out = 24'(40);
			19490: out = 24'(24);
			19491: out = 24'(16);
			19492: out = 24'(8);
			19493: out = 24'(32);
			19494: out = 24'(-36);
			19495: out = 24'(-16);
			19496: out = 24'(4);
			19497: out = 24'(-72);
			19498: out = 24'(-28);
			19499: out = 24'(-60);
			19500: out = 24'(-64);
			19501: out = 24'(-52);
			19502: out = 24'(-104);
			19503: out = 24'(-68);
			19504: out = 24'(-120);
			19505: out = 24'(-84);
			19506: out = 24'(-128);
			19507: out = 24'(-80);
			19508: out = 24'(-164);
			19509: out = 24'(-100);
			19510: out = 24'(-160);
			19511: out = 24'(-116);
			19512: out = 24'(-152);
			19513: out = 24'(-164);
			19514: out = 24'(-184);
			19515: out = 24'(-172);
			19516: out = 24'(-116);
			19517: out = 24'(-244);
			19518: out = 24'(-172);
			19519: out = 24'(-192);
			19520: out = 24'(-196);
			19521: out = 24'(-208);
			19522: out = 24'(-224);
			19523: out = 24'(-220);
			19524: out = 24'(-212);
			19525: out = 24'(-220);
			19526: out = 24'(-196);
			19527: out = 24'(-272);
			19528: out = 24'(-228);
			19529: out = 24'(-220);
			19530: out = 24'(-252);
			19531: out = 24'(-280);
			19532: out = 24'(-244);
			19533: out = 24'(-272);
			19534: out = 24'(-288);
			19535: out = 24'(-296);
			19536: out = 24'(-308);
			19537: out = 24'(-268);
			19538: out = 24'(-332);
			19539: out = 24'(-300);
			19540: out = 24'(-288);
			19541: out = 24'(-316);
			19542: out = 24'(-336);
			19543: out = 24'(-316);
			19544: out = 24'(-320);
			19545: out = 24'(-344);
			19546: out = 24'(-356);
			19547: out = 24'(-368);
			19548: out = 24'(-384);
			19549: out = 24'(-348);
			19550: out = 24'(-380);
			19551: out = 24'(-352);
			19552: out = 24'(-420);
			19553: out = 24'(-344);
			19554: out = 24'(-400);
			19555: out = 24'(-380);
			19556: out = 24'(-416);
			19557: out = 24'(-392);
			19558: out = 24'(-400);
			19559: out = 24'(-416);
			19560: out = 24'(-452);
			19561: out = 24'(-400);
			19562: out = 24'(-448);
			19563: out = 24'(-432);
			19564: out = 24'(-488);
			19565: out = 24'(-420);
			19566: out = 24'(-480);
			19567: out = 24'(-464);
			19568: out = 24'(-468);
			19569: out = 24'(-452);
			19570: out = 24'(-524);
			19571: out = 24'(-448);
			19572: out = 24'(-508);
			19573: out = 24'(-452);
			19574: out = 24'(-508);
			19575: out = 24'(-536);
			19576: out = 24'(-480);
			19577: out = 24'(-524);
			19578: out = 24'(-536);
			19579: out = 24'(-528);
			19580: out = 24'(-528);
			19581: out = 24'(-548);
			19582: out = 24'(-552);
			19583: out = 24'(-548);
			19584: out = 24'(-548);
			19585: out = 24'(-560);
			19586: out = 24'(-580);
			19587: out = 24'(-580);
			19588: out = 24'(-572);
			19589: out = 24'(-600);
			19590: out = 24'(-608);
			19591: out = 24'(-608);
			19592: out = 24'(-624);
			19593: out = 24'(-624);
			19594: out = 24'(-644);
			19595: out = 24'(-628);
			19596: out = 24'(-652);
			19597: out = 24'(-672);
			19598: out = 24'(-664);
			19599: out = 24'(-676);
			19600: out = 24'(-700);
			19601: out = 24'(-692);
			19602: out = 24'(-700);
			19603: out = 24'(-684);
			19604: out = 24'(-696);
			19605: out = 24'(-764);
			19606: out = 24'(-728);
			19607: out = 24'(-720);
			19608: out = 24'(-772);
			19609: out = 24'(-748);
			19610: out = 24'(-760);
			19611: out = 24'(-828);
			19612: out = 24'(-748);
			19613: out = 24'(-820);
			19614: out = 24'(-800);
			19615: out = 24'(-820);
			19616: out = 24'(-860);
			19617: out = 24'(-800);
			19618: out = 24'(-900);
			19619: out = 24'(-844);
			19620: out = 24'(-904);
			19621: out = 24'(-856);
			19622: out = 24'(-908);
			19623: out = 24'(-876);
			19624: out = 24'(-956);
			19625: out = 24'(-880);
			19626: out = 24'(-956);
			19627: out = 24'(-952);
			19628: out = 24'(-972);
			19629: out = 24'(-940);
			19630: out = 24'(-976);
			19631: out = 24'(-980);
			19632: out = 24'(-1000);
			19633: out = 24'(-1000);
			19634: out = 24'(-1004);
			19635: out = 24'(-1068);
			19636: out = 24'(-1016);
			19637: out = 24'(-1092);
			19638: out = 24'(-1052);
			19639: out = 24'(-1060);
			19640: out = 24'(-1084);
			19641: out = 24'(-1044);
			19642: out = 24'(-1128);
			19643: out = 24'(-1052);
			19644: out = 24'(-1128);
			19645: out = 24'(-1084);
			19646: out = 24'(-1104);
			19647: out = 24'(-1160);
			19648: out = 24'(-1116);
			19649: out = 24'(-1120);
			19650: out = 24'(-1152);
			19651: out = 24'(-1144);
			19652: out = 24'(-1116);
			19653: out = 24'(-1184);
			19654: out = 24'(-1164);
			19655: out = 24'(-1168);
			19656: out = 24'(-1144);
			19657: out = 24'(-1216);
			19658: out = 24'(-1188);
			19659: out = 24'(-1192);
			19660: out = 24'(-1200);
			19661: out = 24'(-1200);
			19662: out = 24'(-1224);
			19663: out = 24'(-1208);
			19664: out = 24'(-1220);
			19665: out = 24'(-1220);
			19666: out = 24'(-1240);
			19667: out = 24'(-1216);
			19668: out = 24'(-1248);
			19669: out = 24'(-1256);
			19670: out = 24'(-1252);
			19671: out = 24'(-1200);
			19672: out = 24'(-1264);
			19673: out = 24'(-1256);
			19674: out = 24'(-1232);
			19675: out = 24'(-1264);
			19676: out = 24'(-1296);
			19677: out = 24'(-1240);
			19678: out = 24'(-1272);
			19679: out = 24'(-1284);
			19680: out = 24'(-1252);
			19681: out = 24'(-1292);
			19682: out = 24'(-1284);
			19683: out = 24'(-1268);
			19684: out = 24'(-1288);
			19685: out = 24'(-1268);
			19686: out = 24'(-1260);
			19687: out = 24'(-1316);
			19688: out = 24'(-1288);
			19689: out = 24'(-1292);
			19690: out = 24'(-1296);
			19691: out = 24'(-1268);
			19692: out = 24'(-1332);
			19693: out = 24'(-1292);
			19694: out = 24'(-1280);
			19695: out = 24'(-1300);
			19696: out = 24'(-1292);
			19697: out = 24'(-1312);
			19698: out = 24'(-1280);
			19699: out = 24'(-1292);
			19700: out = 24'(-1332);
			19701: out = 24'(-1284);
			19702: out = 24'(-1296);
			19703: out = 24'(-1312);
			19704: out = 24'(-1312);
			19705: out = 24'(-1316);
			19706: out = 24'(-1308);
			19707: out = 24'(-1336);
			19708: out = 24'(-1304);
			19709: out = 24'(-1320);
			19710: out = 24'(-1328);
			19711: out = 24'(-1312);
			19712: out = 24'(-1292);
			19713: out = 24'(-1328);
			19714: out = 24'(-1328);
			19715: out = 24'(-1316);
			19716: out = 24'(-1272);
			19717: out = 24'(-1316);
			19718: out = 24'(-1340);
			19719: out = 24'(-1284);
			19720: out = 24'(-1308);
			19721: out = 24'(-1280);
			19722: out = 24'(-1348);
			19723: out = 24'(-1316);
			19724: out = 24'(-1252);
			19725: out = 24'(-1332);
			19726: out = 24'(-1316);
			19727: out = 24'(-1280);
			19728: out = 24'(-1284);
			19729: out = 24'(-1332);
			19730: out = 24'(-1292);
			19731: out = 24'(-1280);
			19732: out = 24'(-1320);
			19733: out = 24'(-1304);
			19734: out = 24'(-1288);
			19735: out = 24'(-1320);
			19736: out = 24'(-1280);
			19737: out = 24'(-1312);
			19738: out = 24'(-1280);
			19739: out = 24'(-1296);
			19740: out = 24'(-1312);
			19741: out = 24'(-1256);
			19742: out = 24'(-1284);
			19743: out = 24'(-1272);
			19744: out = 24'(-1284);
			19745: out = 24'(-1288);
			19746: out = 24'(-1296);
			19747: out = 24'(-1268);
			19748: out = 24'(-1284);
			19749: out = 24'(-1304);
			19750: out = 24'(-1236);
			19751: out = 24'(-1308);
			19752: out = 24'(-1236);
			19753: out = 24'(-1272);
			19754: out = 24'(-1256);
			19755: out = 24'(-1252);
			19756: out = 24'(-1264);
			19757: out = 24'(-1240);
			19758: out = 24'(-1220);
			19759: out = 24'(-1304);
			19760: out = 24'(-1236);
			19761: out = 24'(-1204);
			19762: out = 24'(-1284);
			19763: out = 24'(-1252);
			19764: out = 24'(-1220);
			19765: out = 24'(-1252);
			19766: out = 24'(-1240);
			19767: out = 24'(-1224);
			19768: out = 24'(-1240);
			19769: out = 24'(-1220);
			19770: out = 24'(-1192);
			19771: out = 24'(-1280);
			19772: out = 24'(-1236);
			19773: out = 24'(-1196);
			19774: out = 24'(-1244);
			19775: out = 24'(-1152);
			19776: out = 24'(-1264);
			19777: out = 24'(-1192);
			19778: out = 24'(-1188);
			19779: out = 24'(-1200);
			19780: out = 24'(-1196);
			19781: out = 24'(-1188);
			19782: out = 24'(-1200);
			19783: out = 24'(-1148);
			19784: out = 24'(-1192);
			19785: out = 24'(-1200);
			19786: out = 24'(-1152);
			19787: out = 24'(-1152);
			19788: out = 24'(-1184);
			19789: out = 24'(-1164);
			19790: out = 24'(-1144);
			19791: out = 24'(-1144);
			19792: out = 24'(-1172);
			19793: out = 24'(-1132);
			19794: out = 24'(-1144);
			19795: out = 24'(-1132);
			19796: out = 24'(-1140);
			19797: out = 24'(-1108);
			19798: out = 24'(-1092);
			19799: out = 24'(-1100);
			19800: out = 24'(-1132);
			19801: out = 24'(-1076);
			19802: out = 24'(-1116);
			19803: out = 24'(-1092);
			19804: out = 24'(-1064);
			19805: out = 24'(-1104);
			19806: out = 24'(-1092);
			19807: out = 24'(-1032);
			19808: out = 24'(-1048);
			19809: out = 24'(-1064);
			19810: out = 24'(-1044);
			19811: out = 24'(-996);
			19812: out = 24'(-1072);
			19813: out = 24'(-1024);
			19814: out = 24'(-980);
			19815: out = 24'(-1044);
			19816: out = 24'(-1000);
			19817: out = 24'(-1000);
			19818: out = 24'(-988);
			19819: out = 24'(-976);
			19820: out = 24'(-964);
			19821: out = 24'(-964);
			19822: out = 24'(-952);
			19823: out = 24'(-968);
			19824: out = 24'(-876);
			19825: out = 24'(-936);
			19826: out = 24'(-956);
			19827: out = 24'(-884);
			19828: out = 24'(-908);
			19829: out = 24'(-876);
			19830: out = 24'(-900);
			19831: out = 24'(-864);
			19832: out = 24'(-848);
			19833: out = 24'(-860);
			19834: out = 24'(-856);
			19835: out = 24'(-840);
			19836: out = 24'(-828);
			19837: out = 24'(-816);
			19838: out = 24'(-812);
			19839: out = 24'(-796);
			19840: out = 24'(-812);
			19841: out = 24'(-772);
			19842: out = 24'(-788);
			19843: out = 24'(-780);
			19844: out = 24'(-760);
			19845: out = 24'(-788);
			19846: out = 24'(-724);
			19847: out = 24'(-776);
			19848: out = 24'(-716);
			19849: out = 24'(-732);
			19850: out = 24'(-732);
			19851: out = 24'(-712);
			19852: out = 24'(-700);
			19853: out = 24'(-700);
			19854: out = 24'(-688);
			19855: out = 24'(-668);
			19856: out = 24'(-684);
			19857: out = 24'(-652);
			19858: out = 24'(-676);
			19859: out = 24'(-656);
			19860: out = 24'(-600);
			19861: out = 24'(-676);
			19862: out = 24'(-672);
			19863: out = 24'(-572);
			19864: out = 24'(-648);
			19865: out = 24'(-604);
			19866: out = 24'(-608);
			19867: out = 24'(-576);
			19868: out = 24'(-624);
			19869: out = 24'(-572);
			19870: out = 24'(-572);
			19871: out = 24'(-560);
			19872: out = 24'(-540);
			19873: out = 24'(-592);
			19874: out = 24'(-580);
			19875: out = 24'(-496);
			19876: out = 24'(-584);
			19877: out = 24'(-500);
			19878: out = 24'(-524);
			19879: out = 24'(-528);
			19880: out = 24'(-524);
			19881: out = 24'(-484);
			19882: out = 24'(-496);
			19883: out = 24'(-544);
			19884: out = 24'(-476);
			19885: out = 24'(-484);
			19886: out = 24'(-468);
			19887: out = 24'(-492);
			19888: out = 24'(-484);
			19889: out = 24'(-476);
			19890: out = 24'(-412);
			19891: out = 24'(-480);
			19892: out = 24'(-464);
			19893: out = 24'(-436);
			19894: out = 24'(-444);
			19895: out = 24'(-448);
			19896: out = 24'(-412);
			19897: out = 24'(-448);
			19898: out = 24'(-420);
			19899: out = 24'(-396);
			19900: out = 24'(-416);
			19901: out = 24'(-404);
			19902: out = 24'(-368);
			19903: out = 24'(-412);
			19904: out = 24'(-420);
			19905: out = 24'(-380);
			19906: out = 24'(-360);
			19907: out = 24'(-380);
			19908: out = 24'(-416);
			19909: out = 24'(-340);
			19910: out = 24'(-400);
			19911: out = 24'(-324);
			19912: out = 24'(-352);
			19913: out = 24'(-356);
			19914: out = 24'(-352);
			19915: out = 24'(-336);
			19916: out = 24'(-340);
			19917: out = 24'(-320);
			19918: out = 24'(-312);
			19919: out = 24'(-340);
			19920: out = 24'(-316);
			19921: out = 24'(-268);
			19922: out = 24'(-304);
			19923: out = 24'(-292);
			19924: out = 24'(-280);
			19925: out = 24'(-272);
			19926: out = 24'(-296);
			19927: out = 24'(-272);
			19928: out = 24'(-244);
			19929: out = 24'(-272);
			19930: out = 24'(-228);
			19931: out = 24'(-260);
			19932: out = 24'(-192);
			19933: out = 24'(-244);
			19934: out = 24'(-232);
			19935: out = 24'(-208);
			19936: out = 24'(-184);
			19937: out = 24'(-180);
			19938: out = 24'(-216);
			19939: out = 24'(-180);
			19940: out = 24'(-196);
			19941: out = 24'(-148);
			19942: out = 24'(-176);
			19943: out = 24'(-224);
			19944: out = 24'(-144);
			19945: out = 24'(-152);
			19946: out = 24'(-148);
			19947: out = 24'(-148);
			19948: out = 24'(-148);
			19949: out = 24'(-124);
			19950: out = 24'(-152);
			19951: out = 24'(-128);
			19952: out = 24'(-124);
			19953: out = 24'(-136);
			19954: out = 24'(-96);
			19955: out = 24'(-168);
			19956: out = 24'(-84);
			19957: out = 24'(-96);
			19958: out = 24'(-120);
			19959: out = 24'(-88);
			19960: out = 24'(-100);
			19961: out = 24'(-96);
			19962: out = 24'(-80);
			19963: out = 24'(-68);
			19964: out = 24'(-80);
			19965: out = 24'(-88);
			19966: out = 24'(-56);
			19967: out = 24'(-64);
			19968: out = 24'(-72);
			19969: out = 24'(-68);
			19970: out = 24'(-72);
			19971: out = 24'(-16);
			19972: out = 24'(-80);
			19973: out = 24'(-60);
			19974: out = 24'(-20);
			19975: out = 24'(-20);
			19976: out = 24'(-36);
			19977: out = 24'(-20);
			19978: out = 24'(0);
			19979: out = 24'(24);
			19980: out = 24'(-52);
			19981: out = 24'(16);
			19982: out = 24'(20);
			19983: out = 24'(-40);
			19984: out = 24'(4);
			19985: out = 24'(-16);
			19986: out = 24'(56);
			19987: out = 24'(-12);
			19988: out = 24'(12);
			19989: out = 24'(56);
			19990: out = 24'(0);
			19991: out = 24'(32);
			19992: out = 24'(56);
			19993: out = 24'(40);
			19994: out = 24'(60);
			19995: out = 24'(60);
			19996: out = 24'(56);
			19997: out = 24'(48);
			19998: out = 24'(100);
			19999: out = 24'(28);
			20000: out = 24'(52);
			20001: out = 24'(132);
			20002: out = 24'(52);
			20003: out = 24'(72);
			20004: out = 24'(112);
			20005: out = 24'(116);
			20006: out = 24'(88);
			20007: out = 24'(116);
			20008: out = 24'(112);
			20009: out = 24'(96);
			20010: out = 24'(132);
			20011: out = 24'(144);
			20012: out = 24'(120);
			20013: out = 24'(152);
			20014: out = 24'(148);
			20015: out = 24'(160);
			20016: out = 24'(172);
			20017: out = 24'(184);
			20018: out = 24'(172);
			20019: out = 24'(180);
			20020: out = 24'(200);
			20021: out = 24'(204);
			20022: out = 24'(164);
			20023: out = 24'(220);
			20024: out = 24'(212);
			20025: out = 24'(220);
			20026: out = 24'(220);
			20027: out = 24'(232);
			20028: out = 24'(264);
			20029: out = 24'(224);
			20030: out = 24'(272);
			20031: out = 24'(256);
			20032: out = 24'(276);
			20033: out = 24'(248);
			20034: out = 24'(312);
			20035: out = 24'(256);
			20036: out = 24'(308);
			20037: out = 24'(296);
			20038: out = 24'(340);
			20039: out = 24'(320);
			20040: out = 24'(332);
			20041: out = 24'(348);
			20042: out = 24'(348);
			20043: out = 24'(372);
			20044: out = 24'(344);
			20045: out = 24'(368);
			20046: out = 24'(348);
			20047: out = 24'(400);
			20048: out = 24'(380);
			20049: out = 24'(420);
			20050: out = 24'(384);
			20051: out = 24'(436);
			20052: out = 24'(400);
			20053: out = 24'(432);
			20054: out = 24'(448);
			20055: out = 24'(440);
			20056: out = 24'(392);
			20057: out = 24'(488);
			20058: out = 24'(444);
			20059: out = 24'(488);
			20060: out = 24'(452);
			20061: out = 24'(460);
			20062: out = 24'(504);
			20063: out = 24'(484);
			20064: out = 24'(488);
			20065: out = 24'(512);
			20066: out = 24'(524);
			20067: out = 24'(480);
			20068: out = 24'(544);
			20069: out = 24'(516);
			20070: out = 24'(512);
			20071: out = 24'(528);
			20072: out = 24'(556);
			20073: out = 24'(496);
			20074: out = 24'(564);
			20075: out = 24'(564);
			20076: out = 24'(536);
			20077: out = 24'(576);
			20078: out = 24'(508);
			20079: out = 24'(600);
			20080: out = 24'(572);
			20081: out = 24'(580);
			20082: out = 24'(560);
			20083: out = 24'(624);
			20084: out = 24'(584);
			20085: out = 24'(620);
			20086: out = 24'(616);
			20087: out = 24'(584);
			20088: out = 24'(628);
			20089: out = 24'(644);
			20090: out = 24'(572);
			20091: out = 24'(628);
			20092: out = 24'(624);
			20093: out = 24'(628);
			20094: out = 24'(684);
			20095: out = 24'(636);
			20096: out = 24'(620);
			20097: out = 24'(668);
			20098: out = 24'(664);
			20099: out = 24'(668);
			20100: out = 24'(664);
			20101: out = 24'(644);
			20102: out = 24'(664);
			20103: out = 24'(692);
			20104: out = 24'(668);
			20105: out = 24'(680);
			20106: out = 24'(696);
			20107: out = 24'(680);
			20108: out = 24'(696);
			20109: out = 24'(684);
			20110: out = 24'(704);
			20111: out = 24'(656);
			20112: out = 24'(728);
			20113: out = 24'(684);
			20114: out = 24'(704);
			20115: out = 24'(732);
			20116: out = 24'(656);
			20117: out = 24'(712);
			20118: out = 24'(728);
			20119: out = 24'(740);
			20120: out = 24'(728);
			20121: out = 24'(720);
			20122: out = 24'(740);
			20123: out = 24'(720);
			20124: out = 24'(716);
			20125: out = 24'(784);
			20126: out = 24'(688);
			20127: out = 24'(744);
			20128: out = 24'(752);
			20129: out = 24'(752);
			20130: out = 24'(772);
			20131: out = 24'(740);
			20132: out = 24'(764);
			20133: out = 24'(752);
			20134: out = 24'(752);
			20135: out = 24'(776);
			20136: out = 24'(776);
			20137: out = 24'(764);
			20138: out = 24'(784);
			20139: out = 24'(736);
			20140: out = 24'(792);
			20141: out = 24'(768);
			20142: out = 24'(784);
			20143: out = 24'(744);
			20144: out = 24'(796);
			20145: out = 24'(780);
			20146: out = 24'(752);
			20147: out = 24'(780);
			20148: out = 24'(796);
			20149: out = 24'(760);
			20150: out = 24'(816);
			20151: out = 24'(776);
			20152: out = 24'(752);
			20153: out = 24'(808);
			20154: out = 24'(740);
			20155: out = 24'(836);
			20156: out = 24'(732);
			20157: out = 24'(768);
			20158: out = 24'(808);
			20159: out = 24'(784);
			20160: out = 24'(760);
			20161: out = 24'(792);
			20162: out = 24'(784);
			20163: out = 24'(776);
			20164: out = 24'(796);
			20165: out = 24'(752);
			20166: out = 24'(752);
			20167: out = 24'(772);
			20168: out = 24'(776);
			20169: out = 24'(732);
			20170: out = 24'(780);
			20171: out = 24'(768);
			20172: out = 24'(716);
			20173: out = 24'(796);
			20174: out = 24'(760);
			20175: out = 24'(724);
			20176: out = 24'(792);
			20177: out = 24'(724);
			20178: out = 24'(776);
			20179: out = 24'(768);
			20180: out = 24'(716);
			20181: out = 24'(768);
			20182: out = 24'(764);
			20183: out = 24'(732);
			20184: out = 24'(768);
			20185: out = 24'(760);
			20186: out = 24'(724);
			20187: out = 24'(768);
			20188: out = 24'(732);
			20189: out = 24'(752);
			20190: out = 24'(716);
			20191: out = 24'(732);
			20192: out = 24'(748);
			20193: out = 24'(752);
			20194: out = 24'(752);
			20195: out = 24'(696);
			20196: out = 24'(780);
			20197: out = 24'(728);
			20198: out = 24'(732);
			20199: out = 24'(768);
			20200: out = 24'(692);
			20201: out = 24'(716);
			20202: out = 24'(760);
			20203: out = 24'(716);
			20204: out = 24'(740);
			20205: out = 24'(724);
			20206: out = 24'(732);
			20207: out = 24'(724);
			20208: out = 24'(732);
			20209: out = 24'(748);
			20210: out = 24'(740);
			20211: out = 24'(680);
			20212: out = 24'(740);
			20213: out = 24'(732);
			20214: out = 24'(700);
			20215: out = 24'(680);
			20216: out = 24'(732);
			20217: out = 24'(724);
			20218: out = 24'(668);
			20219: out = 24'(712);
			20220: out = 24'(704);
			20221: out = 24'(696);
			20222: out = 24'(692);
			20223: out = 24'(680);
			20224: out = 24'(648);
			20225: out = 24'(676);
			20226: out = 24'(688);
			20227: out = 24'(668);
			20228: out = 24'(656);
			20229: out = 24'(656);
			20230: out = 24'(684);
			20231: out = 24'(672);
			20232: out = 24'(656);
			20233: out = 24'(644);
			20234: out = 24'(668);
			20235: out = 24'(632);
			20236: out = 24'(688);
			20237: out = 24'(632);
			20238: out = 24'(644);
			20239: out = 24'(644);
			20240: out = 24'(596);
			20241: out = 24'(664);
			20242: out = 24'(604);
			20243: out = 24'(628);
			20244: out = 24'(616);
			20245: out = 24'(624);
			20246: out = 24'(632);
			20247: out = 24'(584);
			20248: out = 24'(592);
			20249: out = 24'(608);
			20250: out = 24'(564);
			20251: out = 24'(600);
			20252: out = 24'(572);
			20253: out = 24'(560);
			20254: out = 24'(576);
			20255: out = 24'(556);
			20256: out = 24'(556);
			20257: out = 24'(544);
			20258: out = 24'(552);
			20259: out = 24'(496);
			20260: out = 24'(560);
			20261: out = 24'(492);
			20262: out = 24'(556);
			20263: out = 24'(464);
			20264: out = 24'(476);
			20265: out = 24'(500);
			20266: out = 24'(500);
			20267: out = 24'(460);
			20268: out = 24'(464);
			20269: out = 24'(496);
			20270: out = 24'(440);
			20271: out = 24'(464);
			20272: out = 24'(456);
			20273: out = 24'(408);
			20274: out = 24'(420);
			20275: out = 24'(456);
			20276: out = 24'(408);
			20277: out = 24'(416);
			20278: out = 24'(440);
			20279: out = 24'(396);
			20280: out = 24'(428);
			20281: out = 24'(388);
			20282: out = 24'(420);
			20283: out = 24'(388);
			20284: out = 24'(392);
			20285: out = 24'(368);
			20286: out = 24'(372);
			20287: out = 24'(344);
			20288: out = 24'(392);
			20289: out = 24'(360);
			20290: out = 24'(316);
			20291: out = 24'(348);
			20292: out = 24'(364);
			20293: out = 24'(312);
			20294: out = 24'(336);
			20295: out = 24'(300);
			20296: out = 24'(304);
			20297: out = 24'(312);
			20298: out = 24'(304);
			20299: out = 24'(268);
			20300: out = 24'(300);
			20301: out = 24'(276);
			20302: out = 24'(276);
			20303: out = 24'(308);
			20304: out = 24'(252);
			20305: out = 24'(296);
			20306: out = 24'(216);
			20307: out = 24'(264);
			20308: out = 24'(280);
			20309: out = 24'(228);
			20310: out = 24'(216);
			20311: out = 24'(260);
			20312: out = 24'(248);
			20313: out = 24'(276);
			20314: out = 24'(192);
			20315: out = 24'(228);
			20316: out = 24'(248);
			20317: out = 24'(216);
			20318: out = 24'(184);
			20319: out = 24'(212);
			20320: out = 24'(200);
			20321: out = 24'(208);
			20322: out = 24'(144);
			20323: out = 24'(208);
			20324: out = 24'(152);
			20325: out = 24'(184);
			20326: out = 24'(128);
			20327: out = 24'(196);
			20328: out = 24'(132);
			20329: out = 24'(136);
			20330: out = 24'(160);
			20331: out = 24'(136);
			20332: out = 24'(176);
			20333: out = 24'(88);
			20334: out = 24'(148);
			20335: out = 24'(116);
			20336: out = 24'(160);
			20337: out = 24'(136);
			20338: out = 24'(60);
			20339: out = 24'(156);
			20340: out = 24'(96);
			20341: out = 24'(160);
			20342: out = 24'(56);
			20343: out = 24'(112);
			20344: out = 24'(104);
			20345: out = 24'(128);
			20346: out = 24'(72);
			20347: out = 24'(100);
			20348: out = 24'(112);
			20349: out = 24'(112);
			20350: out = 24'(56);
			20351: out = 24'(68);
			20352: out = 24'(60);
			20353: out = 24'(104);
			20354: out = 24'(12);
			20355: out = 24'(88);
			20356: out = 24'(48);
			20357: out = 24'(28);
			20358: out = 24'(40);
			20359: out = 24'(28);
			20360: out = 24'(48);
			20361: out = 24'(4);
			20362: out = 24'(36);
			20363: out = 24'(28);
			20364: out = 24'(32);
			20365: out = 24'(36);
			20366: out = 24'(-20);
			20367: out = 24'(24);
			20368: out = 24'(24);
			20369: out = 24'(16);
			20370: out = 24'(0);
			20371: out = 24'(-12);
			20372: out = 24'(32);
			20373: out = 24'(-8);
			20374: out = 24'(28);
			20375: out = 24'(-36);
			20376: out = 24'(40);
			20377: out = 24'(-12);
			20378: out = 24'(4);
			20379: out = 24'(16);
			20380: out = 24'(-56);
			20381: out = 24'(-4);
			20382: out = 24'(-20);
			20383: out = 24'(-24);
			20384: out = 24'(-32);
			20385: out = 24'(-52);
			20386: out = 24'(-32);
			20387: out = 24'(-96);
			20388: out = 24'(-16);
			20389: out = 24'(-96);
			20390: out = 24'(-52);
			20391: out = 24'(-88);
			20392: out = 24'(-84);
			20393: out = 24'(-124);
			20394: out = 24'(-108);
			20395: out = 24'(-112);
			20396: out = 24'(-108);
			20397: out = 24'(-144);
			20398: out = 24'(-116);
			20399: out = 24'(-136);
			20400: out = 24'(-148);
			20401: out = 24'(-132);
			20402: out = 24'(-156);
			20403: out = 24'(-180);
			20404: out = 24'(-180);
			20405: out = 24'(-152);
			20406: out = 24'(-148);
			20407: out = 24'(-220);
			20408: out = 24'(-168);
			20409: out = 24'(-196);
			20410: out = 24'(-168);
			20411: out = 24'(-192);
			20412: out = 24'(-216);
			20413: out = 24'(-180);
			20414: out = 24'(-212);
			20415: out = 24'(-228);
			20416: out = 24'(-196);
			20417: out = 24'(-212);
			20418: out = 24'(-216);
			20419: out = 24'(-256);
			20420: out = 24'(-172);
			20421: out = 24'(-268);
			20422: out = 24'(-232);
			20423: out = 24'(-224);
			20424: out = 24'(-276);
			20425: out = 24'(-248);
			20426: out = 24'(-252);
			20427: out = 24'(-252);
			20428: out = 24'(-256);
			20429: out = 24'(-276);
			20430: out = 24'(-260);
			20431: out = 24'(-268);
			20432: out = 24'(-308);
			20433: out = 24'(-292);
			20434: out = 24'(-268);
			20435: out = 24'(-288);
			20436: out = 24'(-312);
			20437: out = 24'(-296);
			20438: out = 24'(-308);
			20439: out = 24'(-340);
			20440: out = 24'(-296);
			20441: out = 24'(-340);
			20442: out = 24'(-316);
			20443: out = 24'(-340);
			20444: out = 24'(-300);
			20445: out = 24'(-324);
			20446: out = 24'(-368);
			20447: out = 24'(-304);
			20448: out = 24'(-344);
			20449: out = 24'(-408);
			20450: out = 24'(-312);
			20451: out = 24'(-368);
			20452: out = 24'(-332);
			20453: out = 24'(-400);
			20454: out = 24'(-364);
			20455: out = 24'(-336);
			20456: out = 24'(-400);
			20457: out = 24'(-384);
			20458: out = 24'(-348);
			20459: out = 24'(-372);
			20460: out = 24'(-404);
			20461: out = 24'(-392);
			20462: out = 24'(-396);
			20463: out = 24'(-380);
			20464: out = 24'(-404);
			20465: out = 24'(-444);
			20466: out = 24'(-416);
			20467: out = 24'(-412);
			20468: out = 24'(-416);
			20469: out = 24'(-460);
			20470: out = 24'(-412);
			20471: out = 24'(-448);
			20472: out = 24'(-412);
			20473: out = 24'(-488);
			20474: out = 24'(-420);
			20475: out = 24'(-456);
			20476: out = 24'(-448);
			20477: out = 24'(-460);
			20478: out = 24'(-504);
			20479: out = 24'(-440);
			20480: out = 24'(-488);
			20481: out = 24'(-456);
			20482: out = 24'(-484);
			20483: out = 24'(-528);
			20484: out = 24'(-480);
			20485: out = 24'(-476);
			20486: out = 24'(-528);
			20487: out = 24'(-508);
			20488: out = 24'(-528);
			20489: out = 24'(-524);
			20490: out = 24'(-500);
			20491: out = 24'(-564);
			20492: out = 24'(-556);
			20493: out = 24'(-512);
			20494: out = 24'(-544);
			20495: out = 24'(-592);
			20496: out = 24'(-548);
			20497: out = 24'(-580);
			20498: out = 24'(-572);
			20499: out = 24'(-584);
			20500: out = 24'(-640);
			20501: out = 24'(-580);
			20502: out = 24'(-592);
			20503: out = 24'(-628);
			20504: out = 24'(-608);
			20505: out = 24'(-644);
			20506: out = 24'(-616);
			20507: out = 24'(-668);
			20508: out = 24'(-636);
			20509: out = 24'(-696);
			20510: out = 24'(-684);
			20511: out = 24'(-668);
			20512: out = 24'(-668);
			20513: out = 24'(-736);
			20514: out = 24'(-688);
			20515: out = 24'(-692);
			20516: out = 24'(-692);
			20517: out = 24'(-740);
			20518: out = 24'(-716);
			20519: out = 24'(-752);
			20520: out = 24'(-740);
			20521: out = 24'(-732);
			20522: out = 24'(-780);
			20523: out = 24'(-748);
			20524: out = 24'(-788);
			20525: out = 24'(-772);
			20526: out = 24'(-816);
			20527: out = 24'(-808);
			20528: out = 24'(-800);
			20529: out = 24'(-792);
			20530: out = 24'(-816);
			20531: out = 24'(-824);
			20532: out = 24'(-828);
			20533: out = 24'(-808);
			20534: out = 24'(-872);
			20535: out = 24'(-824);
			20536: out = 24'(-828);
			20537: out = 24'(-844);
			20538: out = 24'(-892);
			20539: out = 24'(-816);
			20540: out = 24'(-888);
			20541: out = 24'(-900);
			20542: out = 24'(-856);
			20543: out = 24'(-908);
			20544: out = 24'(-888);
			20545: out = 24'(-888);
			20546: out = 24'(-920);
			20547: out = 24'(-904);
			20548: out = 24'(-900);
			20549: out = 24'(-928);
			20550: out = 24'(-916);
			20551: out = 24'(-932);
			20552: out = 24'(-932);
			20553: out = 24'(-960);
			20554: out = 24'(-900);
			20555: out = 24'(-972);
			20556: out = 24'(-932);
			20557: out = 24'(-948);
			20558: out = 24'(-948);
			20559: out = 24'(-920);
			20560: out = 24'(-940);
			20561: out = 24'(-960);
			20562: out = 24'(-968);
			20563: out = 24'(-972);
			20564: out = 24'(-932);
			20565: out = 24'(-976);
			20566: out = 24'(-1016);
			20567: out = 24'(-932);
			20568: out = 24'(-964);
			20569: out = 24'(-972);
			20570: out = 24'(-1012);
			20571: out = 24'(-936);
			20572: out = 24'(-1000);
			20573: out = 24'(-984);
			20574: out = 24'(-996);
			20575: out = 24'(-996);
			20576: out = 24'(-1012);
			20577: out = 24'(-988);
			20578: out = 24'(-1000);
			20579: out = 24'(-988);
			20580: out = 24'(-980);
			20581: out = 24'(-1028);
			20582: out = 24'(-1008);
			20583: out = 24'(-1000);
			20584: out = 24'(-980);
			20585: out = 24'(-988);
			20586: out = 24'(-1052);
			20587: out = 24'(-980);
			20588: out = 24'(-1016);
			20589: out = 24'(-1032);
			20590: out = 24'(-988);
			20591: out = 24'(-1044);
			20592: out = 24'(-1008);
			20593: out = 24'(-1024);
			20594: out = 24'(-980);
			20595: out = 24'(-1020);
			20596: out = 24'(-1004);
			20597: out = 24'(-1028);
			20598: out = 24'(-964);
			20599: out = 24'(-1036);
			20600: out = 24'(-1044);
			20601: out = 24'(-1004);
			20602: out = 24'(-984);
			20603: out = 24'(-1024);
			20604: out = 24'(-1012);
			20605: out = 24'(-984);
			20606: out = 24'(-1004);
			20607: out = 24'(-980);
			20608: out = 24'(-1028);
			20609: out = 24'(-1004);
			20610: out = 24'(-1004);
			20611: out = 24'(-1008);
			20612: out = 24'(-1000);
			20613: out = 24'(-1012);
			20614: out = 24'(-1016);
			20615: out = 24'(-1000);
			20616: out = 24'(-1004);
			20617: out = 24'(-1020);
			20618: out = 24'(-1008);
			20619: out = 24'(-996);
			20620: out = 24'(-1012);
			20621: out = 24'(-1008);
			20622: out = 24'(-1016);
			20623: out = 24'(-1012);
			20624: out = 24'(-1020);
			20625: out = 24'(-976);
			20626: out = 24'(-1036);
			20627: out = 24'(-964);
			20628: out = 24'(-1020);
			20629: out = 24'(-956);
			20630: out = 24'(-1016);
			20631: out = 24'(-988);
			20632: out = 24'(-972);
			20633: out = 24'(-1004);
			20634: out = 24'(-1012);
			20635: out = 24'(-948);
			20636: out = 24'(-1024);
			20637: out = 24'(-1004);
			20638: out = 24'(-980);
			20639: out = 24'(-952);
			20640: out = 24'(-1008);
			20641: out = 24'(-976);
			20642: out = 24'(-940);
			20643: out = 24'(-980);
			20644: out = 24'(-980);
			20645: out = 24'(-976);
			20646: out = 24'(-968);
			20647: out = 24'(-972);
			20648: out = 24'(-960);
			20649: out = 24'(-948);
			20650: out = 24'(-960);
			20651: out = 24'(-964);
			20652: out = 24'(-952);
			20653: out = 24'(-976);
			20654: out = 24'(-920);
			20655: out = 24'(-952);
			20656: out = 24'(-964);
			20657: out = 24'(-936);
			20658: out = 24'(-948);
			20659: out = 24'(-936);
			20660: out = 24'(-968);
			20661: out = 24'(-904);
			20662: out = 24'(-996);
			20663: out = 24'(-932);
			20664: out = 24'(-932);
			20665: out = 24'(-936);
			20666: out = 24'(-920);
			20667: out = 24'(-948);
			20668: out = 24'(-932);
			20669: out = 24'(-916);
			20670: out = 24'(-892);
			20671: out = 24'(-956);
			20672: out = 24'(-892);
			20673: out = 24'(-916);
			20674: out = 24'(-968);
			20675: out = 24'(-864);
			20676: out = 24'(-920);
			20677: out = 24'(-920);
			20678: out = 24'(-888);
			20679: out = 24'(-916);
			20680: out = 24'(-840);
			20681: out = 24'(-936);
			20682: out = 24'(-884);
			20683: out = 24'(-880);
			20684: out = 24'(-856);
			20685: out = 24'(-928);
			20686: out = 24'(-836);
			20687: out = 24'(-904);
			20688: out = 24'(-828);
			20689: out = 24'(-880);
			20690: out = 24'(-888);
			20691: out = 24'(-872);
			20692: out = 24'(-856);
			20693: out = 24'(-840);
			20694: out = 24'(-848);
			20695: out = 24'(-844);
			20696: out = 24'(-836);
			20697: out = 24'(-816);
			20698: out = 24'(-824);
			20699: out = 24'(-840);
			20700: out = 24'(-784);
			20701: out = 24'(-836);
			20702: out = 24'(-788);
			20703: out = 24'(-840);
			20704: out = 24'(-736);
			20705: out = 24'(-792);
			20706: out = 24'(-796);
			20707: out = 24'(-764);
			20708: out = 24'(-776);
			20709: out = 24'(-768);
			20710: out = 24'(-752);
			20711: out = 24'(-760);
			20712: out = 24'(-744);
			20713: out = 24'(-720);
			20714: out = 24'(-768);
			20715: out = 24'(-728);
			20716: out = 24'(-720);
			20717: out = 24'(-736);
			20718: out = 24'(-744);
			20719: out = 24'(-696);
			20720: out = 24'(-704);
			20721: out = 24'(-728);
			20722: out = 24'(-692);
			20723: out = 24'(-688);
			20724: out = 24'(-704);
			20725: out = 24'(-664);
			20726: out = 24'(-684);
			20727: out = 24'(-672);
			20728: out = 24'(-644);
			20729: out = 24'(-644);
			20730: out = 24'(-632);
			20731: out = 24'(-640);
			20732: out = 24'(-656);
			20733: out = 24'(-604);
			20734: out = 24'(-616);
			20735: out = 24'(-628);
			20736: out = 24'(-572);
			20737: out = 24'(-608);
			20738: out = 24'(-592);
			20739: out = 24'(-596);
			20740: out = 24'(-544);
			20741: out = 24'(-592);
			20742: out = 24'(-556);
			20743: out = 24'(-560);
			20744: out = 24'(-516);
			20745: out = 24'(-576);
			20746: out = 24'(-532);
			20747: out = 24'(-532);
			20748: out = 24'(-548);
			20749: out = 24'(-528);
			20750: out = 24'(-492);
			20751: out = 24'(-556);
			20752: out = 24'(-468);
			20753: out = 24'(-564);
			20754: out = 24'(-488);
			20755: out = 24'(-500);
			20756: out = 24'(-532);
			20757: out = 24'(-460);
			20758: out = 24'(-504);
			20759: out = 24'(-468);
			20760: out = 24'(-484);
			20761: out = 24'(-448);
			20762: out = 24'(-476);
			20763: out = 24'(-460);
			20764: out = 24'(-460);
			20765: out = 24'(-480);
			20766: out = 24'(-476);
			20767: out = 24'(-404);
			20768: out = 24'(-476);
			20769: out = 24'(-420);
			20770: out = 24'(-440);
			20771: out = 24'(-408);
			20772: out = 24'(-444);
			20773: out = 24'(-396);
			20774: out = 24'(-408);
			20775: out = 24'(-420);
			20776: out = 24'(-404);
			20777: out = 24'(-384);
			20778: out = 24'(-404);
			20779: out = 24'(-372);
			20780: out = 24'(-388);
			20781: out = 24'(-420);
			20782: out = 24'(-372);
			20783: out = 24'(-400);
			20784: out = 24'(-340);
			20785: out = 24'(-392);
			20786: out = 24'(-384);
			20787: out = 24'(-360);
			20788: out = 24'(-332);
			20789: out = 24'(-332);
			20790: out = 24'(-368);
			20791: out = 24'(-340);
			20792: out = 24'(-324);
			20793: out = 24'(-356);
			20794: out = 24'(-344);
			20795: out = 24'(-324);
			20796: out = 24'(-320);
			20797: out = 24'(-344);
			20798: out = 24'(-332);
			20799: out = 24'(-288);
			20800: out = 24'(-320);
			20801: out = 24'(-300);
			20802: out = 24'(-308);
			20803: out = 24'(-276);
			20804: out = 24'(-308);
			20805: out = 24'(-264);
			20806: out = 24'(-276);
			20807: out = 24'(-300);
			20808: out = 24'(-264);
			20809: out = 24'(-276);
			20810: out = 24'(-288);
			20811: out = 24'(-300);
			20812: out = 24'(-224);
			20813: out = 24'(-268);
			20814: out = 24'(-232);
			20815: out = 24'(-264);
			20816: out = 24'(-208);
			20817: out = 24'(-248);
			20818: out = 24'(-204);
			20819: out = 24'(-244);
			20820: out = 24'(-240);
			20821: out = 24'(-228);
			20822: out = 24'(-172);
			20823: out = 24'(-212);
			20824: out = 24'(-204);
			20825: out = 24'(-200);
			20826: out = 24'(-180);
			20827: out = 24'(-200);
			20828: out = 24'(-208);
			20829: out = 24'(-168);
			20830: out = 24'(-192);
			20831: out = 24'(-160);
			20832: out = 24'(-180);
			20833: out = 24'(-152);
			20834: out = 24'(-136);
			20835: out = 24'(-164);
			20836: out = 24'(-168);
			20837: out = 24'(-160);
			20838: out = 24'(-156);
			20839: out = 24'(-132);
			20840: out = 24'(-124);
			20841: out = 24'(-152);
			20842: out = 24'(-148);
			20843: out = 24'(-108);
			20844: out = 24'(-120);
			20845: out = 24'(-108);
			20846: out = 24'(-132);
			20847: out = 24'(-136);
			20848: out = 24'(-112);
			20849: out = 24'(-80);
			20850: out = 24'(-124);
			20851: out = 24'(-112);
			20852: out = 24'(-84);
			20853: out = 24'(-84);
			20854: out = 24'(-100);
			20855: out = 24'(-72);
			20856: out = 24'(-104);
			20857: out = 24'(-104);
			20858: out = 24'(-80);
			20859: out = 24'(-76);
			20860: out = 24'(-76);
			20861: out = 24'(-84);
			20862: out = 24'(-88);
			20863: out = 24'(-48);
			20864: out = 24'(-84);
			20865: out = 24'(-68);
			20866: out = 24'(-64);
			20867: out = 24'(-32);
			20868: out = 24'(-36);
			20869: out = 24'(-100);
			20870: out = 24'(-32);
			20871: out = 24'(-24);
			20872: out = 24'(-40);
			20873: out = 24'(-52);
			20874: out = 24'(-28);
			20875: out = 24'(-40);
			20876: out = 24'(-36);
			20877: out = 24'(0);
			20878: out = 24'(-60);
			20879: out = 24'(-4);
			20880: out = 24'(-32);
			20881: out = 24'(8);
			20882: out = 24'(-20);
			20883: out = 24'(-32);
			20884: out = 24'(0);
			20885: out = 24'(0);
			20886: out = 24'(-4);
			20887: out = 24'(-28);
			20888: out = 24'(8);
			20889: out = 24'(28);
			20890: out = 24'(-24);
			20891: out = 24'(16);
			20892: out = 24'(40);
			20893: out = 24'(-36);
			20894: out = 24'(76);
			20895: out = 24'(4);
			20896: out = 24'(28);
			20897: out = 24'(20);
			20898: out = 24'(28);
			20899: out = 24'(72);
			20900: out = 24'(24);
			20901: out = 24'(68);
			20902: out = 24'(24);
			20903: out = 24'(96);
			20904: out = 24'(48);
			20905: out = 24'(84);
			20906: out = 24'(84);
			20907: out = 24'(76);
			20908: out = 24'(88);
			20909: out = 24'(80);
			20910: out = 24'(88);
			20911: out = 24'(100);
			20912: out = 24'(104);
			20913: out = 24'(88);
			20914: out = 24'(112);
			20915: out = 24'(112);
			20916: out = 24'(116);
			20917: out = 24'(96);
			20918: out = 24'(128);
			20919: out = 24'(144);
			20920: out = 24'(148);
			20921: out = 24'(144);
			20922: out = 24'(124);
			20923: out = 24'(164);
			20924: out = 24'(152);
			20925: out = 24'(160);
			20926: out = 24'(180);
			20927: out = 24'(152);
			20928: out = 24'(196);
			20929: out = 24'(220);
			20930: out = 24'(180);
			20931: out = 24'(184);
			20932: out = 24'(216);
			20933: out = 24'(252);
			20934: out = 24'(208);
			20935: out = 24'(228);
			20936: out = 24'(256);
			20937: out = 24'(232);
			20938: out = 24'(204);
			20939: out = 24'(296);
			20940: out = 24'(232);
			20941: out = 24'(248);
			20942: out = 24'(260);
			20943: out = 24'(292);
			20944: out = 24'(256);
			20945: out = 24'(280);
			20946: out = 24'(272);
			20947: out = 24'(296);
			20948: out = 24'(272);
			20949: out = 24'(304);
			20950: out = 24'(280);
			20951: out = 24'(336);
			20952: out = 24'(296);
			20953: out = 24'(276);
			20954: out = 24'(356);
			20955: out = 24'(280);
			20956: out = 24'(324);
			20957: out = 24'(336);
			20958: out = 24'(348);
			20959: out = 24'(308);
			20960: out = 24'(340);
			20961: out = 24'(380);
			20962: out = 24'(344);
			20963: out = 24'(356);
			20964: out = 24'(360);
			20965: out = 24'(356);
			20966: out = 24'(380);
			20967: out = 24'(400);
			20968: out = 24'(360);
			20969: out = 24'(388);
			20970: out = 24'(388);
			20971: out = 24'(408);
			20972: out = 24'(408);
			20973: out = 24'(364);
			20974: out = 24'(416);
			20975: out = 24'(420);
			20976: out = 24'(388);
			20977: out = 24'(412);
			20978: out = 24'(404);
			20979: out = 24'(440);
			20980: out = 24'(428);
			20981: out = 24'(404);
			20982: out = 24'(452);
			20983: out = 24'(428);
			20984: out = 24'(432);
			20985: out = 24'(420);
			20986: out = 24'(464);
			20987: out = 24'(432);
			20988: out = 24'(432);
			20989: out = 24'(464);
			20990: out = 24'(436);
			20991: out = 24'(456);
			20992: out = 24'(460);
			20993: out = 24'(460);
			20994: out = 24'(416);
			20995: out = 24'(488);
			20996: out = 24'(452);
			20997: out = 24'(452);
			20998: out = 24'(468);
			20999: out = 24'(468);
			21000: out = 24'(492);
			21001: out = 24'(444);
			21002: out = 24'(500);
			21003: out = 24'(464);
			21004: out = 24'(484);
			21005: out = 24'(480);
			21006: out = 24'(500);
			21007: out = 24'(512);
			21008: out = 24'(468);
			21009: out = 24'(500);
			21010: out = 24'(500);
			21011: out = 24'(500);
			21012: out = 24'(464);
			21013: out = 24'(512);
			21014: out = 24'(476);
			21015: out = 24'(508);
			21016: out = 24'(512);
			21017: out = 24'(468);
			21018: out = 24'(512);
			21019: out = 24'(492);
			21020: out = 24'(532);
			21021: out = 24'(488);
			21022: out = 24'(524);
			21023: out = 24'(508);
			21024: out = 24'(532);
			21025: out = 24'(540);
			21026: out = 24'(484);
			21027: out = 24'(524);
			21028: out = 24'(512);
			21029: out = 24'(564);
			21030: out = 24'(476);
			21031: out = 24'(524);
			21032: out = 24'(532);
			21033: out = 24'(512);
			21034: out = 24'(556);
			21035: out = 24'(484);
			21036: out = 24'(536);
			21037: out = 24'(516);
			21038: out = 24'(576);
			21039: out = 24'(488);
			21040: out = 24'(528);
			21041: out = 24'(536);
			21042: out = 24'(512);
			21043: out = 24'(480);
			21044: out = 24'(564);
			21045: out = 24'(508);
			21046: out = 24'(508);
			21047: out = 24'(540);
			21048: out = 24'(508);
			21049: out = 24'(532);
			21050: out = 24'(512);
			21051: out = 24'(516);
			21052: out = 24'(508);
			21053: out = 24'(468);
			21054: out = 24'(560);
			21055: out = 24'(492);
			21056: out = 24'(484);
			21057: out = 24'(532);
			21058: out = 24'(512);
			21059: out = 24'(500);
			21060: out = 24'(500);
			21061: out = 24'(504);
			21062: out = 24'(500);
			21063: out = 24'(484);
			21064: out = 24'(540);
			21065: out = 24'(496);
			21066: out = 24'(492);
			21067: out = 24'(492);
			21068: out = 24'(528);
			21069: out = 24'(484);
			21070: out = 24'(496);
			21071: out = 24'(464);
			21072: out = 24'(512);
			21073: out = 24'(516);
			21074: out = 24'(484);
			21075: out = 24'(492);
			21076: out = 24'(528);
			21077: out = 24'(512);
			21078: out = 24'(460);
			21079: out = 24'(516);
			21080: out = 24'(496);
			21081: out = 24'(452);
			21082: out = 24'(508);
			21083: out = 24'(460);
			21084: out = 24'(496);
			21085: out = 24'(476);
			21086: out = 24'(488);
			21087: out = 24'(500);
			21088: out = 24'(468);
			21089: out = 24'(496);
			21090: out = 24'(468);
			21091: out = 24'(492);
			21092: out = 24'(488);
			21093: out = 24'(440);
			21094: out = 24'(480);
			21095: out = 24'(468);
			21096: out = 24'(488);
			21097: out = 24'(464);
			21098: out = 24'(488);
			21099: out = 24'(448);
			21100: out = 24'(484);
			21101: out = 24'(480);
			21102: out = 24'(468);
			21103: out = 24'(460);
			21104: out = 24'(488);
			21105: out = 24'(436);
			21106: out = 24'(508);
			21107: out = 24'(444);
			21108: out = 24'(484);
			21109: out = 24'(460);
			21110: out = 24'(452);
			21111: out = 24'(464);
			21112: out = 24'(468);
			21113: out = 24'(440);
			21114: out = 24'(452);
			21115: out = 24'(464);
			21116: out = 24'(448);
			21117: out = 24'(428);
			21118: out = 24'(456);
			21119: out = 24'(448);
			21120: out = 24'(420);
			21121: out = 24'(452);
			21122: out = 24'(432);
			21123: out = 24'(416);
			21124: out = 24'(436);
			21125: out = 24'(440);
			21126: out = 24'(404);
			21127: out = 24'(400);
			21128: out = 24'(392);
			21129: out = 24'(404);
			21130: out = 24'(436);
			21131: out = 24'(392);
			21132: out = 24'(412);
			21133: out = 24'(404);
			21134: out = 24'(392);
			21135: out = 24'(432);
			21136: out = 24'(348);
			21137: out = 24'(380);
			21138: out = 24'(416);
			21139: out = 24'(384);
			21140: out = 24'(396);
			21141: out = 24'(356);
			21142: out = 24'(392);
			21143: out = 24'(380);
			21144: out = 24'(388);
			21145: out = 24'(344);
			21146: out = 24'(352);
			21147: out = 24'(364);
			21148: out = 24'(388);
			21149: out = 24'(320);
			21150: out = 24'(352);
			21151: out = 24'(320);
			21152: out = 24'(368);
			21153: out = 24'(332);
			21154: out = 24'(324);
			21155: out = 24'(320);
			21156: out = 24'(316);
			21157: out = 24'(312);
			21158: out = 24'(300);
			21159: out = 24'(312);
			21160: out = 24'(288);
			21161: out = 24'(308);
			21162: out = 24'(268);
			21163: out = 24'(272);
			21164: out = 24'(260);
			21165: out = 24'(308);
			21166: out = 24'(220);
			21167: out = 24'(256);
			21168: out = 24'(264);
			21169: out = 24'(244);
			21170: out = 24'(244);
			21171: out = 24'(252);
			21172: out = 24'(204);
			21173: out = 24'(228);
			21174: out = 24'(244);
			21175: out = 24'(208);
			21176: out = 24'(192);
			21177: out = 24'(240);
			21178: out = 24'(196);
			21179: out = 24'(200);
			21180: out = 24'(196);
			21181: out = 24'(200);
			21182: out = 24'(220);
			21183: out = 24'(200);
			21184: out = 24'(144);
			21185: out = 24'(200);
			21186: out = 24'(192);
			21187: out = 24'(192);
			21188: out = 24'(196);
			21189: out = 24'(152);
			21190: out = 24'(184);
			21191: out = 24'(168);
			21192: out = 24'(148);
			21193: out = 24'(152);
			21194: out = 24'(132);
			21195: out = 24'(168);
			21196: out = 24'(144);
			21197: out = 24'(160);
			21198: out = 24'(108);
			21199: out = 24'(184);
			21200: out = 24'(112);
			21201: out = 24'(124);
			21202: out = 24'(152);
			21203: out = 24'(84);
			21204: out = 24'(60);
			21205: out = 24'(148);
			21206: out = 24'(88);
			21207: out = 24'(96);
			21208: out = 24'(80);
			21209: out = 24'(108);
			21210: out = 24'(104);
			21211: out = 24'(36);
			21212: out = 24'(96);
			21213: out = 24'(68);
			21214: out = 24'(88);
			21215: out = 24'(52);
			21216: out = 24'(60);
			21217: out = 24'(96);
			21218: out = 24'(56);
			21219: out = 24'(24);
			21220: out = 24'(76);
			21221: out = 24'(32);
			21222: out = 24'(68);
			21223: out = 24'(48);
			21224: out = 24'(20);
			21225: out = 24'(84);
			21226: out = 24'(8);
			21227: out = 24'(24);
			21228: out = 24'(52);
			21229: out = 24'(36);
			21230: out = 24'(-12);
			21231: out = 24'(56);
			21232: out = 24'(16);
			21233: out = 24'(32);
			21234: out = 24'(-4);
			21235: out = 24'(12);
			21236: out = 24'(20);
			21237: out = 24'(0);
			21238: out = 24'(-12);
			21239: out = 24'(20);
			21240: out = 24'(8);
			21241: out = 24'(-24);
			21242: out = 24'(-4);
			21243: out = 24'(20);
			21244: out = 24'(-48);
			21245: out = 24'(12);
			21246: out = 24'(-32);
			21247: out = 24'(-16);
			21248: out = 24'(0);
			21249: out = 24'(-36);
			21250: out = 24'(-16);
			21251: out = 24'(-32);
			21252: out = 24'(-24);
			21253: out = 24'(-4);
			21254: out = 24'(-52);
			21255: out = 24'(-12);
			21256: out = 24'(-40);
			21257: out = 24'(-36);
			21258: out = 24'(-16);
			21259: out = 24'(-36);
			21260: out = 24'(-76);
			21261: out = 24'(-28);
			21262: out = 24'(-36);
			21263: out = 24'(-56);
			21264: out = 24'(-48);
			21265: out = 24'(-64);
			21266: out = 24'(-40);
			21267: out = 24'(-80);
			21268: out = 24'(-56);
			21269: out = 24'(-48);
			21270: out = 24'(-64);
			21271: out = 24'(-88);
			21272: out = 24'(-84);
			21273: out = 24'(-72);
			21274: out = 24'(-64);
			21275: out = 24'(-144);
			21276: out = 24'(-96);
			21277: out = 24'(-88);
			21278: out = 24'(-136);
			21279: out = 24'(-108);
			21280: out = 24'(-96);
			21281: out = 24'(-128);
			21282: out = 24'(-144);
			21283: out = 24'(-132);
			21284: out = 24'(-108);
			21285: out = 24'(-144);
			21286: out = 24'(-132);
			21287: out = 24'(-152);
			21288: out = 24'(-148);
			21289: out = 24'(-136);
			21290: out = 24'(-132);
			21291: out = 24'(-156);
			21292: out = 24'(-152);
			21293: out = 24'(-132);
			21294: out = 24'(-184);
			21295: out = 24'(-124);
			21296: out = 24'(-160);
			21297: out = 24'(-228);
			21298: out = 24'(-132);
			21299: out = 24'(-192);
			21300: out = 24'(-176);
			21301: out = 24'(-184);
			21302: out = 24'(-192);
			21303: out = 24'(-164);
			21304: out = 24'(-232);
			21305: out = 24'(-176);
			21306: out = 24'(-200);
			21307: out = 24'(-196);
			21308: out = 24'(-232);
			21309: out = 24'(-172);
			21310: out = 24'(-224);
			21311: out = 24'(-200);
			21312: out = 24'(-224);
			21313: out = 24'(-212);
			21314: out = 24'(-228);
			21315: out = 24'(-244);
			21316: out = 24'(-216);
			21317: out = 24'(-248);
			21318: out = 24'(-256);
			21319: out = 24'(-268);
			21320: out = 24'(-232);
			21321: out = 24'(-260);
			21322: out = 24'(-268);
			21323: out = 24'(-252);
			21324: out = 24'(-264);
			21325: out = 24'(-252);
			21326: out = 24'(-292);
			21327: out = 24'(-196);
			21328: out = 24'(-316);
			21329: out = 24'(-292);
			21330: out = 24'(-256);
			21331: out = 24'(-292);
			21332: out = 24'(-288);
			21333: out = 24'(-280);
			21334: out = 24'(-260);
			21335: out = 24'(-268);
			21336: out = 24'(-300);
			21337: out = 24'(-288);
			21338: out = 24'(-256);
			21339: out = 24'(-340);
			21340: out = 24'(-268);
			21341: out = 24'(-300);
			21342: out = 24'(-308);
			21343: out = 24'(-292);
			21344: out = 24'(-304);
			21345: out = 24'(-320);
			21346: out = 24'(-292);
			21347: out = 24'(-320);
			21348: out = 24'(-308);
			21349: out = 24'(-332);
			21350: out = 24'(-304);
			21351: out = 24'(-336);
			21352: out = 24'(-332);
			21353: out = 24'(-312);
			21354: out = 24'(-332);
			21355: out = 24'(-356);
			21356: out = 24'(-316);
			21357: out = 24'(-352);
			21358: out = 24'(-392);
			21359: out = 24'(-372);
			21360: out = 24'(-344);
			21361: out = 24'(-360);
			21362: out = 24'(-360);
			21363: out = 24'(-392);
			21364: out = 24'(-364);
			21365: out = 24'(-388);
			21366: out = 24'(-364);
			21367: out = 24'(-348);
			21368: out = 24'(-380);
			21369: out = 24'(-420);
			21370: out = 24'(-356);
			21371: out = 24'(-380);
			21372: out = 24'(-400);
			21373: out = 24'(-400);
			21374: out = 24'(-384);
			21375: out = 24'(-420);
			21376: out = 24'(-396);
			21377: out = 24'(-428);
			21378: out = 24'(-420);
			21379: out = 24'(-428);
			21380: out = 24'(-428);
			21381: out = 24'(-408);
			21382: out = 24'(-456);
			21383: out = 24'(-420);
			21384: out = 24'(-440);
			21385: out = 24'(-444);
			21386: out = 24'(-456);
			21387: out = 24'(-464);
			21388: out = 24'(-460);
			21389: out = 24'(-476);
			21390: out = 24'(-452);
			21391: out = 24'(-468);
			21392: out = 24'(-476);
			21393: out = 24'(-496);
			21394: out = 24'(-480);
			21395: out = 24'(-492);
			21396: out = 24'(-512);
			21397: out = 24'(-532);
			21398: out = 24'(-480);
			21399: out = 24'(-540);
			21400: out = 24'(-512);
			21401: out = 24'(-524);
			21402: out = 24'(-536);
			21403: out = 24'(-508);
			21404: out = 24'(-560);
			21405: out = 24'(-556);
			21406: out = 24'(-552);
			21407: out = 24'(-548);
			21408: out = 24'(-556);
			21409: out = 24'(-608);
			21410: out = 24'(-580);
			21411: out = 24'(-552);
			21412: out = 24'(-592);
			21413: out = 24'(-584);
			21414: out = 24'(-596);
			21415: out = 24'(-576);
			21416: out = 24'(-596);
			21417: out = 24'(-628);
			21418: out = 24'(-580);
			21419: out = 24'(-592);
			21420: out = 24'(-656);
			21421: out = 24'(-608);
			21422: out = 24'(-632);
			21423: out = 24'(-632);
			21424: out = 24'(-640);
			21425: out = 24'(-652);
			21426: out = 24'(-608);
			21427: out = 24'(-656);
			21428: out = 24'(-668);
			21429: out = 24'(-624);
			21430: out = 24'(-664);
			21431: out = 24'(-676);
			21432: out = 24'(-664);
			21433: out = 24'(-672);
			21434: out = 24'(-696);
			21435: out = 24'(-648);
			21436: out = 24'(-696);
			21437: out = 24'(-680);
			21438: out = 24'(-696);
			21439: out = 24'(-704);
			21440: out = 24'(-664);
			21441: out = 24'(-688);
			21442: out = 24'(-744);
			21443: out = 24'(-688);
			21444: out = 24'(-688);
			21445: out = 24'(-684);
			21446: out = 24'(-716);
			21447: out = 24'(-680);
			21448: out = 24'(-736);
			21449: out = 24'(-696);
			21450: out = 24'(-688);
			21451: out = 24'(-764);
			21452: out = 24'(-652);
			21453: out = 24'(-740);
			21454: out = 24'(-736);
			21455: out = 24'(-688);
			21456: out = 24'(-724);
			21457: out = 24'(-740);
			21458: out = 24'(-704);
			21459: out = 24'(-716);
			21460: out = 24'(-724);
			21461: out = 24'(-768);
			21462: out = 24'(-712);
			21463: out = 24'(-744);
			21464: out = 24'(-724);
			21465: out = 24'(-764);
			21466: out = 24'(-728);
			21467: out = 24'(-720);
			21468: out = 24'(-764);
			21469: out = 24'(-732);
			21470: out = 24'(-744);
			21471: out = 24'(-736);
			21472: out = 24'(-760);
			21473: out = 24'(-760);
			21474: out = 24'(-732);
			21475: out = 24'(-736);
			21476: out = 24'(-768);
			21477: out = 24'(-732);
			21478: out = 24'(-740);
			21479: out = 24'(-760);
			21480: out = 24'(-760);
			21481: out = 24'(-772);
			21482: out = 24'(-740);
			21483: out = 24'(-784);
			21484: out = 24'(-764);
			21485: out = 24'(-732);
			21486: out = 24'(-792);
			21487: out = 24'(-740);
			21488: out = 24'(-748);
			21489: out = 24'(-772);
			21490: out = 24'(-740);
			21491: out = 24'(-796);
			21492: out = 24'(-744);
			21493: out = 24'(-736);
			21494: out = 24'(-808);
			21495: out = 24'(-740);
			21496: out = 24'(-736);
			21497: out = 24'(-772);
			21498: out = 24'(-752);
			21499: out = 24'(-752);
			21500: out = 24'(-728);
			21501: out = 24'(-736);
			21502: out = 24'(-796);
			21503: out = 24'(-748);
			21504: out = 24'(-760);
			21505: out = 24'(-764);
			21506: out = 24'(-752);
			21507: out = 24'(-776);
			21508: out = 24'(-740);
			21509: out = 24'(-744);
			21510: out = 24'(-720);
			21511: out = 24'(-792);
			21512: out = 24'(-720);
			21513: out = 24'(-764);
			21514: out = 24'(-784);
			21515: out = 24'(-768);
			21516: out = 24'(-716);
			21517: out = 24'(-752);
			21518: out = 24'(-768);
			21519: out = 24'(-744);
			21520: out = 24'(-728);
			21521: out = 24'(-748);
			21522: out = 24'(-736);
			21523: out = 24'(-752);
			21524: out = 24'(-764);
			21525: out = 24'(-716);
			21526: out = 24'(-764);
			21527: out = 24'(-744);
			21528: out = 24'(-764);
			21529: out = 24'(-760);
			21530: out = 24'(-784);
			21531: out = 24'(-704);
			21532: out = 24'(-776);
			21533: out = 24'(-752);
			21534: out = 24'(-712);
			21535: out = 24'(-768);
			21536: out = 24'(-728);
			21537: out = 24'(-740);
			21538: out = 24'(-748);
			21539: out = 24'(-716);
			21540: out = 24'(-748);
			21541: out = 24'(-728);
			21542: out = 24'(-704);
			21543: out = 24'(-744);
			21544: out = 24'(-724);
			21545: out = 24'(-720);
			21546: out = 24'(-724);
			21547: out = 24'(-724);
			21548: out = 24'(-736);
			21549: out = 24'(-716);
			21550: out = 24'(-728);
			21551: out = 24'(-668);
			21552: out = 24'(-776);
			21553: out = 24'(-712);
			21554: out = 24'(-716);
			21555: out = 24'(-712);
			21556: out = 24'(-712);
			21557: out = 24'(-724);
			21558: out = 24'(-704);
			21559: out = 24'(-696);
			21560: out = 24'(-736);
			21561: out = 24'(-680);
			21562: out = 24'(-724);
			21563: out = 24'(-704);
			21564: out = 24'(-712);
			21565: out = 24'(-692);
			21566: out = 24'(-716);
			21567: out = 24'(-724);
			21568: out = 24'(-652);
			21569: out = 24'(-736);
			21570: out = 24'(-680);
			21571: out = 24'(-700);
			21572: out = 24'(-716);
			21573: out = 24'(-652);
			21574: out = 24'(-724);
			21575: out = 24'(-636);
			21576: out = 24'(-700);
			21577: out = 24'(-684);
			21578: out = 24'(-676);
			21579: out = 24'(-640);
			21580: out = 24'(-656);
			21581: out = 24'(-636);
			21582: out = 24'(-696);
			21583: out = 24'(-636);
			21584: out = 24'(-636);
			21585: out = 24'(-668);
			21586: out = 24'(-644);
			21587: out = 24'(-644);
			21588: out = 24'(-668);
			21589: out = 24'(-608);
			21590: out = 24'(-640);
			21591: out = 24'(-632);
			21592: out = 24'(-644);
			21593: out = 24'(-608);
			21594: out = 24'(-624);
			21595: out = 24'(-632);
			21596: out = 24'(-620);
			21597: out = 24'(-604);
			21598: out = 24'(-616);
			21599: out = 24'(-576);
			21600: out = 24'(-632);
			21601: out = 24'(-592);
			21602: out = 24'(-584);
			21603: out = 24'(-564);
			21604: out = 24'(-600);
			21605: out = 24'(-584);
			21606: out = 24'(-544);
			21607: out = 24'(-540);
			21608: out = 24'(-572);
			21609: out = 24'(-556);
			21610: out = 24'(-532);
			21611: out = 24'(-548);
			21612: out = 24'(-548);
			21613: out = 24'(-524);
			21614: out = 24'(-552);
			21615: out = 24'(-492);
			21616: out = 24'(-528);
			21617: out = 24'(-540);
			21618: out = 24'(-496);
			21619: out = 24'(-552);
			21620: out = 24'(-496);
			21621: out = 24'(-476);
			21622: out = 24'(-532);
			21623: out = 24'(-488);
			21624: out = 24'(-508);
			21625: out = 24'(-444);
			21626: out = 24'(-532);
			21627: out = 24'(-468);
			21628: out = 24'(-464);
			21629: out = 24'(-464);
			21630: out = 24'(-452);
			21631: out = 24'(-492);
			21632: out = 24'(-420);
			21633: out = 24'(-444);
			21634: out = 24'(-448);
			21635: out = 24'(-448);
			21636: out = 24'(-404);
			21637: out = 24'(-428);
			21638: out = 24'(-440);
			21639: out = 24'(-412);
			21640: out = 24'(-432);
			21641: out = 24'(-428);
			21642: out = 24'(-404);
			21643: out = 24'(-444);
			21644: out = 24'(-400);
			21645: out = 24'(-408);
			21646: out = 24'(-412);
			21647: out = 24'(-416);
			21648: out = 24'(-380);
			21649: out = 24'(-436);
			21650: out = 24'(-400);
			21651: out = 24'(-380);
			21652: out = 24'(-392);
			21653: out = 24'(-368);
			21654: out = 24'(-344);
			21655: out = 24'(-408);
			21656: out = 24'(-340);
			21657: out = 24'(-388);
			21658: out = 24'(-336);
			21659: out = 24'(-356);
			21660: out = 24'(-384);
			21661: out = 24'(-372);
			21662: out = 24'(-324);
			21663: out = 24'(-340);
			21664: out = 24'(-344);
			21665: out = 24'(-352);
			21666: out = 24'(-308);
			21667: out = 24'(-316);
			21668: out = 24'(-348);
			21669: out = 24'(-312);
			21670: out = 24'(-332);
			21671: out = 24'(-324);
			21672: out = 24'(-304);
			21673: out = 24'(-316);
			21674: out = 24'(-340);
			21675: out = 24'(-256);
			21676: out = 24'(-324);
			21677: out = 24'(-332);
			21678: out = 24'(-280);
			21679: out = 24'(-292);
			21680: out = 24'(-308);
			21681: out = 24'(-308);
			21682: out = 24'(-308);
			21683: out = 24'(-276);
			21684: out = 24'(-316);
			21685: out = 24'(-280);
			21686: out = 24'(-316);
			21687: out = 24'(-272);
			21688: out = 24'(-272);
			21689: out = 24'(-300);
			21690: out = 24'(-244);
			21691: out = 24'(-268);
			21692: out = 24'(-308);
			21693: out = 24'(-244);
			21694: out = 24'(-256);
			21695: out = 24'(-276);
			21696: out = 24'(-264);
			21697: out = 24'(-260);
			21698: out = 24'(-244);
			21699: out = 24'(-244);
			21700: out = 24'(-252);
			21701: out = 24'(-244);
			21702: out = 24'(-228);
			21703: out = 24'(-240);
			21704: out = 24'(-240);
			21705: out = 24'(-224);
			21706: out = 24'(-240);
			21707: out = 24'(-212);
			21708: out = 24'(-184);
			21709: out = 24'(-224);
			21710: out = 24'(-232);
			21711: out = 24'(-180);
			21712: out = 24'(-196);
			21713: out = 24'(-196);
			21714: out = 24'(-204);
			21715: out = 24'(-192);
			21716: out = 24'(-168);
			21717: out = 24'(-180);
			21718: out = 24'(-208);
			21719: out = 24'(-164);
			21720: out = 24'(-172);
			21721: out = 24'(-216);
			21722: out = 24'(-160);
			21723: out = 24'(-148);
			21724: out = 24'(-216);
			21725: out = 24'(-160);
			21726: out = 24'(-152);
			21727: out = 24'(-172);
			21728: out = 24'(-148);
			21729: out = 24'(-168);
			21730: out = 24'(-120);
			21731: out = 24'(-184);
			21732: out = 24'(-132);
			21733: out = 24'(-160);
			21734: out = 24'(-132);
			21735: out = 24'(-128);
			21736: out = 24'(-148);
			21737: out = 24'(-112);
			21738: out = 24'(-180);
			21739: out = 24'(-100);
			21740: out = 24'(-152);
			21741: out = 24'(-128);
			21742: out = 24'(-120);
			21743: out = 24'(-108);
			21744: out = 24'(-112);
			21745: out = 24'(-112);
			21746: out = 24'(-96);
			21747: out = 24'(-108);
			21748: out = 24'(-108);
			21749: out = 24'(-96);
			21750: out = 24'(-104);
			21751: out = 24'(-96);
			21752: out = 24'(-96);
			21753: out = 24'(-100);
			21754: out = 24'(-108);
			21755: out = 24'(-80);
			21756: out = 24'(-80);
			21757: out = 24'(-128);
			21758: out = 24'(-104);
			21759: out = 24'(-72);
			21760: out = 24'(-88);
			21761: out = 24'(-112);
			21762: out = 24'(-36);
			21763: out = 24'(-104);
			21764: out = 24'(-96);
			21765: out = 24'(-56);
			21766: out = 24'(-76);
			21767: out = 24'(-56);
			21768: out = 24'(-68);
			21769: out = 24'(-88);
			21770: out = 24'(-36);
			21771: out = 24'(-52);
			21772: out = 24'(-56);
			21773: out = 24'(-60);
			21774: out = 24'(-52);
			21775: out = 24'(-28);
			21776: out = 24'(-8);
			21777: out = 24'(-84);
			21778: out = 24'(-36);
			21779: out = 24'(-8);
			21780: out = 24'(-24);
			21781: out = 24'(-36);
			21782: out = 24'(-16);
			21783: out = 24'(-20);
			21784: out = 24'(-48);
			21785: out = 24'(0);
			default: out = 0;
		endcase
	end
endmodule
